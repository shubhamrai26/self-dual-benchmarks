module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 , y20242 , y20243 , y20244 , y20245 , y20246 , y20247 , y20248 , y20249 , y20250 , y20251 , y20252 , y20253 , y20254 , y20255 , y20256 , y20257 , y20258 , y20259 , y20260 , y20261 , y20262 , y20263 , y20264 , y20265 , y20266 , y20267 , y20268 , y20269 , y20270 , y20271 , y20272 , y20273 , y20274 , y20275 , y20276 , y20277 , y20278 , y20279 , y20280 , y20281 , y20282 , y20283 , y20284 , y20285 , y20286 , y20287 , y20288 , y20289 , y20290 , y20291 , y20292 , y20293 , y20294 , y20295 , y20296 , y20297 , y20298 , y20299 , y20300 , y20301 , y20302 , y20303 , y20304 , y20305 , y20306 , y20307 , y20308 , y20309 , y20310 , y20311 , y20312 , y20313 , y20314 , y20315 , y20316 , y20317 , y20318 , y20319 , y20320 , y20321 , y20322 , y20323 , y20324 , y20325 , y20326 , y20327 , y20328 , y20329 , y20330 , y20331 , y20332 , y20333 , y20334 , y20335 , y20336 , y20337 , y20338 , y20339 , y20340 , y20341 , y20342 , y20343 , y20344 , y20345 , y20346 , y20347 , y20348 , y20349 , y20350 , y20351 , y20352 , y20353 , y20354 , y20355 , y20356 , y20357 , y20358 , y20359 , y20360 , y20361 , y20362 , y20363 , y20364 , y20365 , y20366 , y20367 , y20368 , y20369 , y20370 , y20371 , y20372 , y20373 , y20374 , y20375 , y20376 , y20377 , y20378 , y20379 , y20380 , y20381 , y20382 , y20383 , y20384 , y20385 , y20386 , y20387 , y20388 , y20389 , y20390 , y20391 , y20392 , y20393 , y20394 , y20395 , y20396 , y20397 , y20398 , y20399 , y20400 , y20401 , y20402 , y20403 , y20404 , y20405 , y20406 , y20407 , y20408 , y20409 , y20410 , y20411 , y20412 , y20413 , y20414 , y20415 , y20416 , y20417 , y20418 , y20419 , y20420 , y20421 , y20422 , y20423 , y20424 , y20425 , y20426 , y20427 , y20428 , y20429 , y20430 , y20431 , y20432 , y20433 , y20434 , y20435 , y20436 , y20437 , y20438 , y20439 , y20440 , y20441 , y20442 , y20443 , y20444 , y20445 , y20446 , y20447 , y20448 , y20449 , y20450 , y20451 , y20452 , y20453 , y20454 , y20455 , y20456 , y20457 , y20458 , y20459 , y20460 , y20461 , y20462 , y20463 , y20464 , y20465 , y20466 , y20467 , y20468 , y20469 , y20470 , y20471 , y20472 , y20473 , y20474 , y20475 , y20476 , y20477 , y20478 , y20479 , y20480 , y20481 , y20482 , y20483 , y20484 , y20485 , y20486 , y20487 , y20488 , y20489 , y20490 , y20491 , y20492 , y20493 , y20494 , y20495 , y20496 , y20497 , y20498 , y20499 , y20500 , y20501 , y20502 , y20503 , y20504 , y20505 , y20506 , y20507 , y20508 , y20509 , y20510 , y20511 , y20512 , y20513 , y20514 , y20515 , y20516 , y20517 , y20518 , y20519 , y20520 , y20521 , y20522 , y20523 , y20524 , y20525 , y20526 , y20527 , y20528 , y20529 , y20530 , y20531 , y20532 , y20533 , y20534 , y20535 , y20536 , y20537 , y20538 , y20539 , y20540 , y20541 , y20542 , y20543 , y20544 , y20545 , y20546 , y20547 , y20548 , y20549 , y20550 , y20551 , y20552 , y20553 , y20554 , y20555 , y20556 , y20557 , y20558 , y20559 , y20560 , y20561 , y20562 , y20563 , y20564 , y20565 , y20566 , y20567 , y20568 , y20569 , y20570 , y20571 , y20572 , y20573 , y20574 , y20575 , y20576 , y20577 , y20578 , y20579 , y20580 , y20581 , y20582 , y20583 , y20584 , y20585 , y20586 , y20587 , y20588 , y20589 , y20590 , y20591 , y20592 , y20593 , y20594 , y20595 , y20596 , y20597 , y20598 , y20599 , y20600 , y20601 , y20602 , y20603 , y20604 , y20605 , y20606 , y20607 , y20608 , y20609 , y20610 , y20611 , y20612 , y20613 , y20614 , y20615 , y20616 , y20617 , y20618 , y20619 , y20620 , y20621 , y20622 , y20623 , y20624 , y20625 , y20626 , y20627 , y20628 , y20629 , y20630 , y20631 , y20632 , y20633 , y20634 , y20635 , y20636 , y20637 , y20638 , y20639 , y20640 , y20641 , y20642 , y20643 , y20644 , y20645 , y20646 , y20647 , y20648 , y20649 , y20650 , y20651 , y20652 , y20653 , y20654 , y20655 , y20656 , y20657 , y20658 , y20659 , y20660 , y20661 , y20662 , y20663 , y20664 , y20665 , y20666 , y20667 , y20668 , y20669 , y20670 , y20671 , y20672 , y20673 , y20674 , y20675 , y20676 , y20677 , y20678 , y20679 , y20680 , y20681 , y20682 , y20683 , y20684 , y20685 , y20686 , y20687 , y20688 , y20689 , y20690 , y20691 , y20692 , y20693 , y20694 , y20695 , y20696 , y20697 , y20698 , y20699 , y20700 , y20701 , y20702 , y20703 , y20704 , y20705 , y20706 , y20707 , y20708 , y20709 , y20710 , y20711 , y20712 , y20713 , y20714 , y20715 , y20716 , y20717 , y20718 , y20719 , y20720 , y20721 , y20722 , y20723 , y20724 , y20725 , y20726 , y20727 , y20728 , y20729 , y20730 , y20731 , y20732 , y20733 , y20734 , y20735 , y20736 , y20737 , y20738 , y20739 , y20740 , y20741 , y20742 , y20743 , y20744 , y20745 , y20746 , y20747 , y20748 , y20749 , y20750 , y20751 , y20752 , y20753 , y20754 , y20755 , y20756 , y20757 , y20758 , y20759 , y20760 , y20761 , y20762 , y20763 , y20764 , y20765 , y20766 , y20767 , y20768 , y20769 , y20770 , y20771 , y20772 , y20773 , y20774 , y20775 , y20776 , y20777 , y20778 , y20779 , y20780 , y20781 , y20782 , y20783 , y20784 , y20785 , y20786 , y20787 , y20788 , y20789 , y20790 , y20791 , y20792 , y20793 , y20794 , y20795 , y20796 , y20797 , y20798 , y20799 , y20800 , y20801 , y20802 , y20803 , y20804 , y20805 , y20806 , y20807 , y20808 , y20809 , y20810 , y20811 , y20812 , y20813 , y20814 , y20815 , y20816 , y20817 , y20818 , y20819 , y20820 , y20821 , y20822 , y20823 , y20824 , y20825 , y20826 , y20827 , y20828 , y20829 , y20830 , y20831 , y20832 , y20833 , y20834 , y20835 , y20836 , y20837 , y20838 , y20839 , y20840 , y20841 , y20842 , y20843 , y20844 , y20845 , y20846 , y20847 , y20848 , y20849 , y20850 , y20851 , y20852 , y20853 , y20854 , y20855 , y20856 , y20857 , y20858 , y20859 , y20860 , y20861 , y20862 , y20863 , y20864 , y20865 , y20866 , y20867 , y20868 , y20869 , y20870 , y20871 , y20872 , y20873 , y20874 , y20875 , y20876 , y20877 , y20878 , y20879 , y20880 , y20881 , y20882 , y20883 , y20884 , y20885 , y20886 , y20887 , y20888 , y20889 , y20890 , y20891 , y20892 , y20893 , y20894 , y20895 , y20896 , y20897 , y20898 , y20899 , y20900 , y20901 , y20902 , y20903 , y20904 , y20905 , y20906 , y20907 , y20908 , y20909 , y20910 , y20911 , y20912 , y20913 , y20914 , y20915 , y20916 , y20917 , y20918 , y20919 , y20920 , y20921 , y20922 , y20923 , y20924 , y20925 , y20926 , y20927 , y20928 , y20929 , y20930 , y20931 , y20932 , y20933 , y20934 , y20935 , y20936 , y20937 , y20938 , y20939 , y20940 , y20941 , y20942 , y20943 , y20944 , y20945 , y20946 , y20947 , y20948 , y20949 , y20950 , y20951 , y20952 , y20953 , y20954 , y20955 , y20956 , y20957 , y20958 , y20959 , y20960 , y20961 , y20962 , y20963 , y20964 , y20965 , y20966 , y20967 , y20968 , y20969 , y20970 , y20971 , y20972 , y20973 , y20974 , y20975 , y20976 , y20977 , y20978 , y20979 , y20980 , y20981 , y20982 , y20983 , y20984 , y20985 , y20986 , y20987 , y20988 , y20989 , y20990 , y20991 , y20992 , y20993 , y20994 , y20995 , y20996 , y20997 , y20998 , y20999 , y21000 , y21001 , y21002 , y21003 , y21004 , y21005 , y21006 , y21007 , y21008 , y21009 , y21010 , y21011 , y21012 , y21013 , y21014 , y21015 , y21016 , y21017 , y21018 , y21019 , y21020 , y21021 , y21022 , y21023 , y21024 , y21025 , y21026 , y21027 , y21028 , y21029 , y21030 , y21031 , y21032 , y21033 , y21034 , y21035 , y21036 , y21037 , y21038 , y21039 , y21040 , y21041 , y21042 , y21043 , y21044 , y21045 , y21046 , y21047 , y21048 , y21049 , y21050 , y21051 , y21052 , y21053 , y21054 , y21055 , y21056 , y21057 , y21058 , y21059 , y21060 , y21061 , y21062 , y21063 , y21064 , y21065 , y21066 , y21067 , y21068 , y21069 , y21070 , y21071 , y21072 , y21073 , y21074 , y21075 , y21076 , y21077 , y21078 , y21079 , y21080 , y21081 , y21082 , y21083 , y21084 , y21085 , y21086 , y21087 , y21088 , y21089 , y21090 , y21091 , y21092 , y21093 , y21094 , y21095 , y21096 , y21097 , y21098 , y21099 , y21100 , y21101 , y21102 , y21103 , y21104 , y21105 , y21106 , y21107 , y21108 , y21109 , y21110 , y21111 , y21112 , y21113 , y21114 , y21115 , y21116 , y21117 , y21118 , y21119 , y21120 , y21121 , y21122 , y21123 , y21124 , y21125 , y21126 , y21127 , y21128 , y21129 , y21130 , y21131 , y21132 , y21133 , y21134 , y21135 , y21136 , y21137 , y21138 , y21139 , y21140 , y21141 , y21142 , y21143 , y21144 , y21145 , y21146 , y21147 , y21148 , y21149 , y21150 , y21151 , y21152 , y21153 , y21154 , y21155 , y21156 , y21157 , y21158 , y21159 , y21160 , y21161 , y21162 , y21163 , y21164 , y21165 , y21166 , y21167 , y21168 , y21169 , y21170 , y21171 , y21172 , y21173 , y21174 , y21175 , y21176 , y21177 , y21178 , y21179 , y21180 , y21181 , y21182 , y21183 , y21184 , y21185 , y21186 , y21187 , y21188 , y21189 , y21190 , y21191 , y21192 , y21193 , y21194 , y21195 , y21196 , y21197 , y21198 , y21199 , y21200 , y21201 , y21202 , y21203 , y21204 , y21205 , y21206 , y21207 , y21208 , y21209 , y21210 , y21211 , y21212 , y21213 , y21214 , y21215 , y21216 , y21217 , y21218 , y21219 , y21220 , y21221 , y21222 , y21223 , y21224 , y21225 , y21226 , y21227 , y21228 , y21229 , y21230 , y21231 , y21232 , y21233 , y21234 , y21235 , y21236 , y21237 , y21238 , y21239 , y21240 , y21241 , y21242 , y21243 , y21244 , y21245 , y21246 , y21247 , y21248 , y21249 , y21250 , y21251 , y21252 , y21253 , y21254 , y21255 , y21256 , y21257 , y21258 , y21259 , y21260 , y21261 , y21262 , y21263 , y21264 , y21265 , y21266 , y21267 , y21268 , y21269 , y21270 , y21271 , y21272 , y21273 , y21274 , y21275 , y21276 , y21277 , y21278 , y21279 , y21280 , y21281 , y21282 , y21283 , y21284 , y21285 , y21286 , y21287 , y21288 , y21289 , y21290 , y21291 , y21292 , y21293 , y21294 , y21295 , y21296 , y21297 , y21298 , y21299 , y21300 , y21301 , y21302 , y21303 , y21304 , y21305 , y21306 , y21307 , y21308 , y21309 , y21310 , y21311 , y21312 , y21313 , y21314 , y21315 , y21316 , y21317 , y21318 , y21319 , y21320 , y21321 , y21322 , y21323 , y21324 , y21325 , y21326 , y21327 , y21328 , y21329 , y21330 , y21331 , y21332 , y21333 , y21334 , y21335 , y21336 , y21337 , y21338 , y21339 , y21340 , y21341 , y21342 , y21343 , y21344 , y21345 , y21346 , y21347 , y21348 , y21349 , y21350 , y21351 , y21352 , y21353 , y21354 , y21355 , y21356 , y21357 , y21358 , y21359 , y21360 , y21361 , y21362 , y21363 , y21364 , y21365 , y21366 , y21367 , y21368 , y21369 , y21370 , y21371 , y21372 , y21373 , y21374 , y21375 , y21376 , y21377 , y21378 , y21379 , y21380 , y21381 , y21382 , y21383 , y21384 , y21385 , y21386 , y21387 , y21388 , y21389 , y21390 , y21391 , y21392 , y21393 , y21394 , y21395 , y21396 , y21397 , y21398 , y21399 , y21400 , y21401 , y21402 , y21403 , y21404 , y21405 , y21406 , y21407 , y21408 , y21409 , y21410 , y21411 , y21412 , y21413 , y21414 , y21415 , y21416 , y21417 , y21418 , y21419 , y21420 , y21421 , y21422 , y21423 , y21424 , y21425 , y21426 , y21427 , y21428 , y21429 , y21430 , y21431 , y21432 , y21433 , y21434 , y21435 , y21436 , y21437 , y21438 , y21439 , y21440 , y21441 , y21442 , y21443 , y21444 , y21445 , y21446 , y21447 , y21448 , y21449 , y21450 , y21451 , y21452 , y21453 , y21454 , y21455 , y21456 , y21457 , y21458 , y21459 , y21460 , y21461 , y21462 , y21463 , y21464 , y21465 , y21466 , y21467 , y21468 , y21469 , y21470 , y21471 , y21472 , y21473 , y21474 , y21475 , y21476 , y21477 , y21478 , y21479 , y21480 , y21481 , y21482 , y21483 , y21484 , y21485 , y21486 , y21487 , y21488 , y21489 , y21490 , y21491 , y21492 , y21493 , y21494 , y21495 , y21496 , y21497 , y21498 , y21499 , y21500 , y21501 , y21502 , y21503 , y21504 , y21505 , y21506 , y21507 , y21508 , y21509 , y21510 , y21511 , y21512 , y21513 , y21514 , y21515 , y21516 , y21517 , y21518 , y21519 , y21520 , y21521 , y21522 , y21523 , y21524 , y21525 , y21526 , y21527 , y21528 , y21529 , y21530 , y21531 , y21532 , y21533 , y21534 , y21535 , y21536 , y21537 , y21538 , y21539 , y21540 , y21541 , y21542 , y21543 , y21544 , y21545 , y21546 , y21547 , y21548 , y21549 , y21550 , y21551 , y21552 , y21553 , y21554 , y21555 , y21556 , y21557 , y21558 , y21559 , y21560 , y21561 , y21562 , y21563 , y21564 , y21565 , y21566 , y21567 , y21568 , y21569 , y21570 , y21571 , y21572 , y21573 , y21574 , y21575 , y21576 , y21577 , y21578 , y21579 , y21580 , y21581 , y21582 , y21583 , y21584 , y21585 , y21586 , y21587 , y21588 , y21589 , y21590 , y21591 , y21592 , y21593 , y21594 , y21595 , y21596 , y21597 , y21598 , y21599 , y21600 , y21601 , y21602 , y21603 , y21604 , y21605 , y21606 , y21607 , y21608 , y21609 , y21610 , y21611 , y21612 , y21613 , y21614 , y21615 , y21616 , y21617 , y21618 , y21619 , y21620 , y21621 , y21622 , y21623 , y21624 , y21625 , y21626 , y21627 , y21628 , y21629 , y21630 , y21631 , y21632 , y21633 , y21634 , y21635 , y21636 , y21637 , y21638 , y21639 , y21640 , y21641 , y21642 , y21643 , y21644 , y21645 , y21646 , y21647 , y21648 , y21649 , y21650 , y21651 , y21652 , y21653 , y21654 , y21655 , y21656 , y21657 , y21658 , y21659 , y21660 , y21661 , y21662 , y21663 , y21664 , y21665 , y21666 , y21667 , y21668 , y21669 , y21670 , y21671 , y21672 , y21673 , y21674 , y21675 , y21676 , y21677 , y21678 , y21679 , y21680 , y21681 , y21682 , y21683 , y21684 , y21685 , y21686 , y21687 , y21688 , y21689 , y21690 , y21691 , y21692 , y21693 , y21694 , y21695 , y21696 , y21697 , y21698 , y21699 , y21700 , y21701 , y21702 , y21703 , y21704 , y21705 , y21706 , y21707 , y21708 , y21709 , y21710 , y21711 , y21712 , y21713 , y21714 , y21715 , y21716 , y21717 , y21718 , y21719 , y21720 , y21721 , y21722 , y21723 , y21724 , y21725 , y21726 , y21727 , y21728 , y21729 , y21730 , y21731 , y21732 , y21733 , y21734 , y21735 , y21736 , y21737 , y21738 , y21739 , y21740 , y21741 , y21742 , y21743 , y21744 , y21745 , y21746 , y21747 , y21748 , y21749 , y21750 , y21751 , y21752 , y21753 , y21754 , y21755 , y21756 , y21757 , y21758 , y21759 , y21760 , y21761 , y21762 , y21763 , y21764 , y21765 , y21766 , y21767 , y21768 , y21769 , y21770 , y21771 , y21772 , y21773 , y21774 , y21775 , y21776 , y21777 , y21778 , y21779 , y21780 , y21781 , y21782 , y21783 , y21784 , y21785 , y21786 , y21787 , y21788 , y21789 , y21790 , y21791 , y21792 , y21793 , y21794 , y21795 , y21796 , y21797 , y21798 , y21799 , y21800 , y21801 , y21802 , y21803 , y21804 , y21805 , y21806 , y21807 , y21808 , y21809 , y21810 , y21811 , y21812 , y21813 , y21814 , y21815 , y21816 , y21817 , y21818 , y21819 , y21820 , y21821 , y21822 , y21823 , y21824 , y21825 , y21826 , y21827 , y21828 , y21829 , y21830 , y21831 , y21832 , y21833 , y21834 , y21835 , y21836 , y21837 , y21838 , y21839 , y21840 , y21841 , y21842 , y21843 , y21844 , y21845 , y21846 , y21847 , y21848 , y21849 , y21850 , y21851 , y21852 , y21853 , y21854 , y21855 , y21856 , y21857 , y21858 , y21859 , y21860 , y21861 , y21862 , y21863 , y21864 , y21865 , y21866 , y21867 , y21868 , y21869 , y21870 , y21871 , y21872 , y21873 , y21874 , y21875 , y21876 , y21877 , y21878 , y21879 , y21880 , y21881 , y21882 , y21883 , y21884 , y21885 , y21886 , y21887 , y21888 , y21889 , y21890 , y21891 , y21892 , y21893 , y21894 , y21895 , y21896 , y21897 , y21898 , y21899 , y21900 , y21901 , y21902 , y21903 , y21904 , y21905 , y21906 , y21907 , y21908 , y21909 , y21910 , y21911 , y21912 , y21913 , y21914 , y21915 , y21916 , y21917 , y21918 , y21919 , y21920 , y21921 , y21922 , y21923 , y21924 , y21925 , y21926 , y21927 , y21928 , y21929 , y21930 , y21931 , y21932 , y21933 , y21934 , y21935 , y21936 , y21937 , y21938 , y21939 , y21940 , y21941 , y21942 , y21943 , y21944 , y21945 , y21946 , y21947 , y21948 , y21949 , y21950 , y21951 , y21952 , y21953 , y21954 , y21955 , y21956 , y21957 , y21958 , y21959 , y21960 , y21961 , y21962 , y21963 , y21964 , y21965 , y21966 , y21967 , y21968 , y21969 , y21970 , y21971 , y21972 , y21973 , y21974 , y21975 , y21976 , y21977 , y21978 , y21979 , y21980 , y21981 , y21982 , y21983 , y21984 , y21985 , y21986 , y21987 , y21988 , y21989 , y21990 , y21991 , y21992 , y21993 , y21994 , y21995 , y21996 , y21997 , y21998 , y21999 , y22000 , y22001 , y22002 , y22003 , y22004 , y22005 , y22006 , y22007 , y22008 , y22009 , y22010 , y22011 , y22012 , y22013 , y22014 , y22015 , y22016 , y22017 , y22018 , y22019 , y22020 , y22021 , y22022 , y22023 , y22024 , y22025 , y22026 , y22027 , y22028 , y22029 , y22030 , y22031 , y22032 , y22033 , y22034 , y22035 , y22036 , y22037 , y22038 , y22039 , y22040 , y22041 , y22042 , y22043 , y22044 , y22045 , y22046 , y22047 , y22048 , y22049 , y22050 , y22051 , y22052 , y22053 , y22054 , y22055 , y22056 , y22057 , y22058 , y22059 , y22060 , y22061 , y22062 , y22063 , y22064 , y22065 , y22066 , y22067 , y22068 , y22069 , y22070 , y22071 , y22072 , y22073 , y22074 , y22075 , y22076 , y22077 , y22078 , y22079 , y22080 , y22081 , y22082 , y22083 , y22084 , y22085 , y22086 , y22087 , y22088 , y22089 , y22090 , y22091 , y22092 , y22093 , y22094 , y22095 , y22096 , y22097 , y22098 , y22099 , y22100 , y22101 , y22102 , y22103 , y22104 , y22105 , y22106 , y22107 , y22108 , y22109 , y22110 , y22111 , y22112 , y22113 , y22114 , y22115 , y22116 , y22117 , y22118 , y22119 , y22120 , y22121 , y22122 , y22123 , y22124 , y22125 , y22126 , y22127 , y22128 , y22129 , y22130 , y22131 , y22132 , y22133 , y22134 , y22135 , y22136 , y22137 , y22138 , y22139 , y22140 , y22141 , y22142 , y22143 , y22144 , y22145 , y22146 , y22147 , y22148 , y22149 , y22150 , y22151 , y22152 , y22153 , y22154 , y22155 , y22156 , y22157 , y22158 , y22159 , y22160 , y22161 , y22162 , y22163 , y22164 , y22165 , y22166 , y22167 , y22168 , y22169 , y22170 , y22171 , y22172 , y22173 , y22174 , y22175 , y22176 , y22177 , y22178 , y22179 , y22180 , y22181 , y22182 , y22183 , y22184 , y22185 , y22186 , y22187 , y22188 , y22189 , y22190 , y22191 , y22192 , y22193 , y22194 , y22195 , y22196 , y22197 , y22198 , y22199 , y22200 , y22201 , y22202 , y22203 , y22204 , y22205 , y22206 , y22207 , y22208 , y22209 , y22210 , y22211 , y22212 , y22213 , y22214 , y22215 , y22216 , y22217 , y22218 , y22219 , y22220 , y22221 , y22222 , y22223 , y22224 , y22225 , y22226 , y22227 , y22228 , y22229 , y22230 , y22231 , y22232 , y22233 , y22234 , y22235 , y22236 , y22237 , y22238 , y22239 , y22240 , y22241 , y22242 , y22243 , y22244 , y22245 , y22246 , y22247 , y22248 , y22249 , y22250 , y22251 , y22252 , y22253 , y22254 , y22255 , y22256 , y22257 , y22258 , y22259 , y22260 , y22261 , y22262 , y22263 , y22264 , y22265 , y22266 , y22267 , y22268 , y22269 , y22270 , y22271 , y22272 , y22273 , y22274 , y22275 , y22276 , y22277 , y22278 , y22279 , y22280 , y22281 , y22282 , y22283 , y22284 , y22285 , y22286 , y22287 , y22288 , y22289 , y22290 , y22291 , y22292 , y22293 , y22294 , y22295 , y22296 , y22297 , y22298 , y22299 , y22300 , y22301 , y22302 , y22303 , y22304 , y22305 , y22306 , y22307 , y22308 , y22309 , y22310 , y22311 , y22312 , y22313 , y22314 , y22315 , y22316 , y22317 , y22318 , y22319 , y22320 , y22321 , y22322 , y22323 , y22324 , y22325 , y22326 , y22327 , y22328 , y22329 , y22330 , y22331 , y22332 , y22333 , y22334 , y22335 , y22336 , y22337 , y22338 , y22339 , y22340 , y22341 , y22342 , y22343 , y22344 , y22345 , y22346 , y22347 , y22348 , y22349 , y22350 , y22351 , y22352 , y22353 , y22354 , y22355 , y22356 , y22357 , y22358 , y22359 , y22360 , y22361 , y22362 , y22363 , y22364 , y22365 , y22366 , y22367 , y22368 , y22369 , y22370 , y22371 , y22372 , y22373 , y22374 , y22375 , y22376 , y22377 , y22378 , y22379 , y22380 , y22381 , y22382 , y22383 , y22384 , y22385 , y22386 , y22387 , y22388 , y22389 , y22390 , y22391 , y22392 , y22393 , y22394 , y22395 , y22396 , y22397 , y22398 , y22399 , y22400 , y22401 , y22402 , y22403 , y22404 , y22405 , y22406 , y22407 , y22408 , y22409 , y22410 , y22411 , y22412 , y22413 , y22414 , y22415 , y22416 , y22417 , y22418 , y22419 , y22420 , y22421 , y22422 , y22423 , y22424 , y22425 , y22426 , y22427 , y22428 , y22429 , y22430 , y22431 , y22432 , y22433 , y22434 , y22435 , y22436 , y22437 , y22438 , y22439 , y22440 , y22441 , y22442 , y22443 , y22444 , y22445 , y22446 , y22447 , y22448 , y22449 , y22450 , y22451 , y22452 , y22453 , y22454 , y22455 , y22456 , y22457 , y22458 , y22459 , y22460 , y22461 , y22462 , y22463 , y22464 , y22465 , y22466 , y22467 , y22468 , y22469 , y22470 , y22471 , y22472 , y22473 , y22474 , y22475 , y22476 , y22477 , y22478 , y22479 , y22480 , y22481 , y22482 , y22483 , y22484 , y22485 , y22486 , y22487 , y22488 , y22489 , y22490 , y22491 , y22492 , y22493 , y22494 , y22495 , y22496 , y22497 , y22498 , y22499 , y22500 , y22501 , y22502 , y22503 , y22504 , y22505 , y22506 , y22507 , y22508 , y22509 , y22510 , y22511 , y22512 , y22513 , y22514 , y22515 , y22516 , y22517 , y22518 , y22519 , y22520 , y22521 , y22522 , y22523 , y22524 , y22525 , y22526 , y22527 , y22528 , y22529 , y22530 , y22531 , y22532 , y22533 , y22534 , y22535 , y22536 , y22537 , y22538 , y22539 , y22540 , y22541 , y22542 , y22543 , y22544 , y22545 , y22546 , y22547 , y22548 , y22549 , y22550 , y22551 , y22552 , y22553 , y22554 , y22555 , y22556 , y22557 , y22558 , y22559 , y22560 , y22561 , y22562 , y22563 , y22564 , y22565 , y22566 , y22567 , y22568 , y22569 , y22570 , y22571 , y22572 , y22573 , y22574 , y22575 , y22576 , y22577 , y22578 , y22579 , y22580 , y22581 , y22582 , y22583 , y22584 , y22585 , y22586 , y22587 , y22588 , y22589 , y22590 , y22591 , y22592 , y22593 , y22594 , y22595 , y22596 , y22597 , y22598 , y22599 , y22600 , y22601 , y22602 , y22603 , y22604 , y22605 , y22606 , y22607 , y22608 , y22609 , y22610 , y22611 , y22612 , y22613 , y22614 , y22615 , y22616 , y22617 , y22618 , y22619 , y22620 , y22621 , y22622 , y22623 , y22624 , y22625 , y22626 , y22627 , y22628 , y22629 , y22630 , y22631 , y22632 , y22633 , y22634 , y22635 , y22636 , y22637 , y22638 , y22639 , y22640 , y22641 , y22642 , y22643 , y22644 , y22645 , y22646 , y22647 , y22648 , y22649 , y22650 , y22651 , y22652 , y22653 , y22654 , y22655 , y22656 , y22657 , y22658 , y22659 , y22660 , y22661 , y22662 , y22663 , y22664 , y22665 , y22666 , y22667 , y22668 , y22669 , y22670 , y22671 , y22672 , y22673 , y22674 , y22675 , y22676 , y22677 , y22678 , y22679 , y22680 , y22681 , y22682 , y22683 , y22684 , y22685 , y22686 , y22687 , y22688 , y22689 , y22690 , y22691 , y22692 , y22693 , y22694 , y22695 , y22696 , y22697 , y22698 , y22699 , y22700 , y22701 , y22702 , y22703 , y22704 , y22705 , y22706 , y22707 , y22708 , y22709 , y22710 , y22711 , y22712 , y22713 , y22714 , y22715 , y22716 , y22717 , y22718 , y22719 , y22720 , y22721 , y22722 , y22723 , y22724 , y22725 , y22726 , y22727 , y22728 , y22729 , y22730 , y22731 , y22732 , y22733 , y22734 , y22735 , y22736 , y22737 , y22738 , y22739 , y22740 , y22741 , y22742 , y22743 , y22744 , y22745 , y22746 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 , y20242 , y20243 , y20244 , y20245 , y20246 , y20247 , y20248 , y20249 , y20250 , y20251 , y20252 , y20253 , y20254 , y20255 , y20256 , y20257 , y20258 , y20259 , y20260 , y20261 , y20262 , y20263 , y20264 , y20265 , y20266 , y20267 , y20268 , y20269 , y20270 , y20271 , y20272 , y20273 , y20274 , y20275 , y20276 , y20277 , y20278 , y20279 , y20280 , y20281 , y20282 , y20283 , y20284 , y20285 , y20286 , y20287 , y20288 , y20289 , y20290 , y20291 , y20292 , y20293 , y20294 , y20295 , y20296 , y20297 , y20298 , y20299 , y20300 , y20301 , y20302 , y20303 , y20304 , y20305 , y20306 , y20307 , y20308 , y20309 , y20310 , y20311 , y20312 , y20313 , y20314 , y20315 , y20316 , y20317 , y20318 , y20319 , y20320 , y20321 , y20322 , y20323 , y20324 , y20325 , y20326 , y20327 , y20328 , y20329 , y20330 , y20331 , y20332 , y20333 , y20334 , y20335 , y20336 , y20337 , y20338 , y20339 , y20340 , y20341 , y20342 , y20343 , y20344 , y20345 , y20346 , y20347 , y20348 , y20349 , y20350 , y20351 , y20352 , y20353 , y20354 , y20355 , y20356 , y20357 , y20358 , y20359 , y20360 , y20361 , y20362 , y20363 , y20364 , y20365 , y20366 , y20367 , y20368 , y20369 , y20370 , y20371 , y20372 , y20373 , y20374 , y20375 , y20376 , y20377 , y20378 , y20379 , y20380 , y20381 , y20382 , y20383 , y20384 , y20385 , y20386 , y20387 , y20388 , y20389 , y20390 , y20391 , y20392 , y20393 , y20394 , y20395 , y20396 , y20397 , y20398 , y20399 , y20400 , y20401 , y20402 , y20403 , y20404 , y20405 , y20406 , y20407 , y20408 , y20409 , y20410 , y20411 , y20412 , y20413 , y20414 , y20415 , y20416 , y20417 , y20418 , y20419 , y20420 , y20421 , y20422 , y20423 , y20424 , y20425 , y20426 , y20427 , y20428 , y20429 , y20430 , y20431 , y20432 , y20433 , y20434 , y20435 , y20436 , y20437 , y20438 , y20439 , y20440 , y20441 , y20442 , y20443 , y20444 , y20445 , y20446 , y20447 , y20448 , y20449 , y20450 , y20451 , y20452 , y20453 , y20454 , y20455 , y20456 , y20457 , y20458 , y20459 , y20460 , y20461 , y20462 , y20463 , y20464 , y20465 , y20466 , y20467 , y20468 , y20469 , y20470 , y20471 , y20472 , y20473 , y20474 , y20475 , y20476 , y20477 , y20478 , y20479 , y20480 , y20481 , y20482 , y20483 , y20484 , y20485 , y20486 , y20487 , y20488 , y20489 , y20490 , y20491 , y20492 , y20493 , y20494 , y20495 , y20496 , y20497 , y20498 , y20499 , y20500 , y20501 , y20502 , y20503 , y20504 , y20505 , y20506 , y20507 , y20508 , y20509 , y20510 , y20511 , y20512 , y20513 , y20514 , y20515 , y20516 , y20517 , y20518 , y20519 , y20520 , y20521 , y20522 , y20523 , y20524 , y20525 , y20526 , y20527 , y20528 , y20529 , y20530 , y20531 , y20532 , y20533 , y20534 , y20535 , y20536 , y20537 , y20538 , y20539 , y20540 , y20541 , y20542 , y20543 , y20544 , y20545 , y20546 , y20547 , y20548 , y20549 , y20550 , y20551 , y20552 , y20553 , y20554 , y20555 , y20556 , y20557 , y20558 , y20559 , y20560 , y20561 , y20562 , y20563 , y20564 , y20565 , y20566 , y20567 , y20568 , y20569 , y20570 , y20571 , y20572 , y20573 , y20574 , y20575 , y20576 , y20577 , y20578 , y20579 , y20580 , y20581 , y20582 , y20583 , y20584 , y20585 , y20586 , y20587 , y20588 , y20589 , y20590 , y20591 , y20592 , y20593 , y20594 , y20595 , y20596 , y20597 , y20598 , y20599 , y20600 , y20601 , y20602 , y20603 , y20604 , y20605 , y20606 , y20607 , y20608 , y20609 , y20610 , y20611 , y20612 , y20613 , y20614 , y20615 , y20616 , y20617 , y20618 , y20619 , y20620 , y20621 , y20622 , y20623 , y20624 , y20625 , y20626 , y20627 , y20628 , y20629 , y20630 , y20631 , y20632 , y20633 , y20634 , y20635 , y20636 , y20637 , y20638 , y20639 , y20640 , y20641 , y20642 , y20643 , y20644 , y20645 , y20646 , y20647 , y20648 , y20649 , y20650 , y20651 , y20652 , y20653 , y20654 , y20655 , y20656 , y20657 , y20658 , y20659 , y20660 , y20661 , y20662 , y20663 , y20664 , y20665 , y20666 , y20667 , y20668 , y20669 , y20670 , y20671 , y20672 , y20673 , y20674 , y20675 , y20676 , y20677 , y20678 , y20679 , y20680 , y20681 , y20682 , y20683 , y20684 , y20685 , y20686 , y20687 , y20688 , y20689 , y20690 , y20691 , y20692 , y20693 , y20694 , y20695 , y20696 , y20697 , y20698 , y20699 , y20700 , y20701 , y20702 , y20703 , y20704 , y20705 , y20706 , y20707 , y20708 , y20709 , y20710 , y20711 , y20712 , y20713 , y20714 , y20715 , y20716 , y20717 , y20718 , y20719 , y20720 , y20721 , y20722 , y20723 , y20724 , y20725 , y20726 , y20727 , y20728 , y20729 , y20730 , y20731 , y20732 , y20733 , y20734 , y20735 , y20736 , y20737 , y20738 , y20739 , y20740 , y20741 , y20742 , y20743 , y20744 , y20745 , y20746 , y20747 , y20748 , y20749 , y20750 , y20751 , y20752 , y20753 , y20754 , y20755 , y20756 , y20757 , y20758 , y20759 , y20760 , y20761 , y20762 , y20763 , y20764 , y20765 , y20766 , y20767 , y20768 , y20769 , y20770 , y20771 , y20772 , y20773 , y20774 , y20775 , y20776 , y20777 , y20778 , y20779 , y20780 , y20781 , y20782 , y20783 , y20784 , y20785 , y20786 , y20787 , y20788 , y20789 , y20790 , y20791 , y20792 , y20793 , y20794 , y20795 , y20796 , y20797 , y20798 , y20799 , y20800 , y20801 , y20802 , y20803 , y20804 , y20805 , y20806 , y20807 , y20808 , y20809 , y20810 , y20811 , y20812 , y20813 , y20814 , y20815 , y20816 , y20817 , y20818 , y20819 , y20820 , y20821 , y20822 , y20823 , y20824 , y20825 , y20826 , y20827 , y20828 , y20829 , y20830 , y20831 , y20832 , y20833 , y20834 , y20835 , y20836 , y20837 , y20838 , y20839 , y20840 , y20841 , y20842 , y20843 , y20844 , y20845 , y20846 , y20847 , y20848 , y20849 , y20850 , y20851 , y20852 , y20853 , y20854 , y20855 , y20856 , y20857 , y20858 , y20859 , y20860 , y20861 , y20862 , y20863 , y20864 , y20865 , y20866 , y20867 , y20868 , y20869 , y20870 , y20871 , y20872 , y20873 , y20874 , y20875 , y20876 , y20877 , y20878 , y20879 , y20880 , y20881 , y20882 , y20883 , y20884 , y20885 , y20886 , y20887 , y20888 , y20889 , y20890 , y20891 , y20892 , y20893 , y20894 , y20895 , y20896 , y20897 , y20898 , y20899 , y20900 , y20901 , y20902 , y20903 , y20904 , y20905 , y20906 , y20907 , y20908 , y20909 , y20910 , y20911 , y20912 , y20913 , y20914 , y20915 , y20916 , y20917 , y20918 , y20919 , y20920 , y20921 , y20922 , y20923 , y20924 , y20925 , y20926 , y20927 , y20928 , y20929 , y20930 , y20931 , y20932 , y20933 , y20934 , y20935 , y20936 , y20937 , y20938 , y20939 , y20940 , y20941 , y20942 , y20943 , y20944 , y20945 , y20946 , y20947 , y20948 , y20949 , y20950 , y20951 , y20952 , y20953 , y20954 , y20955 , y20956 , y20957 , y20958 , y20959 , y20960 , y20961 , y20962 , y20963 , y20964 , y20965 , y20966 , y20967 , y20968 , y20969 , y20970 , y20971 , y20972 , y20973 , y20974 , y20975 , y20976 , y20977 , y20978 , y20979 , y20980 , y20981 , y20982 , y20983 , y20984 , y20985 , y20986 , y20987 , y20988 , y20989 , y20990 , y20991 , y20992 , y20993 , y20994 , y20995 , y20996 , y20997 , y20998 , y20999 , y21000 , y21001 , y21002 , y21003 , y21004 , y21005 , y21006 , y21007 , y21008 , y21009 , y21010 , y21011 , y21012 , y21013 , y21014 , y21015 , y21016 , y21017 , y21018 , y21019 , y21020 , y21021 , y21022 , y21023 , y21024 , y21025 , y21026 , y21027 , y21028 , y21029 , y21030 , y21031 , y21032 , y21033 , y21034 , y21035 , y21036 , y21037 , y21038 , y21039 , y21040 , y21041 , y21042 , y21043 , y21044 , y21045 , y21046 , y21047 , y21048 , y21049 , y21050 , y21051 , y21052 , y21053 , y21054 , y21055 , y21056 , y21057 , y21058 , y21059 , y21060 , y21061 , y21062 , y21063 , y21064 , y21065 , y21066 , y21067 , y21068 , y21069 , y21070 , y21071 , y21072 , y21073 , y21074 , y21075 , y21076 , y21077 , y21078 , y21079 , y21080 , y21081 , y21082 , y21083 , y21084 , y21085 , y21086 , y21087 , y21088 , y21089 , y21090 , y21091 , y21092 , y21093 , y21094 , y21095 , y21096 , y21097 , y21098 , y21099 , y21100 , y21101 , y21102 , y21103 , y21104 , y21105 , y21106 , y21107 , y21108 , y21109 , y21110 , y21111 , y21112 , y21113 , y21114 , y21115 , y21116 , y21117 , y21118 , y21119 , y21120 , y21121 , y21122 , y21123 , y21124 , y21125 , y21126 , y21127 , y21128 , y21129 , y21130 , y21131 , y21132 , y21133 , y21134 , y21135 , y21136 , y21137 , y21138 , y21139 , y21140 , y21141 , y21142 , y21143 , y21144 , y21145 , y21146 , y21147 , y21148 , y21149 , y21150 , y21151 , y21152 , y21153 , y21154 , y21155 , y21156 , y21157 , y21158 , y21159 , y21160 , y21161 , y21162 , y21163 , y21164 , y21165 , y21166 , y21167 , y21168 , y21169 , y21170 , y21171 , y21172 , y21173 , y21174 , y21175 , y21176 , y21177 , y21178 , y21179 , y21180 , y21181 , y21182 , y21183 , y21184 , y21185 , y21186 , y21187 , y21188 , y21189 , y21190 , y21191 , y21192 , y21193 , y21194 , y21195 , y21196 , y21197 , y21198 , y21199 , y21200 , y21201 , y21202 , y21203 , y21204 , y21205 , y21206 , y21207 , y21208 , y21209 , y21210 , y21211 , y21212 , y21213 , y21214 , y21215 , y21216 , y21217 , y21218 , y21219 , y21220 , y21221 , y21222 , y21223 , y21224 , y21225 , y21226 , y21227 , y21228 , y21229 , y21230 , y21231 , y21232 , y21233 , y21234 , y21235 , y21236 , y21237 , y21238 , y21239 , y21240 , y21241 , y21242 , y21243 , y21244 , y21245 , y21246 , y21247 , y21248 , y21249 , y21250 , y21251 , y21252 , y21253 , y21254 , y21255 , y21256 , y21257 , y21258 , y21259 , y21260 , y21261 , y21262 , y21263 , y21264 , y21265 , y21266 , y21267 , y21268 , y21269 , y21270 , y21271 , y21272 , y21273 , y21274 , y21275 , y21276 , y21277 , y21278 , y21279 , y21280 , y21281 , y21282 , y21283 , y21284 , y21285 , y21286 , y21287 , y21288 , y21289 , y21290 , y21291 , y21292 , y21293 , y21294 , y21295 , y21296 , y21297 , y21298 , y21299 , y21300 , y21301 , y21302 , y21303 , y21304 , y21305 , y21306 , y21307 , y21308 , y21309 , y21310 , y21311 , y21312 , y21313 , y21314 , y21315 , y21316 , y21317 , y21318 , y21319 , y21320 , y21321 , y21322 , y21323 , y21324 , y21325 , y21326 , y21327 , y21328 , y21329 , y21330 , y21331 , y21332 , y21333 , y21334 , y21335 , y21336 , y21337 , y21338 , y21339 , y21340 , y21341 , y21342 , y21343 , y21344 , y21345 , y21346 , y21347 , y21348 , y21349 , y21350 , y21351 , y21352 , y21353 , y21354 , y21355 , y21356 , y21357 , y21358 , y21359 , y21360 , y21361 , y21362 , y21363 , y21364 , y21365 , y21366 , y21367 , y21368 , y21369 , y21370 , y21371 , y21372 , y21373 , y21374 , y21375 , y21376 , y21377 , y21378 , y21379 , y21380 , y21381 , y21382 , y21383 , y21384 , y21385 , y21386 , y21387 , y21388 , y21389 , y21390 , y21391 , y21392 , y21393 , y21394 , y21395 , y21396 , y21397 , y21398 , y21399 , y21400 , y21401 , y21402 , y21403 , y21404 , y21405 , y21406 , y21407 , y21408 , y21409 , y21410 , y21411 , y21412 , y21413 , y21414 , y21415 , y21416 , y21417 , y21418 , y21419 , y21420 , y21421 , y21422 , y21423 , y21424 , y21425 , y21426 , y21427 , y21428 , y21429 , y21430 , y21431 , y21432 , y21433 , y21434 , y21435 , y21436 , y21437 , y21438 , y21439 , y21440 , y21441 , y21442 , y21443 , y21444 , y21445 , y21446 , y21447 , y21448 , y21449 , y21450 , y21451 , y21452 , y21453 , y21454 , y21455 , y21456 , y21457 , y21458 , y21459 , y21460 , y21461 , y21462 , y21463 , y21464 , y21465 , y21466 , y21467 , y21468 , y21469 , y21470 , y21471 , y21472 , y21473 , y21474 , y21475 , y21476 , y21477 , y21478 , y21479 , y21480 , y21481 , y21482 , y21483 , y21484 , y21485 , y21486 , y21487 , y21488 , y21489 , y21490 , y21491 , y21492 , y21493 , y21494 , y21495 , y21496 , y21497 , y21498 , y21499 , y21500 , y21501 , y21502 , y21503 , y21504 , y21505 , y21506 , y21507 , y21508 , y21509 , y21510 , y21511 , y21512 , y21513 , y21514 , y21515 , y21516 , y21517 , y21518 , y21519 , y21520 , y21521 , y21522 , y21523 , y21524 , y21525 , y21526 , y21527 , y21528 , y21529 , y21530 , y21531 , y21532 , y21533 , y21534 , y21535 , y21536 , y21537 , y21538 , y21539 , y21540 , y21541 , y21542 , y21543 , y21544 , y21545 , y21546 , y21547 , y21548 , y21549 , y21550 , y21551 , y21552 , y21553 , y21554 , y21555 , y21556 , y21557 , y21558 , y21559 , y21560 , y21561 , y21562 , y21563 , y21564 , y21565 , y21566 , y21567 , y21568 , y21569 , y21570 , y21571 , y21572 , y21573 , y21574 , y21575 , y21576 , y21577 , y21578 , y21579 , y21580 , y21581 , y21582 , y21583 , y21584 , y21585 , y21586 , y21587 , y21588 , y21589 , y21590 , y21591 , y21592 , y21593 , y21594 , y21595 , y21596 , y21597 , y21598 , y21599 , y21600 , y21601 , y21602 , y21603 , y21604 , y21605 , y21606 , y21607 , y21608 , y21609 , y21610 , y21611 , y21612 , y21613 , y21614 , y21615 , y21616 , y21617 , y21618 , y21619 , y21620 , y21621 , y21622 , y21623 , y21624 , y21625 , y21626 , y21627 , y21628 , y21629 , y21630 , y21631 , y21632 , y21633 , y21634 , y21635 , y21636 , y21637 , y21638 , y21639 , y21640 , y21641 , y21642 , y21643 , y21644 , y21645 , y21646 , y21647 , y21648 , y21649 , y21650 , y21651 , y21652 , y21653 , y21654 , y21655 , y21656 , y21657 , y21658 , y21659 , y21660 , y21661 , y21662 , y21663 , y21664 , y21665 , y21666 , y21667 , y21668 , y21669 , y21670 , y21671 , y21672 , y21673 , y21674 , y21675 , y21676 , y21677 , y21678 , y21679 , y21680 , y21681 , y21682 , y21683 , y21684 , y21685 , y21686 , y21687 , y21688 , y21689 , y21690 , y21691 , y21692 , y21693 , y21694 , y21695 , y21696 , y21697 , y21698 , y21699 , y21700 , y21701 , y21702 , y21703 , y21704 , y21705 , y21706 , y21707 , y21708 , y21709 , y21710 , y21711 , y21712 , y21713 , y21714 , y21715 , y21716 , y21717 , y21718 , y21719 , y21720 , y21721 , y21722 , y21723 , y21724 , y21725 , y21726 , y21727 , y21728 , y21729 , y21730 , y21731 , y21732 , y21733 , y21734 , y21735 , y21736 , y21737 , y21738 , y21739 , y21740 , y21741 , y21742 , y21743 , y21744 , y21745 , y21746 , y21747 , y21748 , y21749 , y21750 , y21751 , y21752 , y21753 , y21754 , y21755 , y21756 , y21757 , y21758 , y21759 , y21760 , y21761 , y21762 , y21763 , y21764 , y21765 , y21766 , y21767 , y21768 , y21769 , y21770 , y21771 , y21772 , y21773 , y21774 , y21775 , y21776 , y21777 , y21778 , y21779 , y21780 , y21781 , y21782 , y21783 , y21784 , y21785 , y21786 , y21787 , y21788 , y21789 , y21790 , y21791 , y21792 , y21793 , y21794 , y21795 , y21796 , y21797 , y21798 , y21799 , y21800 , y21801 , y21802 , y21803 , y21804 , y21805 , y21806 , y21807 , y21808 , y21809 , y21810 , y21811 , y21812 , y21813 , y21814 , y21815 , y21816 , y21817 , y21818 , y21819 , y21820 , y21821 , y21822 , y21823 , y21824 , y21825 , y21826 , y21827 , y21828 , y21829 , y21830 , y21831 , y21832 , y21833 , y21834 , y21835 , y21836 , y21837 , y21838 , y21839 , y21840 , y21841 , y21842 , y21843 , y21844 , y21845 , y21846 , y21847 , y21848 , y21849 , y21850 , y21851 , y21852 , y21853 , y21854 , y21855 , y21856 , y21857 , y21858 , y21859 , y21860 , y21861 , y21862 , y21863 , y21864 , y21865 , y21866 , y21867 , y21868 , y21869 , y21870 , y21871 , y21872 , y21873 , y21874 , y21875 , y21876 , y21877 , y21878 , y21879 , y21880 , y21881 , y21882 , y21883 , y21884 , y21885 , y21886 , y21887 , y21888 , y21889 , y21890 , y21891 , y21892 , y21893 , y21894 , y21895 , y21896 , y21897 , y21898 , y21899 , y21900 , y21901 , y21902 , y21903 , y21904 , y21905 , y21906 , y21907 , y21908 , y21909 , y21910 , y21911 , y21912 , y21913 , y21914 , y21915 , y21916 , y21917 , y21918 , y21919 , y21920 , y21921 , y21922 , y21923 , y21924 , y21925 , y21926 , y21927 , y21928 , y21929 , y21930 , y21931 , y21932 , y21933 , y21934 , y21935 , y21936 , y21937 , y21938 , y21939 , y21940 , y21941 , y21942 , y21943 , y21944 , y21945 , y21946 , y21947 , y21948 , y21949 , y21950 , y21951 , y21952 , y21953 , y21954 , y21955 , y21956 , y21957 , y21958 , y21959 , y21960 , y21961 , y21962 , y21963 , y21964 , y21965 , y21966 , y21967 , y21968 , y21969 , y21970 , y21971 , y21972 , y21973 , y21974 , y21975 , y21976 , y21977 , y21978 , y21979 , y21980 , y21981 , y21982 , y21983 , y21984 , y21985 , y21986 , y21987 , y21988 , y21989 , y21990 , y21991 , y21992 , y21993 , y21994 , y21995 , y21996 , y21997 , y21998 , y21999 , y22000 , y22001 , y22002 , y22003 , y22004 , y22005 , y22006 , y22007 , y22008 , y22009 , y22010 , y22011 , y22012 , y22013 , y22014 , y22015 , y22016 , y22017 , y22018 , y22019 , y22020 , y22021 , y22022 , y22023 , y22024 , y22025 , y22026 , y22027 , y22028 , y22029 , y22030 , y22031 , y22032 , y22033 , y22034 , y22035 , y22036 , y22037 , y22038 , y22039 , y22040 , y22041 , y22042 , y22043 , y22044 , y22045 , y22046 , y22047 , y22048 , y22049 , y22050 , y22051 , y22052 , y22053 , y22054 , y22055 , y22056 , y22057 , y22058 , y22059 , y22060 , y22061 , y22062 , y22063 , y22064 , y22065 , y22066 , y22067 , y22068 , y22069 , y22070 , y22071 , y22072 , y22073 , y22074 , y22075 , y22076 , y22077 , y22078 , y22079 , y22080 , y22081 , y22082 , y22083 , y22084 , y22085 , y22086 , y22087 , y22088 , y22089 , y22090 , y22091 , y22092 , y22093 , y22094 , y22095 , y22096 , y22097 , y22098 , y22099 , y22100 , y22101 , y22102 , y22103 , y22104 , y22105 , y22106 , y22107 , y22108 , y22109 , y22110 , y22111 , y22112 , y22113 , y22114 , y22115 , y22116 , y22117 , y22118 , y22119 , y22120 , y22121 , y22122 , y22123 , y22124 , y22125 , y22126 , y22127 , y22128 , y22129 , y22130 , y22131 , y22132 , y22133 , y22134 , y22135 , y22136 , y22137 , y22138 , y22139 , y22140 , y22141 , y22142 , y22143 , y22144 , y22145 , y22146 , y22147 , y22148 , y22149 , y22150 , y22151 , y22152 , y22153 , y22154 , y22155 , y22156 , y22157 , y22158 , y22159 , y22160 , y22161 , y22162 , y22163 , y22164 , y22165 , y22166 , y22167 , y22168 , y22169 , y22170 , y22171 , y22172 , y22173 , y22174 , y22175 , y22176 , y22177 , y22178 , y22179 , y22180 , y22181 , y22182 , y22183 , y22184 , y22185 , y22186 , y22187 , y22188 , y22189 , y22190 , y22191 , y22192 , y22193 , y22194 , y22195 , y22196 , y22197 , y22198 , y22199 , y22200 , y22201 , y22202 , y22203 , y22204 , y22205 , y22206 , y22207 , y22208 , y22209 , y22210 , y22211 , y22212 , y22213 , y22214 , y22215 , y22216 , y22217 , y22218 , y22219 , y22220 , y22221 , y22222 , y22223 , y22224 , y22225 , y22226 , y22227 , y22228 , y22229 , y22230 , y22231 , y22232 , y22233 , y22234 , y22235 , y22236 , y22237 , y22238 , y22239 , y22240 , y22241 , y22242 , y22243 , y22244 , y22245 , y22246 , y22247 , y22248 , y22249 , y22250 , y22251 , y22252 , y22253 , y22254 , y22255 , y22256 , y22257 , y22258 , y22259 , y22260 , y22261 , y22262 , y22263 , y22264 , y22265 , y22266 , y22267 , y22268 , y22269 , y22270 , y22271 , y22272 , y22273 , y22274 , y22275 , y22276 , y22277 , y22278 , y22279 , y22280 , y22281 , y22282 , y22283 , y22284 , y22285 , y22286 , y22287 , y22288 , y22289 , y22290 , y22291 , y22292 , y22293 , y22294 , y22295 , y22296 , y22297 , y22298 , y22299 , y22300 , y22301 , y22302 , y22303 , y22304 , y22305 , y22306 , y22307 , y22308 , y22309 , y22310 , y22311 , y22312 , y22313 , y22314 , y22315 , y22316 , y22317 , y22318 , y22319 , y22320 , y22321 , y22322 , y22323 , y22324 , y22325 , y22326 , y22327 , y22328 , y22329 , y22330 , y22331 , y22332 , y22333 , y22334 , y22335 , y22336 , y22337 , y22338 , y22339 , y22340 , y22341 , y22342 , y22343 , y22344 , y22345 , y22346 , y22347 , y22348 , y22349 , y22350 , y22351 , y22352 , y22353 , y22354 , y22355 , y22356 , y22357 , y22358 , y22359 , y22360 , y22361 , y22362 , y22363 , y22364 , y22365 , y22366 , y22367 , y22368 , y22369 , y22370 , y22371 , y22372 , y22373 , y22374 , y22375 , y22376 , y22377 , y22378 , y22379 , y22380 , y22381 , y22382 , y22383 , y22384 , y22385 , y22386 , y22387 , y22388 , y22389 , y22390 , y22391 , y22392 , y22393 , y22394 , y22395 , y22396 , y22397 , y22398 , y22399 , y22400 , y22401 , y22402 , y22403 , y22404 , y22405 , y22406 , y22407 , y22408 , y22409 , y22410 , y22411 , y22412 , y22413 , y22414 , y22415 , y22416 , y22417 , y22418 , y22419 , y22420 , y22421 , y22422 , y22423 , y22424 , y22425 , y22426 , y22427 , y22428 , y22429 , y22430 , y22431 , y22432 , y22433 , y22434 , y22435 , y22436 , y22437 , y22438 , y22439 , y22440 , y22441 , y22442 , y22443 , y22444 , y22445 , y22446 , y22447 , y22448 , y22449 , y22450 , y22451 , y22452 , y22453 , y22454 , y22455 , y22456 , y22457 , y22458 , y22459 , y22460 , y22461 , y22462 , y22463 , y22464 , y22465 , y22466 , y22467 , y22468 , y22469 , y22470 , y22471 , y22472 , y22473 , y22474 , y22475 , y22476 , y22477 , y22478 , y22479 , y22480 , y22481 , y22482 , y22483 , y22484 , y22485 , y22486 , y22487 , y22488 , y22489 , y22490 , y22491 , y22492 , y22493 , y22494 , y22495 , y22496 , y22497 , y22498 , y22499 , y22500 , y22501 , y22502 , y22503 , y22504 , y22505 , y22506 , y22507 , y22508 , y22509 , y22510 , y22511 , y22512 , y22513 , y22514 , y22515 , y22516 , y22517 , y22518 , y22519 , y22520 , y22521 , y22522 , y22523 , y22524 , y22525 , y22526 , y22527 , y22528 , y22529 , y22530 , y22531 , y22532 , y22533 , y22534 , y22535 , y22536 , y22537 , y22538 , y22539 , y22540 , y22541 , y22542 , y22543 , y22544 , y22545 , y22546 , y22547 , y22548 , y22549 , y22550 , y22551 , y22552 , y22553 , y22554 , y22555 , y22556 , y22557 , y22558 , y22559 , y22560 , y22561 , y22562 , y22563 , y22564 , y22565 , y22566 , y22567 , y22568 , y22569 , y22570 , y22571 , y22572 , y22573 , y22574 , y22575 , y22576 , y22577 , y22578 , y22579 , y22580 , y22581 , y22582 , y22583 , y22584 , y22585 , y22586 , y22587 , y22588 , y22589 , y22590 , y22591 , y22592 , y22593 , y22594 , y22595 , y22596 , y22597 , y22598 , y22599 , y22600 , y22601 , y22602 , y22603 , y22604 , y22605 , y22606 , y22607 , y22608 , y22609 , y22610 , y22611 , y22612 , y22613 , y22614 , y22615 , y22616 , y22617 , y22618 , y22619 , y22620 , y22621 , y22622 , y22623 , y22624 , y22625 , y22626 , y22627 , y22628 , y22629 , y22630 , y22631 , y22632 , y22633 , y22634 , y22635 , y22636 , y22637 , y22638 , y22639 , y22640 , y22641 , y22642 , y22643 , y22644 , y22645 , y22646 , y22647 , y22648 , y22649 , y22650 , y22651 , y22652 , y22653 , y22654 , y22655 , y22656 , y22657 , y22658 , y22659 , y22660 , y22661 , y22662 , y22663 , y22664 , y22665 , y22666 , y22667 , y22668 , y22669 , y22670 , y22671 , y22672 , y22673 , y22674 , y22675 , y22676 , y22677 , y22678 , y22679 , y22680 , y22681 , y22682 , y22683 , y22684 , y22685 , y22686 , y22687 , y22688 , y22689 , y22690 , y22691 , y22692 , y22693 , y22694 , y22695 , y22696 , y22697 , y22698 , y22699 , y22700 , y22701 , y22702 , y22703 , y22704 , y22705 , y22706 , y22707 , y22708 , y22709 , y22710 , y22711 , y22712 , y22713 , y22714 , y22715 , y22716 , y22717 , y22718 , y22719 , y22720 , y22721 , y22722 , y22723 , y22724 , y22725 , y22726 , y22727 , y22728 , y22729 , y22730 , y22731 , y22732 , y22733 , y22734 , y22735 , y22736 , y22737 , y22738 , y22739 , y22740 , y22741 , y22742 , y22743 , y22744 , y22745 , y22746 ;
  wire n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 ;
  assign n256 = ( x14 & ~x67 ) | ( x14 & x145 ) | ( ~x67 & x145 ) ;
  assign n257 = x145 & x183 ;
  assign n258 = ~x14 & n257 ;
  assign n259 = ( x42 & x253 ) | ( x42 & ~x254 ) | ( x253 & ~x254 ) ;
  assign n260 = x123 & x162 ;
  assign n261 = ~x111 & n260 ;
  assign n262 = x39 & x203 ;
  assign n263 = n261 & n262 ;
  assign n264 = x234 ^ x63 ^ 1'b0 ;
  assign n265 = x63 & n264 ;
  assign n266 = x48 & x163 ;
  assign n267 = ~x102 & n266 ;
  assign n268 = x153 ^ x140 ^ 1'b0 ;
  assign n269 = x17 & n268 ;
  assign n270 = x170 ^ x47 ^ 1'b0 ;
  assign n271 = x70 & n270 ;
  assign n272 = x69 & n271 ;
  assign n273 = ~x77 & n272 ;
  assign n274 = ( x34 & x131 ) | ( x34 & ~x157 ) | ( x131 & ~x157 ) ;
  assign n275 = ( x11 & ~x213 ) | ( x11 & n274 ) | ( ~x213 & n274 ) ;
  assign n276 = x200 ^ x48 ^ 1'b0 ;
  assign n277 = x226 & n276 ;
  assign n278 = x60 & x232 ;
  assign n279 = n278 ^ x136 ^ 1'b0 ;
  assign n280 = x91 ^ x50 ^ 1'b0 ;
  assign n281 = x141 & n280 ;
  assign n282 = x89 & x233 ;
  assign n283 = ~x237 & n282 ;
  assign n284 = ( x46 & x128 ) | ( x46 & ~x140 ) | ( x128 & ~x140 ) ;
  assign n285 = x116 & n284 ;
  assign n286 = n285 ^ x113 ^ 1'b0 ;
  assign n287 = x138 & x158 ;
  assign n288 = ~x238 & n287 ;
  assign n289 = ( x37 & x192 ) | ( x37 & ~x212 ) | ( x192 & ~x212 ) ;
  assign n290 = x53 & x113 ;
  assign n291 = ~x114 & n290 ;
  assign n292 = x12 & ~x101 ;
  assign n293 = x212 & x233 ;
  assign n294 = n293 ^ x66 ^ 1'b0 ;
  assign n295 = x13 & x30 ;
  assign n296 = ~x134 & n295 ;
  assign n297 = x32 & x36 ;
  assign n298 = n297 ^ x168 ^ 1'b0 ;
  assign n299 = ( x143 & ~n296 ) | ( x143 & n298 ) | ( ~n296 & n298 ) ;
  assign n300 = n289 ^ x202 ^ x41 ;
  assign n301 = x176 & ~x187 ;
  assign n302 = x188 ^ x172 ^ 1'b0 ;
  assign n303 = x93 & x114 ;
  assign n304 = ~x197 & n303 ;
  assign n305 = x183 ^ x92 ^ x29 ;
  assign n306 = ( ~x10 & x165 ) | ( ~x10 & x216 ) | ( x165 & x216 ) ;
  assign n307 = x116 & x141 ;
  assign n310 = x176 ^ x103 ^ 1'b0 ;
  assign n311 = x237 & n310 ;
  assign n309 = x48 & x130 ;
  assign n312 = n311 ^ n309 ^ 1'b0 ;
  assign n308 = x133 & ~n274 ;
  assign n313 = n312 ^ n308 ^ 1'b0 ;
  assign n314 = x59 & n313 ;
  assign n315 = x188 ^ x127 ^ x87 ;
  assign n316 = x193 & ~n267 ;
  assign n317 = n316 ^ x22 ^ 1'b0 ;
  assign n318 = x165 & ~n317 ;
  assign n319 = n318 ^ x161 ^ 1'b0 ;
  assign n320 = n283 ^ x122 ^ 1'b0 ;
  assign n321 = x11 & n314 ;
  assign n322 = ~x123 & n321 ;
  assign n323 = x222 ^ x174 ^ x54 ;
  assign n325 = x193 & x198 ;
  assign n326 = n325 ^ x173 ^ 1'b0 ;
  assign n327 = n326 ^ x83 ^ x61 ;
  assign n324 = x154 & x214 ;
  assign n328 = n327 ^ n324 ^ 1'b0 ;
  assign n329 = ( x173 & ~x175 ) | ( x173 & n317 ) | ( ~x175 & n317 ) ;
  assign n330 = x0 & ~n329 ;
  assign n331 = ~x206 & n330 ;
  assign n332 = n305 ^ x235 ^ x8 ;
  assign n333 = n312 ^ n279 ^ x24 ;
  assign n334 = x156 & x243 ;
  assign n335 = n334 ^ x220 ^ 1'b0 ;
  assign n336 = x18 & ~n267 ;
  assign n337 = n336 ^ x238 ^ 1'b0 ;
  assign n338 = n337 ^ x159 ^ 1'b0 ;
  assign n340 = ( x55 & x102 ) | ( x55 & ~x166 ) | ( x102 & ~x166 ) ;
  assign n339 = x16 & x35 ;
  assign n341 = n340 ^ n339 ^ 1'b0 ;
  assign n342 = n341 ^ x221 ^ x190 ;
  assign n343 = x118 ^ x29 ^ 1'b0 ;
  assign n344 = x244 & n343 ;
  assign n345 = ( ~x49 & x67 ) | ( ~x49 & x73 ) | ( x67 & x73 ) ;
  assign n346 = x59 ^ x57 ^ 1'b0 ;
  assign n347 = n345 & n346 ;
  assign n348 = x235 & n347 ;
  assign n349 = ~n344 & n348 ;
  assign n350 = x47 & ~n308 ;
  assign n351 = ~x195 & n350 ;
  assign n353 = ( ~x58 & x122 ) | ( ~x58 & x142 ) | ( x122 & x142 ) ;
  assign n352 = x103 & n345 ;
  assign n354 = n353 ^ n352 ^ 1'b0 ;
  assign n359 = x248 ^ x204 ^ 1'b0 ;
  assign n360 = x244 & n359 ;
  assign n356 = x24 & x252 ;
  assign n357 = n356 ^ x210 ^ 1'b0 ;
  assign n355 = x244 & ~n315 ;
  assign n358 = n357 ^ n355 ^ 1'b0 ;
  assign n361 = n360 ^ n358 ^ x199 ;
  assign n362 = x190 & x211 ;
  assign n363 = ~x109 & n362 ;
  assign n364 = n265 & n344 ;
  assign n365 = n363 & n364 ;
  assign n366 = ( x33 & ~x89 ) | ( x33 & n365 ) | ( ~x89 & n365 ) ;
  assign n367 = x242 ^ x198 ^ x166 ;
  assign n368 = x191 & ~n367 ;
  assign n369 = ~n360 & n368 ;
  assign n370 = x237 & ~n369 ;
  assign n371 = ~x165 & n370 ;
  assign n372 = ( x61 & ~x72 ) | ( x61 & x239 ) | ( ~x72 & x239 ) ;
  assign n373 = x130 & ~n296 ;
  assign n374 = ~x126 & n373 ;
  assign n375 = n340 & ~n374 ;
  assign n376 = ~n372 & n375 ;
  assign n377 = ( ~x96 & x117 ) | ( ~x96 & n376 ) | ( x117 & n376 ) ;
  assign n378 = x64 & x213 ;
  assign n379 = ~x129 & n378 ;
  assign n380 = n379 ^ x78 ^ x61 ;
  assign n381 = n365 ^ n349 ^ x232 ;
  assign n390 = n269 ^ x71 ^ x46 ;
  assign n391 = n390 ^ x144 ^ 1'b0 ;
  assign n392 = x222 & ~n391 ;
  assign n386 = x24 & x143 ;
  assign n387 = ~x111 & n386 ;
  assign n382 = x245 ^ x238 ^ 1'b0 ;
  assign n383 = x212 & n382 ;
  assign n384 = x137 & n383 ;
  assign n385 = n384 ^ n304 ^ 1'b0 ;
  assign n388 = n387 ^ n385 ^ x56 ;
  assign n389 = x91 & n388 ;
  assign n393 = n392 ^ n389 ^ 1'b0 ;
  assign n394 = n353 ^ x135 ^ 1'b0 ;
  assign n395 = x229 & n394 ;
  assign n396 = x76 ^ x41 ^ 1'b0 ;
  assign n397 = ~n393 & n396 ;
  assign n398 = x30 & x146 ;
  assign n399 = n398 ^ n335 ^ 1'b0 ;
  assign n400 = ( ~x42 & x91 ) | ( ~x42 & n335 ) | ( x91 & n335 ) ;
  assign n401 = n347 ^ x252 ^ 1'b0 ;
  assign n402 = x150 ^ x33 ^ x12 ;
  assign n403 = x186 & ~n312 ;
  assign n404 = n403 ^ x197 ^ 1'b0 ;
  assign n405 = ( ~x146 & x159 ) | ( ~x146 & n404 ) | ( x159 & n404 ) ;
  assign n406 = x40 & x49 ;
  assign n407 = ~x63 & n406 ;
  assign n408 = x148 & x157 ;
  assign n409 = n407 & n408 ;
  assign n410 = x56 ^ x30 ^ 1'b0 ;
  assign n411 = ~x171 & n410 ;
  assign n412 = n411 ^ x212 ^ 1'b0 ;
  assign n413 = ~x29 & x198 ;
  assign n414 = x62 & n413 ;
  assign n415 = n414 ^ x30 ^ 1'b0 ;
  assign n416 = x41 & x238 ;
  assign n417 = ~x189 & n416 ;
  assign n418 = x83 & ~n289 ;
  assign n419 = x122 & x127 ;
  assign n420 = ~x99 & n419 ;
  assign n423 = x227 ^ x140 ^ x35 ;
  assign n424 = x39 & ~n423 ;
  assign n425 = n424 ^ x23 ^ 1'b0 ;
  assign n426 = x145 & ~n425 ;
  assign n427 = n426 ^ n320 ^ 1'b0 ;
  assign n422 = x164 & ~n322 ;
  assign n428 = n427 ^ n422 ^ 1'b0 ;
  assign n421 = n347 & ~n367 ;
  assign n429 = n428 ^ n421 ^ 1'b0 ;
  assign n430 = x10 & n429 ;
  assign n431 = n420 & n430 ;
  assign n432 = n267 | n335 ;
  assign n433 = x248 & n344 ;
  assign n434 = ( ~x159 & x224 ) | ( ~x159 & n404 ) | ( x224 & n404 ) ;
  assign n435 = x103 & x127 ;
  assign n436 = n435 ^ x198 ^ 1'b0 ;
  assign n437 = x3 & x84 ;
  assign n438 = ~x13 & n437 ;
  assign n439 = ( x138 & ~x225 ) | ( x138 & n425 ) | ( ~x225 & n425 ) ;
  assign n440 = n438 | n439 ;
  assign n441 = n440 ^ x157 ^ 1'b0 ;
  assign n442 = n271 ^ x144 ^ 1'b0 ;
  assign n443 = ~n387 & n442 ;
  assign n444 = x59 ^ x31 ^ x29 ;
  assign n445 = n444 ^ x63 ^ x11 ;
  assign n446 = ( x214 & ~n443 ) | ( x214 & n445 ) | ( ~n443 & n445 ) ;
  assign n447 = x146 ^ x56 ^ 1'b0 ;
  assign n448 = x138 ^ x51 ^ 1'b0 ;
  assign n449 = x67 & n448 ;
  assign n450 = n274 & ~n425 ;
  assign n451 = n450 ^ x115 ^ 1'b0 ;
  assign n452 = x248 & ~n451 ;
  assign n453 = ~n449 & n452 ;
  assign n454 = x76 & x180 ;
  assign n455 = ~x54 & n454 ;
  assign n456 = ( x130 & x208 ) | ( x130 & n455 ) | ( x208 & n455 ) ;
  assign n458 = ( ~x95 & x109 ) | ( ~x95 & n322 ) | ( x109 & n322 ) ;
  assign n457 = x145 & x247 ;
  assign n459 = n458 ^ n457 ^ 1'b0 ;
  assign n460 = n363 ^ x50 ^ 1'b0 ;
  assign n461 = x158 ^ x48 ^ 1'b0 ;
  assign n462 = n385 & n461 ;
  assign n463 = n288 ^ x221 ^ 1'b0 ;
  assign n464 = x239 & ~n357 ;
  assign n465 = n464 ^ x110 ^ 1'b0 ;
  assign n466 = x240 & ~n465 ;
  assign n467 = n466 ^ x215 ^ 1'b0 ;
  assign n468 = n279 ^ x243 ^ 1'b0 ;
  assign n469 = n256 & ~n468 ;
  assign n470 = n326 ^ x69 ^ 1'b0 ;
  assign n471 = x131 & ~n470 ;
  assign n472 = ( x122 & x247 ) | ( x122 & ~x254 ) | ( x247 & ~x254 ) ;
  assign n473 = ( x74 & x151 ) | ( x74 & ~n472 ) | ( x151 & ~n472 ) ;
  assign n474 = x234 ^ x197 ^ 1'b0 ;
  assign n475 = n265 & n474 ;
  assign n476 = n475 ^ x56 ^ 1'b0 ;
  assign n477 = x246 & n347 ;
  assign n478 = ~x94 & n477 ;
  assign n479 = x179 & n411 ;
  assign n480 = n479 ^ x80 ^ 1'b0 ;
  assign n481 = n480 ^ x69 ^ x33 ;
  assign n482 = n340 ^ x166 ^ x18 ;
  assign n483 = n274 ^ x185 ^ 1'b0 ;
  assign n484 = ~n341 & n483 ;
  assign n485 = ( x34 & ~x179 ) | ( x34 & n472 ) | ( ~x179 & n472 ) ;
  assign n486 = ( x131 & ~x156 ) | ( x131 & x250 ) | ( ~x156 & x250 ) ;
  assign n487 = x221 & n486 ;
  assign n488 = n292 & n487 ;
  assign n489 = n311 ^ x221 ^ 1'b0 ;
  assign n490 = n489 ^ x161 ^ 1'b0 ;
  assign n491 = ( x149 & ~x156 ) | ( x149 & x226 ) | ( ~x156 & x226 ) ;
  assign n492 = n374 ^ x144 ^ 1'b0 ;
  assign n493 = x113 & x239 ;
  assign n494 = ~x241 & n493 ;
  assign n495 = x163 | n494 ;
  assign n496 = x210 & n495 ;
  assign n497 = x188 & ~n496 ;
  assign n498 = n492 & n497 ;
  assign n499 = n498 ^ n317 ^ 1'b0 ;
  assign n500 = x22 & n499 ;
  assign n501 = x84 & x222 ;
  assign n502 = n501 ^ n289 ^ 1'b0 ;
  assign n503 = n502 ^ n443 ^ 1'b0 ;
  assign n504 = n453 | n503 ;
  assign n505 = x9 & ~x34 ;
  assign n506 = ( ~x54 & x85 ) | ( ~x54 & n275 ) | ( x85 & n275 ) ;
  assign n507 = x173 & ~n366 ;
  assign n508 = n507 ^ x159 ^ 1'b0 ;
  assign n509 = n508 ^ n298 ^ x17 ;
  assign n510 = x77 & n344 ;
  assign n511 = n510 ^ x185 ^ 1'b0 ;
  assign n513 = ( x89 & x116 ) | ( x89 & ~x216 ) | ( x116 & ~x216 ) ;
  assign n514 = n513 ^ x128 ^ x45 ;
  assign n515 = n514 ^ x99 ^ 1'b0 ;
  assign n516 = n335 | n515 ;
  assign n512 = ( x68 & x102 ) | ( x68 & ~x158 ) | ( x102 & ~x158 ) ;
  assign n517 = n516 ^ n512 ^ 1'b0 ;
  assign n518 = x182 & ~n517 ;
  assign n519 = ~x60 & x193 ;
  assign n520 = n519 ^ n489 ^ 1'b0 ;
  assign n521 = x50 & n520 ;
  assign n522 = ~x159 & n521 ;
  assign n523 = n432 ^ x49 ^ 1'b0 ;
  assign n524 = x191 & ~n523 ;
  assign n525 = x39 & x105 ;
  assign n526 = n525 ^ n425 ^ 1'b0 ;
  assign n527 = ~x39 & x143 ;
  assign n528 = x63 & x249 ;
  assign n529 = n332 & n528 ;
  assign n536 = x201 ^ x99 ^ x87 ;
  assign n531 = x241 & n326 ;
  assign n532 = x237 & ~n531 ;
  assign n533 = n305 & n532 ;
  assign n534 = x7 & x111 ;
  assign n535 = n533 & n534 ;
  assign n530 = ( x25 & ~x118 ) | ( x25 & x184 ) | ( ~x118 & x184 ) ;
  assign n537 = n536 ^ n535 ^ n530 ;
  assign n538 = n267 ^ x199 ^ x144 ;
  assign n539 = n538 ^ x45 ^ x43 ;
  assign n540 = n539 ^ n395 ^ 1'b0 ;
  assign n541 = n537 | n540 ;
  assign n545 = ( x10 & n308 ) | ( x10 & ~n446 ) | ( n308 & ~n446 ) ;
  assign n542 = x79 ^ x1 ^ 1'b0 ;
  assign n543 = x12 & n542 ;
  assign n544 = n388 & n543 ;
  assign n546 = n545 ^ n544 ^ 1'b0 ;
  assign n547 = x35 & x232 ;
  assign n548 = n498 & n547 ;
  assign n549 = n365 ^ n261 ^ x195 ;
  assign n550 = ~n465 & n549 ;
  assign n551 = x247 & n311 ;
  assign n552 = n551 ^ n277 ^ 1'b0 ;
  assign n553 = ( x13 & n400 ) | ( x13 & n472 ) | ( n400 & n472 ) ;
  assign n554 = n553 ^ x225 ^ 1'b0 ;
  assign n555 = x143 & n554 ;
  assign n556 = x33 & ~n555 ;
  assign n557 = n486 ^ n358 ^ n345 ;
  assign n558 = x236 & n557 ;
  assign n559 = n488 ^ x49 ^ x26 ;
  assign n560 = n559 ^ n279 ^ x166 ;
  assign n561 = x35 & x241 ;
  assign n562 = n273 & n561 ;
  assign n563 = n289 & n562 ;
  assign n564 = n505 ^ x119 ^ 1'b0 ;
  assign n565 = x252 & n564 ;
  assign n566 = x107 & n565 ;
  assign n567 = n566 ^ n512 ^ 1'b0 ;
  assign n568 = x168 & x214 ;
  assign n569 = n405 & n568 ;
  assign n570 = x155 & ~n369 ;
  assign n571 = ( x41 & n569 ) | ( x41 & n570 ) | ( n569 & n570 ) ;
  assign n572 = n377 | n399 ;
  assign n574 = ( x57 & x207 ) | ( x57 & ~x234 ) | ( x207 & ~x234 ) ;
  assign n573 = x214 & n543 ;
  assign n575 = n574 ^ n573 ^ 1'b0 ;
  assign n576 = x36 ^ x11 ^ 1'b0 ;
  assign n577 = ~n390 & n576 ;
  assign n578 = x12 & n577 ;
  assign n579 = ~x1 & n578 ;
  assign n580 = ( x83 & ~x107 ) | ( x83 & x110 ) | ( ~x107 & x110 ) ;
  assign n581 = n580 ^ x173 ^ x90 ;
  assign n582 = x14 & n581 ;
  assign n583 = n582 ^ n328 ^ x79 ;
  assign n584 = ~n579 & n583 ;
  assign n585 = n584 ^ x60 ^ 1'b0 ;
  assign n586 = x120 ^ x69 ^ 1'b0 ;
  assign n587 = ~n363 & n586 ;
  assign n588 = x149 ^ x114 ^ x11 ;
  assign n589 = ~x168 & x210 ;
  assign n590 = n588 & n589 ;
  assign n591 = ( x54 & ~n587 ) | ( x54 & n590 ) | ( ~n587 & n590 ) ;
  assign n592 = n583 ^ n332 ^ n283 ;
  assign n595 = x171 ^ x93 ^ 1'b0 ;
  assign n596 = x33 & n595 ;
  assign n593 = x186 ^ x172 ^ x123 ;
  assign n594 = n593 ^ n433 ^ x139 ;
  assign n597 = n596 ^ n594 ^ n531 ;
  assign n598 = x151 & n574 ;
  assign n599 = x109 & ~n308 ;
  assign n600 = ~x248 & n599 ;
  assign n603 = x5 & x230 ;
  assign n604 = n603 ^ x119 ^ 1'b0 ;
  assign n605 = ( x96 & ~n410 ) | ( x96 & n604 ) | ( ~n410 & n604 ) ;
  assign n601 = ( x5 & ~n512 ) | ( x5 & n565 ) | ( ~n512 & n565 ) ;
  assign n602 = x7 & n601 ;
  assign n606 = n605 ^ n602 ^ 1'b0 ;
  assign n608 = ( x131 & ~x175 ) | ( x131 & x225 ) | ( ~x175 & x225 ) ;
  assign n607 = n345 ^ n326 ^ x162 ;
  assign n609 = n608 ^ n607 ^ 1'b0 ;
  assign n610 = ~n604 & n609 ;
  assign n611 = x153 & x199 ;
  assign n612 = ~n610 & n611 ;
  assign n613 = x93 & ~n291 ;
  assign n614 = ~x146 & n613 ;
  assign n615 = x41 & ~n423 ;
  assign n616 = n614 & n615 ;
  assign n617 = n616 ^ x15 ^ 1'b0 ;
  assign n619 = x87 & ~n329 ;
  assign n620 = ~x44 & n619 ;
  assign n621 = x14 & ~n620 ;
  assign n622 = n621 ^ n357 ^ 1'b0 ;
  assign n623 = n622 ^ x249 ^ x35 ;
  assign n618 = x116 & ~n537 ;
  assign n624 = n623 ^ n618 ^ 1'b0 ;
  assign n627 = n275 ^ x218 ^ 1'b0 ;
  assign n625 = x216 & ~n302 ;
  assign n626 = n625 ^ x177 ^ 1'b0 ;
  assign n628 = n627 ^ n626 ^ 1'b0 ;
  assign n629 = n538 & ~n628 ;
  assign n630 = x72 & x196 ;
  assign n631 = n630 ^ x146 ^ 1'b0 ;
  assign n632 = n631 ^ n608 ^ 1'b0 ;
  assign n633 = n629 & ~n632 ;
  assign n634 = n307 & n633 ;
  assign n635 = n623 ^ x207 ^ x86 ;
  assign n636 = ( x179 & n537 ) | ( x179 & n635 ) | ( n537 & n635 ) ;
  assign n637 = ~x69 & x98 ;
  assign n638 = x56 & x145 ;
  assign n639 = ~x166 & n638 ;
  assign n640 = n639 ^ n329 ^ x85 ;
  assign n641 = n640 ^ x132 ^ 1'b0 ;
  assign n642 = n637 | n641 ;
  assign n643 = n589 ^ n315 ^ x124 ;
  assign n645 = n536 ^ n387 ^ x0 ;
  assign n644 = x129 & ~n541 ;
  assign n646 = n645 ^ n644 ^ 1'b0 ;
  assign n647 = x86 & ~x252 ;
  assign n648 = n647 ^ n296 ^ 1'b0 ;
  assign n649 = x203 & ~n374 ;
  assign n650 = n649 ^ n360 ^ 1'b0 ;
  assign n651 = x102 ^ x39 ^ 1'b0 ;
  assign n652 = x241 & n651 ;
  assign n653 = ~x130 & n652 ;
  assign n654 = ~n305 & n340 ;
  assign n655 = n654 ^ x32 ^ 1'b0 ;
  assign n656 = n655 ^ n298 ^ 1'b0 ;
  assign n657 = n383 & n656 ;
  assign n658 = x101 ^ x59 ^ 1'b0 ;
  assign n659 = n657 & n658 ;
  assign n660 = ( x106 & x132 ) | ( x106 & ~x224 ) | ( x132 & ~x224 ) ;
  assign n661 = n536 & ~n572 ;
  assign n662 = n660 & ~n661 ;
  assign n663 = ~n397 & n662 ;
  assign n664 = x170 & ~n304 ;
  assign n665 = ~x127 & n664 ;
  assign n666 = n543 ^ x100 ^ x15 ;
  assign n673 = n494 ^ x238 ^ 1'b0 ;
  assign n670 = x77 ^ x50 ^ 1'b0 ;
  assign n671 = ~n556 & n670 ;
  assign n668 = ( x131 & ~x144 ) | ( x131 & x194 ) | ( ~x144 & x194 ) ;
  assign n667 = x7 & ~n637 ;
  assign n669 = n668 ^ n667 ^ 1'b0 ;
  assign n672 = n671 ^ n669 ^ 1'b0 ;
  assign n674 = n673 ^ n672 ^ n387 ;
  assign n675 = x239 ^ x215 ^ 1'b0 ;
  assign n676 = n675 ^ x72 ^ 1'b0 ;
  assign n677 = x81 & ~n676 ;
  assign n678 = x183 ^ x51 ^ 1'b0 ;
  assign n679 = x190 & n678 ;
  assign n680 = x22 & n679 ;
  assign n681 = ~x185 & n680 ;
  assign n682 = n433 & ~n516 ;
  assign n683 = n682 ^ x26 ^ 1'b0 ;
  assign n684 = n683 ^ x240 ^ 1'b0 ;
  assign n685 = n681 | n684 ;
  assign n689 = x185 & x246 ;
  assign n690 = n689 ^ x137 ^ 1'b0 ;
  assign n686 = x159 ^ x98 ^ 1'b0 ;
  assign n687 = n634 ^ n413 ^ 1'b0 ;
  assign n688 = n686 & n687 ;
  assign n691 = n690 ^ n688 ^ 1'b0 ;
  assign n692 = n393 | n691 ;
  assign n693 = x187 ^ x137 ^ x134 ;
  assign n694 = x75 & n693 ;
  assign n696 = n390 ^ n283 ^ 1'b0 ;
  assign n697 = ~n417 & n696 ;
  assign n695 = x46 & ~n322 ;
  assign n698 = n697 ^ n695 ^ 1'b0 ;
  assign n699 = n383 & n397 ;
  assign n700 = n699 ^ x92 ^ 1'b0 ;
  assign n701 = x86 & ~n700 ;
  assign n702 = n701 ^ n558 ^ 1'b0 ;
  assign n703 = x216 & ~n400 ;
  assign n704 = n620 & n703 ;
  assign n705 = x55 & n679 ;
  assign n706 = n704 & n705 ;
  assign n707 = ( ~x121 & n360 ) | ( ~x121 & n410 ) | ( n360 & n410 ) ;
  assign n708 = n707 ^ n637 ^ 1'b0 ;
  assign n709 = n412 & ~n708 ;
  assign n710 = x125 & ~n631 ;
  assign n711 = n710 ^ x37 ^ 1'b0 ;
  assign n712 = ~x172 & n570 ;
  assign n713 = ( x96 & ~n306 ) | ( x96 & n712 ) | ( ~n306 & n712 ) ;
  assign n714 = ( ~x47 & x134 ) | ( ~x47 & n514 ) | ( x134 & n514 ) ;
  assign n715 = n433 ^ x225 ^ 1'b0 ;
  assign n716 = n443 & n715 ;
  assign n717 = x16 & n560 ;
  assign n718 = n717 ^ x101 ^ 1'b0 ;
  assign n720 = x116 & n660 ;
  assign n721 = ~x218 & n720 ;
  assign n722 = n627 & ~n721 ;
  assign n723 = ~x12 & n722 ;
  assign n724 = x237 & ~n723 ;
  assign n725 = n724 ^ n647 ^ 1'b0 ;
  assign n726 = x46 & n725 ;
  assign n727 = n726 ^ n411 ^ 1'b0 ;
  assign n719 = n583 ^ n463 ^ n372 ;
  assign n728 = n727 ^ n719 ^ n275 ;
  assign n729 = n304 & ~n728 ;
  assign n730 = n267 | n588 ;
  assign n731 = n730 ^ n390 ^ 1'b0 ;
  assign n732 = n731 ^ x95 ^ 1'b0 ;
  assign n733 = ~x212 & n277 ;
  assign n734 = x246 ^ x132 ^ 1'b0 ;
  assign n735 = n734 ^ x171 ^ 1'b0 ;
  assign n741 = x109 ^ x48 ^ 1'b0 ;
  assign n742 = x203 & n741 ;
  assign n743 = n742 ^ x116 ^ 1'b0 ;
  assign n744 = n743 ^ n669 ^ n417 ;
  assign n737 = n516 ^ x233 ^ x143 ;
  assign n736 = n261 ^ x114 ^ x99 ;
  assign n738 = n737 ^ n736 ^ 1'b0 ;
  assign n739 = ~n549 & n738 ;
  assign n740 = n474 & n739 ;
  assign n745 = n744 ^ n740 ^ 1'b0 ;
  assign n746 = n385 & ~n387 ;
  assign n747 = n746 ^ x94 ^ 1'b0 ;
  assign n748 = n747 ^ n494 ^ 1'b0 ;
  assign n749 = x1 & n748 ;
  assign n750 = x14 & x133 ;
  assign n751 = n750 ^ n407 ^ 1'b0 ;
  assign n752 = n308 & n751 ;
  assign n753 = n458 ^ x227 ^ 1'b0 ;
  assign n754 = n549 ^ n311 ^ 1'b0 ;
  assign n755 = n634 & ~n754 ;
  assign n756 = x57 & n279 ;
  assign n757 = n265 & ~n319 ;
  assign n758 = ~x109 & n757 ;
  assign n759 = ( ~x142 & x200 ) | ( ~x142 & x253 ) | ( x200 & x253 ) ;
  assign n760 = ( x30 & x36 ) | ( x30 & ~n397 ) | ( x36 & ~n397 ) ;
  assign n761 = n760 ^ n377 ^ 1'b0 ;
  assign n762 = n761 ^ n543 ^ x64 ;
  assign n763 = n646 & ~n762 ;
  assign n764 = ~n759 & n763 ;
  assign n765 = n277 & ~n758 ;
  assign n766 = n765 ^ x77 ^ 1'b0 ;
  assign n767 = x140 & ~n562 ;
  assign n768 = ~n660 & n767 ;
  assign n769 = x181 & n520 ;
  assign n770 = n768 & n769 ;
  assign n771 = n372 & ~n770 ;
  assign n772 = ~x154 & n771 ;
  assign n773 = x232 ^ x67 ^ 1'b0 ;
  assign n774 = n545 & n773 ;
  assign n779 = x35 & x218 ;
  assign n780 = n779 ^ x88 ^ 1'b0 ;
  assign n775 = n281 & ~n315 ;
  assign n776 = ~x198 & n775 ;
  assign n777 = x60 & ~n776 ;
  assign n778 = ~x169 & n777 ;
  assign n781 = n780 ^ n778 ^ 1'b0 ;
  assign n782 = n489 ^ x61 ^ 1'b0 ;
  assign n783 = ~n781 & n782 ;
  assign n784 = x88 & n284 ;
  assign n785 = n784 ^ n427 ^ 1'b0 ;
  assign n786 = x175 & ~n785 ;
  assign n787 = n436 & n786 ;
  assign n788 = n669 | n787 ;
  assign n789 = n788 ^ n743 ^ 1'b0 ;
  assign n790 = n429 ^ n351 ^ x53 ;
  assign n791 = n790 ^ n351 ^ n275 ;
  assign n792 = x155 & x231 ;
  assign n793 = ~x179 & n792 ;
  assign n794 = n725 & ~n793 ;
  assign n795 = n794 ^ x159 ^ 1'b0 ;
  assign n796 = n337 | n458 ;
  assign n797 = n796 ^ n600 ^ 1'b0 ;
  assign n798 = ~n506 & n543 ;
  assign n799 = x133 & n372 ;
  assign n800 = ~n327 & n799 ;
  assign n801 = x221 & ~n800 ;
  assign n802 = n801 ^ x44 ^ 1'b0 ;
  assign n803 = n802 ^ x185 ^ x110 ;
  assign n804 = n259 ^ x199 ^ 1'b0 ;
  assign n805 = n458 ^ x210 ^ x196 ;
  assign n806 = x172 & ~n747 ;
  assign n807 = n806 ^ n574 ^ 1'b0 ;
  assign n808 = n805 & n807 ;
  assign n809 = n547 ^ n326 ^ 1'b0 ;
  assign n810 = x170 & ~n647 ;
  assign n811 = ~x110 & n810 ;
  assign n812 = n809 & ~n811 ;
  assign n813 = ~n490 & n812 ;
  assign n814 = n413 ^ x212 ^ 1'b0 ;
  assign n815 = x158 | n814 ;
  assign n816 = n587 ^ x15 ^ 1'b0 ;
  assign n817 = x145 & n816 ;
  assign n818 = x190 & ~n817 ;
  assign n820 = n412 ^ x26 ^ 1'b0 ;
  assign n821 = ~n593 & n820 ;
  assign n819 = x132 & x155 ;
  assign n822 = n821 ^ n819 ^ 1'b0 ;
  assign n823 = n306 & ~n535 ;
  assign n824 = n823 ^ n289 ^ 1'b0 ;
  assign n825 = n756 | n824 ;
  assign n826 = x10 | n825 ;
  assign n827 = ~n315 & n608 ;
  assign n828 = n279 & n827 ;
  assign n829 = x168 & ~n828 ;
  assign n832 = n655 ^ x142 ^ x61 ;
  assign n830 = x201 ^ x110 ^ 1'b0 ;
  assign n831 = x210 & n830 ;
  assign n833 = n832 ^ n831 ^ x148 ;
  assign n834 = n596 & ~n833 ;
  assign n835 = ~n829 & n834 ;
  assign n838 = n743 & ~n828 ;
  assign n839 = n773 & ~n838 ;
  assign n840 = n839 ^ x68 ^ 1'b0 ;
  assign n836 = x5 & ~n535 ;
  assign n837 = x177 & n836 ;
  assign n841 = n840 ^ n837 ^ 1'b0 ;
  assign n842 = x170 & n492 ;
  assign n843 = n842 ^ n496 ^ x98 ;
  assign n844 = x165 & n843 ;
  assign n845 = n844 ^ n423 ^ 1'b0 ;
  assign n853 = x9 & ~n640 ;
  assign n848 = x155 & ~n341 ;
  assign n849 = ~x41 & n848 ;
  assign n850 = n849 ^ n480 ^ 1'b0 ;
  assign n851 = ~n331 & n850 ;
  assign n852 = n851 ^ n753 ^ n567 ;
  assign n846 = x87 & x150 ;
  assign n847 = n846 ^ n369 ^ 1'b0 ;
  assign n854 = n853 ^ n852 ^ n847 ;
  assign n860 = ( x111 & ~x189 ) | ( x111 & x213 ) | ( ~x189 & x213 ) ;
  assign n855 = x136 & ~n263 ;
  assign n856 = n855 ^ x93 ^ 1'b0 ;
  assign n857 = n856 ^ x113 ^ 1'b0 ;
  assign n858 = x195 & ~n857 ;
  assign n859 = x16 & n858 ;
  assign n861 = n860 ^ n859 ^ 1'b0 ;
  assign n862 = x133 & x155 ;
  assign n863 = n862 ^ x82 ^ 1'b0 ;
  assign n864 = x58 & ~n863 ;
  assign n865 = ~n347 & n864 ;
  assign n866 = n361 ^ x236 ^ x207 ;
  assign n867 = n865 | n866 ;
  assign n871 = x162 ^ x23 ^ 1'b0 ;
  assign n868 = x212 ^ x10 ^ 1'b0 ;
  assign n869 = x217 & n868 ;
  assign n870 = x101 & n869 ;
  assign n872 = n871 ^ n870 ^ 1'b0 ;
  assign n873 = n380 ^ x108 ^ 1'b0 ;
  assign n874 = n802 & ~n873 ;
  assign n875 = x129 | n296 ;
  assign n876 = ~x15 & n512 ;
  assign n877 = ~x48 & n876 ;
  assign n878 = n875 | n877 ;
  assign n879 = ( x201 & ~n535 ) | ( x201 & n714 ) | ( ~n535 & n714 ) ;
  assign n880 = n879 ^ n587 ^ n411 ;
  assign n881 = x90 & ~n732 ;
  assign n882 = x67 & x100 ;
  assign n883 = n345 & ~n616 ;
  assign n884 = ~n725 & n883 ;
  assign n885 = x124 & n634 ;
  assign n886 = n885 ^ n759 ^ 1'b0 ;
  assign n887 = ( n882 & ~n884 ) | ( n882 & n886 ) | ( ~n884 & n886 ) ;
  assign n888 = n459 ^ n415 ^ 1'b0 ;
  assign n889 = n569 | n888 ;
  assign n890 = ( x96 & n322 ) | ( x96 & n385 ) | ( n322 & n385 ) ;
  assign n891 = x32 & x82 ;
  assign n892 = ~x254 & n891 ;
  assign n893 = x166 ^ x86 ^ 1'b0 ;
  assign n894 = ~n892 & n893 ;
  assign n895 = x157 & n539 ;
  assign n896 = n895 ^ n774 ^ n665 ;
  assign n897 = n814 ^ x44 ^ 1'b0 ;
  assign n898 = ~x82 & n281 ;
  assign n899 = ~n393 & n520 ;
  assign n900 = n569 & n899 ;
  assign n901 = n898 | n900 ;
  assign n902 = x25 | n901 ;
  assign n903 = x38 & x148 ;
  assign n904 = n903 ^ n488 ^ x29 ;
  assign n905 = n286 ^ n275 ^ x212 ;
  assign n906 = ( x222 & n751 ) | ( x222 & ~n905 ) | ( n751 & ~n905 ) ;
  assign n907 = n735 ^ n583 ^ x203 ;
  assign n908 = n907 ^ n681 ^ n377 ;
  assign n909 = x144 ^ x135 ^ 1'b0 ;
  assign n910 = n332 ^ n281 ^ 1'b0 ;
  assign n911 = x182 & ~n910 ;
  assign n912 = n911 ^ x55 ^ 1'b0 ;
  assign n913 = n909 & n912 ;
  assign n914 = x133 & n652 ;
  assign n915 = n914 ^ x117 ^ 1'b0 ;
  assign n916 = n915 ^ x35 ^ 1'b0 ;
  assign n917 = n913 & ~n916 ;
  assign n918 = n749 & n917 ;
  assign n919 = ~x7 & n488 ;
  assign n920 = n919 ^ n319 ^ 1'b0 ;
  assign n921 = x133 & n920 ;
  assign n922 = ( x35 & ~n277 ) | ( x35 & n529 ) | ( ~n277 & n529 ) ;
  assign n923 = n307 & ~n333 ;
  assign n924 = ~x111 & n923 ;
  assign n925 = n924 ^ x46 ^ 1'b0 ;
  assign n926 = x230 & ~n925 ;
  assign n927 = x13 & n926 ;
  assign n928 = n922 & n927 ;
  assign n929 = n753 & n841 ;
  assign n930 = n620 & n929 ;
  assign n931 = n274 | n930 ;
  assign n932 = n556 ^ x237 ^ x95 ;
  assign n933 = n932 ^ n895 ^ 1'b0 ;
  assign n934 = n933 ^ x74 ^ 1'b0 ;
  assign n935 = n500 & ~n934 ;
  assign n936 = ( x239 & n418 ) | ( x239 & ~n631 ) | ( n418 & ~n631 ) ;
  assign n937 = n936 ^ n723 ^ x69 ;
  assign n938 = n937 ^ n404 ^ 1'b0 ;
  assign n939 = n935 & ~n938 ;
  assign n940 = ( ~n340 & n531 ) | ( ~n340 & n939 ) | ( n531 & n939 ) ;
  assign n941 = x195 & n607 ;
  assign n942 = n941 ^ x145 ^ 1'b0 ;
  assign n943 = n274 & ~n942 ;
  assign n944 = ~x0 & n943 ;
  assign n946 = x128 ^ x104 ^ 1'b0 ;
  assign n945 = n444 | n581 ;
  assign n947 = n946 ^ n945 ^ 1'b0 ;
  assign n948 = n944 & n947 ;
  assign n949 = x186 & n259 ;
  assign n950 = n949 ^ n718 ^ 1'b0 ;
  assign n951 = x83 & n950 ;
  assign n952 = n948 & n951 ;
  assign n953 = n284 & n385 ;
  assign n954 = n953 ^ x233 ^ 1'b0 ;
  assign n955 = n308 ^ x83 ^ 1'b0 ;
  assign n956 = x166 & ~n955 ;
  assign n957 = n956 ^ n433 ^ 1'b0 ;
  assign n958 = n760 ^ n490 ^ 1'b0 ;
  assign n959 = ~n957 & n958 ;
  assign n960 = ( ~n948 & n954 ) | ( ~n948 & n959 ) | ( n954 & n959 ) ;
  assign n961 = n838 ^ n345 ^ 1'b0 ;
  assign n965 = x107 & ~n460 ;
  assign n966 = ~x162 & n965 ;
  assign n962 = x142 & x252 ;
  assign n963 = n962 ^ n338 ^ 1'b0 ;
  assign n964 = n753 | n963 ;
  assign n967 = n966 ^ n964 ^ 1'b0 ;
  assign n968 = n785 ^ n606 ^ x13 ;
  assign n975 = x214 ^ x69 ^ 1'b0 ;
  assign n969 = x186 ^ x139 ^ 1'b0 ;
  assign n970 = x244 & n969 ;
  assign n971 = x80 & n751 ;
  assign n972 = ~n970 & n971 ;
  assign n973 = n783 & ~n972 ;
  assign n974 = ~n883 & n973 ;
  assign n976 = n975 ^ n974 ^ 1'b0 ;
  assign n977 = n527 ^ n505 ^ 1'b0 ;
  assign n978 = n581 | n977 ;
  assign n979 = x144 & n511 ;
  assign n980 = ( x121 & ~n340 ) | ( x121 & n707 ) | ( ~n340 & n707 ) ;
  assign n981 = n980 ^ n417 ^ 1'b0 ;
  assign n982 = ( x14 & n337 ) | ( x14 & ~n981 ) | ( n337 & ~n981 ) ;
  assign n983 = ( n292 & ~n979 ) | ( n292 & n982 ) | ( ~n979 & n982 ) ;
  assign n984 = ( n892 & ~n978 ) | ( n892 & n983 ) | ( ~n978 & n983 ) ;
  assign n985 = ( ~x215 & n399 ) | ( ~x215 & n793 ) | ( n399 & n793 ) ;
  assign n986 = x249 ^ x112 ^ 1'b0 ;
  assign n987 = ~n985 & n986 ;
  assign n988 = ( x202 & n984 ) | ( x202 & n987 ) | ( n984 & n987 ) ;
  assign n989 = n970 ^ x62 ^ 1'b0 ;
  assign n990 = x137 & x163 ;
  assign n991 = n990 ^ x118 ^ 1'b0 ;
  assign n994 = ~x7 & x214 ;
  assign n992 = x252 & ~n785 ;
  assign n993 = ~x229 & n992 ;
  assign n995 = n994 ^ n993 ^ n887 ;
  assign n996 = x250 & n526 ;
  assign n997 = n996 ^ n693 ^ 1'b0 ;
  assign n998 = x120 & ~n997 ;
  assign n1000 = ( n267 & n545 ) | ( n267 & ~n768 ) | ( n545 & ~n768 ) ;
  assign n999 = x122 & ~n626 ;
  assign n1001 = n1000 ^ n999 ^ 1'b0 ;
  assign n1002 = n749 & n791 ;
  assign n1003 = n1002 ^ x189 ^ 1'b0 ;
  assign n1004 = n780 ^ n441 ^ 1'b0 ;
  assign n1005 = x83 & n319 ;
  assign n1006 = x61 & ~n1005 ;
  assign n1007 = n425 ^ x136 ^ 1'b0 ;
  assign n1008 = n261 | n361 ;
  assign n1009 = n1008 ^ x186 ^ 1'b0 ;
  assign n1010 = ~n982 & n1009 ;
  assign n1011 = x110 & n884 ;
  assign n1012 = x200 ^ x90 ^ 1'b0 ;
  assign n1013 = n410 & n1012 ;
  assign n1014 = x221 & n1013 ;
  assign n1015 = ~x19 & n1014 ;
  assign n1016 = n296 | n1015 ;
  assign n1017 = n1016 ^ x41 ^ 1'b0 ;
  assign n1018 = x190 & n1017 ;
  assign n1019 = ~n652 & n1018 ;
  assign n1020 = n894 & ~n1019 ;
  assign n1021 = n1020 ^ n545 ^ 1'b0 ;
  assign n1022 = n413 ^ x237 ^ 1'b0 ;
  assign n1023 = n1022 ^ n492 ^ 1'b0 ;
  assign n1024 = ~n433 & n463 ;
  assign n1025 = ( x193 & ~n488 ) | ( x193 & n972 ) | ( ~n488 & n972 ) ;
  assign n1026 = x88 & n1025 ;
  assign n1027 = x141 ^ x89 ^ 1'b0 ;
  assign n1028 = n706 ^ n549 ^ 1'b0 ;
  assign n1029 = n1027 & n1028 ;
  assign n1030 = ( n256 & n1023 ) | ( n256 & n1029 ) | ( n1023 & n1029 ) ;
  assign n1032 = n539 ^ x233 ^ 1'b0 ;
  assign n1033 = x244 & ~n1032 ;
  assign n1031 = ( n665 & n903 ) | ( n665 & ~n907 ) | ( n903 & ~n907 ) ;
  assign n1034 = n1033 ^ n1031 ^ 1'b0 ;
  assign n1038 = n489 | n616 ;
  assign n1035 = n402 ^ n377 ^ 1'b0 ;
  assign n1036 = x105 & n1035 ;
  assign n1037 = ~x252 & n1036 ;
  assign n1039 = n1038 ^ n1037 ^ 1'b0 ;
  assign n1040 = n385 & ~n1039 ;
  assign n1041 = n994 ^ x85 ^ x28 ;
  assign n1042 = ( x119 & n376 ) | ( x119 & ~n1023 ) | ( n376 & ~n1023 ) ;
  assign n1043 = n755 ^ n645 ^ 1'b0 ;
  assign n1044 = n987 & ~n1043 ;
  assign n1045 = n482 | n963 ;
  assign n1046 = n1045 ^ n902 ^ 1'b0 ;
  assign n1051 = x29 & n399 ;
  assign n1052 = n1051 ^ x120 ^ 1'b0 ;
  assign n1053 = n1052 ^ n895 ^ 1'b0 ;
  assign n1050 = x10 & n289 ;
  assign n1054 = n1053 ^ n1050 ^ 1'b0 ;
  assign n1047 = n652 ^ x101 ^ 1'b0 ;
  assign n1048 = ~n267 & n1047 ;
  assign n1049 = ~x174 & n1048 ;
  assign n1055 = n1054 ^ n1049 ^ x230 ;
  assign n1056 = n494 ^ n488 ^ n337 ;
  assign n1057 = n1048 & ~n1056 ;
  assign n1058 = n1057 ^ n463 ^ 1'b0 ;
  assign n1059 = n485 ^ x220 ^ x147 ;
  assign n1060 = n674 & n1059 ;
  assign n1061 = x242 & n299 ;
  assign n1062 = n1061 ^ x214 ^ 1'b0 ;
  assign n1063 = ( ~x53 & n307 ) | ( ~x53 & n1062 ) | ( n307 & n1062 ) ;
  assign n1065 = x80 & ~n407 ;
  assign n1066 = n1065 ^ x91 ^ 1'b0 ;
  assign n1064 = n514 ^ x140 ^ 1'b0 ;
  assign n1067 = n1066 ^ n1064 ^ x207 ;
  assign n1068 = n1067 ^ x246 ^ 1'b0 ;
  assign n1069 = n994 ^ n478 ^ 1'b0 ;
  assign n1070 = ~n714 & n1069 ;
  assign n1071 = x243 ^ x101 ^ 1'b0 ;
  assign n1072 = ~n563 & n1071 ;
  assign n1073 = n879 & ~n1072 ;
  assign n1074 = n409 | n778 ;
  assign n1075 = x205 | n1074 ;
  assign n1076 = ~n975 & n1075 ;
  assign n1077 = n1076 ^ n397 ^ 1'b0 ;
  assign n1081 = x95 & n1005 ;
  assign n1082 = n854 & ~n1038 ;
  assign n1083 = n462 & ~n1082 ;
  assign n1084 = ~n1081 & n1083 ;
  assign n1078 = x85 & x112 ;
  assign n1079 = ~x53 & n1078 ;
  assign n1080 = n712 | n1079 ;
  assign n1085 = n1084 ^ n1080 ^ 1'b0 ;
  assign n1086 = n1085 ^ n956 ^ n267 ;
  assign n1087 = x140 & x208 ;
  assign n1088 = n1087 ^ n723 ^ 1'b0 ;
  assign n1089 = x74 ^ x7 ^ 1'b0 ;
  assign n1090 = n489 & n1089 ;
  assign n1091 = ( x202 & ~n444 ) | ( x202 & n552 ) | ( ~n444 & n552 ) ;
  assign n1098 = n661 ^ x203 ^ 1'b0 ;
  assign n1092 = x28 & ~n418 ;
  assign n1093 = n1092 ^ x86 ^ 1'b0 ;
  assign n1094 = n366 | n541 ;
  assign n1095 = n1094 ^ n489 ^ 1'b0 ;
  assign n1096 = n1095 ^ n417 ^ x232 ;
  assign n1097 = ( x232 & n1093 ) | ( x232 & n1096 ) | ( n1093 & n1096 ) ;
  assign n1099 = n1098 ^ n1097 ^ 1'b0 ;
  assign n1100 = x144 & n1040 ;
  assign n1101 = n1100 ^ n1070 ^ 1'b0 ;
  assign n1102 = x79 ^ x72 ^ 1'b0 ;
  assign n1103 = ~x23 & n1102 ;
  assign n1107 = ( x158 & ~x177 ) | ( x158 & x196 ) | ( ~x177 & x196 ) ;
  assign n1108 = ~n447 & n1107 ;
  assign n1104 = n512 & n570 ;
  assign n1105 = n267 & n1104 ;
  assign n1106 = n1105 ^ n856 ^ 1'b0 ;
  assign n1109 = n1108 ^ n1106 ^ 1'b0 ;
  assign n1110 = n809 & ~n1109 ;
  assign n1111 = x177 & ~n1110 ;
  assign n1112 = n1022 ^ n407 ^ 1'b0 ;
  assign n1113 = n587 & n1112 ;
  assign n1114 = ~n296 & n1113 ;
  assign n1115 = ~x146 & n1114 ;
  assign n1116 = n1115 ^ n1090 ^ 1'b0 ;
  assign n1117 = n553 & ~n1116 ;
  assign n1118 = n371 | n915 ;
  assign n1119 = n831 | n1118 ;
  assign n1120 = ~x200 & x250 ;
  assign n1121 = n879 & n1027 ;
  assign n1122 = n734 | n1121 ;
  assign n1123 = ~n1101 & n1122 ;
  assign n1124 = n1120 & n1123 ;
  assign n1125 = x180 & ~n589 ;
  assign n1126 = x127 | n1125 ;
  assign n1127 = n728 | n1103 ;
  assign n1128 = n455 | n721 ;
  assign n1129 = n1128 ^ n474 ^ 1'b0 ;
  assign n1130 = n580 & n1129 ;
  assign n1131 = n1072 & n1130 ;
  assign n1132 = ~n1006 & n1131 ;
  assign n1133 = ~x15 & x41 ;
  assign n1134 = ~n491 & n1133 ;
  assign n1135 = x123 & x233 ;
  assign n1136 = n616 & n1135 ;
  assign n1137 = n1136 ^ x100 ^ 1'b0 ;
  assign n1138 = ( n275 & ~n415 ) | ( n275 & n581 ) | ( ~n415 & n581 ) ;
  assign n1139 = n379 ^ n369 ^ 1'b0 ;
  assign n1147 = x126 & ~n505 ;
  assign n1143 = x155 & n599 ;
  assign n1144 = n569 & n1143 ;
  assign n1140 = ( x136 & ~n328 ) | ( x136 & n371 ) | ( ~n328 & n371 ) ;
  assign n1141 = ~n700 & n1140 ;
  assign n1142 = ~n994 & n1141 ;
  assign n1145 = n1144 ^ n1142 ^ n702 ;
  assign n1146 = n583 & n1145 ;
  assign n1148 = n1147 ^ n1146 ^ 1'b0 ;
  assign n1151 = x2 & ~n719 ;
  assign n1149 = x178 & ~n387 ;
  assign n1150 = n1149 ^ n420 ^ 1'b0 ;
  assign n1152 = n1151 ^ n1150 ^ n633 ;
  assign n1153 = x57 & ~n909 ;
  assign n1154 = x160 & ~n1153 ;
  assign n1155 = n1154 ^ n397 ^ 1'b0 ;
  assign n1156 = n1017 ^ x172 ^ x50 ;
  assign n1157 = n467 | n1156 ;
  assign n1158 = x109 | n1157 ;
  assign n1159 = n1158 ^ x235 ^ 1'b0 ;
  assign n1160 = ~n1155 & n1159 ;
  assign n1161 = n574 & ~n579 ;
  assign n1162 = n1161 ^ n344 ^ 1'b0 ;
  assign n1163 = n950 ^ x99 ^ 1'b0 ;
  assign n1164 = ~n605 & n1163 ;
  assign n1165 = x213 & ~n428 ;
  assign n1166 = n1165 ^ n291 ^ 1'b0 ;
  assign n1167 = ~n681 & n1166 ;
  assign n1168 = ~n956 & n1167 ;
  assign n1169 = n298 | n1168 ;
  assign n1170 = n1169 ^ n570 ^ 1'b0 ;
  assign n1171 = ~n811 & n1170 ;
  assign n1172 = n357 & n1171 ;
  assign n1173 = ( n639 & n1164 ) | ( n639 & n1172 ) | ( n1164 & n1172 ) ;
  assign n1181 = ( x120 & ~n589 ) | ( x120 & n882 ) | ( ~n589 & n882 ) ;
  assign n1182 = x251 ^ x155 ^ 1'b0 ;
  assign n1183 = n1182 ^ n1054 ^ 1'b0 ;
  assign n1184 = n1181 & ~n1183 ;
  assign n1174 = n671 ^ n302 ^ 1'b0 ;
  assign n1175 = n690 | n1174 ;
  assign n1176 = ~x19 & x130 ;
  assign n1177 = x219 & ~n413 ;
  assign n1178 = ~n1176 & n1177 ;
  assign n1179 = ~n427 & n1178 ;
  assign n1180 = n1175 & ~n1179 ;
  assign n1185 = n1184 ^ n1180 ^ 1'b0 ;
  assign n1186 = n802 | n1185 ;
  assign n1187 = ( x128 & ~n766 ) | ( x128 & n1172 ) | ( ~n766 & n1172 ) ;
  assign n1188 = n1101 ^ x167 ^ 1'b0 ;
  assign n1189 = n587 ^ n333 ^ 1'b0 ;
  assign n1190 = n809 ^ n805 ^ 1'b0 ;
  assign n1192 = n840 ^ n502 ^ 1'b0 ;
  assign n1191 = x223 ^ x170 ^ x155 ;
  assign n1193 = n1192 ^ n1191 ^ 1'b0 ;
  assign n1194 = n1071 & ~n1193 ;
  assign n1195 = ( ~n342 & n1190 ) | ( ~n342 & n1194 ) | ( n1190 & n1194 ) ;
  assign n1196 = n675 ^ x210 ^ x146 ;
  assign n1197 = n760 ^ n538 ^ n365 ;
  assign n1198 = n1196 & n1197 ;
  assign n1199 = n1198 ^ n995 ^ 1'b0 ;
  assign n1200 = n1066 ^ n768 ^ n653 ;
  assign n1201 = ( x36 & n349 ) | ( x36 & n840 ) | ( n349 & n840 ) ;
  assign n1202 = n273 ^ x109 ^ 1'b0 ;
  assign n1203 = ~n533 & n1202 ;
  assign n1204 = ~n335 & n472 ;
  assign n1205 = n1204 ^ n341 ^ 1'b0 ;
  assign n1206 = x62 ^ x54 ^ 1'b0 ;
  assign n1207 = n1205 & n1206 ;
  assign n1208 = ~n911 & n1207 ;
  assign n1209 = ( ~x5 & x33 ) | ( ~x5 & x197 ) | ( x33 & x197 ) ;
  assign n1210 = n588 & n1209 ;
  assign n1211 = x16 & ~n1210 ;
  assign n1212 = n1211 ^ n716 ^ 1'b0 ;
  assign n1213 = ( n808 & n936 ) | ( n808 & n1049 ) | ( n936 & n1049 ) ;
  assign n1214 = n697 ^ n300 ^ x111 ;
  assign n1216 = n809 ^ n459 ^ 1'b0 ;
  assign n1217 = x253 & n1216 ;
  assign n1215 = n790 ^ x20 ^ 1'b0 ;
  assign n1218 = n1217 ^ n1215 ^ n535 ;
  assign n1219 = n606 & n809 ;
  assign n1220 = n1219 ^ n514 ^ 1'b0 ;
  assign n1221 = n504 ^ n291 ^ 1'b0 ;
  assign n1222 = n821 & n1221 ;
  assign n1223 = n1222 ^ n333 ^ x170 ;
  assign n1224 = n399 & n634 ;
  assign n1225 = n1224 ^ n821 ^ 1'b0 ;
  assign n1226 = n946 & n960 ;
  assign n1227 = n1225 & n1226 ;
  assign n1228 = n663 ^ x131 ^ 1'b0 ;
  assign n1231 = ( x26 & ~x206 ) | ( x26 & n289 ) | ( ~x206 & n289 ) ;
  assign n1229 = x24 & ~n745 ;
  assign n1230 = n1229 ^ n617 ^ 1'b0 ;
  assign n1232 = n1231 ^ n1230 ^ 1'b0 ;
  assign n1233 = n1177 ^ x238 ^ x213 ;
  assign n1234 = x144 | n1233 ;
  assign n1235 = n562 ^ x247 ^ x160 ;
  assign n1236 = x84 & ~n404 ;
  assign n1237 = x181 & ~n1236 ;
  assign n1238 = x234 & n1145 ;
  assign n1239 = n1238 ^ n789 ^ 1'b0 ;
  assign n1240 = n1237 & n1239 ;
  assign n1241 = ~x132 & n1240 ;
  assign n1242 = n614 ^ x176 ^ 1'b0 ;
  assign n1243 = x82 & n1184 ;
  assign n1244 = ~n469 & n1243 ;
  assign n1245 = n1242 & ~n1244 ;
  assign n1246 = n1245 ^ n319 ^ 1'b0 ;
  assign n1247 = n363 ^ n286 ^ 1'b0 ;
  assign n1248 = n675 | n1247 ;
  assign n1249 = x7 | n1248 ;
  assign n1250 = n593 & ~n700 ;
  assign n1251 = n367 | n1250 ;
  assign n1252 = n1251 ^ n445 ^ 1'b0 ;
  assign n1253 = n994 ^ n284 ^ x28 ;
  assign n1254 = n944 & ~n1253 ;
  assign n1255 = n1252 & n1254 ;
  assign n1256 = n993 ^ n640 ^ 1'b0 ;
  assign n1257 = x7 & x78 ;
  assign n1258 = ~x133 & n1257 ;
  assign n1259 = n1258 ^ n411 ^ x26 ;
  assign n1260 = n365 & n1259 ;
  assign n1261 = ( n363 & ~n1129 ) | ( n363 & n1260 ) | ( ~n1129 & n1260 ) ;
  assign n1262 = n1019 ^ n338 ^ 1'b0 ;
  assign n1263 = n1261 | n1262 ;
  assign n1264 = n1263 ^ n527 ^ 1'b0 ;
  assign n1265 = ~x169 & n1117 ;
  assign n1266 = n847 ^ n729 ^ x228 ;
  assign n1267 = n686 ^ x171 ^ 1'b0 ;
  assign n1268 = n275 & n1267 ;
  assign n1269 = n671 ^ n263 ^ 1'b0 ;
  assign n1270 = n1268 & ~n1269 ;
  assign n1271 = ( n590 & n915 ) | ( n590 & ~n1010 ) | ( n915 & ~n1010 ) ;
  assign n1272 = x123 ^ x67 ^ 1'b0 ;
  assign n1273 = ( x232 & n770 ) | ( x232 & ~n1055 ) | ( n770 & ~n1055 ) ;
  assign n1274 = x251 & ~x254 ;
  assign n1275 = n963 ^ n873 ^ n734 ;
  assign n1276 = ~n1142 & n1275 ;
  assign n1277 = n612 & n1276 ;
  assign n1278 = n683 ^ x185 ^ 1'b0 ;
  assign n1279 = n716 ^ n702 ^ x42 ;
  assign n1280 = n1279 ^ n1235 ^ 1'b0 ;
  assign n1281 = ~n545 & n1280 ;
  assign n1284 = n944 ^ n660 ^ x114 ;
  assign n1282 = ~n371 & n392 ;
  assign n1283 = ~n269 & n1282 ;
  assign n1285 = n1284 ^ n1283 ^ n550 ;
  assign n1286 = n1281 & n1285 ;
  assign n1287 = ( x170 & ~x190 ) | ( x170 & n840 ) | ( ~x190 & n840 ) ;
  assign n1288 = ( ~x187 & x198 ) | ( ~x187 & n608 ) | ( x198 & n608 ) ;
  assign n1289 = n404 | n1288 ;
  assign n1290 = ~n957 & n1289 ;
  assign n1291 = n856 & n1290 ;
  assign n1292 = n1287 | n1291 ;
  assign n1293 = n1292 ^ n301 ^ 1'b0 ;
  assign n1294 = x89 ^ x19 ^ 1'b0 ;
  assign n1295 = x61 & n1294 ;
  assign n1296 = x191 & n1295 ;
  assign n1297 = x216 ^ x145 ^ 1'b0 ;
  assign n1298 = n1027 & n1297 ;
  assign n1299 = n301 ^ x104 ^ 1'b0 ;
  assign n1300 = x203 & ~n1299 ;
  assign n1301 = ~n535 & n1300 ;
  assign n1302 = n1301 ^ x20 ^ 1'b0 ;
  assign n1303 = ~n815 & n1197 ;
  assign n1304 = n1303 ^ n500 ^ 1'b0 ;
  assign n1306 = n1096 ^ n858 ^ x56 ;
  assign n1305 = x47 & ~n480 ;
  assign n1307 = n1306 ^ n1305 ^ 1'b0 ;
  assign n1308 = n780 | n1307 ;
  assign n1309 = ~n758 & n1234 ;
  assign n1310 = n1309 ^ n531 ^ 1'b0 ;
  assign n1311 = x169 & x238 ;
  assign n1312 = n787 | n1311 ;
  assign n1313 = ( x205 & n930 ) | ( x205 & n1312 ) | ( n930 & n1312 ) ;
  assign n1314 = n781 & ~n818 ;
  assign n1315 = n1025 ^ n543 ^ 1'b0 ;
  assign n1316 = n273 ^ n265 ^ 1'b0 ;
  assign n1317 = n344 & ~n1316 ;
  assign n1318 = x72 & n1317 ;
  assign n1319 = ~n932 & n1318 ;
  assign n1320 = x1 & ~n1319 ;
  assign n1321 = ~x58 & n1320 ;
  assign n1323 = n500 & n1209 ;
  assign n1324 = n1093 | n1323 ;
  assign n1322 = n995 & n1072 ;
  assign n1325 = n1324 ^ n1322 ^ 1'b0 ;
  assign n1327 = x244 ^ x42 ^ 1'b0 ;
  assign n1326 = n337 | n1059 ;
  assign n1328 = n1327 ^ n1326 ^ 1'b0 ;
  assign n1329 = n832 & ~n1037 ;
  assign n1330 = ~n598 & n1329 ;
  assign n1331 = n752 ^ x15 ^ 1'b0 ;
  assign n1332 = ~n1330 & n1331 ;
  assign n1333 = n1332 ^ n460 ^ 1'b0 ;
  assign n1334 = x70 & ~n1333 ;
  assign n1335 = n639 ^ x193 ^ 1'b0 ;
  assign n1336 = x26 & ~n1335 ;
  assign n1337 = n1336 ^ n617 ^ 1'b0 ;
  assign n1338 = ~n465 & n882 ;
  assign n1339 = ~n1337 & n1338 ;
  assign n1340 = ( x206 & ~x208 ) | ( x206 & n737 ) | ( ~x208 & n737 ) ;
  assign n1341 = x105 & n1340 ;
  assign n1342 = ~n519 & n1341 ;
  assign n1343 = n849 ^ n793 ^ x22 ;
  assign n1344 = n673 ^ n647 ^ 1'b0 ;
  assign n1345 = ~n944 & n1344 ;
  assign n1346 = n1343 & n1345 ;
  assign n1347 = n1346 ^ n688 ^ n371 ;
  assign n1348 = ~n1342 & n1347 ;
  assign n1349 = n1235 ^ n732 ^ 1'b0 ;
  assign n1350 = n446 ^ x79 ^ 1'b0 ;
  assign n1351 = n913 ^ n832 ^ x60 ;
  assign n1352 = n737 & ~n1351 ;
  assign n1353 = n1352 ^ n413 ^ 1'b0 ;
  assign n1354 = x98 ^ x92 ^ 1'b0 ;
  assign n1355 = n1354 ^ n1196 ^ 1'b0 ;
  assign n1356 = ( ~x102 & n980 ) | ( ~x102 & n1355 ) | ( n980 & n1355 ) ;
  assign n1357 = x171 & n652 ;
  assign n1358 = n1357 ^ n513 ^ 1'b0 ;
  assign n1359 = x79 & ~n1358 ;
  assign n1360 = n1359 ^ n530 ^ 1'b0 ;
  assign n1361 = n1085 | n1360 ;
  assign n1362 = n1361 ^ n1027 ^ 1'b0 ;
  assign n1363 = n1036 & ~n1059 ;
  assign n1364 = n1120 & n1363 ;
  assign n1365 = n1364 ^ n818 ^ 1'b0 ;
  assign n1366 = ( x225 & ~x229 ) | ( x225 & n312 ) | ( ~x229 & n312 ) ;
  assign n1367 = n755 & ~n1366 ;
  assign n1368 = ~x169 & n1367 ;
  assign n1369 = ~n1003 & n1266 ;
  assign n1370 = ~x86 & n1369 ;
  assign n1371 = x26 & ~n972 ;
  assign n1372 = n1371 ^ n256 ^ 1'b0 ;
  assign n1373 = n1372 ^ x144 ^ 1'b0 ;
  assign n1377 = ~x195 & n519 ;
  assign n1374 = n1079 ^ x11 ^ 1'b0 ;
  assign n1375 = n942 ^ n485 ^ 1'b0 ;
  assign n1376 = n1374 & ~n1375 ;
  assign n1378 = n1377 ^ n1376 ^ n459 ;
  assign n1379 = x236 & ~n966 ;
  assign n1380 = n1379 ^ n545 ^ 1'b0 ;
  assign n1381 = n1093 ^ n936 ^ n872 ;
  assign n1382 = ~x133 & n1284 ;
  assign n1383 = x220 & ~n1382 ;
  assign n1384 = ~n1310 & n1383 ;
  assign n1385 = n770 | n1306 ;
  assign n1386 = n1385 ^ n666 ^ 1'b0 ;
  assign n1387 = n614 & n829 ;
  assign n1388 = x125 & ~n1387 ;
  assign n1389 = n907 ^ x57 ^ 1'b0 ;
  assign n1390 = n921 & n1389 ;
  assign n1391 = n433 & n1239 ;
  assign n1392 = n1391 ^ n694 ^ 1'b0 ;
  assign n1393 = n983 ^ n311 ^ x32 ;
  assign n1394 = ( x144 & n1023 ) | ( x144 & ~n1393 ) | ( n1023 & ~n1393 ) ;
  assign n1395 = ( ~x151 & x201 ) | ( ~x151 & n764 ) | ( x201 & n764 ) ;
  assign n1396 = x243 ^ x234 ^ x15 ;
  assign n1397 = ( n1098 & n1336 ) | ( n1098 & n1396 ) | ( n1336 & n1396 ) ;
  assign n1399 = x12 & ~n319 ;
  assign n1400 = ~x252 & n1399 ;
  assign n1398 = x31 & n583 ;
  assign n1401 = n1400 ^ n1398 ^ 1'b0 ;
  assign n1402 = n1177 ^ n1097 ^ 1'b0 ;
  assign n1403 = n1401 & n1402 ;
  assign n1404 = ( x65 & ~x229 ) | ( x65 & n298 ) | ( ~x229 & n298 ) ;
  assign n1405 = n431 ^ n258 ^ 1'b0 ;
  assign n1406 = x98 & n1405 ;
  assign n1407 = n1404 & n1406 ;
  assign n1408 = x105 & x254 ;
  assign n1409 = ~n1038 & n1408 ;
  assign n1410 = n1162 | n1409 ;
  assign n1411 = n1407 & ~n1410 ;
  assign n1412 = n960 ^ n877 ^ 1'b0 ;
  assign n1413 = n1247 | n1412 ;
  assign n1414 = x128 & ~n294 ;
  assign n1415 = n1414 ^ n608 ^ 1'b0 ;
  assign n1416 = n1064 | n1415 ;
  assign n1417 = x26 & ~n351 ;
  assign n1418 = n1417 ^ n513 ^ 1'b0 ;
  assign n1419 = ( x183 & ~x254 ) | ( x183 & n1418 ) | ( ~x254 & n1418 ) ;
  assign n1420 = n1419 ^ n363 ^ 1'b0 ;
  assign n1421 = ~n1019 & n1420 ;
  assign n1422 = ~n1416 & n1421 ;
  assign n1423 = n1413 & n1422 ;
  assign n1424 = x179 & n749 ;
  assign n1425 = n1423 & n1424 ;
  assign n1426 = n300 | n661 ;
  assign n1427 = x58 | n1426 ;
  assign n1428 = ~n721 & n1337 ;
  assign n1429 = ~n1427 & n1428 ;
  assign n1430 = ~n498 & n1429 ;
  assign n1431 = n671 & n723 ;
  assign n1432 = ( x15 & ~x133 ) | ( x15 & n1431 ) | ( ~x133 & n1431 ) ;
  assign n1433 = n1406 ^ n926 ^ 1'b0 ;
  assign n1434 = n1433 ^ x95 ^ 1'b0 ;
  assign n1435 = x217 & n1434 ;
  assign n1436 = n732 & ~n797 ;
  assign n1437 = n1436 ^ x50 ^ 1'b0 ;
  assign n1438 = n1437 ^ n895 ^ 1'b0 ;
  assign n1439 = n565 & n1438 ;
  assign n1440 = n643 ^ n606 ^ 1'b0 ;
  assign n1441 = x171 & n1440 ;
  assign n1442 = ~n1439 & n1441 ;
  assign n1443 = ~x177 & n1184 ;
  assign n1444 = n1443 ^ n906 ^ 1'b0 ;
  assign n1450 = n700 ^ n698 ^ n296 ;
  assign n1445 = n614 | n944 ;
  assign n1446 = n1445 ^ n898 ^ 1'b0 ;
  assign n1447 = x200 & ~n1446 ;
  assign n1448 = n1447 ^ n509 ^ 1'b0 ;
  assign n1449 = x101 & n1448 ;
  assign n1451 = n1450 ^ n1449 ^ 1'b0 ;
  assign n1452 = n399 ^ x48 ^ 1'b0 ;
  assign n1453 = n277 & n1452 ;
  assign n1454 = n570 & n1177 ;
  assign n1455 = ~n1453 & n1454 ;
  assign n1456 = n1455 ^ n1360 ^ 1'b0 ;
  assign n1457 = n306 & n1456 ;
  assign n1458 = n939 ^ x118 ^ 1'b0 ;
  assign n1459 = n562 ^ n508 ^ n432 ;
  assign n1460 = n1458 | n1459 ;
  assign n1461 = n451 | n642 ;
  assign n1462 = n1344 | n1461 ;
  assign n1463 = n274 & n860 ;
  assign n1464 = n1463 ^ n1205 ^ 1'b0 ;
  assign n1465 = n1464 ^ n1052 ^ 1'b0 ;
  assign n1466 = ~n492 & n1465 ;
  assign n1467 = x140 & n863 ;
  assign n1468 = ~n785 & n1467 ;
  assign n1469 = ~n1466 & n1468 ;
  assign n1470 = ~x167 & n716 ;
  assign n1471 = x196 & n854 ;
  assign n1472 = n1467 ^ n890 ^ 1'b0 ;
  assign n1475 = n361 & n392 ;
  assign n1476 = n863 ^ n657 ^ 1'b0 ;
  assign n1477 = n832 & ~n1476 ;
  assign n1478 = n1475 & ~n1477 ;
  assign n1479 = n1478 ^ n553 ^ 1'b0 ;
  assign n1473 = ( x253 & ~n404 ) | ( x253 & n1253 ) | ( ~n404 & n1253 ) ;
  assign n1474 = n1473 ^ n879 ^ n657 ;
  assign n1480 = n1479 ^ n1474 ^ 1'b0 ;
  assign n1482 = n351 ^ x253 ^ 1'b0 ;
  assign n1483 = n751 & ~n1482 ;
  assign n1481 = x16 & ~n776 ;
  assign n1484 = n1483 ^ n1481 ^ n300 ;
  assign n1485 = n496 ^ x1 ^ 1'b0 ;
  assign n1486 = x19 & ~n1485 ;
  assign n1487 = ~n1068 & n1486 ;
  assign n1488 = ~n1377 & n1487 ;
  assign n1489 = x7 & n800 ;
  assign n1490 = x15 & n587 ;
  assign n1491 = n443 | n552 ;
  assign n1492 = ~n800 & n1491 ;
  assign n1493 = ~n1490 & n1492 ;
  assign n1494 = n354 & n1017 ;
  assign n1495 = n1494 ^ n1177 ^ 1'b0 ;
  assign n1496 = n1495 ^ n666 ^ n347 ;
  assign n1497 = n1486 & n1496 ;
  assign n1498 = n1497 ^ n563 ^ 1'b0 ;
  assign n1499 = ~n535 & n1498 ;
  assign n1500 = x17 | n533 ;
  assign n1501 = x55 ^ x50 ^ 1'b0 ;
  assign n1502 = n1501 ^ n263 ^ 1'b0 ;
  assign n1503 = n1502 ^ n672 ^ 1'b0 ;
  assign n1504 = ~n1446 & n1503 ;
  assign n1505 = n1504 ^ n314 ^ 1'b0 ;
  assign n1506 = n1500 & n1505 ;
  assign n1507 = n1506 ^ x172 ^ 1'b0 ;
  assign n1508 = n1184 & n1507 ;
  assign n1509 = ~n1365 & n1508 ;
  assign n1512 = x128 ^ x103 ^ x43 ;
  assign n1513 = n900 ^ n447 ^ 1'b0 ;
  assign n1514 = n1512 | n1513 ;
  assign n1510 = x195 ^ x178 ^ x87 ;
  assign n1511 = n1068 | n1510 ;
  assign n1515 = n1514 ^ n1511 ^ 1'b0 ;
  assign n1516 = x215 & ~n341 ;
  assign n1517 = ~x23 & n1516 ;
  assign n1518 = x222 | n1517 ;
  assign n1519 = ( ~n420 & n1082 ) | ( ~n420 & n1182 ) | ( n1082 & n1182 ) ;
  assign n1520 = ~x55 & n809 ;
  assign n1521 = n1415 ^ n520 ^ 1'b0 ;
  assign n1523 = x42 & ~n488 ;
  assign n1524 = n1523 ^ n439 ^ 1'b0 ;
  assign n1522 = n304 | n1413 ;
  assign n1525 = n1524 ^ n1522 ^ 1'b0 ;
  assign n1527 = x91 ^ x54 ^ 1'b0 ;
  assign n1526 = ~x153 & x199 ;
  assign n1528 = n1527 ^ n1526 ^ 1'b0 ;
  assign n1529 = ~n840 & n1295 ;
  assign n1530 = ~n456 & n1529 ;
  assign n1531 = ~n745 & n842 ;
  assign n1532 = n1531 ^ n1311 ^ 1'b0 ;
  assign n1533 = n1137 ^ n407 ^ 1'b0 ;
  assign n1534 = n565 & ~n1132 ;
  assign n1535 = n1534 ^ n1277 ^ 1'b0 ;
  assign n1536 = x242 & ~n294 ;
  assign n1537 = ~n529 & n1536 ;
  assign n1538 = n1537 ^ x243 ^ 1'b0 ;
  assign n1539 = n1365 ^ n1246 ^ 1'b0 ;
  assign n1540 = n1213 & ~n1539 ;
  assign n1541 = n465 ^ n358 ^ n328 ;
  assign n1542 = n1541 ^ n883 ^ 1'b0 ;
  assign n1543 = x194 & ~n1542 ;
  assign n1544 = n530 ^ x48 ^ 1'b0 ;
  assign n1545 = n1543 & n1544 ;
  assign n1546 = n1545 ^ x158 ^ 1'b0 ;
  assign n1547 = n1122 | n1152 ;
  assign n1548 = ( ~x65 & x183 ) | ( ~x65 & n1464 ) | ( x183 & n1464 ) ;
  assign n1549 = x200 & ~n1548 ;
  assign n1550 = n1549 ^ n745 ^ 1'b0 ;
  assign n1551 = ~n734 & n1396 ;
  assign n1552 = n1550 & n1551 ;
  assign n1553 = n1552 ^ n845 ^ 1'b0 ;
  assign n1554 = n946 ^ x2 ^ 1'b0 ;
  assign n1555 = x156 & n1554 ;
  assign n1556 = n1555 ^ n465 ^ 1'b0 ;
  assign n1557 = x7 & ~n1556 ;
  assign n1558 = ( ~x76 & n508 ) | ( ~x76 & n987 ) | ( n508 & n987 ) ;
  assign n1559 = ( x104 & n320 ) | ( x104 & ~n898 ) | ( n320 & ~n898 ) ;
  assign n1560 = n1559 ^ n1446 ^ 1'b0 ;
  assign n1561 = n1558 | n1560 ;
  assign n1562 = x78 & ~n502 ;
  assign n1563 = n1562 ^ n1401 ^ 1'b0 ;
  assign n1564 = n1541 ^ n976 ^ 1'b0 ;
  assign n1565 = n909 ^ x204 ^ 1'b0 ;
  assign n1566 = n1190 ^ x50 ^ 1'b0 ;
  assign n1567 = n970 & n1566 ;
  assign n1568 = n569 ^ n337 ^ 1'b0 ;
  assign n1569 = ~n966 & n1568 ;
  assign n1570 = n1569 ^ n1260 ^ n323 ;
  assign n1571 = n553 ^ x235 ^ 1'b0 ;
  assign n1572 = ( n418 & n1570 ) | ( n418 & n1571 ) | ( n1570 & n1571 ) ;
  assign n1585 = n922 ^ n289 ^ 1'b0 ;
  assign n1580 = ~n537 & n1317 ;
  assign n1581 = n1580 ^ n333 ^ 1'b0 ;
  assign n1573 = x95 & x169 ;
  assign n1574 = ~x224 & n1573 ;
  assign n1575 = n652 ^ n304 ^ x178 ;
  assign n1576 = n1575 ^ n526 ^ 1'b0 ;
  assign n1577 = x245 & n1576 ;
  assign n1578 = ~n1574 & n1577 ;
  assign n1579 = n743 & n1578 ;
  assign n1582 = n1581 ^ n1579 ^ 1'b0 ;
  assign n1583 = n1582 ^ n504 ^ 1'b0 ;
  assign n1584 = n755 & n1583 ;
  assign n1586 = n1585 ^ n1584 ^ 1'b0 ;
  assign n1587 = ~n1572 & n1586 ;
  assign n1593 = n340 ^ x195 ^ x113 ;
  assign n1588 = x108 & ~n1127 ;
  assign n1589 = ~x165 & n1588 ;
  assign n1590 = n686 ^ x12 ^ x1 ;
  assign n1591 = n1590 ^ n933 ^ 1'b0 ;
  assign n1592 = ~n1589 & n1591 ;
  assign n1594 = n1593 ^ n1592 ^ n562 ;
  assign n1595 = n1594 ^ n1298 ^ n354 ;
  assign n1596 = x115 & ~n489 ;
  assign n1597 = n1596 ^ n1390 ^ n880 ;
  assign n1598 = n379 ^ x71 ^ 1'b0 ;
  assign n1599 = x21 & x192 ;
  assign n1600 = n1598 & n1599 ;
  assign n1601 = ~n294 & n536 ;
  assign n1602 = n1601 ^ x38 ^ 1'b0 ;
  assign n1603 = n1288 & n1602 ;
  assign n1604 = n975 & n1603 ;
  assign n1607 = n314 & n443 ;
  assign n1608 = n1607 ^ x59 ^ 1'b0 ;
  assign n1609 = n1608 ^ n338 ^ 1'b0 ;
  assign n1610 = n647 & ~n1609 ;
  assign n1605 = n467 & ~n1263 ;
  assign n1606 = n666 & ~n1605 ;
  assign n1611 = n1610 ^ n1606 ^ 1'b0 ;
  assign n1612 = n327 & n1184 ;
  assign n1613 = n634 & n1232 ;
  assign n1614 = x44 & x96 ;
  assign n1615 = n711 & n1614 ;
  assign n1616 = n1615 ^ n1387 ^ n874 ;
  assign n1617 = n1254 | n1616 ;
  assign n1618 = n1617 ^ n1324 ^ 1'b0 ;
  assign n1619 = ~x237 & n459 ;
  assign n1620 = n438 | n481 ;
  assign n1621 = x120 ^ x112 ^ 1'b0 ;
  assign n1622 = x0 & n1621 ;
  assign n1623 = x64 & x220 ;
  assign n1624 = ~n1622 & n1623 ;
  assign n1625 = ( n1049 & n1620 ) | ( n1049 & n1624 ) | ( n1620 & n1624 ) ;
  assign n1626 = n1625 ^ n1508 ^ 1'b0 ;
  assign n1627 = n393 & n443 ;
  assign n1628 = n327 & n1627 ;
  assign n1629 = ~n643 & n1628 ;
  assign n1630 = n727 | n1629 ;
  assign n1631 = n623 ^ n511 ^ n494 ;
  assign n1632 = n718 ^ n258 ^ 1'b0 ;
  assign n1633 = n1631 & n1632 ;
  assign n1634 = n546 & ~n734 ;
  assign n1635 = ~n1633 & n1634 ;
  assign n1636 = n485 ^ x213 ^ 1'b0 ;
  assign n1637 = n1155 & ~n1636 ;
  assign n1638 = n1136 ^ x234 ^ 1'b0 ;
  assign n1639 = x65 & ~n1638 ;
  assign n1640 = ~n328 & n1639 ;
  assign n1641 = n1640 ^ n968 ^ 1'b0 ;
  assign n1642 = n1641 ^ n256 ^ 1'b0 ;
  assign n1643 = n1637 & ~n1642 ;
  assign n1644 = x135 & ~n1590 ;
  assign n1645 = ~n449 & n1644 ;
  assign n1646 = ( n803 & ~n897 ) | ( n803 & n1645 ) | ( ~n897 & n1645 ) ;
  assign n1647 = x27 & n1046 ;
  assign n1648 = n1647 ^ n462 ^ 1'b0 ;
  assign n1649 = ~n263 & n399 ;
  assign n1650 = n328 & n1649 ;
  assign n1651 = x19 & ~n1650 ;
  assign n1652 = x172 & x229 ;
  assign n1653 = n1652 ^ x31 ^ 1'b0 ;
  assign n1654 = n1653 ^ x105 ^ 1'b0 ;
  assign n1655 = n585 | n1654 ;
  assign n1656 = n805 & ~n1655 ;
  assign n1657 = n963 & n1656 ;
  assign n1658 = n1557 ^ n960 ^ 1'b0 ;
  assign n1659 = x219 ^ x185 ^ 1'b0 ;
  assign n1660 = n277 & n1659 ;
  assign n1661 = n905 ^ n560 ^ 1'b0 ;
  assign n1662 = n1660 & n1661 ;
  assign n1663 = ~x117 & n1662 ;
  assign n1664 = n480 ^ x45 ^ 1'b0 ;
  assign n1665 = x149 & ~n1664 ;
  assign n1666 = n530 ^ n463 ^ 1'b0 ;
  assign n1667 = n1666 ^ x94 ^ 1'b0 ;
  assign n1668 = n1665 & n1667 ;
  assign n1669 = n1668 ^ n1339 ^ 1'b0 ;
  assign n1670 = x200 & ~n1250 ;
  assign n1671 = ~x58 & n1670 ;
  assign n1672 = n292 | n1671 ;
  assign n1673 = n1672 ^ n1069 ^ 1'b0 ;
  assign n1674 = n413 ^ x107 ^ x84 ;
  assign n1675 = n380 & ~n1674 ;
  assign n1676 = n415 | n1022 ;
  assign n1677 = n1676 ^ x61 ^ 1'b0 ;
  assign n1678 = n1677 ^ n1214 ^ n1126 ;
  assign n1679 = n1675 & ~n1678 ;
  assign n1682 = x35 & x175 ;
  assign n1683 = ~n311 & n1682 ;
  assign n1684 = n387 | n1683 ;
  assign n1685 = n1176 & ~n1684 ;
  assign n1686 = n1685 ^ n320 ^ x197 ;
  assign n1680 = ~n548 & n556 ;
  assign n1681 = x169 | n1680 ;
  assign n1687 = n1686 ^ n1681 ^ n900 ;
  assign n1688 = ~n471 & n1687 ;
  assign n1689 = n1075 ^ x106 ^ 1'b0 ;
  assign n1690 = n1689 ^ n957 ^ x212 ;
  assign n1691 = ( n449 & ~n673 ) | ( n449 & n1026 ) | ( ~n673 & n1026 ) ;
  assign n1692 = n1403 | n1691 ;
  assign n1693 = ( x201 & n983 ) | ( x201 & ~n1692 ) | ( n983 & ~n1692 ) ;
  assign n1694 = n429 & ~n1687 ;
  assign n1695 = n952 ^ x251 ^ 1'b0 ;
  assign n1696 = x163 & ~n1000 ;
  assign n1697 = n1696 ^ n443 ^ 1'b0 ;
  assign n1698 = n1697 ^ n1086 ^ x210 ;
  assign n1699 = n698 | n1698 ;
  assign n1700 = n1699 ^ n358 ^ 1'b0 ;
  assign n1701 = ( ~x101 & n1314 ) | ( ~x101 & n1700 ) | ( n1314 & n1700 ) ;
  assign n1702 = n921 ^ n322 ^ 1'b0 ;
  assign n1703 = n1702 ^ n388 ^ 1'b0 ;
  assign n1704 = n760 & n1406 ;
  assign n1705 = n1261 & n1704 ;
  assign n1706 = ( ~n283 & n1144 ) | ( ~n283 & n1705 ) | ( n1144 & n1705 ) ;
  assign n1710 = x159 & n980 ;
  assign n1711 = ~n485 & n1710 ;
  assign n1712 = n1711 ^ n537 ^ n463 ;
  assign n1707 = n471 & ~n751 ;
  assign n1708 = n459 | n706 ;
  assign n1709 = ( n1421 & n1707 ) | ( n1421 & ~n1708 ) | ( n1707 & ~n1708 ) ;
  assign n1713 = n1712 ^ n1709 ^ n768 ;
  assign n1715 = n646 ^ n393 ^ 1'b0 ;
  assign n1714 = ~n486 & n1297 ;
  assign n1716 = n1715 ^ n1714 ^ 1'b0 ;
  assign n1717 = n1354 ^ n1176 ^ 1'b0 ;
  assign n1718 = n739 & ~n1717 ;
  assign n1719 = ~n1716 & n1718 ;
  assign n1720 = n1277 & ~n1474 ;
  assign n1721 = x57 & ~n873 ;
  assign n1722 = n1721 ^ n1358 ^ 1'b0 ;
  assign n1723 = n598 & n1722 ;
  assign n1724 = n889 & n1723 ;
  assign n1725 = n1284 ^ n498 ^ n410 ;
  assign n1726 = ~n279 & n840 ;
  assign n1727 = n1726 ^ x126 ^ 1'b0 ;
  assign n1728 = x78 & ~x202 ;
  assign n1729 = n1728 ^ n1264 ^ 1'b0 ;
  assign n1730 = n1019 ^ n289 ^ 1'b0 ;
  assign n1731 = x10 | n1103 ;
  assign n1732 = n380 & ~n785 ;
  assign n1733 = n1732 ^ n1237 ^ n1210 ;
  assign n1736 = x62 ^ x57 ^ 1'b0 ;
  assign n1734 = x230 & n1457 ;
  assign n1735 = ~n1006 & n1734 ;
  assign n1737 = n1736 ^ n1735 ^ n1528 ;
  assign n1738 = n1686 ^ x243 ^ 1'b0 ;
  assign n1739 = n1091 & ~n1738 ;
  assign n1740 = n1739 ^ x142 ^ 1'b0 ;
  assign n1741 = ~n304 & n1740 ;
  assign n1742 = n1270 ^ n622 ^ 1'b0 ;
  assign n1743 = ~n712 & n1592 ;
  assign n1744 = n1397 & n1743 ;
  assign n1745 = n395 & n874 ;
  assign n1746 = n1745 ^ n787 ^ 1'b0 ;
  assign n1747 = n379 | n1306 ;
  assign n1748 = n1747 ^ n1559 ^ 1'b0 ;
  assign n1754 = n967 ^ n456 ^ 1'b0 ;
  assign n1755 = n1400 | n1754 ;
  assign n1749 = n633 ^ n366 ^ 1'b0 ;
  assign n1750 = n842 & ~n1749 ;
  assign n1751 = n954 | n1302 ;
  assign n1752 = n1751 ^ n627 ^ 1'b0 ;
  assign n1753 = ( x95 & n1750 ) | ( x95 & ~n1752 ) | ( n1750 & ~n1752 ) ;
  assign n1756 = n1755 ^ n1753 ^ 1'b0 ;
  assign n1757 = n1339 | n1756 ;
  assign n1758 = n727 & ~n1241 ;
  assign n1759 = n781 ^ n531 ^ 1'b0 ;
  assign n1760 = n860 & n1759 ;
  assign n1761 = n1760 ^ n1172 ^ 1'b0 ;
  assign n1762 = n1761 ^ n1596 ^ 1'b0 ;
  assign n1763 = ( x23 & ~x56 ) | ( x23 & n1613 ) | ( ~x56 & n1613 ) ;
  assign n1764 = n1033 & ~n1306 ;
  assign n1766 = n259 ^ x155 ^ 1'b0 ;
  assign n1767 = ( x102 & ~n308 ) | ( x102 & n1766 ) | ( ~n308 & n1766 ) ;
  assign n1768 = n1767 ^ n622 ^ 1'b0 ;
  assign n1765 = ~n294 & n1075 ;
  assign n1769 = n1768 ^ n1765 ^ 1'b0 ;
  assign n1770 = n438 | n1098 ;
  assign n1771 = n315 & ~n1770 ;
  assign n1772 = n1771 ^ n1079 ^ x187 ;
  assign n1773 = n1772 ^ n952 ^ 1'b0 ;
  assign n1774 = n1773 ^ n935 ^ 1'b0 ;
  assign n1775 = ~n1769 & n1774 ;
  assign n1776 = x123 & n380 ;
  assign n1777 = n381 & n449 ;
  assign n1778 = x3 & ~n1351 ;
  assign n1779 = n1778 ^ n381 ^ 1'b0 ;
  assign n1780 = x163 & n1779 ;
  assign n1781 = n1780 ^ n591 ^ 1'b0 ;
  assign n1785 = ( x155 & ~x166 ) | ( x155 & n842 ) | ( ~x166 & n842 ) ;
  assign n1786 = n1785 ^ n818 ^ x141 ;
  assign n1782 = ( x86 & x91 ) | ( x86 & n431 ) | ( x91 & n431 ) ;
  assign n1783 = n1782 ^ n679 ^ 1'b0 ;
  assign n1784 = n1783 ^ n719 ^ 1'b0 ;
  assign n1787 = n1786 ^ n1784 ^ 1'b0 ;
  assign n1788 = n322 | n1787 ;
  assign n1789 = x132 | n797 ;
  assign n1790 = n1702 ^ n1009 ^ 1'b0 ;
  assign n1791 = n1144 | n1790 ;
  assign n1792 = n1789 & ~n1791 ;
  assign n1796 = x20 & x123 ;
  assign n1797 = n1796 ^ x248 ^ 1'b0 ;
  assign n1793 = x16 | n723 ;
  assign n1794 = n1070 & n1793 ;
  assign n1795 = n1794 ^ x73 ^ 1'b0 ;
  assign n1798 = n1797 ^ n1795 ^ n1697 ;
  assign n1799 = n781 ^ n570 ^ 1'b0 ;
  assign n1800 = n347 | n1799 ;
  assign n1802 = n274 & ~n441 ;
  assign n1801 = n867 ^ n329 ^ 1'b0 ;
  assign n1803 = n1802 ^ n1801 ^ n622 ;
  assign n1804 = ( n471 & ~n1800 ) | ( n471 & n1803 ) | ( ~n1800 & n1803 ) ;
  assign n1805 = n882 & ~n1567 ;
  assign n1806 = ( ~x22 & n417 ) | ( ~x22 & n987 ) | ( n417 & n987 ) ;
  assign n1807 = n505 & n1618 ;
  assign n1808 = ( x177 & ~x206 ) | ( x177 & n727 ) | ( ~x206 & n727 ) ;
  assign n1809 = ( n597 & ~n1685 ) | ( n597 & n1808 ) | ( ~n1685 & n1808 ) ;
  assign n1810 = x115 & n491 ;
  assign n1811 = n631 & n1810 ;
  assign n1812 = n886 ^ n511 ^ 1'b0 ;
  assign n1813 = ~n1228 & n1812 ;
  assign n1814 = ( n1259 & n1811 ) | ( n1259 & n1813 ) | ( n1811 & n1813 ) ;
  assign n1815 = ~n822 & n1814 ;
  assign n1816 = ~n1809 & n1815 ;
  assign n1817 = n549 ^ x167 ^ 1'b0 ;
  assign n1818 = x158 & n1817 ;
  assign n1819 = n1818 ^ n1722 ^ 1'b0 ;
  assign n1820 = x245 & ~n1056 ;
  assign n1821 = ~n1242 & n1820 ;
  assign n1822 = n1821 ^ n1569 ^ 1'b0 ;
  assign n1823 = n365 & n1256 ;
  assign n1824 = x37 | n1823 ;
  assign n1825 = n1824 ^ n1062 ^ 1'b0 ;
  assign n1826 = ~n1822 & n1825 ;
  assign n1827 = n854 ^ n851 ^ n683 ;
  assign n1828 = ~n476 & n559 ;
  assign n1829 = x222 & n1828 ;
  assign n1830 = n1829 ^ n1598 ^ 1'b0 ;
  assign n1831 = ~n1616 & n1703 ;
  assign n1833 = ~x180 & n411 ;
  assign n1832 = n1115 ^ n970 ^ 1'b0 ;
  assign n1834 = n1833 ^ n1832 ^ 1'b0 ;
  assign n1835 = ~n1464 & n1834 ;
  assign n1836 = ( n709 & ~n1336 ) | ( n709 & n1418 ) | ( ~n1336 & n1418 ) ;
  assign n1837 = n1400 ^ x202 ^ 1'b0 ;
  assign n1838 = n1837 ^ n727 ^ 1'b0 ;
  assign n1839 = x80 & ~n768 ;
  assign n1840 = ~n490 & n1839 ;
  assign n1841 = x12 & ~n1840 ;
  assign n1842 = n1841 ^ n736 ^ 1'b0 ;
  assign n1843 = n399 & ~n1842 ;
  assign n1845 = n1801 ^ n529 ^ 1'b0 ;
  assign n1846 = ~n349 & n1845 ;
  assign n1847 = ( x207 & n650 ) | ( x207 & ~n1069 ) | ( n650 & ~n1069 ) ;
  assign n1848 = n1847 ^ n939 ^ 1'b0 ;
  assign n1849 = n1848 ^ n1832 ^ 1'b0 ;
  assign n1850 = n1846 & n1849 ;
  assign n1844 = n284 & ~n963 ;
  assign n1851 = n1850 ^ n1844 ^ 1'b0 ;
  assign n1852 = n449 & n1783 ;
  assign n1853 = ~n1499 & n1852 ;
  assign n1854 = n1026 | n1277 ;
  assign n1855 = n1297 | n1854 ;
  assign n1856 = n954 ^ n463 ^ 1'b0 ;
  assign n1857 = x56 & ~n1856 ;
  assign n1858 = n1857 ^ x252 ^ 1'b0 ;
  assign n1859 = n1619 ^ n1504 ^ 1'b0 ;
  assign n1860 = ~n1858 & n1859 ;
  assign n1861 = n1270 ^ n1259 ^ 1'b0 ;
  assign n1862 = ~x165 & n1861 ;
  assign n1863 = ( x200 & n261 ) | ( x200 & n1862 ) | ( n261 & n1862 ) ;
  assign n1865 = ( ~n388 & n605 ) | ( ~n388 & n1311 ) | ( n605 & n1311 ) ;
  assign n1864 = x75 & n456 ;
  assign n1866 = n1865 ^ n1864 ^ 1'b0 ;
  assign n1867 = n937 & n988 ;
  assign n1868 = n1867 ^ n1823 ^ 1'b0 ;
  assign n1869 = ( x77 & n822 ) | ( x77 & ~n1136 ) | ( n822 & ~n1136 ) ;
  assign n1870 = n1259 ^ n317 ^ x249 ;
  assign n1871 = n1869 & n1870 ;
  assign n1872 = ( ~x216 & n673 ) | ( ~x216 & n1665 ) | ( n673 & n1665 ) ;
  assign n1873 = n1872 ^ n1354 ^ 1'b0 ;
  assign n1874 = ( x167 & ~n760 ) | ( x167 & n809 ) | ( ~n760 & n809 ) ;
  assign n1875 = n1874 ^ x230 ^ 1'b0 ;
  assign n1876 = n1875 ^ n1370 ^ n972 ;
  assign n1877 = n1797 ^ n1646 ^ n1627 ;
  assign n1878 = ( ~n872 & n1103 ) | ( ~n872 & n1517 ) | ( n1103 & n1517 ) ;
  assign n1879 = n1878 ^ n1427 ^ n760 ;
  assign n1880 = ( ~x224 & n1023 ) | ( ~x224 & n1879 ) | ( n1023 & n1879 ) ;
  assign n1881 = n854 & ~n1099 ;
  assign n1882 = ~n543 & n755 ;
  assign n1883 = n557 | n650 ;
  assign n1884 = n581 & ~n1883 ;
  assign n1885 = n1882 | n1884 ;
  assign n1886 = n1885 ^ n1786 ^ n1678 ;
  assign n1893 = n631 | n1650 ;
  assign n1894 = n1893 ^ n453 ^ 1'b0 ;
  assign n1888 = n590 ^ n518 ^ 1'b0 ;
  assign n1889 = x223 & n1888 ;
  assign n1887 = n307 | n1474 ;
  assign n1890 = n1889 ^ n1887 ^ n635 ;
  assign n1891 = n1190 & ~n1890 ;
  assign n1892 = n1891 ^ n1648 ^ 1'b0 ;
  assign n1895 = n1894 ^ n1892 ^ 1'b0 ;
  assign n1896 = x140 & ~n569 ;
  assign n1897 = n1896 ^ n737 ^ 1'b0 ;
  assign n1898 = n832 ^ x143 ^ 1'b0 ;
  assign n1899 = ~n863 & n1898 ;
  assign n1900 = n527 | n1899 ;
  assign n1901 = x84 & ~n1900 ;
  assign n1902 = n1897 & n1901 ;
  assign n1903 = n832 ^ x106 ^ 1'b0 ;
  assign n1904 = n1903 ^ x192 ^ 1'b0 ;
  assign n1905 = n1626 & ~n1726 ;
  assign n1906 = n301 & n1905 ;
  assign n1907 = ( ~n429 & n1498 ) | ( ~n429 & n1906 ) | ( n1498 & n1906 ) ;
  assign n1908 = n1376 & ~n1495 ;
  assign n1909 = ~n1689 & n1908 ;
  assign n1912 = n1102 ^ n412 ^ x132 ;
  assign n1910 = ( ~n485 & n509 ) | ( ~n485 & n1793 ) | ( n509 & n1793 ) ;
  assign n1911 = n1910 ^ n1856 ^ n489 ;
  assign n1913 = n1912 ^ n1911 ^ 1'b0 ;
  assign n1914 = x16 & ~n1195 ;
  assign n1915 = x34 & n773 ;
  assign n1916 = ~x127 & n1915 ;
  assign n1917 = ( ~n471 & n1677 ) | ( ~n471 & n1916 ) | ( n1677 & n1916 ) ;
  assign n1918 = n1917 ^ n434 ^ 1'b0 ;
  assign n1919 = n513 & n1918 ;
  assign n1920 = ~n1200 & n1919 ;
  assign n1921 = n936 ^ x191 ^ 1'b0 ;
  assign n1922 = ~n458 & n1921 ;
  assign n1923 = n1922 ^ n261 ^ 1'b0 ;
  assign n1924 = n770 | n1923 ;
  assign n1925 = n518 ^ x151 ^ 1'b0 ;
  assign n1926 = ( ~n1608 & n1924 ) | ( ~n1608 & n1925 ) | ( n1924 & n1925 ) ;
  assign n1927 = n411 ^ x38 ^ 1'b0 ;
  assign n1928 = x14 & n1927 ;
  assign n1930 = n1601 ^ n445 ^ n328 ;
  assign n1929 = n742 & n1464 ;
  assign n1931 = n1930 ^ n1929 ^ 1'b0 ;
  assign n1932 = n410 & ~n1931 ;
  assign n1933 = n1928 & n1932 ;
  assign n1934 = ~n744 & n1933 ;
  assign n1935 = n1934 ^ n1247 ^ 1'b0 ;
  assign n1936 = ~n1253 & n1525 ;
  assign n1937 = n1936 ^ n1344 ^ 1'b0 ;
  assign n1938 = n1937 ^ n1200 ^ 1'b0 ;
  assign n1940 = n1686 ^ n1297 ^ n997 ;
  assign n1939 = x132 & n1440 ;
  assign n1941 = n1940 ^ n1939 ^ 1'b0 ;
  assign n1942 = x205 & ~n1941 ;
  assign n1943 = n669 & n1942 ;
  assign n1944 = n1943 ^ x193 ^ 1'b0 ;
  assign n1945 = x36 & x84 ;
  assign n1946 = ~x42 & n1945 ;
  assign n1947 = ~n982 & n1946 ;
  assign n1948 = n1665 & ~n1947 ;
  assign n1949 = n1944 & n1948 ;
  assign n1950 = n1949 ^ n1667 ^ 1'b0 ;
  assign n1951 = n1938 | n1950 ;
  assign n1952 = n1951 ^ n1453 ^ 1'b0 ;
  assign n1953 = n1681 ^ n1213 ^ 1'b0 ;
  assign n1954 = n950 ^ n895 ^ 1'b0 ;
  assign n1955 = x109 & ~n1954 ;
  assign n1958 = n1769 ^ n1705 ^ 1'b0 ;
  assign n1957 = n1641 ^ n813 ^ x60 ;
  assign n1959 = n1958 ^ n1957 ^ x68 ;
  assign n1956 = x161 & ~n1413 ;
  assign n1960 = n1959 ^ n1956 ^ 1'b0 ;
  assign n1961 = x5 | n498 ;
  assign n1962 = ~n335 & n1961 ;
  assign n1963 = n1962 ^ n928 ^ 1'b0 ;
  assign n1964 = n1308 ^ n263 ^ 1'b0 ;
  assign n1965 = ~n379 & n1964 ;
  assign n1966 = n1965 ^ n802 ^ 1'b0 ;
  assign n1967 = n1698 | n1966 ;
  assign n1968 = x174 & n340 ;
  assign n1969 = n1968 ^ n1056 ^ 1'b0 ;
  assign n1970 = n1279 & ~n1969 ;
  assign n1976 = n1023 ^ n587 ^ n374 ;
  assign n1977 = n1976 ^ n1125 ^ 1'b0 ;
  assign n1978 = x19 & n1977 ;
  assign n1971 = n577 & ~n592 ;
  assign n1972 = n723 & n1971 ;
  assign n1973 = n1117 & ~n1972 ;
  assign n1974 = ~n1369 & n1973 ;
  assign n1975 = n1974 ^ n1802 ^ 1'b0 ;
  assign n1979 = n1978 ^ n1975 ^ 1'b0 ;
  assign n1980 = n675 ^ n436 ^ 1'b0 ;
  assign n1981 = n1006 & n1870 ;
  assign n1982 = ~n1739 & n1981 ;
  assign n1983 = n936 | n1429 ;
  assign n1984 = n1750 ^ n1653 ^ x47 ;
  assign n1985 = ( x98 & n399 ) | ( x98 & ~n1984 ) | ( n399 & ~n1984 ) ;
  assign n1986 = x85 & n610 ;
  assign n1987 = n1986 ^ n409 ^ 1'b0 ;
  assign n1988 = n647 | n1987 ;
  assign n1989 = x211 & ~n1988 ;
  assign n1990 = n342 & n1209 ;
  assign n1991 = n1990 ^ x101 ^ 1'b0 ;
  assign n1992 = n1147 | n1991 ;
  assign n1993 = ~n1989 & n1992 ;
  assign n1994 = n1993 ^ n559 ^ 1'b0 ;
  assign n1995 = n1486 & ~n1994 ;
  assign n1996 = x99 & n1156 ;
  assign n1997 = x198 | n704 ;
  assign n1998 = ~n1996 & n1997 ;
  assign n1999 = n760 & n1998 ;
  assign n2000 = ~n432 & n1373 ;
  assign n2001 = n626 | n1444 ;
  assign n2002 = n2000 & ~n2001 ;
  assign n2003 = n989 | n1120 ;
  assign n2004 = n2003 ^ x247 ^ 1'b0 ;
  assign n2005 = n884 | n1384 ;
  assign n2006 = n1506 ^ n445 ^ 1'b0 ;
  assign n2007 = n472 & ~n1703 ;
  assign n2008 = ~n2006 & n2007 ;
  assign n2009 = n904 ^ n661 ^ n478 ;
  assign n2010 = ( ~n1555 & n1762 ) | ( ~n1555 & n2009 ) | ( n1762 & n2009 ) ;
  assign n2011 = n277 ^ x175 ^ 1'b0 ;
  assign n2012 = ( n530 & ~n762 ) | ( n530 & n1418 ) | ( ~n762 & n1418 ) ;
  assign n2013 = n2012 ^ n880 ^ 1'b0 ;
  assign n2014 = n1581 & ~n2013 ;
  assign n2015 = n1795 ^ n840 ^ x132 ;
  assign n2016 = n640 ^ n527 ^ 1'b0 ;
  assign n2017 = n1550 & ~n2016 ;
  assign n2018 = ~n1381 & n1498 ;
  assign n2019 = n2018 ^ n1273 ^ 1'b0 ;
  assign n2020 = n1440 ^ n1209 ^ n612 ;
  assign n2021 = ~n1711 & n2020 ;
  assign n2022 = n2021 ^ n930 ^ 1'b0 ;
  assign n2023 = ( n1577 & ~n1674 ) | ( n1577 & n1681 ) | ( ~n1674 & n1681 ) ;
  assign n2024 = n963 & ~n1212 ;
  assign n2025 = ~n1902 & n2024 ;
  assign n2026 = ~x87 & n2025 ;
  assign n2027 = n1373 | n2026 ;
  assign n2028 = n2023 | n2027 ;
  assign n2029 = ( x139 & ~x225 ) | ( x139 & n462 ) | ( ~x225 & n462 ) ;
  assign n2030 = n1811 ^ n1096 ^ 1'b0 ;
  assign n2031 = n2029 & ~n2030 ;
  assign n2032 = n486 ^ x185 ^ 1'b0 ;
  assign n2033 = x47 & n2032 ;
  assign n2034 = n2033 ^ n1291 ^ n520 ;
  assign n2035 = n1817 & n2034 ;
  assign n2036 = n2035 ^ x68 ^ 1'b0 ;
  assign n2037 = x16 & ~n498 ;
  assign n2038 = ~n742 & n2037 ;
  assign n2039 = n1377 ^ n305 ^ 1'b0 ;
  assign n2040 = n1162 | n2039 ;
  assign n2041 = x108 & ~n1650 ;
  assign n2042 = n333 | n727 ;
  assign n2043 = n444 | n2042 ;
  assign n2044 = n2041 | n2043 ;
  assign n2045 = n1026 | n1106 ;
  assign n2046 = n2044 | n2045 ;
  assign n2047 = ~n1782 & n2046 ;
  assign n2048 = ( n895 & ~n2040 ) | ( n895 & n2047 ) | ( ~n2040 & n2047 ) ;
  assign n2049 = n1996 ^ n713 ^ 1'b0 ;
  assign n2050 = ~n640 & n2049 ;
  assign n2051 = ~n1281 & n2050 ;
  assign n2052 = n1475 ^ n1332 ^ n1101 ;
  assign n2053 = n2052 ^ x246 ^ 1'b0 ;
  assign n2054 = ( x218 & ~n409 ) | ( x218 & n776 ) | ( ~n409 & n776 ) ;
  assign n2055 = n2054 ^ n1259 ^ n1113 ;
  assign n2056 = n1506 & ~n1934 ;
  assign n2057 = n2056 ^ n1258 ^ 1'b0 ;
  assign n2062 = n1250 ^ n332 ^ 1'b0 ;
  assign n2063 = x2 & n2062 ;
  assign n2058 = ~x29 & x185 ;
  assign n2059 = ( x240 & ~n471 ) | ( x240 & n2058 ) | ( ~n471 & n2058 ) ;
  assign n2060 = n760 & n2059 ;
  assign n2061 = ~n1930 & n2060 ;
  assign n2064 = n2063 ^ n2061 ^ 1'b0 ;
  assign n2065 = n2046 ^ n256 ^ x239 ;
  assign n2066 = n472 ^ x222 ^ 1'b0 ;
  assign n2067 = n2066 ^ n1386 ^ n380 ;
  assign n2068 = n1600 ^ n1004 ^ 1'b0 ;
  assign n2069 = n831 & ~n928 ;
  assign n2070 = ~x88 & n2069 ;
  assign n2071 = n646 & ~n1013 ;
  assign n2072 = n360 & n2071 ;
  assign n2073 = ~x206 & n2072 ;
  assign n2074 = n1281 & n2073 ;
  assign n2075 = n1925 ^ x80 ^ 1'b0 ;
  assign n2076 = n436 & n456 ;
  assign n2077 = n1395 ^ n1101 ^ x228 ;
  assign n2078 = n1048 ^ x164 ^ 1'b0 ;
  assign n2079 = n2078 ^ n1231 ^ 1'b0 ;
  assign n2080 = n1324 & n2079 ;
  assign n2081 = ( n1348 & n2077 ) | ( n1348 & n2080 ) | ( n2077 & n2080 ) ;
  assign n2082 = n582 & n2081 ;
  assign n2083 = n516 | n617 ;
  assign n2084 = n2083 ^ n486 ^ 1'b0 ;
  assign n2085 = x97 & n956 ;
  assign n2086 = ~n2084 & n2085 ;
  assign n2087 = ~n484 & n2086 ;
  assign n2088 = x239 & ~n752 ;
  assign n2089 = n2088 ^ x210 ^ 1'b0 ;
  assign n2090 = n1007 ^ n873 ^ 1'b0 ;
  assign n2091 = n921 & n2090 ;
  assign n2092 = ~n647 & n1010 ;
  assign n2093 = n1302 & n2092 ;
  assign n2094 = x30 & ~n2093 ;
  assign n2095 = n1250 & n2094 ;
  assign n2096 = x102 & ~n652 ;
  assign n2097 = ( n1488 & n1569 ) | ( n1488 & n2096 ) | ( n1569 & n2096 ) ;
  assign n2098 = n1527 ^ n1423 ^ 1'b0 ;
  assign n2099 = n624 & n1681 ;
  assign n2100 = n1066 ^ n841 ^ n476 ;
  assign n2101 = x249 & ~n2009 ;
  assign n2102 = n2101 ^ x227 ^ 1'b0 ;
  assign n2103 = n2100 & n2102 ;
  assign n2104 = n1186 ^ n574 ^ 1'b0 ;
  assign n2105 = n2103 | n2104 ;
  assign n2106 = n2105 ^ n747 ^ 1'b0 ;
  assign n2107 = n490 ^ n484 ^ 1'b0 ;
  assign n2108 = n1034 | n2107 ;
  assign n2109 = ~n1641 & n2108 ;
  assign n2117 = n852 ^ x36 ^ 1'b0 ;
  assign n2118 = n491 & ~n2117 ;
  assign n2119 = ~n856 & n2118 ;
  assign n2120 = n2119 ^ x223 ^ 1'b0 ;
  assign n2112 = x20 & x41 ;
  assign n2113 = n2112 ^ n558 ^ 1'b0 ;
  assign n2110 = n1512 ^ n968 ^ 1'b0 ;
  assign n2111 = n1376 & ~n2110 ;
  assign n2114 = n2113 ^ n2111 ^ n1763 ;
  assign n2115 = n1233 ^ n591 ^ 1'b0 ;
  assign n2116 = n2114 | n2115 ;
  assign n2121 = n2120 ^ n2116 ^ 1'b0 ;
  assign n2122 = ~n393 & n2121 ;
  assign n2123 = n1046 & n1498 ;
  assign n2124 = ~n896 & n2123 ;
  assign n2125 = n1266 & n2124 ;
  assign n2126 = x0 & ~n1176 ;
  assign n2127 = n2126 ^ n1095 ^ 1'b0 ;
  assign n2128 = n647 ^ x243 ^ 1'b0 ;
  assign n2129 = n2127 | n2128 ;
  assign n2131 = x163 & ~n1300 ;
  assign n2130 = ~n587 & n821 ;
  assign n2132 = n2131 ^ n2130 ^ 1'b0 ;
  assign n2133 = n1411 & ~n2132 ;
  assign n2134 = n1453 & n2133 ;
  assign n2135 = ( x57 & n376 ) | ( x57 & n679 ) | ( n376 & n679 ) ;
  assign n2136 = ~n458 & n1110 ;
  assign n2137 = n2136 ^ n1115 ^ 1'b0 ;
  assign n2138 = n2137 ^ n652 ^ 1'b0 ;
  assign n2139 = n1013 & n1228 ;
  assign n2140 = n2139 ^ n371 ^ 1'b0 ;
  assign n2141 = ~n826 & n1298 ;
  assign n2143 = n947 & ~n1068 ;
  assign n2144 = n753 & n2143 ;
  assign n2142 = x190 & n512 ;
  assign n2145 = n2144 ^ n2142 ^ 1'b0 ;
  assign n2146 = n1370 | n2145 ;
  assign n2147 = ( x229 & n793 ) | ( x229 & ~n1993 ) | ( n793 & ~n1993 ) ;
  assign n2148 = n2146 & n2147 ;
  assign n2149 = n1575 ^ n1540 ^ 1'b0 ;
  assign n2150 = n1557 & n1626 ;
  assign n2151 = n2150 ^ n865 ^ 1'b0 ;
  assign n2152 = n1263 ^ x110 ^ 1'b0 ;
  assign n2153 = n918 & ~n2152 ;
  assign n2154 = n288 | n872 ;
  assign n2155 = n877 & ~n2154 ;
  assign n2156 = ~n863 & n1295 ;
  assign n2157 = n1527 & ~n2156 ;
  assign n2158 = n2155 & n2157 ;
  assign n2159 = n1222 & n1406 ;
  assign n2160 = n283 & n2159 ;
  assign n2161 = n2160 ^ n294 ^ x107 ;
  assign n2162 = ( n1403 & n1630 ) | ( n1403 & n1906 ) | ( n1630 & n1906 ) ;
  assign n2163 = ~n1648 & n1953 ;
  assign n2164 = n2163 ^ n721 ^ 1'b0 ;
  assign n2165 = ~n944 & n1671 ;
  assign n2166 = n1866 ^ n572 ^ 1'b0 ;
  assign n2167 = x210 & n1166 ;
  assign n2168 = n2167 ^ n936 ^ 1'b0 ;
  assign n2169 = n2168 ^ n400 ^ 1'b0 ;
  assign n2170 = ~n363 & n2169 ;
  assign n2171 = n2170 ^ x231 ^ 1'b0 ;
  assign n2172 = x119 & n1419 ;
  assign n2173 = n2172 ^ n432 ^ 1'b0 ;
  assign n2174 = n736 ^ n686 ^ 1'b0 ;
  assign n2175 = n821 & n1459 ;
  assign n2176 = n2174 & n2175 ;
  assign n2177 = n1004 | n2176 ;
  assign n2178 = n2177 ^ n1688 ^ 1'b0 ;
  assign n2179 = n441 | n753 ;
  assign n2180 = n2179 ^ n1631 ^ x239 ;
  assign n2181 = n1615 ^ n719 ^ n645 ;
  assign n2182 = ( x234 & n2180 ) | ( x234 & ~n2181 ) | ( n2180 & ~n2181 ) ;
  assign n2186 = ( x23 & ~n636 ) | ( x23 & n995 ) | ( ~n636 & n995 ) ;
  assign n2183 = ~x122 & x142 ;
  assign n2184 = n634 | n756 ;
  assign n2185 = ~n2183 & n2184 ;
  assign n2187 = n2186 ^ n2185 ^ 1'b0 ;
  assign n2188 = n319 & ~n2187 ;
  assign n2189 = ~n550 & n1476 ;
  assign n2190 = ~x45 & n2189 ;
  assign n2191 = ( x100 & n735 ) | ( x100 & n1872 ) | ( n735 & n1872 ) ;
  assign n2192 = n2191 ^ n1285 ^ 1'b0 ;
  assign n2193 = n1544 & ~n2192 ;
  assign n2194 = n2190 & n2193 ;
  assign n2195 = n1222 | n2194 ;
  assign n2196 = n555 & ~n1474 ;
  assign n2197 = ~n474 & n2196 ;
  assign n2198 = n390 | n2197 ;
  assign n2199 = n2198 ^ n1829 ^ 1'b0 ;
  assign n2200 = x245 ^ x152 ^ 1'b0 ;
  assign n2201 = x33 & n2200 ;
  assign n2202 = ~n511 & n1225 ;
  assign n2203 = ( n1253 & n2201 ) | ( n1253 & n2202 ) | ( n2201 & n2202 ) ;
  assign n2204 = ( x52 & ~n395 ) | ( x52 & n1258 ) | ( ~n395 & n1258 ) ;
  assign n2205 = n2204 ^ n829 ^ 1'b0 ;
  assign n2206 = n1053 & ~n2205 ;
  assign n2207 = n2206 ^ n829 ^ n659 ;
  assign n2208 = ( ~n500 & n1603 ) | ( ~n500 & n2207 ) | ( n1603 & n2207 ) ;
  assign n2209 = n1170 & n2208 ;
  assign n2210 = n397 & ~n444 ;
  assign n2211 = n749 & n2210 ;
  assign n2212 = n2211 ^ n1009 ^ 1'b0 ;
  assign n2213 = ( n1593 & n1926 ) | ( n1593 & n2212 ) | ( n1926 & n2212 ) ;
  assign n2214 = n2209 | n2213 ;
  assign n2215 = n314 & ~n915 ;
  assign n2216 = n2215 ^ n640 ^ 1'b0 ;
  assign n2217 = n1132 & n2216 ;
  assign n2218 = ~n1069 & n1215 ;
  assign n2219 = n1558 ^ n367 ^ 1'b0 ;
  assign n2220 = n873 | n2219 ;
  assign n2221 = n2218 | n2220 ;
  assign n2222 = n574 ^ n559 ^ 1'b0 ;
  assign n2223 = x94 & n2222 ;
  assign n2224 = ( n1236 & n2101 ) | ( n1236 & ~n2223 ) | ( n2101 & ~n2223 ) ;
  assign n2225 = n1027 | n1241 ;
  assign n2227 = x179 | n647 ;
  assign n2226 = ( x18 & ~x169 ) | ( x18 & x240 ) | ( ~x169 & x240 ) ;
  assign n2228 = n2227 ^ n2226 ^ n536 ;
  assign n2229 = n1540 ^ n579 ^ 1'b0 ;
  assign n2230 = n2228 & ~n2229 ;
  assign n2231 = n2209 & n2230 ;
  assign n2232 = x30 & ~n1824 ;
  assign n2233 = ~n1515 & n2057 ;
  assign n2234 = n1347 & n2233 ;
  assign n2235 = ( x63 & ~n627 ) | ( x63 & n994 ) | ( ~n627 & n994 ) ;
  assign n2236 = n1069 | n1429 ;
  assign n2237 = x40 | n2236 ;
  assign n2238 = n2235 & n2237 ;
  assign n2239 = n2234 & n2238 ;
  assign n2240 = n626 & ~n1897 ;
  assign n2241 = ( x35 & n332 ) | ( x35 & n2240 ) | ( n332 & n2240 ) ;
  assign n2242 = n1213 ^ n1156 ^ 1'b0 ;
  assign n2243 = n2241 & ~n2242 ;
  assign n2244 = n2142 ^ n552 ^ x111 ;
  assign n2245 = ~n747 & n1801 ;
  assign n2246 = n828 & n2245 ;
  assign n2247 = n1023 ^ n956 ^ 1'b0 ;
  assign n2249 = ( x18 & ~n993 ) | ( x18 & n1278 ) | ( ~n993 & n1278 ) ;
  assign n2248 = x149 & ~n768 ;
  assign n2250 = n2249 ^ n2248 ^ n1823 ;
  assign n2251 = x244 | n1261 ;
  assign n2252 = x119 | n2251 ;
  assign n2253 = n1343 ^ n690 ^ x198 ;
  assign n2254 = n1210 ^ n592 ^ 1'b0 ;
  assign n2255 = ~n2253 & n2254 ;
  assign n2256 = n1042 & n2255 ;
  assign n2257 = n2256 ^ n1038 ^ 1'b0 ;
  assign n2259 = n853 ^ n335 ^ 1'b0 ;
  assign n2258 = ( n905 & n1430 ) | ( n905 & ~n1779 ) | ( n1430 & ~n1779 ) ;
  assign n2260 = n2259 ^ n2258 ^ 1'b0 ;
  assign n2261 = ( n1816 & ~n1965 ) | ( n1816 & n2260 ) | ( ~n1965 & n2260 ) ;
  assign n2262 = n2257 & ~n2261 ;
  assign n2263 = n1176 | n1351 ;
  assign n2264 = n2263 ^ n2059 ^ 1'b0 ;
  assign n2265 = n2264 ^ n1430 ^ 1'b0 ;
  assign n2266 = n2262 | n2265 ;
  assign n2267 = x250 & ~n473 ;
  assign n2268 = n716 ^ n341 ^ 1'b0 ;
  assign n2269 = n1961 & ~n2268 ;
  assign n2270 = x197 ^ x169 ^ 1'b0 ;
  assign n2271 = ~n322 & n2270 ;
  assign n2272 = ( n263 & ~n449 ) | ( n263 & n486 ) | ( ~n449 & n486 ) ;
  assign n2273 = n2271 & ~n2272 ;
  assign n2274 = ~n2269 & n2273 ;
  assign n2275 = n351 & ~n723 ;
  assign n2276 = n1252 ^ n926 ^ 1'b0 ;
  assign n2277 = n2276 ^ n2087 ^ 1'b0 ;
  assign n2278 = x54 & n1510 ;
  assign n2279 = n1453 ^ n1409 ^ 1'b0 ;
  assign n2280 = n2279 ^ n331 ^ 1'b0 ;
  assign n2281 = n1184 & n2280 ;
  assign n2282 = ~n1007 & n1833 ;
  assign n2283 = n2282 ^ n693 ^ 1'b0 ;
  assign n2284 = n1358 | n2283 ;
  assign n2285 = n2281 & ~n2284 ;
  assign n2286 = n2140 ^ n1228 ^ n506 ;
  assign n2292 = x218 | n1084 ;
  assign n2287 = n1712 ^ n1683 ^ n1582 ;
  assign n2288 = ~n434 & n677 ;
  assign n2289 = ~n1107 & n2288 ;
  assign n2290 = n1590 | n2289 ;
  assign n2291 = n2287 | n2290 ;
  assign n2293 = n2292 ^ n2291 ^ 1'b0 ;
  assign n2294 = n633 & ~n1974 ;
  assign n2295 = x73 & n1782 ;
  assign n2296 = n2295 ^ n2059 ^ 1'b0 ;
  assign n2297 = n1288 ^ n1081 ^ 1'b0 ;
  assign n2298 = ~n2296 & n2297 ;
  assign n2299 = n1455 | n2298 ;
  assign n2300 = ~n1390 & n2299 ;
  assign n2301 = n267 | n2134 ;
  assign n2302 = n2301 ^ x33 ^ 1'b0 ;
  assign n2303 = n1374 ^ n1215 ^ 1'b0 ;
  assign n2304 = n776 | n2303 ;
  assign n2305 = n1992 | n2304 ;
  assign n2306 = n269 & ~n2305 ;
  assign n2307 = n459 & ~n1661 ;
  assign n2308 = n783 & n1887 ;
  assign n2309 = n2308 ^ n2103 ^ 1'b0 ;
  assign n2310 = n1579 ^ n393 ^ 1'b0 ;
  assign n2311 = n1700 & n2310 ;
  assign n2312 = n1145 ^ n329 ^ 1'b0 ;
  assign n2313 = x58 | n2312 ;
  assign n2314 = n983 ^ n840 ^ 1'b0 ;
  assign n2315 = n1998 ^ x110 ^ 1'b0 ;
  assign n2316 = n2315 ^ n594 ^ 1'b0 ;
  assign n2317 = ~n861 & n2316 ;
  assign n2318 = n1179 ^ n742 ^ 1'b0 ;
  assign n2322 = ( ~x207 & n890 ) | ( ~x207 & n919 ) | ( n890 & n919 ) ;
  assign n2323 = n286 | n2322 ;
  assign n2324 = n2323 ^ x35 ^ 1'b0 ;
  assign n2319 = n279 ^ x10 ^ 1'b0 ;
  assign n2320 = n1949 | n2319 ;
  assign n2321 = n1364 | n2320 ;
  assign n2325 = n2324 ^ n2321 ^ 1'b0 ;
  assign n2326 = n836 & n2325 ;
  assign n2331 = x59 & x123 ;
  assign n2332 = ~x4 & n2331 ;
  assign n2333 = n2332 ^ n942 ^ 1'b0 ;
  assign n2334 = n345 ^ x173 ^ 1'b0 ;
  assign n2335 = n2333 & n2334 ;
  assign n2336 = ~n1164 & n2335 ;
  assign n2337 = n2336 ^ n2259 ^ 1'b0 ;
  assign n2327 = n950 ^ x27 ^ 1'b0 ;
  assign n2328 = x113 & n2327 ;
  assign n2329 = ~x12 & n2328 ;
  assign n2330 = n790 & ~n2329 ;
  assign n2338 = n2337 ^ n2330 ^ 1'b0 ;
  assign n2339 = x211 | n1056 ;
  assign n2340 = n2339 ^ x227 ^ 1'b0 ;
  assign n2341 = ( x103 & n915 ) | ( x103 & ~n2340 ) | ( n915 & ~n2340 ) ;
  assign n2342 = n1319 & ~n2341 ;
  assign n2343 = n605 ^ x108 ^ 1'b0 ;
  assign n2344 = n1932 & ~n2343 ;
  assign n2345 = n1314 | n2344 ;
  assign n2346 = n444 ^ x61 ^ 1'b0 ;
  assign n2347 = n605 | n2346 ;
  assign n2348 = x131 & ~n2347 ;
  assign n2349 = n2348 ^ n753 ^ 1'b0 ;
  assign n2350 = n1192 ^ n518 ^ 1'b0 ;
  assign n2351 = n2350 ^ n1378 ^ n418 ;
  assign n2352 = n2351 ^ n1213 ^ n1075 ;
  assign n2353 = n2352 ^ n635 ^ 1'b0 ;
  assign n2354 = ~x14 & n526 ;
  assign n2355 = n1162 ^ n593 ^ 1'b0 ;
  assign n2356 = n1254 | n1277 ;
  assign n2357 = n1315 | n2356 ;
  assign n2358 = n1764 ^ n1259 ^ 1'b0 ;
  assign n2359 = n753 ^ n315 ^ 1'b0 ;
  assign n2360 = ( n267 & n277 ) | ( n267 & ~n1448 ) | ( n277 & ~n1448 ) ;
  assign n2361 = n1209 ^ n269 ^ 1'b0 ;
  assign n2362 = n1273 & n2361 ;
  assign n2363 = ( n473 & ~n1697 ) | ( n473 & n2362 ) | ( ~n1697 & n2362 ) ;
  assign n2364 = n1009 & n2363 ;
  assign n2365 = n1378 & n2364 ;
  assign n2367 = n797 ^ n617 ^ 1'b0 ;
  assign n2368 = ~n967 & n2367 ;
  assign n2366 = n495 ^ n433 ^ 1'b0 ;
  assign n2369 = n2368 ^ n2366 ^ n1170 ;
  assign n2370 = n1988 ^ n1722 ^ 1'b0 ;
  assign n2371 = n1483 & n2370 ;
  assign n2372 = ~n438 & n747 ;
  assign n2373 = ~n861 & n2372 ;
  assign n2374 = n2373 ^ x251 ^ 1'b0 ;
  assign n2378 = ( n380 & n978 ) | ( n380 & ~n2179 ) | ( n978 & ~n2179 ) ;
  assign n2379 = x197 & n587 ;
  assign n2380 = n2379 ^ x226 ^ 1'b0 ;
  assign n2381 = n631 | n2380 ;
  assign n2382 = n1681 & ~n2381 ;
  assign n2383 = n1444 | n2382 ;
  assign n2384 = n2378 & ~n2383 ;
  assign n2375 = ~n1026 & n1256 ;
  assign n2376 = n2375 ^ n1360 ^ 1'b0 ;
  assign n2377 = n2376 ^ n1068 ^ 1'b0 ;
  assign n2385 = n2384 ^ n2377 ^ 1'b0 ;
  assign n2386 = n315 | n2385 ;
  assign n2387 = n1206 & n1685 ;
  assign n2388 = x249 & ~n2387 ;
  assign n2389 = n2388 ^ n853 ^ 1'b0 ;
  assign n2390 = n1194 ^ x225 ^ 1'b0 ;
  assign n2391 = x127 & ~n798 ;
  assign n2392 = ~n1273 & n2391 ;
  assign n2393 = n1017 & n2392 ;
  assign n2394 = n2393 ^ x71 ^ 1'b0 ;
  assign n2395 = n737 & n1313 ;
  assign n2396 = n2044 ^ x150 ^ 1'b0 ;
  assign n2397 = x78 & n2396 ;
  assign n2398 = n1692 ^ n919 ^ 1'b0 ;
  assign n2399 = x214 & ~n2398 ;
  assign n2400 = n2399 ^ n822 ^ 1'b0 ;
  assign n2401 = n1604 | n2400 ;
  assign n2402 = ( x187 & n1354 ) | ( x187 & n2347 ) | ( n1354 & n2347 ) ;
  assign n2403 = n831 & ~n2402 ;
  assign n2404 = ~n1220 & n2403 ;
  assign n2405 = n2404 ^ n582 ^ 1'b0 ;
  assign n2406 = n2405 ^ n2346 ^ n981 ;
  assign n2407 = ( n400 & n596 ) | ( n400 & ~n911 ) | ( n596 & ~n911 ) ;
  assign n2408 = x236 & ~n1613 ;
  assign n2409 = n1033 & n2408 ;
  assign n2410 = ~n849 & n2341 ;
  assign n2411 = n2410 ^ n1457 ^ 1'b0 ;
  assign n2412 = n1597 ^ n559 ^ 1'b0 ;
  assign n2413 = n2412 ^ n1920 ^ 1'b0 ;
  assign n2414 = n1985 ^ n1480 ^ 1'b0 ;
  assign n2415 = n2000 ^ n617 ^ 1'b0 ;
  assign n2416 = n1027 & n2415 ;
  assign n2417 = ~n729 & n1013 ;
  assign n2418 = ~n558 & n2417 ;
  assign n2419 = n476 & ~n648 ;
  assign n2420 = ( n974 & n2418 ) | ( n974 & ~n2419 ) | ( n2418 & ~n2419 ) ;
  assign n2421 = n2420 ^ n1213 ^ x83 ;
  assign n2422 = n1192 & n2054 ;
  assign n2423 = n1711 ^ n513 ^ 1'b0 ;
  assign n2424 = n2423 ^ n2057 ^ 1'b0 ;
  assign n2425 = n2342 | n2424 ;
  assign n2426 = n1541 ^ n1285 ^ x136 ;
  assign n2427 = n1736 ^ x56 ^ 1'b0 ;
  assign n2428 = ~n550 & n2427 ;
  assign n2429 = ~x7 & n2428 ;
  assign n2430 = n2426 & n2429 ;
  assign n2431 = n1528 ^ n1285 ^ n371 ;
  assign n2432 = n2320 ^ n1995 ^ 1'b0 ;
  assign n2433 = n2431 | n2432 ;
  assign n2435 = x3 & n307 ;
  assign n2436 = n2435 ^ n308 ^ 1'b0 ;
  assign n2437 = ( n594 & n1289 ) | ( n594 & ~n2436 ) | ( n1289 & ~n2436 ) ;
  assign n2434 = n349 & n1096 ;
  assign n2438 = n2437 ^ n2434 ^ 1'b0 ;
  assign n2439 = x6 & ~n928 ;
  assign n2440 = n2439 ^ n939 ^ 1'b0 ;
  assign n2441 = ~n677 & n1835 ;
  assign n2442 = n2169 ^ n972 ^ 1'b0 ;
  assign n2443 = ~n942 & n1543 ;
  assign n2444 = n2443 ^ n1156 ^ 1'b0 ;
  assign n2447 = x215 | n1339 ;
  assign n2445 = ( n404 & n453 ) | ( n404 & n773 ) | ( n453 & n773 ) ;
  assign n2446 = n1284 & ~n2445 ;
  assign n2448 = n2447 ^ n2446 ^ 1'b0 ;
  assign n2449 = x117 & ~n2448 ;
  assign n2450 = n2067 ^ n1688 ^ 1'b0 ;
  assign n2451 = n444 | n2340 ;
  assign n2452 = n2451 ^ n1162 ^ 1'b0 ;
  assign n2453 = n714 ^ x180 ^ 1'b0 ;
  assign n2454 = n1829 | n2453 ;
  assign n2455 = ( ~x64 & n349 ) | ( ~x64 & n1024 ) | ( n349 & n1024 ) ;
  assign n2456 = n1009 & ~n2455 ;
  assign n2457 = n1007 & n2456 ;
  assign n2458 = n1824 ^ n1471 ^ 1'b0 ;
  assign n2459 = ~n2457 & n2458 ;
  assign n2460 = ( n650 & n1732 ) | ( n650 & ~n1881 ) | ( n1732 & ~n1881 ) ;
  assign n2461 = n1708 ^ n1311 ^ 1'b0 ;
  assign n2462 = n2460 | n2461 ;
  assign n2463 = n1275 ^ n1070 ^ 1'b0 ;
  assign n2464 = x219 & x232 ;
  assign n2465 = n2464 ^ n550 ^ 1'b0 ;
  assign n2466 = ( n1486 & n2034 ) | ( n1486 & ~n2465 ) | ( n2034 & ~n2465 ) ;
  assign n2467 = n2463 | n2466 ;
  assign n2468 = ( n420 & n541 ) | ( n420 & ~n2467 ) | ( n541 & ~n2467 ) ;
  assign n2469 = n1350 | n2111 ;
  assign n2470 = x184 & n1665 ;
  assign n2471 = n1695 ^ n1105 ^ n591 ;
  assign n2472 = ~n1514 & n1801 ;
  assign n2473 = n2471 & n2472 ;
  assign n2474 = ~n702 & n2048 ;
  assign n2475 = ~n866 & n2474 ;
  assign n2476 = x126 & ~x194 ;
  assign n2485 = n1222 & ~n1510 ;
  assign n2486 = n2485 ^ x37 ^ 1'b0 ;
  assign n2487 = n328 | n2486 ;
  assign n2488 = n2487 ^ x151 ^ 1'b0 ;
  assign n2478 = x198 ^ x97 ^ 1'b0 ;
  assign n2479 = x144 & n2478 ;
  assign n2480 = ( x53 & n331 ) | ( x53 & ~n2479 ) | ( n331 & ~n2479 ) ;
  assign n2481 = n2480 ^ n617 ^ n385 ;
  assign n2482 = n589 & ~n2481 ;
  assign n2483 = n2482 ^ n1237 ^ 1'b0 ;
  assign n2484 = ( n596 & n1055 ) | ( n596 & n2483 ) | ( n1055 & n2483 ) ;
  assign n2477 = n967 | n1337 ;
  assign n2489 = n2488 ^ n2484 ^ n2477 ;
  assign n2490 = n2187 ^ n1615 ^ 1'b0 ;
  assign n2491 = n694 | n1124 ;
  assign n2492 = n1477 & ~n2491 ;
  assign n2493 = n2492 ^ n1848 ^ 1'b0 ;
  assign n2494 = ~n1657 & n1981 ;
  assign n2495 = n331 & n2494 ;
  assign n2497 = n1633 ^ x46 ^ 1'b0 ;
  assign n2498 = n358 ^ x153 ^ 1'b0 ;
  assign n2499 = x20 & n2498 ;
  assign n2500 = ( x177 & ~n1182 ) | ( x177 & n2499 ) | ( ~n1182 & n2499 ) ;
  assign n2501 = ( n1755 & ~n2497 ) | ( n1755 & n2500 ) | ( ~n2497 & n2500 ) ;
  assign n2496 = n740 & ~n2061 ;
  assign n2502 = n2501 ^ n2496 ^ 1'b0 ;
  assign n2503 = ( n1327 & n2212 ) | ( n1327 & ~n2502 ) | ( n2212 & ~n2502 ) ;
  assign n2504 = n2503 ^ n2346 ^ 1'b0 ;
  assign n2505 = x86 & n909 ;
  assign n2506 = ~n918 & n2505 ;
  assign n2507 = ( n932 & n1321 ) | ( n932 & n2239 ) | ( n1321 & n2239 ) ;
  assign n2508 = n1164 & ~n1227 ;
  assign n2509 = n2508 ^ x127 ^ 1'b0 ;
  assign n2510 = n843 & n1975 ;
  assign n2511 = n2509 & n2510 ;
  assign n2517 = n892 ^ n367 ^ 1'b0 ;
  assign n2518 = n2517 ^ n2387 ^ n323 ;
  assign n2512 = n1946 ^ n358 ^ 1'b0 ;
  assign n2513 = n2512 ^ n441 ^ 1'b0 ;
  assign n2514 = n302 & ~n756 ;
  assign n2515 = n2513 & ~n2514 ;
  assign n2516 = ~x6 & n2515 ;
  assign n2519 = n2518 ^ n2516 ^ n1726 ;
  assign n2520 = n1162 ^ x85 ^ 1'b0 ;
  assign n2521 = n2519 & ~n2520 ;
  assign n2522 = n1475 ^ n669 ^ 1'b0 ;
  assign n2527 = ~n594 & n931 ;
  assign n2523 = n1270 ^ n1062 ^ 1'b0 ;
  assign n2524 = ( n596 & n989 ) | ( n596 & n1136 ) | ( n989 & n1136 ) ;
  assign n2525 = n2524 ^ n1285 ^ n593 ;
  assign n2526 = n2523 & n2525 ;
  assign n2528 = n2527 ^ n2526 ^ 1'b0 ;
  assign n2529 = ( n1772 & n2522 ) | ( n1772 & ~n2528 ) | ( n2522 & ~n2528 ) ;
  assign n2530 = ( n811 & n2190 ) | ( n811 & n2216 ) | ( n2190 & n2216 ) ;
  assign n2531 = ~n1829 & n2530 ;
  assign n2532 = n2171 & ~n2531 ;
  assign n2533 = n772 ^ n612 ^ 1'b0 ;
  assign n2534 = ~n692 & n2533 ;
  assign n2535 = x133 ^ x38 ^ 1'b0 ;
  assign n2536 = ~n963 & n2535 ;
  assign n2537 = x178 & n508 ;
  assign n2538 = n1140 | n2340 ;
  assign n2539 = n449 & ~n545 ;
  assign n2541 = n1885 & n2260 ;
  assign n2540 = n1892 & n2004 ;
  assign n2542 = n2541 ^ n2540 ^ 1'b0 ;
  assign n2543 = n516 ^ x147 ^ 1'b0 ;
  assign n2544 = ~n288 & n2543 ;
  assign n2545 = n1843 & ~n2544 ;
  assign n2546 = n2545 ^ n1233 ^ 1'b0 ;
  assign n2548 = n1129 & ~n1736 ;
  assign n2549 = ~n2418 & n2548 ;
  assign n2547 = n2492 ^ n1090 ^ x55 ;
  assign n2550 = n2549 ^ n2547 ^ n2272 ;
  assign n2551 = n1453 ^ x189 ^ 1'b0 ;
  assign n2552 = ~n954 & n2551 ;
  assign n2553 = n2480 & n2552 ;
  assign n2554 = n449 & ~n1003 ;
  assign n2555 = n1208 & n2554 ;
  assign n2556 = ( x199 & n1967 ) | ( x199 & ~n2555 ) | ( n1967 & ~n2555 ) ;
  assign n2557 = n333 ^ x92 ^ 1'b0 ;
  assign n2558 = n1443 & n1620 ;
  assign n2559 = n2557 & n2558 ;
  assign n2560 = n2559 ^ n1863 ^ 1'b0 ;
  assign n2561 = n2358 & n2560 ;
  assign n2562 = ~n317 & n489 ;
  assign n2563 = n2562 ^ n950 ^ 1'b0 ;
  assign n2564 = n2563 ^ n2306 ^ 1'b0 ;
  assign n2565 = n455 ^ x40 ^ 1'b0 ;
  assign n2566 = n2051 | n2565 ;
  assign n2567 = n1274 & ~n1712 ;
  assign n2568 = x178 | n631 ;
  assign n2569 = n1959 | n2568 ;
  assign n2570 = ~n787 & n2569 ;
  assign n2571 = n1705 & n2570 ;
  assign n2572 = n1496 ^ n571 ^ 1'b0 ;
  assign n2573 = ~n665 & n2572 ;
  assign n2574 = n1992 & n2063 ;
  assign n2575 = n2573 & ~n2574 ;
  assign n2576 = n1622 & n1767 ;
  assign n2577 = n2575 & n2576 ;
  assign n2583 = n2169 ^ x177 ^ 1'b0 ;
  assign n2584 = n1200 & n2583 ;
  assign n2578 = n553 & ~n884 ;
  assign n2579 = x27 & n753 ;
  assign n2580 = ~n2578 & n2579 ;
  assign n2581 = n2580 ^ n1115 ^ 1'b0 ;
  assign n2582 = n2581 ^ n668 ^ 1'b0 ;
  assign n2585 = n2584 ^ n2582 ^ x10 ;
  assign n2586 = n1268 ^ x60 ^ 1'b0 ;
  assign n2587 = ~x60 & n2586 ;
  assign n2588 = n2587 ^ n1223 ^ n530 ;
  assign n2589 = ~n1166 & n1643 ;
  assign n2590 = n2588 & n2589 ;
  assign n2594 = n500 & ~n770 ;
  assign n2595 = ~x73 & n2594 ;
  assign n2591 = n2248 & ~n2434 ;
  assign n2592 = n2591 ^ n1780 ^ 1'b0 ;
  assign n2593 = x137 & ~n2592 ;
  assign n2596 = n2595 ^ n2593 ^ 1'b0 ;
  assign n2597 = n2207 ^ x171 ^ 1'b0 ;
  assign n2598 = n2597 ^ n2005 ^ 1'b0 ;
  assign n2599 = n1762 ^ n556 ^ 1'b0 ;
  assign n2600 = n506 & n2599 ;
  assign n2601 = n2600 ^ n441 ^ 1'b0 ;
  assign n2602 = n2601 ^ n1651 ^ 1'b0 ;
  assign n2603 = n2598 & n2602 ;
  assign n2608 = ~n524 & n2503 ;
  assign n2605 = n2486 ^ n434 ^ 1'b0 ;
  assign n2606 = n2605 ^ n1493 ^ 1'b0 ;
  assign n2607 = n413 & ~n2606 ;
  assign n2609 = n2608 ^ n2607 ^ 1'b0 ;
  assign n2604 = n858 & ~n1253 ;
  assign n2610 = n2609 ^ n2604 ^ 1'b0 ;
  assign n2611 = n995 & n1536 ;
  assign n2612 = ( n409 & ~n1462 ) | ( n409 & n2611 ) | ( ~n1462 & n2611 ) ;
  assign n2613 = ( ~n1170 & n2592 ) | ( ~n1170 & n2612 ) | ( n2592 & n2612 ) ;
  assign n2614 = n1800 ^ n367 ^ 1'b0 ;
  assign n2615 = x81 | n1961 ;
  assign n2616 = n1762 ^ n1739 ^ 1'b0 ;
  assign n2617 = x232 & ~n2616 ;
  assign n2618 = n1997 ^ n1547 ^ 1'b0 ;
  assign n2619 = n983 ^ n861 ^ x63 ;
  assign n2620 = n2252 ^ n2243 ^ 1'b0 ;
  assign n2621 = ~n2619 & n2620 ;
  assign n2622 = n390 | n1430 ;
  assign n2623 = n2622 ^ n2431 ^ 1'b0 ;
  assign n2625 = x100 & n805 ;
  assign n2626 = n2625 ^ x176 ^ 1'b0 ;
  assign n2624 = n451 & n853 ;
  assign n2627 = n2626 ^ n2624 ^ 1'b0 ;
  assign n2628 = ~n2368 & n2627 ;
  assign n2629 = n645 | n2628 ;
  assign n2630 = n2629 ^ n1593 ^ 1'b0 ;
  assign n2631 = n2630 ^ n1096 ^ 1'b0 ;
  assign n2632 = n731 | n2631 ;
  assign n2633 = n2623 | n2632 ;
  assign n2634 = n1797 & ~n2633 ;
  assign n2635 = n2634 ^ n1038 ^ 1'b0 ;
  assign n2636 = ~n661 & n1213 ;
  assign n2637 = n2636 ^ n2201 ^ n505 ;
  assign n2638 = n1029 & ~n1597 ;
  assign n2639 = n2638 ^ n1336 ^ 1'b0 ;
  assign n2640 = n2481 | n2639 ;
  assign n2641 = n2640 ^ n1339 ^ n1024 ;
  assign n2642 = n2628 ^ n1277 ^ 1'b0 ;
  assign n2643 = n1776 & n2642 ;
  assign n2644 = n1683 & n2643 ;
  assign n2645 = n1791 & n2012 ;
  assign n2646 = n1060 & n1448 ;
  assign n2647 = n2646 ^ n2080 ^ 1'b0 ;
  assign n2648 = n2647 ^ n1862 ^ 1'b0 ;
  assign n2649 = n2264 ^ n498 ^ 1'b0 ;
  assign n2650 = ( n811 & n1563 ) | ( n811 & ~n2649 ) | ( n1563 & ~n2649 ) ;
  assign n2651 = n2314 ^ n1603 ^ 1'b0 ;
  assign n2652 = n2463 ^ n1851 ^ 1'b0 ;
  assign n2653 = ~x68 & n1235 ;
  assign n2654 = n1650 ^ n679 ^ 1'b0 ;
  assign n2655 = n2652 ^ n1831 ^ 1'b0 ;
  assign n2656 = n428 | n2655 ;
  assign n2657 = n1724 ^ n1615 ^ 1'b0 ;
  assign n2658 = n804 & n2657 ;
  assign n2659 = ~n562 & n1158 ;
  assign n2660 = n2659 ^ n657 ^ x217 ;
  assign n2661 = n1103 & ~n2660 ;
  assign n2662 = n686 & ~n2661 ;
  assign n2663 = n1086 & n2662 ;
  assign n2666 = n395 & ~n863 ;
  assign n2667 = n2666 ^ n513 ^ 1'b0 ;
  assign n2668 = ( n1237 & ~n1247 ) | ( n1237 & n2667 ) | ( ~n1247 & n2667 ) ;
  assign n2664 = n1315 ^ n1176 ^ 1'b0 ;
  assign n2665 = n2080 & ~n2664 ;
  assign n2669 = n2668 ^ n2665 ^ 1'b0 ;
  assign n2670 = n1870 & ~n2669 ;
  assign n2671 = n436 ^ n433 ^ 1'b0 ;
  assign n2672 = n1102 & ~n2671 ;
  assign n2673 = n271 & ~n2672 ;
  assign n2674 = n2673 ^ n2279 ^ 1'b0 ;
  assign n2675 = n2674 ^ n2507 ^ 1'b0 ;
  assign n2676 = n1476 ^ n413 ^ x15 ;
  assign n2677 = n2676 ^ x36 ^ 1'b0 ;
  assign n2678 = ~n1413 & n2677 ;
  assign n2679 = ~n1772 & n1987 ;
  assign n2680 = ~x46 & n2679 ;
  assign n2681 = n2680 ^ n761 ^ 1'b0 ;
  assign n2682 = n2681 ^ n1967 ^ 1'b0 ;
  assign n2683 = n1584 ^ x169 ^ 1'b0 ;
  assign n2684 = ~n2682 & n2683 ;
  assign n2685 = ( n397 & ~n2058 ) | ( n397 & n2287 ) | ( ~n2058 & n2287 ) ;
  assign n2686 = n2685 ^ n2298 ^ 1'b0 ;
  assign n2687 = n635 & ~n2686 ;
  assign n2688 = ( x69 & n2207 ) | ( x69 & ~n2687 ) | ( n2207 & ~n2687 ) ;
  assign n2689 = n1256 ^ x133 ^ 1'b0 ;
  assign n2690 = x39 & n1298 ;
  assign n2691 = n2689 & n2690 ;
  assign n2692 = n2691 ^ n1615 ^ 1'b0 ;
  assign n2693 = n1122 ^ n734 ^ 1'b0 ;
  assign n2694 = n1608 | n2693 ;
  assign n2695 = n1590 ^ n1194 ^ 1'b0 ;
  assign n2696 = n2694 | n2695 ;
  assign n2697 = n2573 ^ x241 ^ 1'b0 ;
  assign n2698 = n513 ^ x216 ^ x158 ;
  assign n2699 = n2698 ^ n516 ^ 1'b0 ;
  assign n2700 = n2699 ^ n1067 ^ 1'b0 ;
  assign n2701 = n2697 & ~n2700 ;
  assign n2702 = ~n835 & n2701 ;
  assign n2703 = ( ~n1526 & n2652 ) | ( ~n1526 & n2702 ) | ( n2652 & n2702 ) ;
  assign n2704 = ( ~n1328 & n1914 ) | ( ~n1328 & n2469 ) | ( n1914 & n2469 ) ;
  assign n2706 = x76 & x132 ;
  assign n2705 = n425 | n2231 ;
  assign n2707 = n2706 ^ n2705 ^ 1'b0 ;
  assign n2708 = n2362 ^ n1430 ^ n663 ;
  assign n2709 = n2708 ^ n1297 ^ 1'b0 ;
  assign n2710 = n2709 ^ n516 ^ n372 ;
  assign n2711 = n2710 ^ n1575 ^ x200 ;
  assign n2712 = n2711 ^ n1871 ^ 1'b0 ;
  assign n2713 = ~n1356 & n2540 ;
  assign n2714 = n361 ^ n340 ^ 1'b0 ;
  assign n2723 = n308 | n388 ;
  assign n2715 = n663 ^ x235 ^ 1'b0 ;
  assign n2717 = x125 & ~n1702 ;
  assign n2718 = n2717 ^ n976 ^ 1'b0 ;
  assign n2719 = n2718 ^ n502 ^ 1'b0 ;
  assign n2720 = n2719 ^ n2661 ^ n1876 ;
  assign n2716 = n1481 & n1963 ;
  assign n2721 = n2720 ^ n2716 ^ 1'b0 ;
  assign n2722 = n2715 & ~n2721 ;
  assign n2724 = n2723 ^ n2722 ^ 1'b0 ;
  assign n2725 = n994 & ~n2724 ;
  assign n2726 = n1177 | n1228 ;
  assign n2727 = n2726 ^ x254 ^ x56 ;
  assign n2737 = ( x76 & ~n1152 ) | ( x76 & n1254 ) | ( ~n1152 & n1254 ) ;
  assign n2734 = n418 | n712 ;
  assign n2735 = n2734 ^ n563 ^ 1'b0 ;
  assign n2733 = ~n462 & n1206 ;
  assign n2736 = n2735 ^ n2733 ^ 1'b0 ;
  assign n2728 = ~n1421 & n2339 ;
  assign n2729 = n795 | n1139 ;
  assign n2730 = n2728 & ~n2729 ;
  assign n2731 = n1544 & ~n2730 ;
  assign n2732 = n2667 & n2731 ;
  assign n2738 = n2737 ^ n2736 ^ n2732 ;
  assign n2739 = n1972 ^ x52 ^ 1'b0 ;
  assign n2740 = n441 & ~n2739 ;
  assign n2741 = n2740 ^ n476 ^ 1'b0 ;
  assign n2742 = n2741 ^ n1404 ^ 1'b0 ;
  assign n2743 = n485 & ~n2742 ;
  assign n2744 = n478 ^ x218 ^ 1'b0 ;
  assign n2745 = n2744 ^ n1101 ^ 1'b0 ;
  assign n2746 = n574 & ~n2745 ;
  assign n2747 = ~n1244 & n2746 ;
  assign n2748 = ~x203 & n2747 ;
  assign n2749 = n2748 ^ n273 ^ 1'b0 ;
  assign n2750 = n1535 & n2749 ;
  assign n2751 = ~n2600 & n2750 ;
  assign n2752 = n2751 ^ n2038 ^ n1095 ;
  assign n2753 = n1548 ^ n1295 ^ 1'b0 ;
  assign n2754 = n1017 & ~n2753 ;
  assign n2755 = x187 & ~n2754 ;
  assign n2756 = x31 & ~n1394 ;
  assign n2757 = n1889 ^ n937 ^ n562 ;
  assign n2758 = n1038 | n1319 ;
  assign n2759 = n2758 ^ x43 ^ 1'b0 ;
  assign n2760 = n2759 ^ n1390 ^ 1'b0 ;
  assign n2761 = n2134 | n2760 ;
  assign n2762 = n2054 ^ x159 ^ 1'b0 ;
  assign n2763 = ( x224 & ~n292 ) | ( x224 & n2253 ) | ( ~n292 & n2253 ) ;
  assign n2764 = x124 & n2522 ;
  assign n2765 = ~n2763 & n2764 ;
  assign n2766 = n2762 | n2765 ;
  assign n2772 = ~x149 & x249 ;
  assign n2771 = ~n322 & n2276 ;
  assign n2773 = n2772 ^ n2771 ^ 1'b0 ;
  assign n2770 = ( n1275 & ~n1783 ) | ( n1275 & n2183 ) | ( ~n1783 & n2183 ) ;
  assign n2767 = x150 & n1036 ;
  assign n2768 = ~n1768 & n2767 ;
  assign n2769 = n2768 ^ x128 ^ 1'b0 ;
  assign n2774 = n2773 ^ n2770 ^ n2769 ;
  assign n2775 = ( x147 & n1062 ) | ( x147 & n1821 ) | ( n1062 & n1821 ) ;
  assign n2776 = n411 & n1688 ;
  assign n2777 = n2776 ^ n2384 ^ 1'b0 ;
  assign n2778 = ~n1553 & n2777 ;
  assign n2779 = n2190 ^ n936 ^ 1'b0 ;
  assign n2780 = n1506 & ~n2779 ;
  assign n2781 = ~n752 & n1253 ;
  assign n2782 = ~n776 & n2781 ;
  assign n2783 = n2782 ^ n488 ^ 1'b0 ;
  assign n2785 = n2148 ^ n1233 ^ n570 ;
  assign n2784 = n1295 & ~n1947 ;
  assign n2786 = n2785 ^ n2784 ^ 1'b0 ;
  assign n2787 = ( n798 & n882 ) | ( n798 & ~n1349 ) | ( n882 & ~n1349 ) ;
  assign n2788 = n331 | n1720 ;
  assign n2789 = n2788 ^ n2548 ^ 1'b0 ;
  assign n2790 = n1831 & ~n2789 ;
  assign n2791 = n991 & n2790 ;
  assign n2792 = n1592 ^ n281 ^ 1'b0 ;
  assign n2793 = ~n778 & n2792 ;
  assign n2794 = n2793 ^ n1760 ^ n570 ;
  assign n2795 = n2794 ^ n1780 ^ n1387 ;
  assign n2796 = ( n2543 & n2746 ) | ( n2543 & ~n2795 ) | ( n2746 & ~n2795 ) ;
  assign n2797 = n1064 ^ x49 ^ 1'b0 ;
  assign n2798 = n981 & n2797 ;
  assign n2799 = ~n847 & n2798 ;
  assign n2800 = ~x30 & n1555 ;
  assign n2801 = n383 | n1368 ;
  assign n2802 = n2801 ^ n2164 ^ 1'b0 ;
  assign n2803 = n601 ^ x253 ^ 1'b0 ;
  assign n2804 = x118 & n2803 ;
  assign n2805 = n2285 & n2804 ;
  assign n2806 = n2805 ^ n1113 ^ 1'b0 ;
  assign n2807 = n1382 ^ n1254 ^ x175 ;
  assign n2808 = x162 | n2807 ;
  assign n2809 = n732 & ~n2694 ;
  assign n2810 = ~n560 & n2809 ;
  assign n2811 = ( n332 & n1789 ) | ( n332 & n2289 ) | ( n1789 & n2289 ) ;
  assign n2812 = ( n587 & n2473 ) | ( n587 & n2811 ) | ( n2473 & n2811 ) ;
  assign n2813 = n327 & n392 ;
  assign n2814 = n335 & n2813 ;
  assign n2815 = n527 | n557 ;
  assign n2816 = ( n989 & n2814 ) | ( n989 & ~n2815 ) | ( n2814 & ~n2815 ) ;
  assign n2817 = n612 | n2816 ;
  assign n2818 = ~n1084 & n1312 ;
  assign n2819 = ( n1949 & n2344 ) | ( n1949 & ~n2818 ) | ( n2344 & ~n2818 ) ;
  assign n2820 = x29 & n903 ;
  assign n2821 = n302 & n2820 ;
  assign n2822 = n2557 & ~n2821 ;
  assign n2823 = ~n411 & n2822 ;
  assign n2824 = n2823 ^ n2202 ^ n512 ;
  assign n2825 = n869 & n2399 ;
  assign n2826 = n2824 & n2825 ;
  assign n2827 = n643 ^ n607 ^ x94 ;
  assign n2828 = ~n776 & n1166 ;
  assign n2829 = ~x42 & n2828 ;
  assign n2830 = n2829 ^ n1605 ^ 1'b0 ;
  assign n2831 = n1459 & ~n2830 ;
  assign n2832 = n358 | n2831 ;
  assign n2833 = n2827 | n2832 ;
  assign n2839 = n1484 ^ n1323 ^ 1'b0 ;
  assign n2834 = n2689 ^ n1469 ^ x173 ;
  assign n2835 = n2834 ^ n976 ^ 1'b0 ;
  assign n2836 = n526 & ~n2835 ;
  assign n2837 = ~n1291 & n2836 ;
  assign n2838 = n2837 ^ n633 ^ 1'b0 ;
  assign n2840 = n2839 ^ n2838 ^ 1'b0 ;
  assign n2841 = n773 & n2840 ;
  assign n2842 = n907 & n1575 ;
  assign n2843 = ~n1855 & n2842 ;
  assign n2844 = x147 & ~n2843 ;
  assign n2845 = n1693 ^ n1528 ^ 1'b0 ;
  assign n2846 = n2844 & ~n2845 ;
  assign n2847 = x179 & n1415 ;
  assign n2848 = ~n1912 & n2847 ;
  assign n2849 = n2332 & n2848 ;
  assign n2850 = n2849 ^ n587 ^ 1'b0 ;
  assign n2852 = ~x56 & x172 ;
  assign n2851 = n1996 ^ n647 ^ 1'b0 ;
  assign n2853 = n2852 ^ n2851 ^ n1611 ;
  assign n2854 = x34 & ~x90 ;
  assign n2855 = n2672 ^ n1052 ^ n660 ;
  assign n2856 = ( n342 & ~n1121 ) | ( n342 & n2855 ) | ( ~n1121 & n2855 ) ;
  assign n2857 = n1551 & n2856 ;
  assign n2858 = n2857 ^ x91 ^ 1'b0 ;
  assign n2859 = x21 & ~n2858 ;
  assign n2860 = x178 & n2859 ;
  assign n2861 = n1220 ^ x236 ^ 1'b0 ;
  assign n2862 = x227 & n2861 ;
  assign n2863 = n395 & n2527 ;
  assign n2864 = n2863 ^ x38 ^ 1'b0 ;
  assign n2865 = n702 | n948 ;
  assign n2866 = n2864 & ~n2865 ;
  assign n2867 = n1965 & ~n2866 ;
  assign n2868 = ~n2862 & n2867 ;
  assign n2869 = n865 & n2437 ;
  assign n2870 = n2869 ^ x29 ^ 1'b0 ;
  assign n2871 = n2870 ^ n1858 ^ n545 ;
  assign n2872 = x127 & n2871 ;
  assign n2873 = n2872 ^ n1793 ^ 1'b0 ;
  assign n2874 = x13 & n1192 ;
  assign n2875 = n2874 ^ n538 ^ 1'b0 ;
  assign n2876 = n2048 & ~n2875 ;
  assign n2877 = n2876 ^ n663 ^ 1'b0 ;
  assign n2878 = n1746 & n2877 ;
  assign n2879 = ~n2217 & n2878 ;
  assign n2880 = n1269 & ~n2879 ;
  assign n2881 = n2880 ^ n481 ^ 1'b0 ;
  assign n2882 = n2455 & n2697 ;
  assign n2883 = n1987 ^ n1612 ^ 1'b0 ;
  assign n2884 = ( ~n704 & n1421 ) | ( ~n704 & n1851 ) | ( n1421 & n1851 ) ;
  assign n2885 = n939 ^ n582 ^ 1'b0 ;
  assign n2886 = n1959 & n2885 ;
  assign n2887 = n1707 & n2886 ;
  assign n2888 = n2887 ^ n256 ^ 1'b0 ;
  assign n2889 = n2888 ^ n2692 ^ 1'b0 ;
  assign n2890 = n2281 & n2889 ;
  assign n2891 = n2122 & ~n2483 ;
  assign n2892 = n2891 ^ x164 ^ 1'b0 ;
  assign n2893 = n2873 ^ n2783 ^ 1'b0 ;
  assign n2894 = n854 & n1880 ;
  assign n2895 = ~n879 & n2894 ;
  assign n2896 = n902 ^ n861 ^ 1'b0 ;
  assign n2897 = n1053 & ~n2896 ;
  assign n2898 = n2269 ^ n745 ^ 1'b0 ;
  assign n2899 = n2793 ^ n1470 ^ 1'b0 ;
  assign n2900 = ~x72 & n1013 ;
  assign n2901 = x209 & n983 ;
  assign n2902 = n2901 ^ n2347 ^ 1'b0 ;
  assign n2903 = ( ~n2635 & n2641 ) | ( ~n2635 & n2902 ) | ( n2641 & n2902 ) ;
  assign n2904 = n645 | n1356 ;
  assign n2905 = n2904 ^ n1601 ^ 1'b0 ;
  assign n2906 = ~n491 & n2905 ;
  assign n2907 = n2906 ^ n410 ^ 1'b0 ;
  assign n2908 = n2070 ^ n2033 ^ 1'b0 ;
  assign n2909 = n2011 & ~n2908 ;
  assign n2910 = n772 | n2909 ;
  assign n2912 = n277 ^ x182 ^ 1'b0 ;
  assign n2913 = n413 & n2912 ;
  assign n2911 = ~n322 & n1130 ;
  assign n2914 = n2913 ^ n2911 ^ 1'b0 ;
  assign n2915 = n2914 ^ n2630 ^ n2248 ;
  assign n2916 = ~n1055 & n2915 ;
  assign n2920 = n759 & ~n954 ;
  assign n2921 = n2920 ^ n456 ^ 1'b0 ;
  assign n2917 = n1186 | n2067 ;
  assign n2918 = n2230 | n2917 ;
  assign n2919 = ~n2855 & n2918 ;
  assign n2922 = n2921 ^ n2919 ^ 1'b0 ;
  assign n2923 = ~x15 & n1348 ;
  assign n2924 = n2923 ^ n985 ^ 1'b0 ;
  assign n2925 = ( n1798 & ~n1981 ) | ( n1798 & n2924 ) | ( ~n1981 & n2924 ) ;
  assign n2926 = n593 | n2067 ;
  assign n2927 = n2926 ^ x50 ^ 1'b0 ;
  assign n2928 = n1555 ^ n340 ^ 1'b0 ;
  assign n2929 = x96 & n2928 ;
  assign n2930 = n1924 ^ n471 ^ 1'b0 ;
  assign n2931 = n2929 & n2930 ;
  assign n2932 = n2931 ^ n2913 ^ 1'b0 ;
  assign n2934 = n622 & n1571 ;
  assign n2935 = ~n520 & n2934 ;
  assign n2933 = x74 & ~n1314 ;
  assign n2936 = n2935 ^ n2933 ^ 1'b0 ;
  assign n2937 = n683 ^ x17 ^ 1'b0 ;
  assign n2938 = n1637 & n2587 ;
  assign n2939 = n2938 ^ n1261 ^ 1'b0 ;
  assign n2940 = ~n867 & n2939 ;
  assign n2941 = n2940 ^ n1311 ^ 1'b0 ;
  assign n2942 = n2941 ^ x159 ^ x2 ;
  assign n2943 = n1874 ^ n791 ^ 1'b0 ;
  assign n2944 = n842 ^ n600 ^ 1'b0 ;
  assign n2945 = x2 & ~n2944 ;
  assign n2946 = n2943 & ~n2945 ;
  assign n2947 = n1377 ^ x185 ^ 1'b0 ;
  assign n2948 = n1027 & ~n1387 ;
  assign n2949 = n2948 ^ n1096 ^ 1'b0 ;
  assign n2950 = ( n453 & ~n1085 ) | ( n453 & n2949 ) | ( ~n1085 & n2949 ) ;
  assign n2951 = n2950 ^ n2051 ^ x56 ;
  assign n2952 = ~n2550 & n2951 ;
  assign n2953 = ( x62 & ~x130 ) | ( x62 & n706 ) | ( ~x130 & n706 ) ;
  assign n2955 = n785 ^ n520 ^ 1'b0 ;
  assign n2956 = n2955 ^ n1281 ^ x31 ;
  assign n2954 = n1349 & n1728 ;
  assign n2957 = n2956 ^ n2954 ^ n2250 ;
  assign n2958 = n2296 ^ n1689 ^ x121 ;
  assign n2959 = n2958 ^ n1337 ^ 1'b0 ;
  assign n2960 = n1750 ^ n1011 ^ 1'b0 ;
  assign n2961 = ( n1003 & ~n2959 ) | ( n1003 & n2960 ) | ( ~n2959 & n2960 ) ;
  assign n2964 = x216 & n946 ;
  assign n2965 = n2964 ^ x29 ^ 1'b0 ;
  assign n2966 = n2965 ^ n1633 ^ x39 ;
  assign n2963 = n905 ^ n727 ^ x148 ;
  assign n2967 = n2966 ^ n2963 ^ 1'b0 ;
  assign n2962 = n1315 & ~n1633 ;
  assign n2968 = n2967 ^ n2962 ^ 1'b0 ;
  assign n2970 = n2118 ^ n438 ^ x87 ;
  assign n2969 = n462 & ~n498 ;
  assign n2971 = n2970 ^ n2969 ^ n1937 ;
  assign n2972 = ( ~n1425 & n1527 ) | ( ~n1425 & n1702 ) | ( n1527 & n1702 ) ;
  assign n2973 = ~x241 & n2972 ;
  assign n2975 = ~n1004 & n1217 ;
  assign n2974 = x105 & ~n582 ;
  assign n2976 = n2975 ^ n2974 ^ 1'b0 ;
  assign n2978 = n480 | n944 ;
  assign n2979 = n456 | n2978 ;
  assign n2980 = n2690 ^ n286 ^ 1'b0 ;
  assign n2981 = n2979 & ~n2980 ;
  assign n2977 = n1533 | n1706 ;
  assign n2982 = n2981 ^ n2977 ^ 1'b0 ;
  assign n2983 = ( x71 & n1067 ) | ( x71 & n1900 ) | ( n1067 & n1900 ) ;
  assign n2984 = n2759 ^ x254 ^ 1'b0 ;
  assign n2985 = n935 & ~n2207 ;
  assign n2986 = n2985 ^ x172 ^ 1'b0 ;
  assign n2987 = n1685 | n2986 ;
  assign n2988 = n1459 | n2987 ;
  assign n2989 = ( n849 & n852 ) | ( n849 & n2988 ) | ( n852 & n2988 ) ;
  assign n2990 = n2118 | n2989 ;
  assign n2991 = ( n505 & ~n1152 ) | ( n505 & n2402 ) | ( ~n1152 & n2402 ) ;
  assign n2992 = n884 ^ n417 ^ 1'b0 ;
  assign n2993 = n2991 & n2992 ;
  assign n2994 = n267 | n1073 ;
  assign n2995 = n2994 ^ n335 ^ 1'b0 ;
  assign n2996 = ~n1106 & n2224 ;
  assign n2997 = n1548 ^ n1158 ^ 1'b0 ;
  assign n2998 = x27 & n2997 ;
  assign n2999 = n863 ^ x94 ^ 1'b0 ;
  assign n3000 = x210 & ~n2999 ;
  assign n3001 = ( n1419 & ~n2937 ) | ( n1419 & n3000 ) | ( ~n2937 & n3000 ) ;
  assign n3002 = n2244 ^ n1709 ^ x81 ;
  assign n3003 = n1626 ^ n711 ^ n335 ;
  assign n3004 = n1021 & ~n3003 ;
  assign n3005 = n1462 & n3004 ;
  assign n3007 = ~n2131 & n2194 ;
  assign n3008 = ( x88 & ~n1789 ) | ( x88 & n3007 ) | ( ~n1789 & n3007 ) ;
  assign n3009 = n2664 ^ n2513 ^ 1'b0 ;
  assign n3010 = n3008 & n3009 ;
  assign n3006 = x112 & ~n1395 ;
  assign n3011 = n3010 ^ n3006 ^ 1'b0 ;
  assign n3012 = ~n729 & n1323 ;
  assign n3013 = ~n560 & n3012 ;
  assign n3014 = n3013 ^ n2298 ^ 1'b0 ;
  assign n3015 = n3014 ^ n2871 ^ 1'b0 ;
  assign n3016 = n2277 & n3015 ;
  assign n3017 = n659 & n1038 ;
  assign n3018 = n261 & n3017 ;
  assign n3019 = n572 ^ x117 ^ 1'b0 ;
  assign n3020 = x208 & ~n3019 ;
  assign n3021 = n3020 ^ x82 ^ 1'b0 ;
  assign n3022 = n2012 ^ n271 ^ 1'b0 ;
  assign n3023 = ~n3021 & n3022 ;
  assign n3024 = n3023 ^ n1317 ^ n258 ;
  assign n3025 = ( n993 & n3018 ) | ( n993 & n3024 ) | ( n3018 & n3024 ) ;
  assign n3026 = n3025 ^ n1651 ^ 1'b0 ;
  assign n3027 = n3016 | n3026 ;
  assign n3028 = n2518 | n3027 ;
  assign n3029 = n3028 ^ n548 ^ 1'b0 ;
  assign n3034 = x244 & ~n2426 ;
  assign n3030 = n486 & n2015 ;
  assign n3031 = n3030 ^ n538 ^ 1'b0 ;
  assign n3032 = ~n1394 & n3031 ;
  assign n3033 = ~n2630 & n3032 ;
  assign n3035 = n3034 ^ n3033 ^ 1'b0 ;
  assign n3037 = x145 & n385 ;
  assign n3038 = n2272 & n3037 ;
  assign n3039 = ( n858 & n2574 ) | ( n858 & n3038 ) | ( n2574 & n3038 ) ;
  assign n3036 = n1996 ^ x149 ^ 1'b0 ;
  assign n3040 = n3039 ^ n3036 ^ n1416 ;
  assign n3041 = x195 | n2074 ;
  assign n3042 = n3041 ^ n1214 ^ 1'b0 ;
  assign n3043 = n2856 & n3042 ;
  assign n3044 = n694 ^ x164 ^ 1'b0 ;
  assign n3045 = n3043 & ~n3044 ;
  assign n3047 = n482 & n1975 ;
  assign n3046 = n1692 & n1866 ;
  assign n3048 = n3047 ^ n3046 ^ 1'b0 ;
  assign n3049 = ~n1069 & n2979 ;
  assign n3050 = ~n2181 & n3049 ;
  assign n3051 = n2853 ^ n1708 ^ 1'b0 ;
  assign n3052 = x206 & ~n2971 ;
  assign n3053 = ~x90 & n587 ;
  assign n3054 = ~n1595 & n3053 ;
  assign n3055 = n798 & n3054 ;
  assign n3056 = n3055 ^ n2512 ^ 1'b0 ;
  assign n3057 = n639 ^ x7 ^ 1'b0 ;
  assign n3058 = n2409 | n3057 ;
  assign n3059 = n894 & n2597 ;
  assign n3060 = n3059 ^ x246 ^ 1'b0 ;
  assign n3061 = ( x84 & n275 ) | ( x84 & ~n481 ) | ( n275 & ~n481 ) ;
  assign n3062 = n3061 ^ n1912 ^ 1'b0 ;
  assign n3063 = n718 ^ n455 ^ 1'b0 ;
  assign n3064 = n3063 ^ n1658 ^ n840 ;
  assign n3065 = x76 & n1113 ;
  assign n3066 = n3065 ^ n661 ^ 1'b0 ;
  assign n3067 = ~n2345 & n3066 ;
  assign n3068 = n585 & ~n1418 ;
  assign n3069 = x214 & n2298 ;
  assign n3070 = n3069 ^ n269 ^ 1'b0 ;
  assign n3071 = n2806 & ~n3070 ;
  assign n3072 = n1358 ^ x163 ^ 1'b0 ;
  assign n3073 = ( n269 & ~n755 ) | ( n269 & n3072 ) | ( ~n755 & n3072 ) ;
  assign n3074 = n3073 ^ n867 ^ 1'b0 ;
  assign n3076 = n3000 ^ n2380 ^ 1'b0 ;
  assign n3077 = n1823 | n3076 ;
  assign n3075 = n572 | n1823 ;
  assign n3078 = n3077 ^ n3075 ^ 1'b0 ;
  assign n3079 = n1373 | n1926 ;
  assign n3080 = n1871 & n2558 ;
  assign n3081 = n3080 ^ n366 ^ 1'b0 ;
  assign n3082 = n3021 | n3081 ;
  assign n3083 = n3079 & n3082 ;
  assign n3084 = ~n2178 & n3083 ;
  assign n3085 = n2882 ^ x133 ^ 1'b0 ;
  assign n3086 = n1036 & n2902 ;
  assign n3087 = n2380 & n3086 ;
  assign n3088 = ( n291 & n1027 ) | ( n291 & ~n1832 ) | ( n1027 & ~n1832 ) ;
  assign n3089 = n3088 ^ n379 ^ 1'b0 ;
  assign n3090 = n3089 ^ n2260 ^ 1'b0 ;
  assign n3091 = n1645 | n2918 ;
  assign n3092 = n686 & ~n1917 ;
  assign n3093 = n3092 ^ x76 ^ 1'b0 ;
  assign n3094 = n1739 ^ n516 ^ x222 ;
  assign n3095 = ~n861 & n3094 ;
  assign n3096 = ~n1013 & n1889 ;
  assign n3097 = n3096 ^ n930 ^ 1'b0 ;
  assign n3098 = ~n759 & n3097 ;
  assign n3099 = n3098 ^ n707 ^ x134 ;
  assign n3100 = ( ~x69 & n2335 ) | ( ~x69 & n3099 ) | ( n2335 & n3099 ) ;
  assign n3101 = x126 & n2201 ;
  assign n3102 = n3101 ^ n1378 ^ 1'b0 ;
  assign n3103 = n3102 ^ n1925 ^ 1'b0 ;
  assign n3104 = ( n1340 & n2203 ) | ( n1340 & ~n3103 ) | ( n2203 & ~n3103 ) ;
  assign n3105 = ~n593 & n2778 ;
  assign n3106 = n3105 ^ n2610 ^ 1'b0 ;
  assign n3107 = ( ~n915 & n1917 ) | ( ~n915 & n2008 ) | ( n1917 & n2008 ) ;
  assign n3108 = n755 & ~n3107 ;
  assign n3109 = n3108 ^ n2148 ^ 1'b0 ;
  assign n3110 = n2047 & ~n2623 ;
  assign n3111 = n3110 ^ n1106 ^ 1'b0 ;
  assign n3112 = n2002 ^ n327 ^ 1'b0 ;
  assign n3113 = n2230 ^ n1160 ^ 1'b0 ;
  assign n3114 = ~n1717 & n3113 ;
  assign n3115 = n3114 ^ n614 ^ 1'b0 ;
  assign n3116 = n1648 ^ n332 ^ 1'b0 ;
  assign n3117 = n1439 ^ n1024 ^ 1'b0 ;
  assign n3118 = x184 & n3117 ;
  assign n3119 = ~n2224 & n3118 ;
  assign n3120 = n3119 ^ n1027 ^ 1'b0 ;
  assign n3121 = n2577 ^ n2536 ^ 1'b0 ;
  assign n3122 = n946 & ~n1709 ;
  assign n3123 = n3122 ^ n2255 ^ 1'b0 ;
  assign n3124 = x170 | n3123 ;
  assign n3125 = ~n1541 & n2004 ;
  assign n3126 = n3125 ^ n648 ^ 1'b0 ;
  assign n3127 = x143 ^ x69 ^ x7 ;
  assign n3128 = n890 | n3127 ;
  assign n3129 = ( x225 & n3126 ) | ( x225 & ~n3128 ) | ( n3126 & ~n3128 ) ;
  assign n3130 = x70 & x181 ;
  assign n3131 = ~n265 & n3130 ;
  assign n3132 = ~n1038 & n2100 ;
  assign n3133 = n3131 | n3132 ;
  assign n3134 = ( x196 & ~n2421 ) | ( x196 & n2871 ) | ( ~n2421 & n2871 ) ;
  assign n3137 = n365 | n480 ;
  assign n3138 = n3137 ^ n1780 ^ 1'b0 ;
  assign n3135 = ( n535 & ~n635 ) | ( n535 & n805 ) | ( ~n635 & n805 ) ;
  assign n3136 = n3135 ^ n2548 ^ n1064 ;
  assign n3139 = n3138 ^ n3136 ^ n1462 ;
  assign n3140 = n1702 & ~n3139 ;
  assign n3141 = ( ~n2237 & n2368 ) | ( ~n2237 & n3140 ) | ( n2368 & n3140 ) ;
  assign n3143 = n1259 & n1737 ;
  assign n3144 = n3143 ^ n1210 ^ 1'b0 ;
  assign n3142 = ( n598 & n742 ) | ( n598 & ~n1814 ) | ( n742 & ~n1814 ) ;
  assign n3145 = n3144 ^ n3142 ^ 1'b0 ;
  assign n3146 = n405 & n2006 ;
  assign n3147 = ~n2797 & n3146 ;
  assign n3148 = n956 ^ n905 ^ n405 ;
  assign n3149 = n3148 ^ n2627 ^ 1'b0 ;
  assign n3150 = n3149 ^ x174 ^ 1'b0 ;
  assign n3151 = n1885 | n3150 ;
  assign n3152 = n1530 & ~n3151 ;
  assign n3153 = ( ~n1477 & n3147 ) | ( ~n1477 & n3152 ) | ( n3147 & n3152 ) ;
  assign n3154 = n508 | n1122 ;
  assign n3155 = n3154 ^ n1882 ^ 1'b0 ;
  assign n3156 = n2512 | n3155 ;
  assign n3157 = n1880 ^ n826 ^ 1'b0 ;
  assign n3158 = x18 & ~n3157 ;
  assign n3160 = ~n948 & n2935 ;
  assign n3159 = n761 & ~n1729 ;
  assign n3161 = n3160 ^ n3159 ^ 1'b0 ;
  assign n3162 = n596 & n3161 ;
  assign n3163 = ~n1147 & n3162 ;
  assign n3164 = n2311 & ~n2853 ;
  assign n3169 = ~x235 & n706 ;
  assign n3170 = n1203 | n3169 ;
  assign n3165 = n597 ^ n491 ^ 1'b0 ;
  assign n3166 = n860 & n3165 ;
  assign n3167 = ~n502 & n3166 ;
  assign n3168 = ~x6 & n3167 ;
  assign n3171 = n3170 ^ n3168 ^ 1'b0 ;
  assign n3173 = n522 | n1711 ;
  assign n3174 = n1150 | n3173 ;
  assign n3172 = ( n1060 & n1535 ) | ( n1060 & ~n1725 ) | ( n1535 & ~n1725 ) ;
  assign n3175 = n3174 ^ n3172 ^ n600 ;
  assign n3176 = ~n998 & n3175 ;
  assign n3177 = n2070 | n2732 ;
  assign n3178 = n3177 ^ n2140 ^ 1'b0 ;
  assign n3179 = n2580 ^ x176 ^ 1'b0 ;
  assign n3180 = n3178 & ~n3179 ;
  assign n3184 = n967 ^ n365 ^ 1'b0 ;
  assign n3185 = n2224 & n3184 ;
  assign n3181 = x137 & ~n365 ;
  assign n3182 = n3181 ^ n1354 ^ 1'b0 ;
  assign n3183 = n3182 ^ n1608 ^ n1162 ;
  assign n3186 = n3185 ^ n3183 ^ 1'b0 ;
  assign n3187 = x169 & n3186 ;
  assign n3193 = n1044 ^ x94 ^ 1'b0 ;
  assign n3194 = n3193 ^ n3038 ^ 1'b0 ;
  assign n3195 = n952 | n3194 ;
  assign n3188 = ~n471 & n1998 ;
  assign n3189 = ~n543 & n3188 ;
  assign n3190 = n1932 & ~n3189 ;
  assign n3191 = n3190 ^ n2448 ^ 1'b0 ;
  assign n3192 = n505 & n3191 ;
  assign n3196 = n3195 ^ n3192 ^ 1'b0 ;
  assign n3197 = n541 | n1593 ;
  assign n3198 = n351 & ~n3197 ;
  assign n3199 = n3198 ^ n1462 ^ 1'b0 ;
  assign n3200 = x112 & n2024 ;
  assign n3201 = ~n1741 & n3200 ;
  assign n3202 = x121 & n1894 ;
  assign n3203 = n3202 ^ n1223 ^ x193 ;
  assign n3204 = n1416 & ~n3021 ;
  assign n3205 = n721 ^ x47 ^ 1'b0 ;
  assign n3206 = n2746 & ~n3205 ;
  assign n3207 = n963 & n3206 ;
  assign n3208 = ~n1152 & n1733 ;
  assign n3209 = n3208 ^ x123 ^ 1'b0 ;
  assign n3210 = n3209 ^ n1693 ^ n860 ;
  assign n3211 = x40 & n2651 ;
  assign n3212 = n3211 ^ n835 ^ 1'b0 ;
  assign n3213 = n1275 & ~n3212 ;
  assign n3222 = n840 & n1040 ;
  assign n3214 = n2282 ^ n847 ^ 1'b0 ;
  assign n3215 = n2617 & n3214 ;
  assign n3216 = ( n1373 & ~n2327 ) | ( n1373 & n3215 ) | ( ~n2327 & n3215 ) ;
  assign n3217 = n1003 | n2171 ;
  assign n3218 = n935 | n3217 ;
  assign n3219 = ~x244 & n3218 ;
  assign n3220 = n3216 & n3219 ;
  assign n3221 = n2895 | n3220 ;
  assign n3223 = n3222 ^ n3221 ^ 1'b0 ;
  assign n3224 = n1416 ^ n984 ^ 1'b0 ;
  assign n3225 = n3097 & n3224 ;
  assign n3226 = n1184 & ~n1890 ;
  assign n3227 = n1330 & n3226 ;
  assign n3228 = n3227 ^ n1075 ^ 1'b0 ;
  assign n3229 = n1360 ^ n982 ^ n940 ;
  assign n3230 = ( n3225 & n3228 ) | ( n3225 & ~n3229 ) | ( n3228 & ~n3229 ) ;
  assign n3231 = ( ~x101 & n1095 ) | ( ~x101 & n2664 ) | ( n1095 & n2664 ) ;
  assign n3232 = n3231 ^ n441 ^ 1'b0 ;
  assign n3233 = n3232 ^ n2768 ^ x210 ;
  assign n3234 = ~n301 & n2102 ;
  assign n3235 = n2969 & n3234 ;
  assign n3236 = n1653 ^ n439 ^ 1'b0 ;
  assign n3237 = n2968 & ~n3236 ;
  assign n3238 = n2292 ^ n1629 ^ 1'b0 ;
  assign n3239 = ~n1067 & n3238 ;
  assign n3240 = n924 & n3239 ;
  assign n3241 = n1155 ^ n707 ^ 1'b0 ;
  assign n3243 = x26 & x194 ;
  assign n3244 = n3243 ^ n2247 ^ 1'b0 ;
  assign n3245 = ( ~n1058 & n2637 ) | ( ~n1058 & n3244 ) | ( n2637 & n3244 ) ;
  assign n3246 = n2989 & n3245 ;
  assign n3247 = n2709 ^ n1579 ^ 1'b0 ;
  assign n3248 = n3246 | n3247 ;
  assign n3242 = ( n344 & n1384 ) | ( n344 & ~n2575 ) | ( n1384 & ~n2575 ) ;
  assign n3249 = n3248 ^ n3242 ^ x200 ;
  assign n3253 = n1570 | n1594 ;
  assign n3254 = n3253 ^ n2164 ^ x102 ;
  assign n3250 = n1062 & n3229 ;
  assign n3251 = ~n1752 & n3250 ;
  assign n3252 = n665 | n3251 ;
  assign n3255 = n3254 ^ n3252 ^ 1'b0 ;
  assign n3256 = ( n387 & n2431 ) | ( n387 & n3067 ) | ( n2431 & n3067 ) ;
  assign n3257 = n2169 ^ x103 ^ 1'b0 ;
  assign n3258 = ~n1353 & n3257 ;
  assign n3259 = n3258 ^ n1624 ^ 1'b0 ;
  assign n3260 = n2022 & n3259 ;
  assign n3261 = n3260 ^ n629 ^ 1'b0 ;
  assign n3262 = n1033 ^ n956 ^ 1'b0 ;
  assign n3263 = ~n3261 & n3262 ;
  assign n3264 = ( n2404 & ~n2413 ) | ( n2404 & n3263 ) | ( ~n2413 & n3263 ) ;
  assign n3265 = n2647 ^ n1474 ^ 1'b0 ;
  assign n3266 = x219 & ~n2155 ;
  assign n3267 = n3266 ^ n1728 ^ 1'b0 ;
  assign n3270 = x190 & ~n887 ;
  assign n3271 = ~n2450 & n3270 ;
  assign n3268 = x75 & n2443 ;
  assign n3269 = n3268 ^ n256 ^ 1'b0 ;
  assign n3272 = n3271 ^ n3269 ^ 1'b0 ;
  assign n3273 = x64 & ~n2450 ;
  assign n3274 = n3230 ^ x111 ^ 1'b0 ;
  assign n3278 = x29 & n2513 ;
  assign n3279 = n3278 ^ x239 ^ 1'b0 ;
  assign n3280 = n3279 ^ n3024 ^ 1'b0 ;
  assign n3281 = ~n3232 & n3280 ;
  assign n3275 = n349 | n935 ;
  assign n3276 = n1627 ^ x77 ^ 1'b0 ;
  assign n3277 = n3275 & n3276 ;
  assign n3282 = n3281 ^ n3277 ^ 1'b0 ;
  assign n3285 = n1785 & n2237 ;
  assign n3286 = n648 & n3285 ;
  assign n3287 = n560 & n3286 ;
  assign n3288 = n2362 & ~n3287 ;
  assign n3283 = n319 ^ x74 ^ 1'b0 ;
  assign n3284 = n832 & ~n3283 ;
  assign n3289 = n3288 ^ n3284 ^ 1'b0 ;
  assign n3290 = n601 & ~n1031 ;
  assign n3291 = n3290 ^ x219 ^ 1'b0 ;
  assign n3292 = ~n863 & n3291 ;
  assign n3293 = ( n686 & n828 ) | ( n686 & n1527 ) | ( n828 & n1527 ) ;
  assign n3294 = ( ~x59 & n1827 ) | ( ~x59 & n3293 ) | ( n1827 & n3293 ) ;
  assign n3295 = ( x122 & n304 ) | ( x122 & n322 ) | ( n304 & n322 ) ;
  assign n3296 = n3295 ^ x142 ^ 1'b0 ;
  assign n3297 = n1356 | n3279 ;
  assign n3298 = x188 & ~n753 ;
  assign n3299 = n1512 & n3298 ;
  assign n3300 = n3299 ^ n1444 ^ 1'b0 ;
  assign n3301 = ( ~n822 & n2935 ) | ( ~n822 & n3300 ) | ( n2935 & n3300 ) ;
  assign n3302 = n306 & n3301 ;
  assign n3303 = n838 | n1127 ;
  assign n3304 = n3303 ^ n431 ^ 1'b0 ;
  assign n3305 = n3304 ^ n2040 ^ 1'b0 ;
  assign n3306 = n3305 ^ n2636 ^ 1'b0 ;
  assign n3307 = ( n587 & n944 ) | ( n587 & ~n2885 ) | ( n944 & ~n2885 ) ;
  assign n3308 = n3307 ^ n2274 ^ n1786 ;
  assign n3309 = x184 ^ x74 ^ 1'b0 ;
  assign n3310 = ~n2156 & n3309 ;
  assign n3311 = n3310 ^ n1484 ^ n718 ;
  assign n3312 = n2799 & ~n3311 ;
  assign n3313 = n395 & ~n2925 ;
  assign n3314 = n1791 ^ n490 ^ 1'b0 ;
  assign n3315 = n1726 | n3314 ;
  assign n3316 = n856 & ~n3315 ;
  assign n3317 = ~n3287 & n3316 ;
  assign n3318 = n2527 ^ n872 ^ n367 ;
  assign n3319 = x83 & ~n2955 ;
  assign n3320 = ~n854 & n3319 ;
  assign n3321 = n3320 ^ n2279 ^ 1'b0 ;
  assign n3322 = ( ~x212 & x247 ) | ( ~x212 & n3321 ) | ( x247 & n3321 ) ;
  assign n3323 = n2725 ^ n712 ^ 1'b0 ;
  assign n3324 = n878 | n3323 ;
  assign n3325 = n1110 | n1877 ;
  assign n3326 = ( n2573 & ~n2618 ) | ( n2573 & n2674 ) | ( ~n2618 & n2674 ) ;
  assign n3327 = n1246 & n3166 ;
  assign n3328 = ~n1813 & n3327 ;
  assign n3329 = x128 & ~n3328 ;
  assign n3330 = n3329 ^ n2573 ^ 1'b0 ;
  assign n3331 = n1079 | n3330 ;
  assign n3332 = n2547 | n3331 ;
  assign n3333 = ~x176 & n2276 ;
  assign n3334 = n3333 ^ n2465 ^ 1'b0 ;
  assign n3335 = n831 ^ n327 ^ 1'b0 ;
  assign n3336 = x3 & n3335 ;
  assign n3337 = n1538 | n2097 ;
  assign n3338 = n3336 | n3337 ;
  assign n3339 = n3338 ^ n2207 ^ 1'b0 ;
  assign n3340 = n2637 | n3339 ;
  assign n3341 = n2851 ^ n273 ^ 1'b0 ;
  assign n3342 = n516 | n3341 ;
  assign n3343 = ( ~x83 & n1917 ) | ( ~x83 & n2050 ) | ( n1917 & n2050 ) ;
  assign n3344 = ( x114 & n2782 ) | ( x114 & ~n3343 ) | ( n2782 & ~n3343 ) ;
  assign n3345 = n1650 & ~n2467 ;
  assign n3346 = n1462 & n3345 ;
  assign n3347 = ~n1587 & n3346 ;
  assign n3348 = x19 & n3347 ;
  assign n3349 = ~n685 & n2517 ;
  assign n3350 = ~n3138 & n3349 ;
  assign n3351 = n2575 ^ n1330 ^ 1'b0 ;
  assign n3352 = ~n3350 & n3351 ;
  assign n3353 = n1355 | n1777 ;
  assign n3354 = n3353 ^ n778 ^ 1'b0 ;
  assign n3359 = ( n399 & n634 ) | ( n399 & ~n1260 ) | ( n634 & ~n1260 ) ;
  assign n3356 = ~n681 & n2009 ;
  assign n3357 = n1957 & n3356 ;
  assign n3358 = x92 & ~n3357 ;
  assign n3360 = n3359 ^ n3358 ^ 1'b0 ;
  assign n3355 = n1308 | n2630 ;
  assign n3361 = n3360 ^ n3355 ^ 1'b0 ;
  assign n3362 = ( n2247 & n2974 ) | ( n2247 & n3361 ) | ( n2974 & n3361 ) ;
  assign n3363 = n2525 ^ n1884 ^ 1'b0 ;
  assign n3364 = ~n1993 & n2736 ;
  assign n3365 = n2097 & n3364 ;
  assign n3366 = n3363 & ~n3365 ;
  assign n3367 = ( n1620 & n2626 ) | ( n1620 & ~n2775 ) | ( n2626 & ~n2775 ) ;
  assign n3368 = n286 | n1115 ;
  assign n3369 = x82 | n3368 ;
  assign n3372 = x34 & x72 ;
  assign n3373 = n3372 ^ n1558 ^ 1'b0 ;
  assign n3370 = x0 & ~n675 ;
  assign n3371 = n3370 ^ n1470 ^ 1'b0 ;
  assign n3374 = n3373 ^ n3371 ^ 1'b0 ;
  assign n3375 = n1853 & ~n3374 ;
  assign n3376 = n3375 ^ n1695 ^ 1'b0 ;
  assign n3377 = n2223 ^ n1904 ^ 1'b0 ;
  assign n3378 = ~n1724 & n3377 ;
  assign n3379 = n277 & n2046 ;
  assign n3380 = n1873 & n3379 ;
  assign n3381 = n3380 ^ n3223 ^ 1'b0 ;
  assign n3382 = ~x149 & n2925 ;
  assign n3383 = n514 & n936 ;
  assign n3384 = ~n733 & n813 ;
  assign n3385 = x26 & n1665 ;
  assign n3386 = n3385 ^ n1287 ^ 1'b0 ;
  assign n3387 = n3386 ^ n1261 ^ 1'b0 ;
  assign n3388 = n455 | n3387 ;
  assign n3389 = n3388 ^ n2582 ^ 1'b0 ;
  assign n3390 = n1059 | n3389 ;
  assign n3391 = n3384 & ~n3390 ;
  assign n3392 = n2253 ^ n1970 ^ 1'b0 ;
  assign n3393 = n3392 ^ n2890 ^ 1'b0 ;
  assign n3394 = ~n755 & n931 ;
  assign n3395 = n1972 | n2093 ;
  assign n3396 = n909 | n3135 ;
  assign n3397 = ~n1564 & n3396 ;
  assign n3398 = n3395 & n3397 ;
  assign n3399 = n629 & ~n2557 ;
  assign n3400 = n3399 ^ n2376 ^ 1'b0 ;
  assign n3401 = x15 & ~n3400 ;
  assign n3402 = n2269 ^ x4 ^ 1'b0 ;
  assign n3403 = n2393 | n3402 ;
  assign n3404 = ( x221 & n1201 ) | ( x221 & ~n3403 ) | ( n1201 & ~n3403 ) ;
  assign n3405 = ( ~x168 & n3172 ) | ( ~x168 & n3404 ) | ( n3172 & n3404 ) ;
  assign n3406 = x20 & ~n1263 ;
  assign n3407 = n3098 ^ n1084 ^ 1'b0 ;
  assign n3408 = n3406 & n3407 ;
  assign n3409 = n2564 & n3408 ;
  assign n3410 = ~n1907 & n3409 ;
  assign n3414 = n314 & n1144 ;
  assign n3411 = x117 & n2421 ;
  assign n3412 = ~n1319 & n3411 ;
  assign n3413 = n3412 ^ n752 ^ 1'b0 ;
  assign n3415 = n3414 ^ n3413 ^ n283 ;
  assign n3416 = n700 | n762 ;
  assign n3417 = n909 | n3416 ;
  assign n3418 = ~n900 & n3417 ;
  assign n3419 = n3418 ^ n539 ^ 1'b0 ;
  assign n3420 = ~n1489 & n3419 ;
  assign n3421 = ( n1093 & n1215 ) | ( n1093 & n3420 ) | ( n1215 & n3420 ) ;
  assign n3422 = n2841 ^ n2230 ^ 1'b0 ;
  assign n3423 = ( ~n585 & n2452 ) | ( ~n585 & n2601 ) | ( n2452 & n2601 ) ;
  assign n3430 = n1369 | n1372 ;
  assign n3424 = n332 & n1627 ;
  assign n3425 = ( n1350 & n1961 ) | ( n1350 & n3424 ) | ( n1961 & n3424 ) ;
  assign n3426 = n2864 ^ n1355 ^ 1'b0 ;
  assign n3427 = x25 & n3426 ;
  assign n3428 = ~n3425 & n3427 ;
  assign n3429 = n1833 & n3428 ;
  assign n3431 = n3430 ^ n3429 ^ 1'b0 ;
  assign n3432 = n749 & ~n2921 ;
  assign n3433 = n3027 & n3432 ;
  assign n3436 = n1453 ^ n1298 ^ n1129 ;
  assign n3437 = n1703 ^ n522 ^ 1'b0 ;
  assign n3438 = n3436 & n3437 ;
  assign n3435 = ~n725 & n907 ;
  assign n3434 = n1374 ^ n326 ^ 1'b0 ;
  assign n3439 = n3438 ^ n3435 ^ n3434 ;
  assign n3440 = n2692 ^ x20 ^ 1'b0 ;
  assign n3441 = n1315 & n3440 ;
  assign n3442 = n2405 ^ n2372 ^ 1'b0 ;
  assign n3443 = n3441 & n3442 ;
  assign n3444 = x70 & n3161 ;
  assign n3445 = n3444 ^ n1411 ^ 1'b0 ;
  assign n3446 = x248 ^ x138 ^ 1'b0 ;
  assign n3447 = n3068 & n3446 ;
  assign n3449 = n1574 ^ n998 ^ x222 ;
  assign n3448 = n3103 ^ n2571 ^ 1'b0 ;
  assign n3450 = n3449 ^ n3448 ^ x247 ;
  assign n3451 = n3041 ^ n3035 ^ 1'b0 ;
  assign n3452 = n1058 | n1526 ;
  assign n3453 = n427 | n3452 ;
  assign n3454 = ( ~n1369 & n1618 ) | ( ~n1369 & n2228 ) | ( n1618 & n2228 ) ;
  assign n3455 = n3454 ^ n1403 ^ 1'b0 ;
  assign n3456 = ~n1458 & n3455 ;
  assign n3458 = x135 & n1722 ;
  assign n3459 = ~x206 & n3458 ;
  assign n3457 = n1166 & ~n1594 ;
  assign n3460 = n3459 ^ n3457 ^ 1'b0 ;
  assign n3461 = n3460 ^ x225 ^ 1'b0 ;
  assign n3462 = n3456 & n3461 ;
  assign n3463 = ~n428 & n2357 ;
  assign n3464 = n3463 ^ n3048 ^ 1'b0 ;
  assign n3465 = n3464 ^ n1062 ^ 1'b0 ;
  assign n3466 = n1558 ^ n1033 ^ 1'b0 ;
  assign n3467 = ( n1296 & n3296 ) | ( n1296 & n3466 ) | ( n3296 & n3466 ) ;
  assign n3470 = n1430 ^ n388 ^ 1'b0 ;
  assign n3471 = n3470 ^ n2981 ^ 1'b0 ;
  assign n3472 = ~n366 & n3471 ;
  assign n3468 = n1980 ^ n1780 ^ n463 ;
  assign n3469 = ( ~n1827 & n2957 ) | ( ~n1827 & n3468 ) | ( n2957 & n3468 ) ;
  assign n3473 = n3472 ^ n3469 ^ n1629 ;
  assign n3474 = n2363 ^ n2228 ^ 1'b0 ;
  assign n3475 = n3474 ^ n3002 ^ 1'b0 ;
  assign n3476 = ( n991 & n1380 ) | ( n991 & ~n3316 ) | ( n1380 & ~n3316 ) ;
  assign n3477 = n2823 ^ n1217 ^ 1'b0 ;
  assign n3478 = n3477 ^ n1203 ^ 1'b0 ;
  assign n3479 = x144 & n3478 ;
  assign n3480 = n2664 ^ n1520 ^ n332 ;
  assign n3481 = n1140 | n1394 ;
  assign n3482 = n535 | n3481 ;
  assign n3483 = n3482 ^ n2609 ^ 1'b0 ;
  assign n3484 = n3483 ^ n2580 ^ 1'b0 ;
  assign n3485 = n3480 & ~n3484 ;
  assign n3486 = n3485 ^ n2000 ^ n642 ;
  assign n3487 = x20 & n1037 ;
  assign n3488 = ~n1702 & n3487 ;
  assign n3489 = ~n345 & n3488 ;
  assign n3492 = n2575 | n3384 ;
  assign n3490 = ~x23 & x223 ;
  assign n3491 = n2492 | n3490 ;
  assign n3493 = n3492 ^ n3491 ^ 1'b0 ;
  assign n3494 = n524 ^ x59 ^ 1'b0 ;
  assign n3495 = ~n315 & n3494 ;
  assign n3496 = n3024 & n3495 ;
  assign n3497 = n3496 ^ n2759 ^ 1'b0 ;
  assign n3498 = n982 ^ n451 ^ 1'b0 ;
  assign n3503 = ~n800 & n1300 ;
  assign n3504 = ~n1295 & n3503 ;
  assign n3501 = x192 ^ x183 ^ 1'b0 ;
  assign n3502 = n3501 ^ n2124 ^ 1'b0 ;
  assign n3505 = n3504 ^ n3502 ^ n1686 ;
  assign n3500 = n894 & n2118 ;
  assign n3506 = n3505 ^ n3500 ^ 1'b0 ;
  assign n3499 = ( n886 & n1711 ) | ( n886 & n2346 ) | ( n1711 & n2346 ) ;
  assign n3507 = n3506 ^ n3499 ^ 1'b0 ;
  assign n3508 = n2654 & ~n3282 ;
  assign n3509 = n1088 | n2490 ;
  assign n3510 = n2431 ^ n1166 ^ 1'b0 ;
  assign n3511 = n1126 | n3510 ;
  assign n3512 = n972 | n1683 ;
  assign n3513 = n1209 | n3512 ;
  assign n3514 = n1695 | n3513 ;
  assign n3515 = n3514 ^ n1403 ^ 1'b0 ;
  assign n3516 = n1095 ^ n392 ^ 1'b0 ;
  assign n3517 = n3516 ^ n2965 ^ 1'b0 ;
  assign n3518 = n527 & n1788 ;
  assign n3519 = n3007 ^ n1011 ^ 1'b0 ;
  assign n3520 = n3518 & ~n3519 ;
  assign n3521 = ~n3517 & n3520 ;
  assign n3522 = x228 & n1903 ;
  assign n3523 = ~x191 & n3522 ;
  assign n3524 = n2134 & ~n3523 ;
  assign n3525 = ~n2720 & n2890 ;
  assign n3526 = ( ~n1106 & n2925 ) | ( ~n1106 & n3525 ) | ( n2925 & n3525 ) ;
  assign n3527 = x11 & n299 ;
  assign n3528 = ~x111 & n3527 ;
  assign n3529 = x247 & ~n3528 ;
  assign n3530 = n3529 ^ n1295 ^ 1'b0 ;
  assign n3531 = n3530 ^ n1541 ^ 1'b0 ;
  assign n3533 = n3166 ^ n2710 ^ n2113 ;
  assign n3532 = n2654 & n3060 ;
  assign n3534 = n3533 ^ n3532 ^ 1'b0 ;
  assign n3535 = ~n2495 & n2913 ;
  assign n3536 = n3534 & n3535 ;
  assign n3537 = n3531 & ~n3536 ;
  assign n3538 = n600 & n3537 ;
  assign n3539 = n3222 ^ n1380 ^ 1'b0 ;
  assign n3540 = n1557 & ~n3539 ;
  assign n3541 = n1658 | n1712 ;
  assign n3542 = n3541 ^ x15 ^ 1'b0 ;
  assign n3543 = n2075 | n3542 ;
  assign n3544 = n2719 | n3543 ;
  assign n3545 = n3544 ^ x11 ^ 1'b0 ;
  assign n3546 = ( ~x71 & n805 ) | ( ~x71 & n3545 ) | ( n805 & n3545 ) ;
  assign n3547 = x220 | n1134 ;
  assign n3548 = x112 & ~n2555 ;
  assign n3549 = n3548 ^ n2558 ^ 1'b0 ;
  assign n3550 = n2546 & n3549 ;
  assign n3551 = n2834 ^ n1194 ^ 1'b0 ;
  assign n3552 = n2389 ^ n1296 ^ 1'b0 ;
  assign n3553 = n2517 ^ n2249 ^ 1'b0 ;
  assign n3554 = ~n1475 & n3553 ;
  assign n3555 = n301 & n3406 ;
  assign n3556 = x17 & n3555 ;
  assign n3557 = n3556 ^ n1027 ^ 1'b0 ;
  assign n3558 = n3557 ^ x171 ^ 1'b0 ;
  assign n3559 = ~n886 & n2586 ;
  assign n3560 = ~n1610 & n3559 ;
  assign n3561 = n668 & n866 ;
  assign n3562 = ~n489 & n3561 ;
  assign n3563 = n2486 | n3562 ;
  assign n3564 = n3560 & ~n3563 ;
  assign n3565 = x169 & ~n3564 ;
  assign n3566 = ~n2888 & n3565 ;
  assign n3571 = x203 & n950 ;
  assign n3572 = n3571 ^ n519 ^ 1'b0 ;
  assign n3573 = n2224 & n3572 ;
  assign n3567 = n624 & n2068 ;
  assign n3568 = n3567 ^ n1252 ^ 1'b0 ;
  assign n3569 = n2860 | n3568 ;
  assign n3570 = n3569 ^ n548 ^ 1'b0 ;
  assign n3574 = n3573 ^ n3570 ^ 1'b0 ;
  assign n3575 = n1881 & n3574 ;
  assign n3576 = n2949 & n3575 ;
  assign n3577 = n1203 & n1358 ;
  assign n3578 = n3577 ^ n1803 ^ 1'b0 ;
  assign n3579 = n1462 & ~n3578 ;
  assign n3580 = n3579 ^ n369 ^ 1'b0 ;
  assign n3581 = ~n1370 & n3580 ;
  assign n3584 = n2345 ^ n2320 ^ 1'b0 ;
  assign n3582 = n1795 & n2047 ;
  assign n3583 = ~n2540 & n3582 ;
  assign n3585 = n3584 ^ n3583 ^ 1'b0 ;
  assign n3586 = n3581 & n3585 ;
  assign n3587 = n2448 ^ n1919 ^ 1'b0 ;
  assign n3588 = n883 ^ x226 ^ 1'b0 ;
  assign n3595 = n2378 ^ n2292 ^ 1'b0 ;
  assign n3589 = n2991 ^ x55 ^ 1'b0 ;
  assign n3590 = x135 & n3589 ;
  assign n3591 = x167 & n3590 ;
  assign n3592 = n1488 & n3591 ;
  assign n3593 = n3592 ^ n2952 ^ 1'b0 ;
  assign n3594 = x76 & n3593 ;
  assign n3596 = n3595 ^ n3594 ^ 1'b0 ;
  assign n3597 = n1233 ^ x5 ^ 1'b0 ;
  assign n3598 = n3597 ^ n1746 ^ n1724 ;
  assign n3599 = ( ~n1472 & n2523 ) | ( ~n1472 & n3598 ) | ( n2523 & n3598 ) ;
  assign n3600 = ~n978 & n3599 ;
  assign n3601 = n2548 ^ n2516 ^ n650 ;
  assign n3602 = ~n3343 & n3601 ;
  assign n3603 = n3602 ^ n2827 ^ 1'b0 ;
  assign n3604 = x54 & ~n3603 ;
  assign n3605 = n3604 ^ n533 ^ 1'b0 ;
  assign n3606 = n3600 & n3605 ;
  assign n3607 = ~n2409 & n2804 ;
  assign n3608 = n3607 ^ n2250 ^ 1'b0 ;
  assign n3609 = n1548 | n3608 ;
  assign n3610 = n3609 ^ x104 ^ 1'b0 ;
  assign n3611 = n2006 ^ n1930 ^ 1'b0 ;
  assign n3616 = n392 & n1273 ;
  assign n3617 = n3616 ^ n1404 ^ 1'b0 ;
  assign n3614 = n814 ^ x52 ^ 1'b0 ;
  assign n3615 = n1206 & ~n3614 ;
  assign n3612 = n3490 ^ n2988 ^ 1'b0 ;
  assign n3613 = n1701 | n3612 ;
  assign n3618 = n3617 ^ n3615 ^ n3613 ;
  assign n3619 = n1023 | n2914 ;
  assign n3620 = n1000 & ~n3619 ;
  assign n3621 = n3090 ^ n2412 ^ 1'b0 ;
  assign n3622 = n3620 | n3621 ;
  assign n3623 = n629 & n2264 ;
  assign n3624 = n3623 ^ n380 ^ 1'b0 ;
  assign n3625 = ~n1416 & n3624 ;
  assign n3626 = ~n326 & n2955 ;
  assign n3627 = ~n3625 & n3626 ;
  assign n3628 = n1813 ^ n425 ^ 1'b0 ;
  assign n3629 = n2611 & ~n3628 ;
  assign n3630 = n795 & n3629 ;
  assign n3631 = n347 & n1374 ;
  assign n3632 = n1882 & n3631 ;
  assign n3633 = n3632 ^ n2303 ^ 1'b0 ;
  assign n3634 = ~n2669 & n3633 ;
  assign n3635 = n3630 & n3634 ;
  assign n3640 = ~x128 & n836 ;
  assign n3641 = ( x94 & ~n874 ) | ( x94 & n3640 ) | ( ~n874 & n3640 ) ;
  assign n3642 = ( n634 & n1416 ) | ( n634 & n3641 ) | ( n1416 & n3641 ) ;
  assign n3637 = n608 & ~n2040 ;
  assign n3638 = n3637 ^ n1258 ^ 1'b0 ;
  assign n3636 = ~n569 & n2517 ;
  assign n3639 = n3638 ^ n3636 ^ 1'b0 ;
  assign n3643 = n3642 ^ n3639 ^ 1'b0 ;
  assign n3644 = n755 | n1259 ;
  assign n3645 = n3644 ^ n2765 ^ 1'b0 ;
  assign n3646 = n1344 ^ n884 ^ n331 ;
  assign n3647 = n3646 ^ n2361 ^ 1'b0 ;
  assign n3648 = n3647 ^ n1935 ^ 1'b0 ;
  assign n3649 = n1103 ^ n488 ^ 1'b0 ;
  assign n3650 = n2523 & ~n3649 ;
  assign n3651 = ( n903 & n1085 ) | ( n903 & ~n3650 ) | ( n1085 & ~n3650 ) ;
  assign n3652 = ( x175 & ~n2782 ) | ( x175 & n3055 ) | ( ~n2782 & n3055 ) ;
  assign n3653 = n3045 ^ n1368 ^ n1234 ;
  assign n3654 = n1785 ^ n685 ^ n432 ;
  assign n3656 = n344 & n1349 ;
  assign n3657 = ~n3579 & n3656 ;
  assign n3658 = n3657 ^ n1247 ^ n367 ;
  assign n3659 = n2125 & n3658 ;
  assign n3655 = n1386 & ~n2457 ;
  assign n3660 = n3659 ^ n3655 ^ 1'b0 ;
  assign n3661 = n1296 & ~n1319 ;
  assign n3662 = n1419 & n3661 ;
  assign n3663 = n2058 ^ n1958 ^ 1'b0 ;
  assign n3664 = ~n3662 & n3663 ;
  assign n3665 = ~n1066 & n2715 ;
  assign n3666 = ~n3203 & n3665 ;
  assign n3667 = n2836 ^ n465 ^ 1'b0 ;
  assign n3670 = n1928 | n2219 ;
  assign n3671 = ( n766 & ~n800 ) | ( n766 & n3670 ) | ( ~n800 & n3670 ) ;
  assign n3668 = ( ~n756 & n948 ) | ( ~n756 & n1353 ) | ( n948 & n1353 ) ;
  assign n3669 = n3267 & ~n3668 ;
  assign n3672 = n3671 ^ n3669 ^ 1'b0 ;
  assign n3673 = n3111 ^ n1138 ^ 1'b0 ;
  assign n3674 = n558 & n660 ;
  assign n3675 = ~x108 & n3674 ;
  assign n3676 = n1177 | n3675 ;
  assign n3677 = n672 & n1081 ;
  assign n3678 = ~n2264 & n3677 ;
  assign n3679 = n1506 & ~n3678 ;
  assign n3680 = n2748 & n3679 ;
  assign n3681 = n446 ^ n404 ^ x17 ;
  assign n3682 = n3681 ^ n1145 ^ 1'b0 ;
  assign n3683 = ~n1369 & n3682 ;
  assign n3684 = n3126 ^ x30 ^ 1'b0 ;
  assign n3685 = ~n3683 & n3684 ;
  assign n3686 = n2053 & n3144 ;
  assign n3687 = n939 | n1934 ;
  assign n3688 = x17 & n1210 ;
  assign n3689 = n3687 | n3688 ;
  assign n3690 = n1478 ^ n1404 ^ 1'b0 ;
  assign n3691 = n1001 & n2065 ;
  assign n3692 = n3402 ^ n1960 ^ 1'b0 ;
  assign n3693 = n3692 ^ n2746 ^ 1'b0 ;
  assign n3694 = n2345 & ~n3693 ;
  assign n3695 = n1892 ^ n597 ^ 1'b0 ;
  assign n3696 = n3399 & n3695 ;
  assign n3697 = n3696 ^ n749 ^ 1'b0 ;
  assign n3698 = ( ~n617 & n1212 ) | ( ~n617 & n2759 ) | ( n1212 & n2759 ) ;
  assign n3699 = n1009 & n3698 ;
  assign n3700 = n3699 ^ n2549 ^ 1'b0 ;
  assign n3701 = n2752 ^ n1525 ^ n1142 ;
  assign n3705 = x180 | n1680 ;
  assign n3703 = n1711 ^ n968 ^ 1'b0 ;
  assign n3704 = n634 & ~n3703 ;
  assign n3702 = ~n308 & n2214 ;
  assign n3706 = n3705 ^ n3704 ^ n3702 ;
  assign n3707 = n366 | n380 ;
  assign n3708 = n3707 ^ n1339 ^ n681 ;
  assign n3709 = n311 | n718 ;
  assign n3710 = n2203 & ~n3709 ;
  assign n3711 = ( n581 & n2468 ) | ( n581 & ~n3710 ) | ( n2468 & ~n3710 ) ;
  assign n3712 = ~n1571 & n3009 ;
  assign n3713 = n1819 | n3712 ;
  assign n3714 = n3711 & ~n3713 ;
  assign n3715 = n2127 ^ n1922 ^ 1'b0 ;
  assign n3716 = n2227 & ~n3715 ;
  assign n3717 = ~n298 & n1090 ;
  assign n3718 = n3717 ^ n2181 ^ 1'b0 ;
  assign n3719 = n3718 ^ n1289 ^ 1'b0 ;
  assign n3720 = n3716 & ~n3719 ;
  assign n3721 = n546 & ~n1850 ;
  assign n3722 = x180 & n2855 ;
  assign n3723 = n3722 ^ n1557 ^ 1'b0 ;
  assign n3724 = x196 & n608 ;
  assign n3725 = n3724 ^ n1489 ^ 1'b0 ;
  assign n3726 = n2893 ^ n1666 ^ 1'b0 ;
  assign n3727 = n2320 ^ n861 ^ 1'b0 ;
  assign n3728 = n3727 ^ n385 ^ 1'b0 ;
  assign n3729 = ~n3726 & n3728 ;
  assign n3730 = ~n3725 & n3729 ;
  assign n3731 = n3723 & n3730 ;
  assign n3732 = n3731 ^ n3216 ^ x26 ;
  assign n3733 = n3687 ^ n814 ^ 1'b0 ;
  assign n3734 = ( n2361 & ~n2661 ) | ( n2361 & n3733 ) | ( ~n2661 & n3733 ) ;
  assign n3743 = n3615 ^ n2483 ^ n562 ;
  assign n3736 = ~n993 & n1192 ;
  assign n3737 = n3736 ^ n898 ^ 1'b0 ;
  assign n3738 = n3737 ^ n460 ^ 1'b0 ;
  assign n3739 = n3738 ^ n904 ^ 1'b0 ;
  assign n3740 = n1912 | n3739 ;
  assign n3741 = ~n1277 & n3740 ;
  assign n3735 = n2065 | n2516 ;
  assign n3742 = n3741 ^ n3735 ^ 1'b0 ;
  assign n3744 = n3743 ^ n3742 ^ n2569 ;
  assign n3745 = n1164 ^ n1113 ^ 1'b0 ;
  assign n3746 = n3154 & n3745 ;
  assign n3747 = n1836 & ~n1912 ;
  assign n3748 = n597 & ~n1389 ;
  assign n3749 = ~n3747 & n3748 ;
  assign n3750 = n304 | n1501 ;
  assign n3751 = n1486 & n1693 ;
  assign n3752 = x192 & n3751 ;
  assign n3753 = x216 & ~n3334 ;
  assign n3754 = n3752 & n3753 ;
  assign n3755 = ( n575 & n2118 ) | ( n575 & ~n3754 ) | ( n2118 & ~n3754 ) ;
  assign n3756 = n3430 ^ n2573 ^ 1'b0 ;
  assign n3757 = ~n2332 & n3756 ;
  assign n3758 = n1525 & ~n3757 ;
  assign n3759 = n1991 & n3758 ;
  assign n3760 = n1075 & n2794 ;
  assign n3761 = n1450 & n3760 ;
  assign n3762 = n3545 ^ n1059 ^ 1'b0 ;
  assign n3763 = n3082 & ~n3762 ;
  assign n3764 = ( n972 & n1527 ) | ( n972 & ~n3011 ) | ( n1527 & ~n3011 ) ;
  assign n3765 = ( ~n2160 & n2870 ) | ( ~n2160 & n3764 ) | ( n2870 & n3764 ) ;
  assign n3766 = n3490 ^ n663 ^ 1'b0 ;
  assign n3767 = ~n3434 & n3766 ;
  assign n3768 = n2959 ^ n2142 ^ 1'b0 ;
  assign n3769 = n2988 & n3768 ;
  assign n3770 = ( n365 & ~n605 ) | ( n365 & n2172 ) | ( ~n605 & n2172 ) ;
  assign n3771 = n2619 ^ n983 ^ 1'b0 ;
  assign n3772 = ~n3770 & n3771 ;
  assign n3773 = n2649 ^ n2272 ^ 1'b0 ;
  assign n3774 = n329 | n1836 ;
  assign n3775 = n3773 | n3774 ;
  assign n3776 = n2534 & n3775 ;
  assign n3777 = ( n737 & n756 ) | ( n737 & ~n2294 ) | ( n756 & ~n2294 ) ;
  assign n3778 = n3777 ^ n737 ^ 1'b0 ;
  assign n3779 = ( ~n2560 & n3485 ) | ( ~n2560 & n3778 ) | ( n3485 & n3778 ) ;
  assign n3780 = n3776 & ~n3779 ;
  assign n3781 = n3780 ^ n3216 ^ 1'b0 ;
  assign n3782 = ( n335 & n2299 ) | ( n335 & n3781 ) | ( n2299 & n3781 ) ;
  assign n3783 = n2696 ^ n2052 ^ n1706 ;
  assign n3784 = n1716 & n3783 ;
  assign n3785 = ~n546 & n3784 ;
  assign n3786 = n3168 ^ x189 ^ 1'b0 ;
  assign n3787 = n2181 ^ n1881 ^ 1'b0 ;
  assign n3788 = n3787 ^ n1214 ^ 1'b0 ;
  assign n3789 = n3013 | n3343 ;
  assign n3790 = n749 | n3789 ;
  assign n3791 = n3790 ^ n1140 ^ 1'b0 ;
  assign n3792 = n1474 ^ x7 ^ 1'b0 ;
  assign n3793 = n3791 & ~n3792 ;
  assign n3794 = n1055 | n1612 ;
  assign n3795 = n3794 ^ n2024 ^ 1'b0 ;
  assign n3796 = n1038 | n3795 ;
  assign n3797 = n590 & n2648 ;
  assign n3798 = n3797 ^ n2437 ^ 1'b0 ;
  assign n3799 = n3668 ^ n3261 ^ 1'b0 ;
  assign n3800 = ~n1247 & n3799 ;
  assign n3801 = n994 ^ n780 ^ x234 ;
  assign n3802 = n3039 & n3128 ;
  assign n3803 = n3802 ^ n787 ^ 1'b0 ;
  assign n3804 = ( n3371 & n3801 ) | ( n3371 & ~n3803 ) | ( n3801 & ~n3803 ) ;
  assign n3805 = n259 & ~n3646 ;
  assign n3806 = n3804 & n3805 ;
  assign n3813 = n1081 & ~n2647 ;
  assign n3814 = ~n3477 & n3813 ;
  assign n3811 = n2296 ^ n1147 ^ 1'b0 ;
  assign n3807 = ~n3307 & n3495 ;
  assign n3808 = ~x83 & n3807 ;
  assign n3809 = n3533 ^ n728 ^ 1'b0 ;
  assign n3810 = ~n3808 & n3809 ;
  assign n3812 = n3811 ^ n3810 ^ 1'b0 ;
  assign n3815 = n3814 ^ n3812 ^ n349 ;
  assign n3816 = n3317 ^ n1555 ^ 1'b0 ;
  assign n3817 = ~n645 & n3816 ;
  assign n3818 = ~n269 & n1782 ;
  assign n3819 = n3818 ^ n3245 ^ 1'b0 ;
  assign n3820 = x55 & ~n1394 ;
  assign n3821 = ~n2250 & n3820 ;
  assign n3822 = ( n1217 & n2972 ) | ( n1217 & n3821 ) | ( n2972 & n3821 ) ;
  assign n3826 = n854 ^ x15 ^ 1'b0 ;
  assign n3823 = n289 & ~n593 ;
  assign n3824 = n3823 ^ n555 ^ 1'b0 ;
  assign n3825 = ( ~n1085 & n3676 ) | ( ~n1085 & n3824 ) | ( n3676 & n3824 ) ;
  assign n3827 = n3826 ^ n3825 ^ 1'b0 ;
  assign n3828 = n1618 ^ n1491 ^ 1'b0 ;
  assign n3829 = ~n793 & n3828 ;
  assign n3830 = ( n880 & n2587 ) | ( n880 & n3829 ) | ( n2587 & n3829 ) ;
  assign n3831 = n3830 ^ n3126 ^ n322 ;
  assign n3832 = n2718 ^ n1194 ^ 1'b0 ;
  assign n3833 = n3832 ^ n2893 ^ 1'b0 ;
  assign n3834 = n1236 ^ n549 ^ n363 ;
  assign n3835 = n3834 ^ n2497 ^ n1902 ;
  assign n3836 = ~n669 & n3835 ;
  assign n3837 = ~n2466 & n3836 ;
  assign n3838 = n2737 ^ x93 ^ 1'b0 ;
  assign n3839 = x125 & n3838 ;
  assign n3840 = n1720 ^ n1387 ^ 1'b0 ;
  assign n3841 = n3839 & n3840 ;
  assign n3842 = n1697 | n2171 ;
  assign n3843 = n1317 & n3842 ;
  assign n3844 = n3843 ^ n3015 ^ 1'b0 ;
  assign n3845 = n2667 ^ n2497 ^ x25 ;
  assign n3846 = n3845 ^ n3801 ^ 1'b0 ;
  assign n3847 = n2995 | n3846 ;
  assign n3848 = n3265 ^ n1288 ^ x7 ;
  assign n3849 = x210 & ~n863 ;
  assign n3850 = n3849 ^ x200 ^ 1'b0 ;
  assign n3851 = n924 | n3253 ;
  assign n3852 = n3850 & ~n3851 ;
  assign n3853 = n2178 & n3852 ;
  assign n3854 = n2382 ^ n1934 ^ n552 ;
  assign n3857 = ~x77 & n3336 ;
  assign n3855 = n1569 ^ n446 ^ 1'b0 ;
  assign n3856 = n269 & n3855 ;
  assign n3858 = n3857 ^ n3856 ^ 1'b0 ;
  assign n3859 = n3854 & ~n3858 ;
  assign n3860 = n3145 ^ n2523 ^ 1'b0 ;
  assign n3861 = n2426 | n3860 ;
  assign n3862 = n3861 ^ n557 ^ 1'b0 ;
  assign n3863 = n3112 & ~n3862 ;
  assign n3864 = n3863 ^ n2495 ^ 1'b0 ;
  assign n3868 = n806 ^ n776 ^ 1'b0 ;
  assign n3865 = ~n579 & n1209 ;
  assign n3866 = n1173 & n3865 ;
  assign n3867 = n1030 & ~n3866 ;
  assign n3869 = n3868 ^ n3867 ^ 1'b0 ;
  assign n3870 = n2924 & n3869 ;
  assign n3871 = n3870 ^ n1067 ^ 1'b0 ;
  assign n3872 = n3794 ^ n2050 ^ 1'b0 ;
  assign n3873 = n2601 | n3872 ;
  assign n3874 = n3873 ^ n2359 ^ 1'b0 ;
  assign n3875 = n2452 ^ x220 ^ 1'b0 ;
  assign n3876 = n829 & n2479 ;
  assign n3877 = ~n1731 & n3876 ;
  assign n3878 = n3877 ^ n2057 ^ 1'b0 ;
  assign n3879 = ( n1650 & n3875 ) | ( n1650 & n3878 ) | ( n3875 & n3878 ) ;
  assign n3880 = n1145 & n2644 ;
  assign n3881 = n789 & n1504 ;
  assign n3882 = n3881 ^ n3366 ^ n674 ;
  assign n3883 = n911 & ~n2617 ;
  assign n3884 = n3883 ^ n1236 ^ 1'b0 ;
  assign n3885 = n982 & n2071 ;
  assign n3886 = ~n1358 & n1587 ;
  assign n3887 = n3886 ^ n852 ^ 1'b0 ;
  assign n3888 = n2636 ^ n833 ^ 1'b0 ;
  assign n3889 = n3888 ^ n3499 ^ 1'b0 ;
  assign n3890 = x169 & n337 ;
  assign n3891 = ( ~n1001 & n3704 ) | ( ~n1001 & n3890 ) | ( n3704 & n3890 ) ;
  assign n3892 = n2756 & ~n3891 ;
  assign n3893 = n3892 ^ n3336 ^ 1'b0 ;
  assign n3894 = n2151 ^ x15 ^ 1'b0 ;
  assign n3897 = ~x13 & n1269 ;
  assign n3898 = n3897 ^ n1168 ^ 1'b0 ;
  assign n3895 = ~n2208 & n2935 ;
  assign n3896 = n2389 | n3895 ;
  assign n3899 = n3898 ^ n3896 ^ 1'b0 ;
  assign n3900 = ~n1232 & n2970 ;
  assign n3901 = ~n2519 & n3900 ;
  assign n3902 = x166 & ~n605 ;
  assign n3903 = n3902 ^ n1181 ^ 1'b0 ;
  assign n3904 = n1362 ^ n591 ^ n429 ;
  assign n3905 = n3903 & ~n3904 ;
  assign n3906 = n2897 ^ n1476 ^ 1'b0 ;
  assign n3907 = n3905 & n3906 ;
  assign n3908 = n1362 & ~n2418 ;
  assign n3909 = n1258 ^ n648 ^ n502 ;
  assign n3910 = n3909 ^ n1525 ^ n1044 ;
  assign n3911 = n1735 ^ n1175 ^ 1'b0 ;
  assign n3912 = n3911 ^ n2939 ^ 1'b0 ;
  assign n3913 = ( n3908 & n3910 ) | ( n3908 & ~n3912 ) | ( n3910 & ~n3912 ) ;
  assign n3914 = n3737 & ~n3913 ;
  assign n3915 = ~n3907 & n3914 ;
  assign n3916 = ~n1372 & n2366 ;
  assign n3917 = ~x203 & n3916 ;
  assign n3918 = n3504 ^ n2862 ^ n2216 ;
  assign n3919 = ( ~n1995 & n2955 ) | ( ~n1995 & n3918 ) | ( n2955 & n3918 ) ;
  assign n3920 = n3919 ^ n539 ^ 1'b0 ;
  assign n3921 = n3917 & n3920 ;
  assign n3922 = n2057 ^ n1960 ^ 1'b0 ;
  assign n3923 = n729 ^ n332 ^ 1'b0 ;
  assign n3924 = n3922 | n3923 ;
  assign n3928 = n404 & n1466 ;
  assign n3929 = ~n383 & n3928 ;
  assign n3934 = ~n498 & n911 ;
  assign n3935 = ~x237 & n3934 ;
  assign n3931 = n1090 & ~n1532 ;
  assign n3932 = ~n1886 & n3931 ;
  assign n3930 = ~n1086 & n1506 ;
  assign n3933 = n3932 ^ n3930 ^ 1'b0 ;
  assign n3936 = n3935 ^ n3933 ^ 1'b0 ;
  assign n3937 = n3929 | n3936 ;
  assign n3926 = n706 | n909 ;
  assign n3925 = x188 & ~n3511 ;
  assign n3927 = n3926 ^ n3925 ^ 1'b0 ;
  assign n3938 = n3937 ^ n3927 ^ n2329 ;
  assign n3939 = n1430 | n2762 ;
  assign n3940 = n3939 ^ n3422 ^ n3413 ;
  assign n3941 = n2022 ^ x42 ^ 1'b0 ;
  assign n3942 = n2499 & n3941 ;
  assign n3943 = ( n2274 & n2372 ) | ( n2274 & n3942 ) | ( n2372 & n3942 ) ;
  assign n3944 = n3943 ^ n913 ^ 1'b0 ;
  assign n3945 = n1890 | n2124 ;
  assign n3946 = n3944 & ~n3945 ;
  assign n3947 = x169 & ~n3443 ;
  assign n3948 = n2818 ^ n2778 ^ 1'b0 ;
  assign n3949 = n762 | n3948 ;
  assign n3950 = x57 & n635 ;
  assign n3951 = n3949 & n3950 ;
  assign n3952 = n1947 ^ n553 ^ 1'b0 ;
  assign n3953 = n269 & ~n3952 ;
  assign n3954 = n3720 ^ n3492 ^ 1'b0 ;
  assign n3955 = n3954 ^ n1451 ^ 1'b0 ;
  assign n3956 = ~n579 & n2466 ;
  assign n3957 = ~n1984 & n3956 ;
  assign n3958 = n3957 ^ n1842 ^ x40 ;
  assign n3959 = n3099 ^ n2694 ^ 1'b0 ;
  assign n3960 = n3959 ^ n1368 ^ 1'b0 ;
  assign n3961 = n2335 ^ n1932 ^ n1179 ;
  assign n3962 = ~n2457 & n3961 ;
  assign n3963 = n492 | n2697 ;
  assign n3964 = n2091 & ~n3963 ;
  assign n3965 = ~x67 & n3964 ;
  assign n3966 = n3307 ^ n1733 ^ 1'b0 ;
  assign n3967 = n3966 ^ n3912 ^ 1'b0 ;
  assign n3968 = n2521 & ~n3967 ;
  assign n3969 = n1930 ^ n495 ^ 1'b0 ;
  assign n3970 = n1158 & ~n3969 ;
  assign n3971 = ~n718 & n2804 ;
  assign n3972 = n2387 & n3971 ;
  assign n3973 = n3970 & n3972 ;
  assign n3974 = x92 & ~n3770 ;
  assign n3975 = ~n472 & n3974 ;
  assign n3978 = x15 & ~x242 ;
  assign n3979 = n731 & n3978 ;
  assign n3976 = ( ~n307 & n909 ) | ( ~n307 & n2574 ) | ( n909 & n2574 ) ;
  assign n3977 = n2490 & n3976 ;
  assign n3980 = n3979 ^ n3977 ^ 1'b0 ;
  assign n3981 = ~n2093 & n3980 ;
  assign n3982 = x87 ^ x16 ^ 1'b0 ;
  assign n3983 = n3982 ^ n3749 ^ 1'b0 ;
  assign n3984 = n1590 | n2870 ;
  assign n3985 = n3984 ^ n592 ^ 1'b0 ;
  assign n3986 = ~n884 & n3691 ;
  assign n3987 = n1992 ^ n1115 ^ 1'b0 ;
  assign n3988 = n3010 & ~n3987 ;
  assign n3991 = x216 & ~n692 ;
  assign n3992 = n3991 ^ n2953 ^ 1'b0 ;
  assign n3989 = n302 & n1850 ;
  assign n3990 = ~n1979 & n3989 ;
  assign n3993 = n3992 ^ n3990 ^ 1'b0 ;
  assign n3994 = n3988 & ~n3993 ;
  assign n3995 = n3994 ^ n2895 ^ 1'b0 ;
  assign n3996 = n1885 | n3995 ;
  assign n3997 = n3996 ^ n1233 ^ 1'b0 ;
  assign n3998 = ( x105 & n659 ) | ( x105 & n1139 ) | ( n659 & n1139 ) ;
  assign n3999 = ~n3543 & n3998 ;
  assign n4000 = n3999 ^ n314 ^ 1'b0 ;
  assign n4001 = n2473 & n2839 ;
  assign n4002 = x65 & ~n1589 ;
  assign n4003 = n3095 ^ n886 ^ 1'b0 ;
  assign n4004 = n4002 & ~n4003 ;
  assign n4005 = ( x173 & n972 ) | ( x173 & n2823 ) | ( n972 & n2823 ) ;
  assign n4006 = n4005 ^ n3439 ^ 1'b0 ;
  assign n4007 = n3909 & ~n4006 ;
  assign n4008 = ~n1241 & n2744 ;
  assign n4009 = n1480 & n4008 ;
  assign n4017 = n312 ^ x43 ^ 1'b0 ;
  assign n4018 = n1541 | n4017 ;
  assign n4014 = n835 ^ n372 ^ 1'b0 ;
  assign n4015 = n2207 | n4014 ;
  assign n4010 = n2543 ^ n1354 ^ n265 ;
  assign n4011 = n1234 & n4010 ;
  assign n4012 = n4011 ^ n1685 ^ 1'b0 ;
  assign n4013 = ~n3232 & n4012 ;
  assign n4016 = n4015 ^ n4013 ^ 1'b0 ;
  assign n4019 = n4018 ^ n4016 ^ n1683 ;
  assign n4020 = n4009 & ~n4019 ;
  assign n4023 = n3530 ^ n3254 ^ 1'b0 ;
  assign n4021 = ( ~x143 & n905 ) | ( ~x143 & n2208 ) | ( n905 & n2208 ) ;
  assign n4022 = n2680 | n4021 ;
  assign n4024 = n4023 ^ n4022 ^ 1'b0 ;
  assign n4025 = ~n1346 & n2686 ;
  assign n4026 = n2158 & n4025 ;
  assign n4027 = n2009 | n3365 ;
  assign n4028 = n4026 | n4027 ;
  assign n4029 = n4024 & ~n4028 ;
  assign n4031 = x79 & n1237 ;
  assign n4032 = n1612 & n4031 ;
  assign n4033 = n2253 & n4032 ;
  assign n4034 = ( ~n329 & n2212 ) | ( ~n329 & n4033 ) | ( n2212 & n4033 ) ;
  assign n4030 = n3917 ^ x185 ^ 1'b0 ;
  assign n4035 = n4034 ^ n4030 ^ n665 ;
  assign n4036 = n2443 ^ n560 ^ 1'b0 ;
  assign n4037 = ~n1192 & n4036 ;
  assign n4038 = ~n1070 & n2969 ;
  assign n4039 = n1760 & ~n3817 ;
  assign n4041 = n764 ^ x125 ^ 1'b0 ;
  assign n4042 = n1906 & ~n4041 ;
  assign n4043 = ( ~n1491 & n1733 ) | ( ~n1491 & n4042 ) | ( n1733 & n4042 ) ;
  assign n4044 = n1351 | n4043 ;
  assign n4045 = n4044 ^ x246 ^ 1'b0 ;
  assign n4040 = ~n1382 & n2428 ;
  assign n4046 = n4045 ^ n4040 ^ 1'b0 ;
  assign n4047 = n3917 ^ n1145 ^ 1'b0 ;
  assign n4048 = n4047 ^ n2547 ^ 1'b0 ;
  assign n4053 = x188 & x227 ;
  assign n4054 = n4053 ^ n1897 ^ 1'b0 ;
  assign n4049 = x72 & ~n449 ;
  assign n4050 = ( n653 & n1767 ) | ( n653 & ~n4049 ) | ( n1767 & ~n4049 ) ;
  assign n4051 = n3239 & n4050 ;
  assign n4052 = n3334 & n4051 ;
  assign n4055 = n4054 ^ n4052 ^ 1'b0 ;
  assign n4056 = n3336 & ~n3472 ;
  assign n4057 = ~n950 & n3517 ;
  assign n4058 = n3769 | n4057 ;
  assign n4059 = n4058 ^ n2654 ^ 1'b0 ;
  assign n4060 = n1716 ^ n438 ^ x247 ;
  assign n4061 = n4060 ^ n3721 ^ 1'b0 ;
  assign n4062 = n3108 & n4061 ;
  assign n4063 = n3336 ^ n2855 ^ 1'b0 ;
  assign n4064 = n1624 ^ n612 ^ x218 ;
  assign n4065 = n513 & ~n1865 ;
  assign n4066 = x157 | n1330 ;
  assign n4067 = n4065 & ~n4066 ;
  assign n4068 = n4064 & n4067 ;
  assign n4069 = n1458 ^ n392 ^ 1'b0 ;
  assign n4070 = n2144 | n4069 ;
  assign n4071 = ~n1306 & n2394 ;
  assign n4072 = ~n1279 & n4071 ;
  assign n4073 = ( n671 & n875 ) | ( n671 & n4072 ) | ( n875 & n4072 ) ;
  assign n4074 = n3924 | n4073 ;
  assign n4075 = n1886 & ~n4074 ;
  assign n4076 = n4070 & n4075 ;
  assign n4077 = n626 ^ n585 ^ 1'b0 ;
  assign n4078 = n3705 ^ n1941 ^ n764 ;
  assign n4079 = n4078 ^ n2271 ^ 1'b0 ;
  assign n4080 = n1239 & ~n4079 ;
  assign n4081 = n1275 & n4080 ;
  assign n4082 = n909 & n4081 ;
  assign n4083 = n4082 ^ x19 ^ 1'b0 ;
  assign n4084 = n4083 ^ x118 ^ 1'b0 ;
  assign n4085 = n2352 & ~n4084 ;
  assign n4086 = ~n4077 & n4085 ;
  assign n4087 = x247 & ~n3018 ;
  assign n4088 = n2005 ^ n1490 ^ 1'b0 ;
  assign n4089 = n3725 | n4088 ;
  assign n4090 = n1814 & ~n3692 ;
  assign n4091 = n4089 & n4090 ;
  assign n4092 = n3189 | n4091 ;
  assign n4093 = n1564 & ~n4092 ;
  assign n4094 = ~n395 & n2959 ;
  assign n4095 = ~n982 & n4094 ;
  assign n4096 = n1527 & ~n3275 ;
  assign n4097 = n4096 ^ n3985 ^ 1'b0 ;
  assign n4098 = ~n800 & n4097 ;
  assign n4099 = ~n344 & n4098 ;
  assign n4100 = n1164 ^ x23 ^ 1'b0 ;
  assign n4101 = n455 & ~n2721 ;
  assign n4102 = n4101 ^ n358 ^ 1'b0 ;
  assign n4103 = n2943 & ~n4102 ;
  assign n4104 = ~n4100 & n4103 ;
  assign n4105 = n3481 ^ x11 ^ 1'b0 ;
  assign n4107 = n1871 & ~n2630 ;
  assign n4108 = ~x28 & n4107 ;
  assign n4106 = x67 & ~n1404 ;
  assign n4109 = n4108 ^ n4106 ^ 1'b0 ;
  assign n4110 = ( n693 & n4105 ) | ( n693 & n4109 ) | ( n4105 & n4109 ) ;
  assign n4111 = n998 ^ n480 ^ 1'b0 ;
  assign n4112 = ~n2797 & n4111 ;
  assign n4113 = ~n4110 & n4112 ;
  assign n4114 = n4113 ^ n2532 ^ 1'b0 ;
  assign n4115 = n2036 & ~n2064 ;
  assign n4116 = n1360 | n2040 ;
  assign n4117 = n4116 ^ n2085 ^ 1'b0 ;
  assign n4118 = n4117 ^ n2518 ^ 1'b0 ;
  assign n4119 = n311 & ~n4118 ;
  assign n4120 = n4115 & n4119 ;
  assign n4125 = x212 & x246 ;
  assign n4126 = n4125 ^ n516 ^ 1'b0 ;
  assign n4123 = n3278 ^ n766 ^ 1'b0 ;
  assign n4124 = n4123 ^ n1354 ^ 1'b0 ;
  assign n4127 = n4126 ^ n4124 ^ 1'b0 ;
  assign n4122 = n306 & ~n1685 ;
  assign n4128 = n4127 ^ n4122 ^ 1'b0 ;
  assign n4121 = n911 & ~n3131 ;
  assign n4129 = n4128 ^ n4121 ^ 1'b0 ;
  assign n4131 = n947 & ~n1202 ;
  assign n4132 = n4131 ^ n2053 ^ 1'b0 ;
  assign n4133 = x125 & ~n1572 ;
  assign n4134 = n4132 & n4133 ;
  assign n4135 = n1585 & n4134 ;
  assign n4130 = n304 | n3583 ;
  assign n4136 = n4135 ^ n4130 ^ 1'b0 ;
  assign n4137 = n304 ^ x211 ^ 1'b0 ;
  assign n4138 = n4137 ^ n1069 ^ 1'b0 ;
  assign n4139 = n326 | n4138 ;
  assign n4140 = x220 & ~n1344 ;
  assign n4141 = n4139 | n4140 ;
  assign n4142 = n471 | n4141 ;
  assign n4143 = n4142 ^ n3001 ^ 1'b0 ;
  assign n4144 = n1835 & ~n4143 ;
  assign n4145 = ( n1142 & ~n1418 ) | ( n1142 & n3270 ) | ( ~n1418 & n3270 ) ;
  assign n4146 = n4145 ^ n2907 ^ n838 ;
  assign n4147 = n1005 & ~n2997 ;
  assign n4148 = ( ~n1054 & n1757 ) | ( ~n1054 & n2595 ) | ( n1757 & n2595 ) ;
  assign n4149 = n1500 & ~n4148 ;
  assign n4150 = n1873 & n4149 ;
  assign n4151 = n4150 ^ n3878 ^ 1'b0 ;
  assign n4152 = n1698 | n4151 ;
  assign n4153 = n1813 ^ n574 ^ 1'b0 ;
  assign n4156 = n2335 ^ n1528 ^ n317 ;
  assign n4157 = n4156 ^ n3809 ^ n1358 ;
  assign n4154 = n3009 ^ n2252 ^ 1'b0 ;
  assign n4155 = ~n3422 & n4154 ;
  assign n4158 = n4157 ^ n4155 ^ 1'b0 ;
  assign n4159 = n922 | n2628 ;
  assign n4160 = n1871 | n4159 ;
  assign n4161 = x235 & ~n535 ;
  assign n4162 = n275 ^ x146 ^ 1'b0 ;
  assign n4163 = x23 & n4162 ;
  assign n4164 = n1140 ^ n776 ^ 1'b0 ;
  assign n4165 = n4163 & ~n4164 ;
  assign n4166 = n4161 & n4165 ;
  assign n4167 = n4166 ^ n1813 ^ 1'b0 ;
  assign n4168 = n1725 & n3903 ;
  assign n4169 = n1553 | n4168 ;
  assign n4170 = n883 ^ n511 ^ 1'b0 ;
  assign n4171 = n4083 ^ n395 ^ 1'b0 ;
  assign n4172 = ~n4170 & n4171 ;
  assign n4173 = n2036 ^ x7 ^ 1'b0 ;
  assign n4177 = n1651 ^ n1425 ^ n1152 ;
  assign n4178 = n4083 ^ x41 ^ 1'b0 ;
  assign n4179 = n4177 | n4178 ;
  assign n4174 = n2431 ^ n1215 ^ n1203 ;
  assign n4175 = n1166 | n2471 ;
  assign n4176 = n4174 & ~n4175 ;
  assign n4180 = n4179 ^ n4176 ^ 1'b0 ;
  assign n4184 = n2023 & ~n2091 ;
  assign n4182 = ( n2814 & n3533 ) | ( n2814 & n4080 ) | ( n3533 & n4080 ) ;
  assign n4181 = n2173 & ~n3714 ;
  assign n4183 = n4182 ^ n4181 ^ 1'b0 ;
  assign n4185 = n4184 ^ n4183 ^ 1'b0 ;
  assign n4186 = n3378 & n4185 ;
  assign n4187 = n2289 ^ n1120 ^ 1'b0 ;
  assign n4188 = n742 & ~n1037 ;
  assign n4189 = n4188 ^ n821 ^ 1'b0 ;
  assign n4190 = n4189 ^ n1877 ^ 1'b0 ;
  assign n4191 = n2358 & n4190 ;
  assign n4192 = ~x17 & x112 ;
  assign n4193 = n4191 | n4192 ;
  assign n4194 = n1295 & n4023 ;
  assign n4195 = n286 & n1782 ;
  assign n4196 = n4115 ^ n1783 ^ 1'b0 ;
  assign n4197 = n4196 ^ n1155 ^ 1'b0 ;
  assign n4198 = n4026 | n4197 ;
  assign n4199 = x115 & n956 ;
  assign n4200 = n4199 ^ n1175 ^ 1'b0 ;
  assign n4201 = n4200 ^ n2649 ^ n2630 ;
  assign n4202 = n790 & ~n4201 ;
  assign n4203 = n1041 & n4202 ;
  assign n4204 = n1795 ^ x88 ^ 1'b0 ;
  assign n4205 = n1011 | n4204 ;
  assign n4206 = n4126 ^ n631 ^ 1'b0 ;
  assign n4207 = n557 | n4206 ;
  assign n4208 = n4207 ^ n4124 ^ x218 ;
  assign n4209 = n1792 & ~n3841 ;
  assign n4210 = ( ~n4205 & n4208 ) | ( ~n4205 & n4209 ) | ( n4208 & n4209 ) ;
  assign n4211 = n3381 ^ n3361 ^ x230 ;
  assign n4212 = ( ~n768 & n1758 ) | ( ~n768 & n2434 ) | ( n1758 & n2434 ) ;
  assign n4213 = n4212 ^ n308 ^ x230 ;
  assign n4214 = n526 & ~n4213 ;
  assign n4215 = n4214 ^ n456 ^ 1'b0 ;
  assign n4216 = n4215 ^ n2660 ^ 1'b0 ;
  assign n4217 = n2566 ^ n537 ^ 1'b0 ;
  assign n4218 = ~n3937 & n4217 ;
  assign n4219 = x16 & x61 ;
  assign n4220 = ~n311 & n4219 ;
  assign n4221 = n3328 | n3688 ;
  assign n4222 = n4221 ^ n1095 ^ 1'b0 ;
  assign n4223 = n1031 | n4222 ;
  assign n4224 = ( n2596 & ~n4220 ) | ( n2596 & n4223 ) | ( ~n4220 & n4223 ) ;
  assign n4225 = n4224 ^ n2772 ^ 1'b0 ;
  assign n4226 = n4218 & n4225 ;
  assign n4227 = ~n1715 & n4226 ;
  assign n4228 = n4216 & n4227 ;
  assign n4229 = n2378 ^ n1215 ^ 1'b0 ;
  assign n4230 = ~n502 & n1319 ;
  assign n4231 = ~n2232 & n4230 ;
  assign n4232 = n4231 ^ n1769 ^ 1'b0 ;
  assign n4233 = ~n1546 & n2243 ;
  assign n4234 = n4233 ^ n2346 ^ 1'b0 ;
  assign n4235 = ( n1483 & ~n4232 ) | ( n1483 & n4234 ) | ( ~n4232 & n4234 ) ;
  assign n4241 = n279 & ~n1882 ;
  assign n4238 = n1122 ^ n1041 ^ n650 ;
  assign n4239 = n2101 | n4238 ;
  assign n4240 = n4239 ^ x22 ^ 1'b0 ;
  assign n4242 = n4241 ^ n4240 ^ 1'b0 ;
  assign n4243 = n3072 | n4242 ;
  assign n4244 = n4243 ^ n2668 ^ n2084 ;
  assign n4245 = n323 & ~n4244 ;
  assign n4236 = n970 | n1625 ;
  assign n4237 = ~n3692 & n4236 ;
  assign n4246 = n4245 ^ n4237 ^ 1'b0 ;
  assign n4247 = n3138 & ~n3227 ;
  assign n4252 = n1348 & n2132 ;
  assign n4248 = n932 ^ x247 ^ 1'b0 ;
  assign n4249 = n869 & n4248 ;
  assign n4250 = n4249 ^ n2347 ^ 1'b0 ;
  assign n4251 = n2253 | n4250 ;
  assign n4253 = n4252 ^ n4251 ^ 1'b0 ;
  assign n4254 = n2463 ^ x247 ^ 1'b0 ;
  assign n4255 = n3147 | n4254 ;
  assign n4256 = n4255 ^ n2144 ^ n1798 ;
  assign n4257 = n1926 ^ n1493 ^ 1'b0 ;
  assign n4258 = n1764 & ~n2521 ;
  assign n4259 = n2360 ^ n550 ^ 1'b0 ;
  assign n4260 = n599 | n1126 ;
  assign n4261 = n4260 ^ n744 ^ 1'b0 ;
  assign n4262 = n2956 & ~n3732 ;
  assign n4263 = ~n4261 & n4262 ;
  assign n4266 = n1691 ^ x88 ^ 1'b0 ;
  assign n4264 = n2648 | n3150 ;
  assign n4265 = x2 & ~n4264 ;
  assign n4267 = n4266 ^ n4265 ^ 1'b0 ;
  assign n4268 = ( x118 & n852 ) | ( x118 & ~n1907 ) | ( n852 & ~n1907 ) ;
  assign n4269 = n1448 ^ n552 ^ 1'b0 ;
  assign n4270 = ~n863 & n4269 ;
  assign n4271 = n4270 ^ n1657 ^ 1'b0 ;
  assign n4272 = n4271 ^ n327 ^ 1'b0 ;
  assign n4273 = n4268 & ~n4272 ;
  assign n4274 = n4273 ^ n3523 ^ 1'b0 ;
  assign n4275 = n4062 & ~n4274 ;
  assign n4278 = n3434 ^ n560 ^ 1'b0 ;
  assign n4276 = n449 | n634 ;
  assign n4277 = n4182 & n4276 ;
  assign n4279 = n4278 ^ n4277 ^ 1'b0 ;
  assign n4280 = x137 | n1976 ;
  assign n4281 = n4280 ^ n4207 ^ n420 ;
  assign n4282 = x124 & ~x140 ;
  assign n4283 = ( n1006 & ~n4281 ) | ( n1006 & n4282 ) | ( ~n4281 & n4282 ) ;
  assign n4288 = x147 & ~n1548 ;
  assign n4289 = n4288 ^ n1733 ^ 1'b0 ;
  assign n4284 = n1176 ^ n511 ^ n376 ;
  assign n4285 = ~n1941 & n4284 ;
  assign n4286 = ~n513 & n4285 ;
  assign n4287 = n2849 | n4286 ;
  assign n4290 = n4289 ^ n4287 ^ n1063 ;
  assign n4291 = ~n593 & n1601 ;
  assign n4292 = n4280 & n4291 ;
  assign n4293 = n1963 ^ x112 ^ 1'b0 ;
  assign n4294 = n2261 | n3246 ;
  assign n4295 = n4293 & ~n4294 ;
  assign n4296 = n4295 ^ n377 ^ 1'b0 ;
  assign n4302 = x231 ^ x225 ^ 1'b0 ;
  assign n4297 = n1958 & ~n3868 ;
  assign n4298 = n4297 ^ n1889 ^ 1'b0 ;
  assign n4299 = n4298 ^ n2561 ^ 1'b0 ;
  assign n4300 = n597 & n4299 ;
  assign n4301 = n3289 & n4300 ;
  assign n4303 = n4302 ^ n4301 ^ 1'b0 ;
  assign n4304 = n1000 ^ x41 ^ 1'b0 ;
  assign n4305 = n315 | n4304 ;
  assign n4306 = n4305 ^ n2942 ^ 1'b0 ;
  assign n4307 = n1179 | n3150 ;
  assign n4308 = n4307 ^ n2668 ^ 1'b0 ;
  assign n4309 = n2850 ^ n2765 ^ x88 ;
  assign n4310 = ~n344 & n1850 ;
  assign n4311 = n2168 | n3881 ;
  assign n4312 = n563 & ~n4311 ;
  assign n4313 = ~n3209 & n3415 ;
  assign n4314 = x186 & ~n4313 ;
  assign n4315 = ~x202 & n4314 ;
  assign n4316 = n574 & ~n1442 ;
  assign n4317 = n4316 ^ n2586 ^ 1'b0 ;
  assign n4318 = ~n1819 & n3738 ;
  assign n4319 = n4318 ^ n856 ^ 1'b0 ;
  assign n4320 = n4317 & n4319 ;
  assign n4321 = ~n1232 & n2285 ;
  assign n4322 = n4320 & n4321 ;
  assign n4323 = n4322 ^ n3790 ^ n449 ;
  assign n4324 = ~n2528 & n4160 ;
  assign n4325 = n3920 & n4324 ;
  assign n4326 = n1805 & ~n4325 ;
  assign n4327 = n4326 ^ n727 ^ 1'b0 ;
  assign n4328 = n3598 & ~n4327 ;
  assign n4332 = n1285 | n2204 ;
  assign n4333 = n4332 ^ x167 ^ 1'b0 ;
  assign n4329 = ~n928 & n2648 ;
  assign n4330 = n4329 ^ n269 ^ 1'b0 ;
  assign n4331 = n836 & ~n4330 ;
  assign n4334 = n4333 ^ n4331 ^ 1'b0 ;
  assign n4335 = n1702 & ~n1894 ;
  assign n4337 = n2970 ^ n1256 ^ 1'b0 ;
  assign n4338 = n2612 & n4337 ;
  assign n4336 = ~n1179 & n3166 ;
  assign n4339 = n4338 ^ n4336 ^ 1'b0 ;
  assign n4340 = ( n2946 & n4335 ) | ( n2946 & n4339 ) | ( n4335 & n4339 ) ;
  assign n4341 = n1633 ^ x5 ^ 1'b0 ;
  assign n4342 = n847 & n4341 ;
  assign n4343 = n2660 | n4342 ;
  assign n4344 = n429 & ~n4343 ;
  assign n4345 = ~n2538 & n4344 ;
  assign n4346 = n4345 ^ n2965 ^ 1'b0 ;
  assign n4347 = n3638 ^ n1804 ^ 1'b0 ;
  assign n4348 = n674 & ~n1777 ;
  assign n4349 = n2124 & n4348 ;
  assign n4350 = n519 & ~n4349 ;
  assign n4351 = n3617 & n4350 ;
  assign n4352 = n4351 ^ n3502 ^ n2536 ;
  assign n4353 = n2149 ^ n1374 ^ x0 ;
  assign n4354 = n4353 ^ n3709 ^ n3431 ;
  assign n4357 = ~n2640 & n3475 ;
  assign n4358 = n267 & n4357 ;
  assign n4355 = n2810 ^ n1788 ^ 1'b0 ;
  assign n4356 = n4355 ^ n706 ^ 1'b0 ;
  assign n4359 = n4358 ^ n4356 ^ n1000 ;
  assign n4361 = ~n2192 & n2463 ;
  assign n4362 = n4361 ^ n344 ^ 1'b0 ;
  assign n4363 = n917 & ~n4362 ;
  assign n4360 = n1395 | n1717 ;
  assign n4364 = n4363 ^ n4360 ^ 1'b0 ;
  assign n4365 = n2829 ^ n354 ^ 1'b0 ;
  assign n4366 = n926 & n4365 ;
  assign n4367 = ~n432 & n4366 ;
  assign n4368 = ~n1218 & n4367 ;
  assign n4369 = n3016 ^ n2441 ^ n666 ;
  assign n4370 = n1431 ^ n902 ^ 1'b0 ;
  assign n4371 = n4370 ^ n2085 ^ 1'b0 ;
  assign n4372 = n1601 & ~n3222 ;
  assign n4373 = ~x1 & n4372 ;
  assign n4374 = n4373 ^ n4338 ^ 1'b0 ;
  assign n4375 = n3818 & ~n4374 ;
  assign n4376 = n1199 & ~n1579 ;
  assign n4377 = n380 & ~n1446 ;
  assign n4378 = ~n4376 & n4377 ;
  assign n4379 = ( n2467 & n3779 ) | ( n2467 & ~n4378 ) | ( n3779 & ~n4378 ) ;
  assign n4380 = n4126 ^ n2573 ^ n867 ;
  assign n4381 = n907 & n1559 ;
  assign n4382 = ~n1752 & n4381 ;
  assign n4383 = ( n735 & n4380 ) | ( n735 & n4382 ) | ( n4380 & n4382 ) ;
  assign n4384 = n1347 ^ n1308 ^ 1'b0 ;
  assign n4385 = n1182 & n4384 ;
  assign n4386 = n332 | n4385 ;
  assign n4387 = n381 | n4386 ;
  assign n4388 = x15 & ~n4387 ;
  assign n4389 = x15 & ~n1991 ;
  assign n4390 = ~n3639 & n4389 ;
  assign n4391 = n4388 & n4390 ;
  assign n4393 = n1369 & n1874 ;
  assign n4394 = n4393 ^ n858 ^ 1'b0 ;
  assign n4392 = n459 & n4010 ;
  assign n4395 = n4394 ^ n4392 ^ 1'b0 ;
  assign n4396 = n4395 ^ n668 ^ 1'b0 ;
  assign n4398 = n4242 ^ n2362 ^ x204 ;
  assign n4399 = n1440 & n4398 ;
  assign n4400 = n4399 ^ n605 ^ 1'b0 ;
  assign n4397 = n1213 & ~n2544 ;
  assign n4401 = n4400 ^ n4397 ^ 1'b0 ;
  assign n4402 = n4320 | n4401 ;
  assign n4403 = x38 & x253 ;
  assign n4404 = ~n2240 & n4403 ;
  assign n4405 = n4404 ^ n4126 ^ n1225 ;
  assign n4406 = n3926 ^ n1728 ^ 1'b0 ;
  assign n4407 = n890 & n2707 ;
  assign n4408 = n530 & n3225 ;
  assign n4409 = ~n3417 & n4408 ;
  assign n4410 = ( x72 & x235 ) | ( x72 & n1172 ) | ( x235 & n1172 ) ;
  assign n4411 = n1838 & ~n3282 ;
  assign n4412 = n1797 & n4411 ;
  assign n4413 = n4412 ^ n4405 ^ 1'b0 ;
  assign n4414 = n4410 | n4413 ;
  assign n4415 = n4409 & ~n4414 ;
  assign n4416 = n1168 | n2116 ;
  assign n4417 = n4416 ^ n410 ^ 1'b0 ;
  assign n4418 = n4417 ^ x132 ^ 1'b0 ;
  assign n4419 = ~n1472 & n3003 ;
  assign n4420 = n2500 & n4419 ;
  assign n4421 = n610 & n4420 ;
  assign n4422 = ~n2151 & n2335 ;
  assign n4423 = n1350 ^ n648 ^ 1'b0 ;
  assign n4424 = n4422 & n4423 ;
  assign n4425 = ~n1138 & n4424 ;
  assign n4426 = ~n645 & n1618 ;
  assign n4428 = n354 & n2276 ;
  assign n4427 = n847 & ~n1991 ;
  assign n4429 = n4428 ^ n4427 ^ 1'b0 ;
  assign n4430 = n1881 & n4429 ;
  assign n4431 = n4052 | n4430 ;
  assign n4432 = n4431 ^ n2208 ^ 1'b0 ;
  assign n4433 = n481 & n2959 ;
  assign n4434 = n469 ^ n443 ^ 1'b0 ;
  assign n4435 = n1263 | n2160 ;
  assign n4436 = ( ~x2 & n4434 ) | ( ~x2 & n4435 ) | ( n4434 & n4435 ) ;
  assign n4437 = ~n1613 & n2281 ;
  assign n4438 = ~n1386 & n4437 ;
  assign n4439 = n781 | n4438 ;
  assign n4440 = n349 & ~n4439 ;
  assign n4441 = n4440 ^ n1666 ^ 1'b0 ;
  assign n4442 = ~n4436 & n4441 ;
  assign n4443 = n3909 ^ n712 ^ 1'b0 ;
  assign n4444 = x233 & ~n4443 ;
  assign n4445 = ~x153 & n4444 ;
  assign n4446 = ~x17 & n1786 ;
  assign n4447 = n4446 ^ n1635 ^ 1'b0 ;
  assign n4448 = ( ~n732 & n903 ) | ( ~n732 & n4447 ) | ( n903 & n4447 ) ;
  assign n4449 = ~x7 & n4448 ;
  assign n4450 = ~n725 & n4449 ;
  assign n4451 = n1980 | n3413 ;
  assign n4452 = n4451 ^ n2080 ^ 1'b0 ;
  assign n4453 = n932 & n3302 ;
  assign n4454 = ~n3980 & n4453 ;
  assign n4455 = x130 & n3734 ;
  assign n4456 = n2970 ^ n1567 ^ 1'b0 ;
  assign n4457 = n4456 ^ n2057 ^ 1'b0 ;
  assign n4461 = x85 & ~n2131 ;
  assign n4462 = n4461 ^ n3459 ^ 1'b0 ;
  assign n4463 = ~x190 & n4462 ;
  assign n4464 = n302 & ~n4463 ;
  assign n4458 = n256 | n2694 ;
  assign n4459 = x12 & n2230 ;
  assign n4460 = ~n4458 & n4459 ;
  assign n4465 = n4464 ^ n4460 ^ 1'b0 ;
  assign n4466 = n2667 | n4465 ;
  assign n4467 = n2179 ^ x123 ^ 1'b0 ;
  assign n4468 = n1988 | n4305 ;
  assign n4469 = ( ~x220 & n2637 ) | ( ~x220 & n2882 ) | ( n2637 & n2882 ) ;
  assign n4470 = n4469 ^ n2228 ^ 1'b0 ;
  assign n4471 = ~n1258 & n1978 ;
  assign n4472 = ~n4470 & n4471 ;
  assign n4473 = n4472 ^ n2300 ^ 1'b0 ;
  assign n4474 = n3557 ^ n2523 ^ 1'b0 ;
  assign n4475 = ~n288 & n520 ;
  assign n4476 = n4475 ^ n805 ^ 1'b0 ;
  assign n4477 = ( x114 & n2873 ) | ( x114 & ~n4476 ) | ( n2873 & ~n4476 ) ;
  assign n4478 = n791 ^ n605 ^ 1'b0 ;
  assign n4479 = n3141 | n4478 ;
  assign n4480 = x241 & ~n3866 ;
  assign n4481 = ~x38 & n4333 ;
  assign n4482 = n4480 | n4481 ;
  assign n4483 = n4482 ^ n592 ^ 1'b0 ;
  assign n4484 = n2772 ^ n637 ^ 1'b0 ;
  assign n4485 = n2689 & ~n4484 ;
  assign n4486 = x85 & ~n1346 ;
  assign n4487 = ~n4353 & n4486 ;
  assign n4488 = n3708 ^ n2990 ^ n2685 ;
  assign n4489 = n2900 ^ n1194 ^ 1'b0 ;
  assign n4490 = n1184 & n4489 ;
  assign n4491 = n4490 ^ n2113 ^ 1'b0 ;
  assign n4492 = ~n1726 & n2436 ;
  assign n4493 = n4492 ^ n1247 ^ 1'b0 ;
  assign n4494 = ~x111 & n4493 ;
  assign n4495 = n939 & n4494 ;
  assign n4496 = ~n2160 & n2225 ;
  assign n4497 = ( n1822 & ~n3731 ) | ( n1822 & n4406 ) | ( ~n3731 & n4406 ) ;
  assign n4498 = n640 ^ n592 ^ 1'b0 ;
  assign n4499 = n3456 ^ n2737 ^ n2008 ;
  assign n4500 = n2815 | n4499 ;
  assign n4501 = n4450 & n4500 ;
  assign n4502 = n756 ^ x160 ^ 1'b0 ;
  assign n4503 = n2621 & ~n4502 ;
  assign n4504 = x76 & ~n648 ;
  assign n4505 = ~n1230 & n4504 ;
  assign n4506 = n3078 & ~n4505 ;
  assign n4507 = n4506 ^ n4382 ^ 1'b0 ;
  assign n4508 = n1767 & n3901 ;
  assign n4509 = x4 | n2619 ;
  assign n4510 = n3193 ^ n2426 ^ n1166 ;
  assign n4511 = n4509 | n4510 ;
  assign n4512 = n3932 ^ n2728 ^ 1'b0 ;
  assign n4513 = ~n3741 & n4512 ;
  assign n4514 = ~n3229 & n4161 ;
  assign n4515 = n1742 & ~n2253 ;
  assign n4516 = n4515 ^ n666 ^ 1'b0 ;
  assign n4517 = n728 | n4516 ;
  assign n4518 = n539 | n4517 ;
  assign n4519 = n4514 | n4518 ;
  assign n4520 = n4513 | n4519 ;
  assign n4523 = n886 ^ n420 ^ 1'b0 ;
  assign n4524 = x155 & n4523 ;
  assign n4525 = n4524 ^ n2935 ^ n320 ;
  assign n4526 = n2363 & ~n4525 ;
  assign n4521 = n1494 ^ n1337 ^ 1'b0 ;
  assign n4522 = n2287 & n4521 ;
  assign n4527 = n4526 ^ n4522 ^ 1'b0 ;
  assign n4528 = n4527 ^ n3809 ^ 1'b0 ;
  assign n4529 = n2766 ^ n538 ^ 1'b0 ;
  assign n4530 = ~n1085 & n3338 ;
  assign n4531 = n1411 & n4530 ;
  assign n4532 = n3055 ^ n1646 ^ n1464 ;
  assign n4533 = ~n2490 & n3098 ;
  assign n4534 = x81 & ~n4533 ;
  assign n4535 = n1680 ^ n841 ^ 1'b0 ;
  assign n4536 = ~n1719 & n4535 ;
  assign n4537 = n2101 & n4536 ;
  assign n4538 = n1188 ^ x111 ^ 1'b0 ;
  assign n4539 = n4346 & ~n4538 ;
  assign n4540 = n3721 & n4539 ;
  assign n4541 = n2775 ^ n666 ^ 1'b0 ;
  assign n4542 = n541 | n4541 ;
  assign n4543 = n4174 ^ n1473 ^ 1'b0 ;
  assign n4544 = n3843 & n4543 ;
  assign n4545 = n4542 | n4544 ;
  assign n4546 = ~n341 & n2972 ;
  assign n4547 = n4546 ^ n2444 ^ 1'b0 ;
  assign n4548 = ( n770 & ~n781 ) | ( n770 & n4547 ) | ( ~n781 & n4547 ) ;
  assign n4549 = ( x116 & n1673 ) | ( x116 & n1850 ) | ( n1673 & n1850 ) ;
  assign n4550 = n2902 ^ x217 ^ 1'b0 ;
  assign n4552 = n928 & ~n1715 ;
  assign n4551 = n755 | n2991 ;
  assign n4553 = n4552 ^ n4551 ^ 1'b0 ;
  assign n4554 = ~n492 & n2352 ;
  assign n4555 = n3425 & n4554 ;
  assign n4556 = n4555 ^ n4466 ^ n275 ;
  assign n4557 = n2471 | n4397 ;
  assign n4558 = n739 ^ n610 ^ 1'b0 ;
  assign n4559 = n4558 ^ n1851 ^ 1'b0 ;
  assign n4560 = ~n1685 & n4559 ;
  assign n4561 = n4560 ^ n636 ^ 1'b0 ;
  assign n4562 = n3917 ^ n1571 ^ 1'b0 ;
  assign n4563 = ( n3752 & n3908 ) | ( n3752 & n4562 ) | ( n3908 & n4562 ) ;
  assign n4564 = n4563 ^ n2067 ^ 1'b0 ;
  assign n4565 = ~n957 & n4564 ;
  assign n4566 = n4565 ^ n1324 ^ 1'b0 ;
  assign n4567 = ~n1777 & n4566 ;
  assign n4568 = x44 & ~n1594 ;
  assign n4569 = ~n1295 & n4568 ;
  assign n4570 = n4386 ^ n1660 ^ x119 ;
  assign n4571 = ( n2774 & n4569 ) | ( n2774 & n4570 ) | ( n4569 & n4570 ) ;
  assign n4572 = ~n1272 & n1887 ;
  assign n4573 = n1232 & n4572 ;
  assign n4574 = n1925 & ~n4573 ;
  assign n4575 = n843 & ~n1206 ;
  assign n4576 = ( n4571 & ~n4574 ) | ( n4571 & n4575 ) | ( ~n4574 & n4575 ) ;
  assign n4577 = n2932 | n3560 ;
  assign n4578 = n1900 & ~n4577 ;
  assign n4579 = ( x173 & ~n1072 ) | ( x173 & n4578 ) | ( ~n1072 & n4578 ) ;
  assign n4580 = x141 | n1175 ;
  assign n4581 = n4246 ^ n3909 ^ 1'b0 ;
  assign n4582 = n1192 | n4581 ;
  assign n4583 = n1192 | n1716 ;
  assign n4584 = ( ~n709 & n2194 ) | ( ~n709 & n3386 ) | ( n2194 & n3386 ) ;
  assign n4585 = n4463 ^ n2443 ^ 1'b0 ;
  assign n4586 = n305 | n4585 ;
  assign n4587 = n4586 ^ n3039 ^ 1'b0 ;
  assign n4588 = n3126 ^ x208 ^ 1'b0 ;
  assign n4589 = n445 & n4588 ;
  assign n4590 = ~n1170 & n4589 ;
  assign n4591 = n2204 ^ n1450 ^ 1'b0 ;
  assign n4592 = n4591 ^ n1984 ^ n1716 ;
  assign n4593 = n4592 ^ n4145 ^ n3172 ;
  assign n4594 = n3375 ^ n1155 ^ x175 ;
  assign n4595 = n3750 & ~n4594 ;
  assign n4596 = n405 & ~n3011 ;
  assign n4597 = n2991 & n4596 ;
  assign n4598 = n4597 ^ n874 ^ 1'b0 ;
  assign n4599 = n1725 & ~n4598 ;
  assign n4600 = n2560 ^ n2376 ^ n329 ;
  assign n4601 = x15 | n1732 ;
  assign n4602 = ( x26 & n412 ) | ( x26 & ~n4601 ) | ( n412 & ~n4601 ) ;
  assign n4603 = n762 | n4410 ;
  assign n4604 = n4603 ^ n3174 ^ 1'b0 ;
  assign n4605 = n4604 ^ n3483 ^ 1'b0 ;
  assign n4606 = n624 & n4605 ;
  assign n4607 = n3803 & ~n4606 ;
  assign n4608 = n2390 ^ n577 ^ 1'b0 ;
  assign n4609 = n2124 ^ n911 ^ 1'b0 ;
  assign n4610 = n572 | n4609 ;
  assign n4611 = ( n2991 & n4608 ) | ( n2991 & n4610 ) | ( n4608 & n4610 ) ;
  assign n4612 = n1235 & ~n3140 ;
  assign n4613 = ~n2959 & n4612 ;
  assign n4614 = n4613 ^ n3785 ^ 1'b0 ;
  assign n4615 = x16 & n1233 ;
  assign n4616 = n4615 ^ n3056 ^ 1'b0 ;
  assign n4617 = ~n1897 & n2945 ;
  assign n4618 = n4617 ^ n822 ^ 1'b0 ;
  assign n4619 = ~n4015 & n4618 ;
  assign n4620 = ~n2022 & n4619 ;
  assign n4621 = n1563 | n4620 ;
  assign n4622 = n4621 ^ n2149 ^ 1'b0 ;
  assign n4625 = n1435 & n4618 ;
  assign n4626 = n4625 ^ n1033 ^ 1'b0 ;
  assign n4623 = n2680 ^ n847 ^ 1'b0 ;
  assign n4624 = n1073 | n4623 ;
  assign n4627 = n4626 ^ n4624 ^ 1'b0 ;
  assign n4628 = n3133 ^ n404 ^ 1'b0 ;
  assign n4629 = n4628 ^ n1989 ^ 1'b0 ;
  assign n4630 = n2667 | n4629 ;
  assign n4631 = n2586 ^ n2109 ^ n1077 ;
  assign n4632 = ~n1347 & n1953 ;
  assign n4633 = ~n4631 & n4632 ;
  assign n4634 = n1205 & ~n4633 ;
  assign n4638 = ~n2910 & n2972 ;
  assign n4635 = n2344 ^ n871 ^ 1'b0 ;
  assign n4636 = n1489 & n4635 ;
  assign n4637 = n471 & n4636 ;
  assign n4639 = n4638 ^ n4637 ^ 1'b0 ;
  assign n4641 = n1392 & ~n2571 ;
  assign n4640 = ~n755 & n3182 ;
  assign n4642 = n4641 ^ n4640 ^ 1'b0 ;
  assign n4643 = n4639 & ~n4642 ;
  assign n4644 = ~n1164 & n2169 ;
  assign n4645 = n4447 ^ n2028 ^ 1'b0 ;
  assign n4646 = n4644 & n4645 ;
  assign n4647 = ~n1935 & n4646 ;
  assign n4648 = ( n1509 & ~n2127 ) | ( n1509 & n4647 ) | ( ~n2127 & n4647 ) ;
  assign n4649 = n395 & ~n3322 ;
  assign n4650 = n4649 ^ n634 ^ 1'b0 ;
  assign n4651 = n2068 | n4428 ;
  assign n4655 = n420 & n679 ;
  assign n4656 = n4655 ^ x184 ^ 1'b0 ;
  assign n4653 = ~n326 & n4240 ;
  assign n4654 = ~n869 & n4653 ;
  assign n4657 = n4656 ^ n4654 ^ 1'b0 ;
  assign n4652 = ( n875 & n3229 ) | ( n875 & ~n4325 ) | ( n3229 & ~n4325 ) ;
  assign n4658 = n4657 ^ n4652 ^ 1'b0 ;
  assign n4659 = n1498 & n3059 ;
  assign n4660 = n259 & ~n1176 ;
  assign n4661 = ~x53 & n4660 ;
  assign n4662 = ( n3883 & n4370 ) | ( n3883 & ~n4661 ) | ( n4370 & ~n4661 ) ;
  assign n4663 = n4659 & n4662 ;
  assign n4664 = n4663 ^ n2095 ^ 1'b0 ;
  assign n4665 = n2070 ^ n1176 ^ 1'b0 ;
  assign n4666 = n4664 & n4665 ;
  assign n4669 = ~x241 & n1913 ;
  assign n4670 = n4669 ^ x7 ^ 1'b0 ;
  assign n4667 = n4148 ^ x43 ^ 1'b0 ;
  assign n4668 = n2279 | n4667 ;
  assign n4671 = n4670 ^ n4668 ^ 1'b0 ;
  assign n4672 = n1863 | n4671 ;
  assign n4673 = n1846 ^ x184 ^ 1'b0 ;
  assign n4674 = n2324 & ~n2531 ;
  assign n4675 = ~n363 & n574 ;
  assign n4676 = n4675 ^ n817 ^ 1'b0 ;
  assign n4677 = n342 & ~n4676 ;
  assign n4678 = n3676 & n4677 ;
  assign n4679 = n4678 ^ n677 ^ 1'b0 ;
  assign n4680 = n4679 ^ n518 ^ 1'b0 ;
  assign n4681 = n2720 & ~n4680 ;
  assign n4682 = n1514 ^ n1415 ^ 1'b0 ;
  assign n4683 = n1980 & n4682 ;
  assign n4684 = ~n3088 & n4683 ;
  assign n4685 = n1055 | n2127 ;
  assign n4686 = n1608 & ~n4685 ;
  assign n4687 = n3468 & ~n3668 ;
  assign n4688 = n1757 & n4687 ;
  assign n4689 = n4686 & ~n4688 ;
  assign n4690 = n3228 ^ n312 ^ 1'b0 ;
  assign n4691 = n4689 | n4690 ;
  assign n4692 = n420 | n4043 ;
  assign n4693 = n4692 ^ n4031 ^ 1'b0 ;
  assign n4694 = n1760 ^ n987 ^ 1'b0 ;
  assign n4695 = ~n3135 & n4694 ;
  assign n4696 = n4473 & n4695 ;
  assign n4700 = n1380 & n1860 ;
  assign n4701 = n4700 ^ n3333 ^ 1'b0 ;
  assign n4702 = x171 & ~n4701 ;
  assign n4703 = ~n1284 & n4702 ;
  assign n4697 = n1249 & n4137 ;
  assign n4698 = n4697 ^ n1700 ^ 1'b0 ;
  assign n4699 = n4698 ^ n1430 ^ 1'b0 ;
  assign n4704 = n4703 ^ n4699 ^ 1'b0 ;
  assign n4705 = n4704 ^ n1885 ^ 1'b0 ;
  assign n4706 = ~n2901 & n3161 ;
  assign n4707 = n4706 ^ x15 ^ 1'b0 ;
  assign n4710 = n2897 & ~n3328 ;
  assign n4708 = n4338 ^ n3322 ^ 1'b0 ;
  assign n4709 = ~n1729 & n4708 ;
  assign n4711 = n4710 ^ n4709 ^ n4187 ;
  assign n4712 = x136 & n683 ;
  assign n4713 = n4033 & n4712 ;
  assign n4714 = n860 ^ n719 ^ 1'b0 ;
  assign n4715 = n1064 ^ n652 ^ 1'b0 ;
  assign n4716 = n4715 ^ n1312 ^ 1'b0 ;
  assign n4717 = n1949 | n2728 ;
  assign n4718 = n4717 ^ n1147 ^ 1'b0 ;
  assign n4719 = n4718 ^ n1665 ^ n449 ;
  assign n4720 = n1278 | n2320 ;
  assign n4721 = n624 | n4720 ;
  assign n4722 = n4721 ^ n1166 ^ x143 ;
  assign n4723 = n2973 ^ n1860 ^ 1'b0 ;
  assign n4724 = n1469 & ~n2314 ;
  assign n4729 = n2028 & n4505 ;
  assign n4726 = n3088 & n3465 ;
  assign n4727 = n4726 ^ n731 ^ 1'b0 ;
  assign n4725 = ~n381 & n3166 ;
  assign n4728 = n4727 ^ n4725 ^ 1'b0 ;
  assign n4730 = n4729 ^ n4728 ^ 1'b0 ;
  assign n4731 = ~n4724 & n4730 ;
  assign n4732 = ~n1512 & n3888 ;
  assign n4733 = ~n1199 & n2012 ;
  assign n4734 = n4733 ^ n2182 ^ 1'b0 ;
  assign n4735 = ( n2786 & n4732 ) | ( n2786 & ~n4734 ) | ( n4732 & ~n4734 ) ;
  assign n4736 = n1024 & ~n4735 ;
  assign n4737 = n3809 ^ n3740 ^ 1'b0 ;
  assign n4738 = n3556 & ~n4737 ;
  assign n4739 = n1199 & ~n4517 ;
  assign n4740 = n4738 & ~n4739 ;
  assign n4741 = n4740 ^ n933 ^ 1'b0 ;
  assign n4742 = ~n2160 & n4383 ;
  assign n4743 = n4513 ^ n2337 ^ 1'b0 ;
  assign n4744 = n4743 ^ x208 ^ 1'b0 ;
  assign n4745 = n4331 ^ n2087 ^ 1'b0 ;
  assign n4746 = n1657 | n4745 ;
  assign n4747 = n2481 | n4746 ;
  assign n4748 = n1679 | n4747 ;
  assign n4749 = n4386 & n4748 ;
  assign n4750 = n3777 & n3970 ;
  assign n4751 = n4750 ^ n2735 ^ 1'b0 ;
  assign n4752 = x185 & n354 ;
  assign n4753 = ( x11 & n604 ) | ( x11 & n3164 ) | ( n604 & n3164 ) ;
  assign n4754 = n3035 | n4753 ;
  assign n4758 = x189 | n1766 ;
  assign n4759 = n704 ^ n415 ^ n284 ;
  assign n4760 = n4759 ^ n1741 ^ 1'b0 ;
  assign n4761 = ( n2708 & ~n4758 ) | ( n2708 & n4760 ) | ( ~n4758 & n4760 ) ;
  assign n4755 = ~n305 & n1626 ;
  assign n4756 = ~n1792 & n4755 ;
  assign n4757 = ( ~n822 & n4422 ) | ( ~n822 & n4756 ) | ( n4422 & n4756 ) ;
  assign n4762 = n4761 ^ n4757 ^ n4467 ;
  assign n4763 = n537 | n1884 ;
  assign n4764 = n4763 ^ n1889 ^ 1'b0 ;
  assign n4765 = n1887 & n4764 ;
  assign n4766 = n4123 ^ n3782 ^ n3490 ;
  assign n4767 = n4765 & n4766 ;
  assign n4768 = ( ~n897 & n970 ) | ( ~n897 & n2173 ) | ( n970 & n2173 ) ;
  assign n4769 = n4768 ^ n571 ^ 1'b0 ;
  assign n4770 = n4769 ^ n1493 ^ 1'b0 ;
  assign n4771 = n4042 ^ n3586 ^ 1'b0 ;
  assign n4772 = n731 | n4771 ;
  assign n4773 = ( n1559 & n4770 ) | ( n1559 & n4772 ) | ( n4770 & n4772 ) ;
  assign n4774 = ( n2217 & ~n3175 ) | ( n2217 & n4773 ) | ( ~n3175 & n4773 ) ;
  assign n4775 = n1878 ^ n449 ^ 1'b0 ;
  assign n4777 = n1817 ^ n1558 ^ n492 ;
  assign n4776 = ~n405 & n3600 ;
  assign n4778 = n4777 ^ n4776 ^ x16 ;
  assign n4779 = n692 | n1023 ;
  assign n4780 = n504 | n4779 ;
  assign n4781 = n1665 & n2991 ;
  assign n4782 = n4781 ^ n506 ^ 1'b0 ;
  assign n4783 = ~n4780 & n4782 ;
  assign n4786 = n1177 ^ x45 ^ 1'b0 ;
  assign n4787 = n659 & n4786 ;
  assign n4788 = ~n4289 & n4787 ;
  assign n4789 = n3770 & n4788 ;
  assign n4784 = n2207 ^ n1202 ^ 1'b0 ;
  assign n4785 = ~n1600 & n4784 ;
  assign n4790 = n4789 ^ n4785 ^ 1'b0 ;
  assign n4791 = n3419 ^ n1166 ^ 1'b0 ;
  assign n4792 = ~n3584 & n4791 ;
  assign n4793 = n707 & n1223 ;
  assign n4794 = n345 & n4793 ;
  assign n4795 = n4794 ^ n1944 ^ 1'b0 ;
  assign n4796 = n2955 | n4795 ;
  assign n4797 = ~n1176 & n4796 ;
  assign n4798 = n832 & ~n1124 ;
  assign n4799 = n1600 & n4798 ;
  assign n4800 = n535 & ~n4799 ;
  assign n4801 = n535 ^ x133 ^ 1'b0 ;
  assign n4802 = n2755 | n4801 ;
  assign n4803 = n4802 ^ n3222 ^ n791 ;
  assign n4804 = n1544 ^ x139 ^ 1'b0 ;
  assign n4805 = n2623 | n4804 ;
  assign n4806 = n1981 | n4805 ;
  assign n4807 = x112 | n4049 ;
  assign n4808 = n1648 ^ n1255 ^ n545 ;
  assign n4809 = ( ~n4286 & n4807 ) | ( ~n4286 & n4808 ) | ( n4807 & n4808 ) ;
  assign n4810 = n4809 ^ n3310 ^ n1732 ;
  assign n4811 = n4174 ^ n3750 ^ 1'b0 ;
  assign n4812 = ~n1067 & n4811 ;
  assign n4813 = n2303 | n4724 ;
  assign n4814 = n1225 & ~n4813 ;
  assign n4815 = n2171 & n4814 ;
  assign n4816 = ~x7 & n2249 ;
  assign n4817 = n1081 | n4816 ;
  assign n4818 = n3373 & n4817 ;
  assign n4819 = ~x176 & n740 ;
  assign n4820 = n4819 ^ n2244 ^ 1'b0 ;
  assign n4821 = n4137 ^ n1446 ^ 1'b0 ;
  assign n4822 = n1253 | n1258 ;
  assign n4823 = n2423 & ~n4822 ;
  assign n4824 = n4823 ^ n731 ^ 1'b0 ;
  assign n4825 = n4821 | n4824 ;
  assign n4826 = n1228 & ~n4825 ;
  assign n4829 = x132 & n3131 ;
  assign n4827 = x23 & ~n622 ;
  assign n4828 = ( x21 & ~n764 ) | ( x21 & n4827 ) | ( ~n764 & n4827 ) ;
  assign n4830 = n4829 ^ n4828 ^ 1'b0 ;
  assign n4831 = n418 | n4252 ;
  assign n4832 = n4831 ^ n924 ^ 1'b0 ;
  assign n4838 = n3150 ^ n1423 ^ 1'b0 ;
  assign n4839 = n2651 & n4838 ;
  assign n4833 = n527 ^ x78 ^ 1'b0 ;
  assign n4834 = n2521 & n4833 ;
  assign n4835 = n4834 ^ x230 ^ 1'b0 ;
  assign n4836 = ~n4514 & n4835 ;
  assign n4837 = ~n4140 & n4836 ;
  assign n4840 = n4839 ^ n4837 ^ 1'b0 ;
  assign n4841 = n306 ^ x194 ^ 1'b0 ;
  assign n4842 = n1879 & n4841 ;
  assign n4843 = ~n1515 & n3097 ;
  assign n4844 = ~n3421 & n4843 ;
  assign n4845 = ( n482 & n1115 ) | ( n482 & ~n1228 ) | ( n1115 & ~n1228 ) ;
  assign n4846 = n4845 ^ n4729 ^ 1'b0 ;
  assign n4847 = n882 & ~n4505 ;
  assign n4848 = n2765 & n4847 ;
  assign n4849 = ~n3384 & n4848 ;
  assign n4850 = n4047 ^ n1579 ^ 1'b0 ;
  assign n4853 = x175 | n436 ;
  assign n4851 = n1783 ^ n265 ^ 1'b0 ;
  assign n4852 = ~n617 & n4851 ;
  assign n4854 = n4853 ^ n4852 ^ 1'b0 ;
  assign n4855 = n2523 & n4854 ;
  assign n4856 = ~n718 & n4855 ;
  assign n4857 = ~n790 & n4856 ;
  assign n4858 = n4857 ^ n522 ^ 1'b0 ;
  assign n4859 = ( n874 & n1024 ) | ( n874 & ~n2943 ) | ( n1024 & ~n2943 ) ;
  assign n4860 = ~n259 & n2956 ;
  assign n4861 = n3419 & ~n4860 ;
  assign n4862 = n4861 ^ n2378 ^ 1'b0 ;
  assign n4863 = n4859 & n4862 ;
  assign n4864 = ~n803 & n4863 ;
  assign n4865 = n4864 ^ n3402 ^ n2854 ;
  assign n4866 = ~n1023 & n1767 ;
  assign n4867 = n4866 ^ x126 ^ 1'b0 ;
  assign n4868 = n4867 ^ n1272 ^ 1'b0 ;
  assign n4869 = n1289 ^ x120 ^ 1'b0 ;
  assign n4870 = ~n3071 & n4869 ;
  assign n4871 = n580 & n1722 ;
  assign n4872 = n4871 ^ n539 ^ 1'b0 ;
  assign n4873 = n4872 ^ n4638 ^ n2063 ;
  assign n4875 = ~n1703 & n2241 ;
  assign n4876 = n267 & n4875 ;
  assign n4877 = n4876 ^ n2363 ^ 1'b0 ;
  assign n4878 = n1040 & ~n4877 ;
  assign n4874 = ~n365 & n3687 ;
  assign n4879 = n4878 ^ n4874 ^ 1'b0 ;
  assign n4880 = n4879 ^ n4583 ^ n1746 ;
  assign n4881 = ~n2434 & n3689 ;
  assign n4882 = n1192 & ~n2081 ;
  assign n4889 = n2719 ^ n1777 ^ x81 ;
  assign n4883 = n4220 ^ n2282 ^ 1'b0 ;
  assign n4884 = n1681 | n4883 ;
  assign n4885 = n4884 ^ n3434 ^ n1126 ;
  assign n4886 = n4885 ^ n1965 ^ 1'b0 ;
  assign n4887 = n577 & n4886 ;
  assign n4888 = n3843 & n4887 ;
  assign n4890 = n4889 ^ n4888 ^ 1'b0 ;
  assign n4896 = n589 ^ x213 ^ 1'b0 ;
  assign n4891 = n1340 ^ n869 ^ n439 ;
  assign n4892 = n300 & n4891 ;
  assign n4893 = ~n639 & n4892 ;
  assign n4894 = n1378 & n4893 ;
  assign n4895 = n4894 ^ n1526 ^ n365 ;
  assign n4897 = n4896 ^ n4895 ^ 1'b0 ;
  assign n4898 = ~n2100 & n4897 ;
  assign n4899 = ( ~n4654 & n4750 ) | ( ~n4654 & n4898 ) | ( n4750 & n4898 ) ;
  assign n4900 = n4899 ^ n3000 ^ 1'b0 ;
  assign n4901 = n335 & ~n1917 ;
  assign n4902 = n1819 | n1882 ;
  assign n4903 = ~n778 & n4902 ;
  assign n4904 = n4903 ^ n4642 ^ 1'b0 ;
  assign n4905 = n4901 & n4904 ;
  assign n4906 = n2674 ^ n527 ^ 1'b0 ;
  assign n4907 = x1 & ~n4906 ;
  assign n4910 = ( n281 & n1058 ) | ( n281 & ~n1603 ) | ( n1058 & ~n1603 ) ;
  assign n4908 = n843 & ~n4686 ;
  assign n4909 = n4908 ^ n527 ^ 1'b0 ;
  assign n4911 = n4910 ^ n4909 ^ n1475 ;
  assign n4912 = n1244 & n4911 ;
  assign n4913 = ~n1134 & n2826 ;
  assign n4914 = n3752 | n4505 ;
  assign n4915 = n3709 & ~n4914 ;
  assign n4916 = n1403 ^ n1110 ^ 1'b0 ;
  assign n4917 = n1138 & n4916 ;
  assign n4918 = ( n737 & n1631 ) | ( n737 & ~n4917 ) | ( n1631 & ~n4917 ) ;
  assign n4919 = n4585 ^ n694 ^ 1'b0 ;
  assign n4920 = x84 & ~n4919 ;
  assign n4921 = n4920 ^ n3330 ^ n549 ;
  assign n4922 = n4921 ^ n2567 ^ 1'b0 ;
  assign n4923 = n4918 & ~n4922 ;
  assign n4924 = n1692 ^ n1571 ^ 1'b0 ;
  assign n4925 = ~n4923 & n4924 ;
  assign n4926 = n3008 ^ x10 ^ 1'b0 ;
  assign n4927 = n4926 ^ n4146 ^ n2101 ;
  assign n4928 = n3829 ^ n2640 ^ 1'b0 ;
  assign n4929 = n686 & ~n4928 ;
  assign n4931 = ( n2264 & ~n3716 ) | ( n2264 & n4585 ) | ( ~n3716 & n4585 ) ;
  assign n4932 = ~n1801 & n4819 ;
  assign n4933 = n2218 ^ n1527 ^ 1'b0 ;
  assign n4934 = ~n4932 & n4933 ;
  assign n4935 = n939 & n4934 ;
  assign n4936 = ~n4931 & n4935 ;
  assign n4930 = n3239 & ~n4027 ;
  assign n4937 = n4936 ^ n4930 ^ 1'b0 ;
  assign n4938 = n2678 ^ n905 ^ 1'b0 ;
  assign n4939 = n3696 ^ n288 ^ 1'b0 ;
  assign n4940 = n4938 & n4939 ;
  assign n4941 = n2614 & n4940 ;
  assign n4942 = n729 ^ n583 ^ 1'b0 ;
  assign n4943 = n2302 & ~n4942 ;
  assign n4944 = ~n4941 & n4943 ;
  assign n4945 = ~n2050 & n4944 ;
  assign n4946 = x29 & n3182 ;
  assign n4947 = ~x74 & n4946 ;
  assign n4948 = ( x36 & ~n1823 ) | ( x36 & n4947 ) | ( ~n1823 & n4947 ) ;
  assign n4949 = ~n781 & n4948 ;
  assign n4950 = n3552 & n4949 ;
  assign n4951 = n322 & ~n1832 ;
  assign n4952 = x116 & x251 ;
  assign n4953 = n4952 ^ x213 ^ 1'b0 ;
  assign n4954 = n4953 ^ n4881 ^ n1472 ;
  assign n4959 = n531 | n924 ;
  assign n4956 = n1052 ^ n472 ^ 1'b0 ;
  assign n4955 = n1289 & n3118 ;
  assign n4957 = n4956 ^ n4955 ^ 1'b0 ;
  assign n4958 = n1007 | n4957 ;
  assign n4960 = n4959 ^ n4958 ^ 1'b0 ;
  assign n4961 = n3399 ^ n1308 ^ 1'b0 ;
  assign n4962 = ~n640 & n4961 ;
  assign n4963 = n1026 | n1909 ;
  assign n4964 = x207 | n4963 ;
  assign n4965 = n4964 ^ n1179 ^ 1'b0 ;
  assign n4966 = n984 & ~n4965 ;
  assign n4967 = ~x195 & n4966 ;
  assign n4968 = n2597 | n4967 ;
  assign n4969 = n4962 | n4968 ;
  assign n4970 = n721 & n4428 ;
  assign n4971 = n2525 & ~n4970 ;
  assign n4972 = n3170 & ~n4220 ;
  assign n4973 = ~n1928 & n4972 ;
  assign n4974 = n998 | n2682 ;
  assign n4975 = n1780 & ~n4974 ;
  assign n4976 = n4973 | n4975 ;
  assign n4977 = n4976 ^ n4674 ^ 1'b0 ;
  assign n4978 = n1764 & ~n2659 ;
  assign n4980 = ( x234 & n338 ) | ( x234 & ~n1275 ) | ( n338 & ~n1275 ) ;
  assign n4979 = n1313 & n4160 ;
  assign n4981 = n4980 ^ n4979 ^ 1'b0 ;
  assign n4982 = n1871 | n4981 ;
  assign n4989 = ~n315 & n988 ;
  assign n4990 = ~n2151 & n4989 ;
  assign n4983 = x136 & n1097 ;
  assign n4984 = ~n3978 & n4983 ;
  assign n4985 = n1261 | n4984 ;
  assign n4986 = n1010 & ~n4985 ;
  assign n4987 = n4986 ^ n449 ^ 1'b0 ;
  assign n4988 = ~n2433 & n4987 ;
  assign n4991 = n4990 ^ n4988 ^ 1'b0 ;
  assign n4992 = x178 & ~n3089 ;
  assign n4993 = n4992 ^ n2076 ^ 1'b0 ;
  assign n4994 = n1455 & n4993 ;
  assign n4995 = n718 ^ n358 ^ n294 ;
  assign n4996 = n1760 ^ x35 ^ 1'b0 ;
  assign n4997 = n690 | n4404 ;
  assign n4998 = n2212 & ~n4997 ;
  assign n4999 = n4996 | n4998 ;
  assign n5000 = ~n4023 & n4870 ;
  assign n5001 = n1707 & n5000 ;
  assign n5002 = n4156 ^ n4076 ^ 1'b0 ;
  assign n5003 = x194 & ~n5002 ;
  assign n5004 = ~n1019 & n3232 ;
  assign n5005 = n1520 | n5004 ;
  assign n5006 = n856 & ~n5005 ;
  assign n5007 = n371 ^ x243 ^ 1'b0 ;
  assign n5008 = x48 & ~n5007 ;
  assign n5009 = ~n1716 & n5008 ;
  assign n5010 = n2967 ^ n2902 ^ 1'b0 ;
  assign n5011 = n5010 ^ n311 ^ 1'b0 ;
  assign n5012 = n2481 | n3132 ;
  assign n5013 = n5012 ^ n4661 ^ 1'b0 ;
  assign n5014 = n5013 ^ n3131 ^ 1'b0 ;
  assign n5015 = x76 & ~n2595 ;
  assign n5016 = ~n3345 & n5015 ;
  assign n5017 = n5014 | n5016 ;
  assign n5018 = n441 & ~n840 ;
  assign n5019 = ~n2255 & n5018 ;
  assign n5020 = n1737 | n5019 ;
  assign n5021 = n2684 | n4364 ;
  assign n5022 = ( n393 & ~n1113 ) | ( n393 & n3183 ) | ( ~n1113 & n3183 ) ;
  assign n5023 = x243 & n511 ;
  assign n5024 = n610 | n3223 ;
  assign n5025 = n3842 & ~n5024 ;
  assign n5026 = x15 | n612 ;
  assign n5027 = n5025 & ~n5026 ;
  assign n5028 = ( n1431 & n2827 ) | ( n1431 & ~n4585 ) | ( n2827 & ~n4585 ) ;
  assign n5029 = n4379 | n5028 ;
  assign n5030 = n686 & n4532 ;
  assign n5031 = n5030 ^ n2637 ^ 1'b0 ;
  assign n5032 = ~n1924 & n2959 ;
  assign n5033 = n5032 ^ n397 ^ 1'b0 ;
  assign n5034 = n3419 & ~n5033 ;
  assign n5035 = n5034 ^ n5010 ^ 1'b0 ;
  assign n5036 = n3289 & n5035 ;
  assign n5037 = n288 | n1575 ;
  assign n5038 = n5037 ^ n2738 ^ 1'b0 ;
  assign n5039 = n5038 ^ n3388 ^ n2253 ;
  assign n5040 = ( n1889 & ~n2761 ) | ( n1889 & n4255 ) | ( ~n2761 & n4255 ) ;
  assign n5042 = n1546 ^ n415 ^ 1'b0 ;
  assign n5041 = ~n900 & n1692 ;
  assign n5043 = n5042 ^ n5041 ^ 1'b0 ;
  assign n5044 = n5040 & n5043 ;
  assign n5045 = n5044 ^ n1547 ^ 1'b0 ;
  assign n5046 = n1678 ^ x247 ^ 1'b0 ;
  assign n5047 = n3367 | n3641 ;
  assign n5048 = n4021 ^ n3755 ^ n2965 ;
  assign n5049 = n1230 & n4395 ;
  assign n5050 = n5049 ^ n2826 ^ n1250 ;
  assign n5051 = ( n2830 & n3490 ) | ( n2830 & n4655 ) | ( n3490 & n4655 ) ;
  assign n5052 = ( ~n904 & n1739 ) | ( ~n904 & n5051 ) | ( n1739 & n5051 ) ;
  assign n5053 = x15 | n1127 ;
  assign n5054 = n4284 ^ n3592 ^ n527 ;
  assign n5055 = n526 ^ n485 ^ 1'b0 ;
  assign n5056 = ~n2644 & n5055 ;
  assign n5057 = ~x125 & n1409 ;
  assign n5058 = n1486 & n2871 ;
  assign n5059 = ~n817 & n5058 ;
  assign n5060 = n5059 ^ n4137 ^ 1'b0 ;
  assign n5061 = n5060 ^ n1622 ^ 1'b0 ;
  assign n5062 = n4580 ^ n3218 ^ 1'b0 ;
  assign n5063 = n4026 | n5062 ;
  assign n5064 = ~x17 & n2981 ;
  assign n5065 = n4982 ^ n4096 ^ 1'b0 ;
  assign n5066 = n2648 & n5065 ;
  assign n5067 = n5066 ^ n858 ^ 1'b0 ;
  assign n5068 = ~n1536 & n5023 ;
  assign n5069 = n2830 & n3043 ;
  assign n5070 = ~n2690 & n5069 ;
  assign n5071 = n3972 ^ n1876 ^ n1275 ;
  assign n5072 = n2305 | n5071 ;
  assign n5073 = ~n1538 & n3441 ;
  assign n5074 = n5073 ^ n3696 ^ n2320 ;
  assign n5075 = n1416 & n2477 ;
  assign n5076 = x254 & ~n873 ;
  assign n5077 = ~x123 & n5076 ;
  assign n5078 = n5077 ^ n631 ^ 1'b0 ;
  assign n5079 = x73 & n5078 ;
  assign n5080 = ~n3261 & n4323 ;
  assign n5081 = ~n5079 & n5080 ;
  assign n5082 = n921 & n4077 ;
  assign n5083 = n5082 ^ n1253 ^ 1'b0 ;
  assign n5084 = n5083 ^ n1860 ^ n1111 ;
  assign n5085 = ~n1334 & n1866 ;
  assign n5086 = n5085 ^ n2382 ^ 1'b0 ;
  assign n5087 = ~n3832 & n5086 ;
  assign n5088 = n1525 ^ n372 ^ 1'b0 ;
  assign n5089 = ~n3778 & n5088 ;
  assign n5090 = ~n5087 & n5089 ;
  assign n5091 = n2221 ^ x164 ^ 1'b0 ;
  assign n5092 = x62 & n3672 ;
  assign n5093 = ~x104 & n3082 ;
  assign n5094 = n860 ^ n553 ^ 1'b0 ;
  assign n5095 = n1666 & ~n5094 ;
  assign n5096 = n2956 & ~n5095 ;
  assign n5097 = n1308 ^ x101 ^ 1'b0 ;
  assign n5098 = n5096 & n5097 ;
  assign n5099 = n5098 ^ n4921 ^ n2726 ;
  assign n5100 = n1295 ^ n296 ^ 1'b0 ;
  assign n5101 = x143 & ~n3903 ;
  assign n5102 = n5100 & n5101 ;
  assign n5103 = n2586 ^ n690 ^ 1'b0 ;
  assign n5104 = n5103 ^ n5006 ^ 1'b0 ;
  assign n5105 = ~n1404 & n5104 ;
  assign n5107 = n2970 ^ n967 ^ n729 ;
  assign n5106 = n1610 & n2294 ;
  assign n5108 = n5107 ^ n5106 ^ 1'b0 ;
  assign n5109 = n5108 ^ n1122 ^ 1'b0 ;
  assign n5110 = ~n780 & n5109 ;
  assign n5111 = n2527 & n3208 ;
  assign n5112 = ~n4618 & n5111 ;
  assign n5113 = n833 & ~n5112 ;
  assign n5115 = ( n852 & ~n1347 ) | ( n852 & n1903 ) | ( ~n1347 & n1903 ) ;
  assign n5114 = n1479 & n3686 ;
  assign n5116 = n5115 ^ n5114 ^ n2667 ;
  assign n5117 = x6 & n2736 ;
  assign n5121 = ( x239 & n1358 ) | ( x239 & ~n2160 ) | ( n1358 & ~n2160 ) ;
  assign n5118 = ~n781 & n1555 ;
  assign n5119 = n5118 ^ n1168 ^ 1'b0 ;
  assign n5120 = ~n1943 & n5119 ;
  assign n5122 = n5121 ^ n5120 ^ 1'b0 ;
  assign n5123 = n5122 ^ n2349 ^ 1'b0 ;
  assign n5124 = ~n1139 & n5123 ;
  assign n5125 = n1582 ^ n626 ^ 1'b0 ;
  assign n5126 = n2340 | n5125 ;
  assign n5127 = n4478 & ~n5126 ;
  assign n5128 = n4987 ^ n2885 ^ 1'b0 ;
  assign n5129 = ~n5127 & n5128 ;
  assign n5130 = n5129 ^ n3714 ^ 1'b0 ;
  assign n5131 = n5130 ^ n2962 ^ n740 ;
  assign n5132 = ( n387 & n677 ) | ( n387 & ~n4638 ) | ( n677 & ~n4638 ) ;
  assign n5133 = n5132 ^ n3409 ^ 1'b0 ;
  assign n5134 = n294 & ~n2664 ;
  assign n5135 = n1354 & ~n1771 ;
  assign n5136 = n5135 ^ n2201 ^ x170 ;
  assign n5137 = n5136 ^ n2431 ^ n967 ;
  assign n5138 = n3557 & ~n5137 ;
  assign n5139 = n5138 ^ n2866 ^ n1766 ;
  assign n5140 = ~x26 & n284 ;
  assign n5141 = n4418 | n5140 ;
  assign n5142 = n4500 ^ x81 ^ 1'b0 ;
  assign n5143 = ( x15 & n947 ) | ( x15 & ~n4212 ) | ( n947 & ~n4212 ) ;
  assign n5144 = n840 & ~n2674 ;
  assign n5145 = n5144 ^ n4549 ^ n1060 ;
  assign n5148 = n2561 | n3169 ;
  assign n5149 = n1500 | n5148 ;
  assign n5146 = x32 | n1126 ;
  assign n5147 = n5146 ^ n1486 ^ 1'b0 ;
  assign n5150 = n5149 ^ n5147 ^ n4881 ;
  assign n5151 = n3208 ^ n3007 ^ 1'b0 ;
  assign n5152 = ~n3227 & n5151 ;
  assign n5153 = n5152 ^ n2875 ^ 1'b0 ;
  assign n5154 = ~n2950 & n5153 ;
  assign n5155 = ( x120 & ~x195 ) | ( x120 & n2548 ) | ( ~x195 & n2548 ) ;
  assign n5156 = n5155 ^ n2852 ^ 1'b0 ;
  assign n5157 = n1105 | n5156 ;
  assign n5158 = n5157 ^ n3152 ^ 1'b0 ;
  assign n5159 = n1369 & n5158 ;
  assign n5160 = n5159 ^ n3133 ^ 1'b0 ;
  assign n5161 = n2020 ^ n633 ^ 1'b0 ;
  assign n5162 = n1593 ^ n1129 ^ n418 ;
  assign n5163 = n5161 & n5162 ;
  assign n5164 = n5163 ^ n473 ^ 1'b0 ;
  assign n5165 = x221 ^ x3 ^ 1'b0 ;
  assign n5166 = n3854 & n5165 ;
  assign n5167 = n5166 ^ n1829 ^ 1'b0 ;
  assign n5168 = n2339 & n3555 ;
  assign n5169 = n5168 ^ x91 ^ 1'b0 ;
  assign n5170 = n5169 ^ n2974 ^ x239 ;
  assign n5171 = n5170 ^ n4245 ^ 1'b0 ;
  assign n5172 = n3087 | n5171 ;
  assign n5173 = n4864 ^ n2897 ^ 1'b0 ;
  assign n5174 = n2618 ^ n1906 ^ 1'b0 ;
  assign n5175 = n3598 & ~n5174 ;
  assign n5176 = n1233 | n5175 ;
  assign n5177 = ( ~n1233 & n2573 ) | ( ~n1233 & n3198 ) | ( n2573 & n3198 ) ;
  assign n5178 = n5177 ^ n3658 ^ 1'b0 ;
  assign n5182 = ( x123 & x170 ) | ( x123 & ~x254 ) | ( x170 & ~x254 ) ;
  assign n5183 = n2259 & n5182 ;
  assign n5184 = n2289 & n5183 ;
  assign n5179 = n4910 ^ n481 ^ 1'b0 ;
  assign n5180 = n4677 & n5179 ;
  assign n5181 = n3979 & n5180 ;
  assign n5185 = n5184 ^ n5181 ^ 1'b0 ;
  assign n5186 = ~n954 & n1260 ;
  assign n5187 = n698 & n5186 ;
  assign n5188 = n5187 ^ n2101 ^ 1'b0 ;
  assign n5189 = n1101 | n5188 ;
  assign n5190 = n2714 & ~n5189 ;
  assign n5191 = n3307 ^ n2849 ^ 1'b0 ;
  assign n5192 = n1177 & n5191 ;
  assign n5193 = n1283 & n5192 ;
  assign n5194 = n4573 ^ n1486 ^ 1'b0 ;
  assign n5195 = n5194 ^ n993 ^ x71 ;
  assign n5196 = n4817 & ~n5195 ;
  assign n5197 = n5196 ^ n2768 ^ 1'b0 ;
  assign n5198 = ~n5193 & n5197 ;
  assign n5199 = n3185 ^ n481 ^ 1'b0 ;
  assign n5200 = n5198 & ~n5199 ;
  assign n5201 = x20 & ~n4035 ;
  assign n5202 = ~x10 & n5201 ;
  assign n5203 = n3183 & ~n5202 ;
  assign n5204 = n2603 ^ n1645 ^ 1'b0 ;
  assign n5205 = n733 | n5204 ;
  assign n5206 = n4015 ^ n2686 ^ 1'b0 ;
  assign n5207 = n2085 & ~n5206 ;
  assign n5208 = n5207 ^ n1970 ^ 1'b0 ;
  assign n5209 = ~n847 & n3547 ;
  assign n5210 = n1603 | n2187 ;
  assign n5211 = ~n3905 & n5210 ;
  assign n5212 = x253 & n2248 ;
  assign n5213 = n5212 ^ n1499 ^ 1'b0 ;
  assign n5214 = n5213 ^ n3208 ^ 1'b0 ;
  assign n5215 = n5211 & ~n5214 ;
  assign n5216 = ~n5209 & n5215 ;
  assign n5218 = n317 & ~n1148 ;
  assign n5217 = n1319 & n1692 ;
  assign n5219 = n5218 ^ n5217 ^ n2483 ;
  assign n5220 = ~n3769 & n5219 ;
  assign n5221 = n4280 ^ n776 ^ 1'b0 ;
  assign n5222 = n5221 ^ n4373 ^ 1'b0 ;
  assign n5223 = n5220 & ~n5222 ;
  assign n5224 = n3638 ^ n2709 ^ 1'b0 ;
  assign n5225 = n5224 ^ n3919 ^ 1'b0 ;
  assign n5229 = n2882 ^ n2031 ^ 1'b0 ;
  assign n5226 = n1017 ^ x83 ^ 1'b0 ;
  assign n5227 = n5226 ^ n3921 ^ n3104 ;
  assign n5228 = n976 & n5227 ;
  assign n5230 = n5229 ^ n5228 ^ n2287 ;
  assign n5231 = x106 & ~n4463 ;
  assign n5232 = n1766 ^ n718 ^ 1'b0 ;
  assign n5233 = ( ~n441 & n3725 ) | ( ~n441 & n5232 ) | ( n3725 & n5232 ) ;
  assign n5234 = n3881 ^ n583 ^ 1'b0 ;
  assign n5235 = n5233 | n5234 ;
  assign n5240 = ~n562 & n2521 ;
  assign n5241 = n1582 & n5240 ;
  assign n5237 = n267 | n2452 ;
  assign n5238 = n1315 | n5237 ;
  assign n5239 = n668 & n5238 ;
  assign n5242 = n5241 ^ n5239 ^ 1'b0 ;
  assign n5236 = n2871 & n4986 ;
  assign n5243 = n5242 ^ n5236 ^ 1'b0 ;
  assign n5244 = n5243 ^ n4444 ^ n3275 ;
  assign n5245 = n1601 & n1786 ;
  assign n5246 = ~n1284 & n5245 ;
  assign n5247 = n4015 & ~n5246 ;
  assign n5248 = n5247 ^ n4934 ^ n3860 ;
  assign n5249 = x56 & x242 ;
  assign n5250 = ~x124 & n5249 ;
  assign n5251 = n337 | n5250 ;
  assign n5252 = n5251 ^ n2442 ^ 1'b0 ;
  assign n5253 = n4655 ^ n2949 ^ 1'b0 ;
  assign n5254 = n2225 & ~n4846 ;
  assign n5255 = n5254 ^ x16 ^ 1'b0 ;
  assign n5256 = n3050 ^ n2884 ^ n2706 ;
  assign n5257 = ( n1439 & n1453 ) | ( n1439 & n2419 ) | ( n1453 & n2419 ) ;
  assign n5258 = n4597 ^ x94 ^ 1'b0 ;
  assign n5259 = n5257 | n5258 ;
  assign n5262 = ( x152 & n1212 ) | ( x152 & ~n1666 ) | ( n1212 & ~n1666 ) ;
  assign n5263 = n5262 ^ n1142 ^ 1'b0 ;
  assign n5260 = n2315 ^ n428 ^ 1'b0 ;
  assign n5261 = n4898 & n5260 ;
  assign n5264 = n5263 ^ n5261 ^ n5155 ;
  assign n5265 = ~n814 & n5130 ;
  assign n5266 = ~n5264 & n5265 ;
  assign n5267 = n1937 ^ n1274 ^ 1'b0 ;
  assign n5268 = n1730 & n2397 ;
  assign n5269 = n5267 & n5268 ;
  assign n5270 = ~n1136 & n2226 ;
  assign n5271 = n5019 & n5270 ;
  assign n5272 = n2830 & ~n5271 ;
  assign n5273 = n3301 ^ n806 ^ 1'b0 ;
  assign n5274 = n3738 & n5273 ;
  assign n5275 = n5272 & n5274 ;
  assign n5276 = n5275 ^ n5114 ^ 1'b0 ;
  assign n5277 = n3883 ^ n1488 ^ 1'b0 ;
  assign n5278 = n2252 ^ n1943 ^ 1'b0 ;
  assign n5279 = n5278 ^ n2942 ^ 1'b0 ;
  assign n5280 = ~n5177 & n5279 ;
  assign n5281 = n5277 & n5280 ;
  assign n5282 = ( n761 & n4565 ) | ( n761 & n5281 ) | ( n4565 & n5281 ) ;
  assign n5283 = ~n753 & n3801 ;
  assign n5284 = n4450 ^ n3875 ^ 1'b0 ;
  assign n5285 = ~n4210 & n5284 ;
  assign n5286 = n2930 ^ n495 ^ 1'b0 ;
  assign n5287 = x4 & n1295 ;
  assign n5288 = n5287 ^ x52 ^ 1'b0 ;
  assign n5289 = ( ~n648 & n822 ) | ( ~n648 & n5288 ) | ( n822 & n5288 ) ;
  assign n5290 = n5289 ^ n607 ^ 1'b0 ;
  assign n5291 = n4144 & n5290 ;
  assign n5292 = n5291 ^ n2871 ^ 1'b0 ;
  assign n5294 = ( n944 & n2144 ) | ( n944 & ~n2296 ) | ( n2144 & ~n2296 ) ;
  assign n5295 = n3363 | n5294 ;
  assign n5293 = ~x235 & n271 ;
  assign n5296 = n5295 ^ n5293 ^ 1'b0 ;
  assign n5297 = ~n4123 & n4768 ;
  assign n5298 = n5297 ^ n291 ^ 1'b0 ;
  assign n5299 = n2300 ^ n451 ^ 1'b0 ;
  assign n5300 = n4280 | n5299 ;
  assign n5301 = n2632 | n5300 ;
  assign n5302 = n5301 ^ n4982 ^ 1'b0 ;
  assign n5303 = ( x108 & n3308 ) | ( x108 & n5302 ) | ( n3308 & n5302 ) ;
  assign n5304 = n4627 ^ n363 ^ 1'b0 ;
  assign n5305 = x42 & ~n4567 ;
  assign n5306 = n4175 ^ x227 ^ x108 ;
  assign n5307 = n4043 ^ x137 ^ 1'b0 ;
  assign n5308 = n1763 | n5307 ;
  assign n5309 = n5306 & ~n5308 ;
  assign n5310 = n5305 & n5309 ;
  assign n5314 = n2097 ^ n1188 ^ 1'b0 ;
  assign n5311 = ( ~n299 & n579 ) | ( ~n299 & n2169 ) | ( n579 & n2169 ) ;
  assign n5312 = n3508 & n5311 ;
  assign n5313 = ( n1980 & ~n4713 ) | ( n1980 & n5312 ) | ( ~n4713 & n5312 ) ;
  assign n5315 = n5314 ^ n5313 ^ n2261 ;
  assign n5316 = n4812 ^ n2452 ^ 1'b0 ;
  assign n5317 = n5315 & ~n5316 ;
  assign n5318 = n2249 & ~n4876 ;
  assign n5319 = n5318 ^ n2054 ^ 1'b0 ;
  assign n5320 = n982 | n2667 ;
  assign n5321 = n1015 & ~n5320 ;
  assign n5322 = n1021 & n3008 ;
  assign n5323 = n5321 & n5322 ;
  assign n5324 = n5323 ^ n3240 ^ 1'b0 ;
  assign n5325 = ( n337 & n1025 ) | ( n337 & ~n2303 ) | ( n1025 & ~n2303 ) ;
  assign n5326 = n5325 ^ n3283 ^ x210 ;
  assign n5327 = x87 & ~n3043 ;
  assign n5328 = ( ~n438 & n538 ) | ( ~n438 & n5327 ) | ( n538 & n5327 ) ;
  assign n5329 = ~n5326 & n5328 ;
  assign n5331 = x8 & n697 ;
  assign n5332 = ( n429 & n1010 ) | ( n429 & ~n1732 ) | ( n1010 & ~n1732 ) ;
  assign n5333 = n4574 & n5332 ;
  assign n5334 = ~n5247 & n5333 ;
  assign n5335 = n5331 & ~n5334 ;
  assign n5336 = n5335 ^ n2074 ^ 1'b0 ;
  assign n5337 = ~n2055 & n5336 ;
  assign n5338 = n5337 ^ n791 ^ 1'b0 ;
  assign n5330 = n1360 ^ x17 ^ 1'b0 ;
  assign n5339 = n5338 ^ n5330 ^ 1'b0 ;
  assign n5349 = n317 | n418 ;
  assign n5350 = n5349 ^ n376 ^ 1'b0 ;
  assign n5351 = n2465 ^ n1103 ^ 1'b0 ;
  assign n5352 = n5350 | n5351 ;
  assign n5347 = n3000 ^ n472 ^ 1'b0 ;
  assign n5348 = n5347 ^ n1779 ^ n331 ;
  assign n5353 = n5352 ^ n5348 ^ 1'b0 ;
  assign n5354 = ~n2171 & n5353 ;
  assign n5340 = n2017 ^ n956 ^ 1'b0 ;
  assign n5341 = n1323 & n5340 ;
  assign n5342 = n3809 ^ n1951 ^ 1'b0 ;
  assign n5343 = n1499 & ~n5342 ;
  assign n5344 = n3796 | n3860 ;
  assign n5345 = n5343 | n5344 ;
  assign n5346 = n5341 & n5345 ;
  assign n5355 = n5354 ^ n5346 ^ 1'b0 ;
  assign n5356 = n5355 ^ n5055 ^ n1340 ;
  assign n5357 = n3824 & ~n5321 ;
  assign n5358 = n3051 ^ n2722 ^ 1'b0 ;
  assign n5359 = n3995 & n5358 ;
  assign n5360 = n5357 & n5359 ;
  assign n5361 = ~n1478 & n5360 ;
  assign n5362 = n1987 ^ n404 ^ 1'b0 ;
  assign n5363 = ~n1944 & n5362 ;
  assign n5364 = n3791 ^ n3039 ^ 1'b0 ;
  assign n5365 = n1735 | n5364 ;
  assign n5366 = n2029 ^ x187 ^ 1'b0 ;
  assign n5367 = n5366 ^ n3398 ^ 1'b0 ;
  assign n5368 = ~n5365 & n5367 ;
  assign n5369 = n5368 ^ n2054 ^ 1'b0 ;
  assign n5370 = n4806 ^ n3282 ^ 1'b0 ;
  assign n5371 = n3594 ^ n3267 ^ 1'b0 ;
  assign n5372 = x195 & n5371 ;
  assign n5373 = ( x194 & ~n2066 ) | ( x194 & n2702 ) | ( ~n2066 & n2702 ) ;
  assign n5374 = ~n1313 & n5373 ;
  assign n5375 = n1561 & n5374 ;
  assign n5376 = n2369 & ~n5375 ;
  assign n5377 = n2617 ^ n753 ^ 1'b0 ;
  assign n5378 = n2153 & n5377 ;
  assign n5379 = ~n390 & n1059 ;
  assign n5380 = n5378 & n5379 ;
  assign n5381 = n1070 | n3794 ;
  assign n5382 = n1048 & ~n2065 ;
  assign n5383 = n5382 ^ n2023 ^ 1'b0 ;
  assign n5384 = n1969 & n5383 ;
  assign n5385 = ( x179 & ~n5257 ) | ( x179 & n5384 ) | ( ~n5257 & n5384 ) ;
  assign n5386 = n4691 ^ n4112 ^ n543 ;
  assign n5387 = n2719 ^ n1401 ^ 1'b0 ;
  assign n5388 = n2298 ^ n1984 ^ n1574 ;
  assign n5389 = ~n4902 & n5388 ;
  assign n5390 = n2082 ^ x185 ^ 1'b0 ;
  assign n5391 = n5389 & n5390 ;
  assign n5392 = x246 & ~n2673 ;
  assign n5393 = n5392 ^ n4150 ^ 1'b0 ;
  assign n5394 = n755 & n2282 ;
  assign n5395 = n5394 ^ n1376 ^ 1'b0 ;
  assign n5396 = ( n2720 & ~n2932 ) | ( n2720 & n5395 ) | ( ~n2932 & n5395 ) ;
  assign n5397 = n5393 & n5396 ;
  assign n5398 = n1831 & ~n5397 ;
  assign n5399 = n575 | n1145 ;
  assign n5400 = n5399 ^ x24 ^ 1'b0 ;
  assign n5401 = x56 & ~n2002 ;
  assign n5402 = ~n3336 & n5401 ;
  assign n5403 = n790 & ~n3743 ;
  assign n5404 = n2530 & n5403 ;
  assign n5405 = n5393 & ~n5404 ;
  assign n5406 = ~n2285 & n5405 ;
  assign n5407 = n3803 ^ x247 ^ 1'b0 ;
  assign n5408 = n790 & n5407 ;
  assign n5411 = n1695 ^ x95 ^ 1'b0 ;
  assign n5409 = n2178 & ~n4074 ;
  assign n5410 = n3059 & n5409 ;
  assign n5412 = n5411 ^ n5410 ^ 1'b0 ;
  assign n5413 = ( ~n2275 & n3091 ) | ( ~n2275 & n3363 ) | ( n3091 & n3363 ) ;
  assign n5414 = n727 & n3557 ;
  assign n5415 = n3399 & ~n4241 ;
  assign n5416 = n2807 | n5415 ;
  assign n5417 = n5416 ^ n3626 ^ 1'b0 ;
  assign n5420 = ~n1250 & n2382 ;
  assign n5418 = n1188 ^ n840 ^ 1'b0 ;
  assign n5419 = ~n5311 & n5418 ;
  assign n5421 = n5420 ^ n5419 ^ 1'b0 ;
  assign n5422 = ~n727 & n1093 ;
  assign n5423 = ( n1258 & ~n1629 ) | ( n1258 & n2118 ) | ( ~n1629 & n2118 ) ;
  assign n5424 = n5422 & n5423 ;
  assign n5425 = n4170 & n5424 ;
  assign n5426 = n5425 ^ n3752 ^ n1001 ;
  assign n5427 = n1176 | n3523 ;
  assign n5428 = n5427 ^ n1514 ^ 1'b0 ;
  assign n5429 = n5338 ^ n2276 ^ 1'b0 ;
  assign n5430 = ~n5428 & n5429 ;
  assign n5431 = ~n2468 & n3096 ;
  assign n5432 = n4505 ^ n4182 ^ n453 ;
  assign n5433 = n5432 ^ n4817 ^ 1'b0 ;
  assign n5434 = n5433 ^ n2887 ^ 1'b0 ;
  assign n5435 = ~n5431 & n5434 ;
  assign n5436 = n5435 ^ n2107 ^ 1'b0 ;
  assign n5437 = n1372 | n5436 ;
  assign n5438 = n3778 ^ n2341 ^ 1'b0 ;
  assign n5439 = n489 & ~n5438 ;
  assign n5440 = n1829 ^ n445 ^ 1'b0 ;
  assign n5441 = n593 | n5440 ;
  assign n5442 = n3517 & ~n3778 ;
  assign n5443 = n5441 & n5442 ;
  assign n5444 = n3097 & ~n5443 ;
  assign n5445 = n5444 ^ n4296 ^ 1'b0 ;
  assign n5446 = n2026 ^ x141 ^ 1'b0 ;
  assign n5447 = n2276 | n4802 ;
  assign n5448 = n5447 ^ n4458 ^ 1'b0 ;
  assign n5449 = n2450 ^ n539 ^ 1'b0 ;
  assign n5450 = n5027 ^ n4826 ^ 1'b0 ;
  assign n5451 = n2368 & n5450 ;
  assign n5452 = n2023 ^ n1817 ^ n1026 ;
  assign n5453 = n5452 ^ n1987 ^ 1'b0 ;
  assign n5454 = n5453 ^ n455 ^ 1'b0 ;
  assign n5455 = ~n2645 & n5454 ;
  assign n5459 = n1972 ^ n1327 ^ 1'b0 ;
  assign n5460 = x61 & ~n5459 ;
  assign n5456 = n1279 & n4698 ;
  assign n5457 = n5456 ^ n4975 ^ 1'b0 ;
  assign n5458 = n259 & n5457 ;
  assign n5461 = n5460 ^ n5458 ^ 1'b0 ;
  assign n5462 = ( n960 & n2300 ) | ( n960 & ~n3554 ) | ( n2300 & ~n3554 ) ;
  assign n5464 = n4105 ^ n529 ^ n434 ;
  assign n5463 = n2276 ^ n1633 ^ n1182 ;
  assign n5465 = n5464 ^ n5463 ^ 1'b0 ;
  assign n5466 = n3383 | n5465 ;
  assign n5467 = n5466 ^ n3872 ^ 1'b0 ;
  assign n5468 = ( ~n4722 & n5462 ) | ( ~n4722 & n5467 ) | ( n5462 & n5467 ) ;
  assign n5472 = n2004 & ~n2808 ;
  assign n5473 = ~n2218 & n5472 ;
  assign n5474 = ( x130 & ~n2134 ) | ( x130 & n3678 ) | ( ~n2134 & n3678 ) ;
  assign n5475 = ~n5473 & n5474 ;
  assign n5476 = n5475 ^ n3133 ^ 1'b0 ;
  assign n5469 = ( n781 & n2945 ) | ( n781 & ~n3231 ) | ( n2945 & ~n3231 ) ;
  assign n5470 = n443 & ~n4435 ;
  assign n5471 = n5469 & n5470 ;
  assign n5477 = n5476 ^ n5471 ^ n2352 ;
  assign n5478 = n5477 ^ n5001 ^ 1'b0 ;
  assign n5479 = ( n2531 & ~n3723 ) | ( n2531 & n3912 ) | ( ~n3723 & n3912 ) ;
  assign n5480 = ~n721 & n3524 ;
  assign n5481 = ~n360 & n5480 ;
  assign n5482 = x42 | n5481 ;
  assign n5483 = n5482 ^ n3702 ^ 1'b0 ;
  assign n5484 = x67 & n637 ;
  assign n5485 = n5484 ^ n2499 ^ 1'b0 ;
  assign n5486 = n5485 ^ n3495 ^ 1'b0 ;
  assign n5487 = n1955 & n5486 ;
  assign n5489 = n420 & n3008 ;
  assign n5490 = ( ~n3666 & n4104 ) | ( ~n3666 & n5489 ) | ( n4104 & n5489 ) ;
  assign n5488 = x117 & ~n3671 ;
  assign n5491 = n5490 ^ n5488 ^ 1'b0 ;
  assign n5492 = n5491 ^ x211 ^ 1'b0 ;
  assign n5493 = n5487 & n5492 ;
  assign n5494 = n686 ^ x187 ^ 1'b0 ;
  assign n5495 = n1892 & ~n5494 ;
  assign n5496 = n5495 ^ n3436 ^ n299 ;
  assign n5497 = n5496 ^ n3477 ^ n2968 ;
  assign n5498 = x235 | n1917 ;
  assign n5499 = n340 | n5498 ;
  assign n5500 = n3567 ^ n374 ^ 1'b0 ;
  assign n5501 = n538 & n5500 ;
  assign n5502 = n365 | n5298 ;
  assign n5503 = n1773 & n2097 ;
  assign n5504 = ~n1188 & n5503 ;
  assign n5505 = n723 | n4436 ;
  assign n5506 = n333 & ~n5505 ;
  assign n5507 = n3018 ^ n2768 ^ x129 ;
  assign n5508 = n548 ^ n327 ^ 1'b0 ;
  assign n5509 = ( ~n922 & n5507 ) | ( ~n922 & n5508 ) | ( n5507 & n5508 ) ;
  assign n5510 = ( n5339 & n5506 ) | ( n5339 & ~n5509 ) | ( n5506 & ~n5509 ) ;
  assign n5511 = n2527 & ~n5370 ;
  assign n5512 = n3804 ^ n2237 ^ 1'b0 ;
  assign n5513 = n5512 ^ n4829 ^ n3504 ;
  assign n5514 = n5513 ^ n2214 ^ 1'b0 ;
  assign n5515 = n3111 ^ n2774 ^ x134 ;
  assign n5516 = n2703 & n4433 ;
  assign n5517 = n5516 ^ n3556 ^ 1'b0 ;
  assign n5518 = n5515 & ~n5517 ;
  assign n5519 = n3738 ^ n2103 ^ 1'b0 ;
  assign n5520 = n5519 ^ n2218 ^ 1'b0 ;
  assign n5521 = n4093 | n5520 ;
  assign n5522 = ~n3696 & n5521 ;
  assign n5523 = n3825 ^ n2206 ^ 1'b0 ;
  assign n5524 = n2164 & ~n2674 ;
  assign n5525 = n5524 ^ n2746 ^ 1'b0 ;
  assign n5526 = x25 & x84 ;
  assign n5527 = n5526 ^ n2744 ^ 1'b0 ;
  assign n5528 = n5527 ^ n1842 ^ n653 ;
  assign n5529 = n3895 ^ n1847 ^ 1'b0 ;
  assign n5530 = n1151 & ~n4941 ;
  assign n5531 = ~n4274 & n5530 ;
  assign n5533 = ~n2289 & n4281 ;
  assign n5534 = n5533 ^ n2191 ^ 1'b0 ;
  assign n5532 = ( ~n434 & n884 ) | ( ~n434 & n1264 ) | ( n884 & n1264 ) ;
  assign n5535 = n5534 ^ n5532 ^ 1'b0 ;
  assign n5536 = ( n1490 & n1793 ) | ( n1490 & n4860 ) | ( n1793 & n4860 ) ;
  assign n5537 = ( n2772 & n4000 ) | ( n2772 & n4679 ) | ( n4000 & n4679 ) ;
  assign n5539 = ~n1343 & n2519 ;
  assign n5540 = x15 & n5539 ;
  assign n5538 = n2694 ^ n2102 ^ n395 ;
  assign n5541 = n5540 ^ n5538 ^ 1'b0 ;
  assign n5542 = ( x121 & n1209 ) | ( x121 & ~n2028 ) | ( n1209 & ~n2028 ) ;
  assign n5543 = n5542 ^ n626 ^ x59 ;
  assign n5545 = n5115 ^ n1587 ^ 1'b0 ;
  assign n5546 = n265 & n5545 ;
  assign n5544 = x72 & ~n580 ;
  assign n5547 = n5546 ^ n5544 ^ 1'b0 ;
  assign n5548 = n5547 ^ n1033 ^ 1'b0 ;
  assign n5549 = n5543 & n5548 ;
  assign n5550 = n5549 ^ n4772 ^ 1'b0 ;
  assign n5551 = n524 & n3577 ;
  assign n5552 = ~n5550 & n5551 ;
  assign n5553 = n1775 & ~n2040 ;
  assign n5554 = n5553 ^ n4905 ^ 1'b0 ;
  assign n5555 = n5554 ^ n5264 ^ 1'b0 ;
  assign n5556 = n3942 & ~n5555 ;
  assign n5557 = ~n1685 & n4643 ;
  assign n5558 = ~n4168 & n5557 ;
  assign n5559 = x181 & ~n4951 ;
  assign n5560 = ~n259 & n5559 ;
  assign n5565 = n1470 ^ n1125 ^ 1'b0 ;
  assign n5563 = n2164 ^ n1788 ^ 1'b0 ;
  assign n5564 = x108 & ~n5563 ;
  assign n5561 = n3163 ^ n733 ^ 1'b0 ;
  assign n5562 = n3708 & n5561 ;
  assign n5566 = n5565 ^ n5564 ^ n5562 ;
  assign n5567 = n3521 | n5566 ;
  assign n5568 = n1400 & ~n4286 ;
  assign n5569 = ( n1712 & ~n3126 ) | ( n1712 & n5154 ) | ( ~n3126 & n5154 ) ;
  assign n5570 = n2746 ^ n1443 ^ 1'b0 ;
  assign n5571 = n887 & ~n5570 ;
  assign n5572 = n5571 ^ n1228 ^ n634 ;
  assign n5573 = ~n5221 & n5572 ;
  assign n5574 = x153 & n2368 ;
  assign n5575 = n5574 ^ n3557 ^ 1'b0 ;
  assign n5576 = n3728 & n5575 ;
  assign n5577 = ~n2081 & n4677 ;
  assign n5578 = n1575 ^ n610 ^ 1'b0 ;
  assign n5579 = n3485 ^ n3291 ^ n3015 ;
  assign n5580 = ~n822 & n5579 ;
  assign n5581 = n2386 & n5580 ;
  assign n5582 = n4905 ^ n1323 ^ 1'b0 ;
  assign n5583 = ~n418 & n1106 ;
  assign n5584 = n2762 ^ n1941 ^ x97 ;
  assign n5585 = ~n3850 & n5584 ;
  assign n5586 = n2547 & n5585 ;
  assign n5587 = x119 & n4591 ;
  assign n5588 = n5587 ^ x128 ^ 1'b0 ;
  assign n5589 = n5586 & ~n5588 ;
  assign n5590 = n1823 ^ n1081 ^ n538 ;
  assign n5591 = n2699 ^ n1735 ^ 1'b0 ;
  assign n5593 = n3829 ^ n2608 ^ 1'b0 ;
  assign n5594 = x28 & ~n5593 ;
  assign n5592 = n791 & n1266 ;
  assign n5595 = n5594 ^ n5592 ^ 1'b0 ;
  assign n5596 = n5591 & n5595 ;
  assign n5597 = n2188 & n2239 ;
  assign n5598 = n5597 ^ x218 ^ 1'b0 ;
  assign n5599 = x224 & n954 ;
  assign n5600 = ( n690 & n1592 ) | ( n690 & ~n1620 ) | ( n1592 & ~n1620 ) ;
  assign n5601 = n3010 & ~n5600 ;
  assign n5602 = n1048 ^ x140 ^ 1'b0 ;
  assign n5603 = n587 & n5602 ;
  assign n5604 = x20 & n5603 ;
  assign n5605 = n5604 ^ n1473 ^ 1'b0 ;
  assign n5606 = n5051 | n5605 ;
  assign n5607 = n5606 ^ n3548 ^ 1'b0 ;
  assign n5608 = n1425 ^ n1374 ^ 1'b0 ;
  assign n5612 = ~n2257 & n2797 ;
  assign n5613 = ~n671 & n5612 ;
  assign n5611 = n557 | n1258 ;
  assign n5614 = n5613 ^ n5611 ^ 1'b0 ;
  assign n5615 = n2801 & n2925 ;
  assign n5616 = n5614 & n5615 ;
  assign n5609 = n1558 ^ n572 ^ 1'b0 ;
  assign n5610 = ~n4033 & n5609 ;
  assign n5617 = n5616 ^ n5610 ^ x22 ;
  assign n5618 = n4294 ^ n3493 ^ 1'b0 ;
  assign n5619 = ~n3564 & n4887 ;
  assign n5620 = n2019 & n5619 ;
  assign n5621 = n2155 ^ n948 ^ 1'b0 ;
  assign n5622 = ~n1208 & n1527 ;
  assign n5623 = n5622 ^ n813 ^ 1'b0 ;
  assign n5629 = x22 & ~n1235 ;
  assign n5624 = n3406 ^ n1382 ^ 1'b0 ;
  assign n5625 = n5366 ^ n1577 ^ 1'b0 ;
  assign n5626 = ~n5624 & n5625 ;
  assign n5627 = n5626 ^ n1882 ^ 1'b0 ;
  assign n5628 = n1940 & ~n5627 ;
  assign n5630 = n5629 ^ n5628 ^ n2445 ;
  assign n5631 = ~n3712 & n5630 ;
  assign n5632 = n5631 ^ n3949 ^ 1'b0 ;
  assign n5633 = n5632 ^ n4373 ^ 1'b0 ;
  assign n5634 = n2838 | n5633 ;
  assign n5635 = ( n1691 & n2797 ) | ( n1691 & ~n5634 ) | ( n2797 & ~n5634 ) ;
  assign n5636 = ( n3806 & n5623 ) | ( n3806 & ~n5635 ) | ( n5623 & ~n5635 ) ;
  assign n5637 = n580 & n1779 ;
  assign n5638 = n1726 ^ n1122 ^ 1'b0 ;
  assign n5639 = n1218 & n2582 ;
  assign n5640 = x133 & n401 ;
  assign n5641 = n5640 ^ n751 ^ 1'b0 ;
  assign n5642 = n5641 ^ n5517 ^ 1'b0 ;
  assign n5643 = n2371 & ~n5642 ;
  assign n5644 = n4047 ^ n281 ^ 1'b0 ;
  assign n5645 = n5644 ^ n3518 ^ n1527 ;
  assign n5646 = n5645 ^ n3875 ^ n3501 ;
  assign n5647 = n5646 ^ n3911 ^ 1'b0 ;
  assign n5648 = n2973 & n3453 ;
  assign n5649 = n571 & ~n4644 ;
  assign n5650 = n2640 | n2991 ;
  assign n5651 = n3429 ^ n815 ^ 1'b0 ;
  assign n5652 = x140 & n5651 ;
  assign n5653 = ~n1894 & n5652 ;
  assign n5654 = n5653 ^ x30 ^ 1'b0 ;
  assign n5655 = n5650 & n5654 ;
  assign n5658 = n1920 ^ n1622 ^ n744 ;
  assign n5656 = n4405 ^ n411 ^ 1'b0 ;
  assign n5657 = n5656 ^ n567 ^ n413 ;
  assign n5659 = n5658 ^ n5657 ^ 1'b0 ;
  assign n5660 = n2942 & ~n5659 ;
  assign n5661 = x83 & ~n3373 ;
  assign n5662 = n5661 ^ n2054 ^ 1'b0 ;
  assign n5663 = x115 & n5662 ;
  assign n5664 = x139 & n2993 ;
  assign n5665 = ~x209 & n5664 ;
  assign n5666 = n5663 & ~n5665 ;
  assign n5667 = ( ~n3705 & n5469 ) | ( ~n3705 & n5666 ) | ( n5469 & n5666 ) ;
  assign n5668 = n3731 ^ n1929 ^ n1007 ;
  assign n5669 = n5668 ^ n1960 ^ n273 ;
  assign n5670 = n2998 & n3210 ;
  assign n5671 = n5670 ^ n2600 ^ x32 ;
  assign n5672 = n5671 ^ n785 ^ 1'b0 ;
  assign n5673 = n5522 ^ n2893 ^ x76 ;
  assign n5674 = n4830 ^ n4323 ^ n2692 ;
  assign n5675 = ( n2059 & n2689 ) | ( n2059 & n4538 ) | ( n2689 & n4538 ) ;
  assign n5676 = n5675 ^ n1344 ^ 1'b0 ;
  assign n5677 = n3716 ^ x231 ^ 1'b0 ;
  assign n5678 = n5031 ^ n3244 ^ 1'b0 ;
  assign n5679 = ~n319 & n643 ;
  assign n5680 = n1390 & n5679 ;
  assign n5681 = n5187 ^ n4540 ^ 1'b0 ;
  assign n5682 = n1996 | n2910 ;
  assign n5683 = n5682 ^ n2942 ^ 1'b0 ;
  assign n5684 = n2536 & n3690 ;
  assign n5685 = n5684 ^ n5414 ^ n3523 ;
  assign n5686 = n427 & n3228 ;
  assign n5687 = n5686 ^ n4541 ^ 1'b0 ;
  assign n5688 = n1484 & ~n5687 ;
  assign n5689 = ( n1148 & n1266 ) | ( n1148 & ~n2224 ) | ( n1266 & ~n2224 ) ;
  assign n5690 = n5689 ^ n2669 ^ 1'b0 ;
  assign n5691 = n3611 & ~n4145 ;
  assign n5692 = n4215 | n4469 ;
  assign n5693 = n2481 & ~n5692 ;
  assign n5694 = x57 | n308 ;
  assign n5695 = ( n380 & ~n1639 ) | ( n380 & n5694 ) | ( ~n1639 & n5694 ) ;
  assign n5696 = n2156 | n5695 ;
  assign n5697 = n548 & ~n5696 ;
  assign n5698 = ~n5693 & n5697 ;
  assign n5699 = ~n549 & n5008 ;
  assign n5700 = ~n3770 & n3926 ;
  assign n5701 = n5700 ^ n536 ^ 1'b0 ;
  assign n5702 = n877 | n1976 ;
  assign n5703 = n3547 | n5702 ;
  assign n5704 = n817 & n2612 ;
  assign n5705 = ~n2957 & n5704 ;
  assign n5706 = n1698 | n2199 ;
  assign n5707 = n5706 ^ n1073 ^ 1'b0 ;
  assign n5708 = n4207 ^ n3096 ^ 1'b0 ;
  assign n5709 = n5708 ^ n865 ^ 1'b0 ;
  assign n5710 = n5707 | n5709 ;
  assign n5711 = x46 & n863 ;
  assign n5713 = n1701 ^ n1106 ^ 1'b0 ;
  assign n5712 = n3430 & n4833 ;
  assign n5714 = n5713 ^ n5712 ^ 1'b0 ;
  assign n5715 = n5538 & n5714 ;
  assign n5716 = n5711 & n5715 ;
  assign n5717 = n1098 ^ x93 ^ 1'b0 ;
  assign n5718 = n4657 & ~n5717 ;
  assign n5719 = x176 & ~n3804 ;
  assign n5720 = n5719 ^ n2903 ^ n1766 ;
  assign n5721 = n1970 & ~n2651 ;
  assign n5722 = n2506 ^ x150 ^ 1'b0 ;
  assign n5723 = n1881 & ~n4679 ;
  assign n5724 = n5723 ^ n2091 ^ 1'b0 ;
  assign n5725 = n502 & ~n5724 ;
  assign n5726 = n5722 | n5725 ;
  assign n5727 = n1196 & n2959 ;
  assign n5728 = n2125 & n5727 ;
  assign n5732 = n1140 & n2660 ;
  assign n5733 = n5732 ^ n433 ^ 1'b0 ;
  assign n5734 = n5733 ^ n1604 ^ 1'b0 ;
  assign n5735 = n2363 & ~n5734 ;
  assign n5729 = x114 & n1190 ;
  assign n5730 = n5366 & ~n5729 ;
  assign n5731 = n2073 | n5730 ;
  assign n5736 = n5735 ^ n5731 ^ 1'b0 ;
  assign n5737 = n5736 ^ n2635 ^ 1'b0 ;
  assign n5738 = n5728 | n5737 ;
  assign n5739 = n3021 ^ n2174 ^ n2057 ;
  assign n5740 = n5739 ^ n2350 ^ 1'b0 ;
  assign n5741 = n5740 ^ n4580 ^ x33 ;
  assign n5742 = n1855 & n3852 ;
  assign n5743 = n650 | n4436 ;
  assign n5744 = n5743 ^ n458 ^ 1'b0 ;
  assign n5745 = n1761 | n5744 ;
  assign n5746 = n5745 ^ n456 ^ 1'b0 ;
  assign n5747 = n3782 ^ n655 ^ 1'b0 ;
  assign n5748 = n3782 & ~n5747 ;
  assign n5749 = n5748 ^ n887 ^ 1'b0 ;
  assign n5750 = n5746 & n5749 ;
  assign n5751 = n3245 ^ n2387 ^ 1'b0 ;
  assign n5752 = n2397 ^ n2286 ^ 1'b0 ;
  assign n5753 = x109 & ~n4388 ;
  assign n5754 = n5753 ^ n1648 ^ 1'b0 ;
  assign n5755 = n5754 ^ n4192 ^ x80 ;
  assign n5756 = n1225 | n2549 ;
  assign n5757 = n5756 ^ n2653 ^ 1'b0 ;
  assign n5758 = ( x225 & ~n1272 ) | ( x225 & n5757 ) | ( ~n1272 & n5757 ) ;
  assign n5759 = ( n1789 & n3590 ) | ( n1789 & ~n5758 ) | ( n3590 & ~n5758 ) ;
  assign n5760 = ( ~n286 & n635 ) | ( ~n286 & n3036 ) | ( n635 & n3036 ) ;
  assign n5761 = n2454 | n2711 ;
  assign n5762 = n2061 & ~n5761 ;
  assign n5763 = ( ~x62 & n1140 ) | ( ~x62 & n1925 ) | ( n1140 & n1925 ) ;
  assign n5764 = n2749 & n5763 ;
  assign n5765 = n5762 & n5764 ;
  assign n5766 = x195 & n3270 ;
  assign n5767 = ~n5765 & n5766 ;
  assign n5768 = n3894 ^ n3847 ^ 1'b0 ;
  assign n5769 = n1574 ^ n1256 ^ 1'b0 ;
  assign n5770 = n5769 ^ n529 ^ 1'b0 ;
  assign n5771 = n5770 ^ n2888 ^ 1'b0 ;
  assign n5772 = n4807 | n5771 ;
  assign n5773 = n4481 ^ n2530 ^ 1'b0 ;
  assign n5774 = n5042 ^ n997 ^ 1'b0 ;
  assign n5775 = n5772 | n5774 ;
  assign n5776 = n1358 ^ n979 ^ 1'b0 ;
  assign n5777 = n815 | n5776 ;
  assign n5778 = n5777 ^ x22 ^ 1'b0 ;
  assign n5783 = n2524 | n4124 ;
  assign n5784 = n2539 & n5783 ;
  assign n5785 = n5784 ^ n3625 ^ 1'b0 ;
  assign n5779 = n3135 ^ n3098 ^ 1'b0 ;
  assign n5780 = n513 & ~n5779 ;
  assign n5781 = ~n802 & n5780 ;
  assign n5782 = n4807 & n5781 ;
  assign n5786 = n5785 ^ n5782 ^ 1'b0 ;
  assign n5787 = ~n1442 & n4031 ;
  assign n5788 = n1514 & n5787 ;
  assign n5789 = n3779 | n4772 ;
  assign n5790 = n3335 & ~n5789 ;
  assign n5791 = ( n3912 & n4460 ) | ( n3912 & ~n5790 ) | ( n4460 & ~n5790 ) ;
  assign n5792 = ~n802 & n3940 ;
  assign n5793 = n4622 & n5792 ;
  assign n5794 = n2968 | n3530 ;
  assign n5795 = n2413 | n5794 ;
  assign n5796 = n1064 | n3958 ;
  assign n5797 = n5589 & ~n5796 ;
  assign n5798 = n917 | n1166 ;
  assign n5799 = n558 & n2954 ;
  assign n5800 = ( n2080 & ~n4644 ) | ( n2080 & n5799 ) | ( ~n4644 & n5799 ) ;
  assign n5801 = n922 & ~n4029 ;
  assign n5802 = n3756 ^ n3720 ^ 1'b0 ;
  assign n5803 = n3150 ^ x227 ^ 1'b0 ;
  assign n5804 = n2324 & ~n5803 ;
  assign n5805 = n5804 ^ n1677 ^ x110 ;
  assign n5806 = n3227 | n5805 ;
  assign n5807 = n5250 ^ n3310 ^ n1269 ;
  assign n5808 = n607 & ~n3837 ;
  assign n5809 = ~n5807 & n5808 ;
  assign n5810 = n2773 & n4126 ;
  assign n5811 = n5810 ^ n4557 ^ 1'b0 ;
  assign n5812 = ( n1453 & ~n5809 ) | ( n1453 & n5811 ) | ( ~n5809 & n5811 ) ;
  assign n5813 = n2543 | n3085 ;
  assign n5814 = n3909 & ~n5019 ;
  assign n5815 = ~n405 & n1610 ;
  assign n5816 = n5815 ^ n3978 ^ 1'b0 ;
  assign n5817 = n915 & ~n5816 ;
  assign n5818 = n5817 ^ n4748 ^ 1'b0 ;
  assign n5819 = ~n3359 & n3485 ;
  assign n5820 = n683 & n5819 ;
  assign n5821 = n4509 ^ n1376 ^ 1'b0 ;
  assign n5822 = ~n3434 & n5821 ;
  assign n5823 = ~n2885 & n5822 ;
  assign n5824 = n1811 & n5823 ;
  assign n5825 = ~n677 & n5546 ;
  assign n5826 = n5825 ^ n3413 ^ 1'b0 ;
  assign n5827 = ~n4280 & n4405 ;
  assign n5828 = n5827 ^ n3296 ^ 1'b0 ;
  assign n5829 = ( ~n4579 & n5531 ) | ( ~n4579 & n5828 ) | ( n5531 & n5828 ) ;
  assign n5830 = n5829 ^ n5491 ^ 1'b0 ;
  assign n5831 = n1980 ^ n1571 ^ 1'b0 ;
  assign n5832 = ~n840 & n5831 ;
  assign n5833 = ( n3233 & n3708 ) | ( n3233 & ~n3854 ) | ( n3708 & ~n3854 ) ;
  assign n5834 = n1373 | n2100 ;
  assign n5835 = n5605 ^ n2945 ^ x15 ;
  assign n5836 = n5835 ^ n1084 ^ 1'b0 ;
  assign n5837 = n4509 ^ n331 ^ 1'b0 ;
  assign n5838 = x159 & ~n326 ;
  assign n5839 = ( n5836 & ~n5837 ) | ( n5836 & n5838 ) | ( ~n5837 & n5838 ) ;
  assign n5840 = n5670 ^ n3708 ^ 1'b0 ;
  assign n5841 = n4099 ^ n3000 ^ 1'b0 ;
  assign n5842 = n2366 ^ n1234 ^ 1'b0 ;
  assign n5843 = ~n2402 & n5842 ;
  assign n5844 = ~n1639 & n5843 ;
  assign n5845 = n5283 | n5844 ;
  assign n5846 = n5845 ^ x222 ^ 1'b0 ;
  assign n5847 = n4996 ^ n4984 ^ 1'b0 ;
  assign n5848 = n972 | n5847 ;
  assign n5849 = ~n548 & n5848 ;
  assign n5850 = ~n3018 & n3122 ;
  assign n5851 = ( ~n1203 & n2127 ) | ( ~n1203 & n5850 ) | ( n2127 & n5850 ) ;
  assign n5852 = n1932 ^ n1907 ^ 1'b0 ;
  assign n5853 = n2777 ^ n946 ^ 1'b0 ;
  assign n5854 = n5853 ^ n4267 ^ 1'b0 ;
  assign n5855 = n3256 | n5854 ;
  assign n5863 = n815 | n2733 ;
  assign n5864 = x106 | n5863 ;
  assign n5856 = n296 | n1258 ;
  assign n5857 = n5856 ^ n772 ^ 1'b0 ;
  assign n5858 = ( x55 & ~n1213 ) | ( x55 & n5857 ) | ( ~n1213 & n5857 ) ;
  assign n5859 = ( n2685 & n5042 ) | ( n2685 & ~n5858 ) | ( n5042 & ~n5858 ) ;
  assign n5860 = n4339 | n5859 ;
  assign n5861 = n5860 ^ n1044 ^ 1'b0 ;
  assign n5862 = ~n681 & n5861 ;
  assign n5865 = n5864 ^ n5862 ^ 1'b0 ;
  assign n5866 = n1567 & ~n4158 ;
  assign n5867 = n4168 & n4434 ;
  assign n5868 = n690 & n5867 ;
  assign n5869 = ~n4128 & n4300 ;
  assign n5870 = n3311 & ~n4435 ;
  assign n5871 = n2488 & n3825 ;
  assign n5872 = n5871 ^ n2613 ^ 1'b0 ;
  assign n5873 = n4524 & n5872 ;
  assign n5874 = n982 & n5873 ;
  assign n5875 = n1762 & ~n1769 ;
  assign n5876 = ( n3884 & ~n4404 ) | ( n3884 & n5875 ) | ( ~n4404 & n5875 ) ;
  assign n5877 = ( ~n963 & n1177 ) | ( ~n963 & n1409 ) | ( n1177 & n1409 ) ;
  assign n5878 = n737 & n5877 ;
  assign n5879 = n5878 ^ n4157 ^ 1'b0 ;
  assign n5880 = ( n924 & n2905 ) | ( n924 & ~n5660 ) | ( n2905 & ~n5660 ) ;
  assign n5881 = n1585 | n5880 ;
  assign n5882 = n3686 | n5881 ;
  assign n5883 = n5879 & n5882 ;
  assign n5884 = n5698 & n5883 ;
  assign n5885 = n460 & n854 ;
  assign n5886 = n942 | n5885 ;
  assign n5887 = n5886 ^ n1735 ^ 1'b0 ;
  assign n5888 = n5887 ^ n3084 ^ n2437 ;
  assign n5889 = n2915 ^ n1427 ^ 1'b0 ;
  assign n5890 = n2807 | n5889 ;
  assign n5891 = n2344 & n5780 ;
  assign n5892 = n5891 ^ n2395 ^ 1'b0 ;
  assign n5893 = n4764 & n5892 ;
  assign n5894 = n5579 & n5893 ;
  assign n5895 = n5890 & n5894 ;
  assign n5896 = ( n924 & ~n1085 ) | ( n924 & n2884 ) | ( ~n1085 & n2884 ) ;
  assign n5897 = n1000 & n5896 ;
  assign n5898 = ~n4839 & n5897 ;
  assign n5899 = n5898 ^ n1209 ^ 1'b0 ;
  assign n5900 = n4792 ^ n548 ^ 1'b0 ;
  assign n5901 = n4593 & ~n5900 ;
  assign n5902 = n4428 & n5040 ;
  assign n5903 = n5902 ^ n3043 ^ 1'b0 ;
  assign n5904 = n314 & ~n5903 ;
  assign n5905 = n1830 & n5904 ;
  assign n5906 = ~n3811 & n4870 ;
  assign n5907 = n5906 ^ x29 ^ 1'b0 ;
  assign n5908 = n471 & ~n5907 ;
  assign n5909 = n5905 & n5908 ;
  assign n5910 = ~n420 & n3782 ;
  assign n5911 = n444 | n1227 ;
  assign n5912 = n1709 | n5911 ;
  assign n5913 = n1725 & n5912 ;
  assign n5914 = n5913 ^ x61 ^ 1'b0 ;
  assign n5915 = n1340 | n5914 ;
  assign n5916 = n5915 ^ n2052 ^ 1'b0 ;
  assign n5917 = n2943 & n4317 ;
  assign n5918 = ~x224 & n5917 ;
  assign n5919 = n5673 ^ n3325 ^ 1'b0 ;
  assign n5920 = x82 & ~n5919 ;
  assign n5921 = n3646 | n4753 ;
  assign n5922 = n2991 ^ n1404 ^ n1308 ;
  assign n5923 = n5922 ^ n4234 ^ n3254 ;
  assign n5924 = ~n1795 & n3895 ;
  assign n5925 = n4173 | n5797 ;
  assign n5926 = n5924 & ~n5925 ;
  assign n5927 = n4378 ^ n2527 ^ 1'b0 ;
  assign n5928 = n5840 ^ x58 ^ 1'b0 ;
  assign n5929 = ~n1650 & n5928 ;
  assign n5930 = n4395 ^ x12 ^ 1'b0 ;
  assign n5931 = n5930 ^ n2941 ^ n2298 ;
  assign n5932 = n4761 ^ n1919 ^ n673 ;
  assign n5933 = n2615 ^ x221 ^ 1'b0 ;
  assign n5934 = n5932 & ~n5933 ;
  assign n5935 = n3556 & n5934 ;
  assign n5936 = ~n5934 & n5935 ;
  assign n5937 = n2276 | n5936 ;
  assign n5938 = n2895 & ~n3251 ;
  assign n5939 = n5938 ^ n5769 ^ 1'b0 ;
  assign n5940 = n5937 & n5939 ;
  assign n5941 = ~n5931 & n5940 ;
  assign n5942 = n2113 ^ n826 ^ 1'b0 ;
  assign n5943 = n5942 ^ n5170 ^ n4593 ;
  assign n5944 = n2374 ^ n1782 ^ 1'b0 ;
  assign n5945 = n5944 ^ n4976 ^ n4726 ;
  assign n5951 = n2452 ^ x229 ^ 1'b0 ;
  assign n5952 = n1924 | n5951 ;
  assign n5947 = ~n1766 & n2519 ;
  assign n5948 = n4373 ^ n1328 ^ 1'b0 ;
  assign n5949 = n3760 | n5948 ;
  assign n5950 = n5947 & ~n5949 ;
  assign n5953 = n5952 ^ n5950 ^ 1'b0 ;
  assign n5946 = n4252 ^ n2224 ^ n2068 ;
  assign n5954 = n5953 ^ n5946 ^ n5312 ;
  assign n5955 = n2781 | n3958 ;
  assign n5956 = n5955 ^ n2454 ^ 1'b0 ;
  assign n5957 = n3712 ^ n1944 ^ 1'b0 ;
  assign n5958 = ~n3312 & n5957 ;
  assign n5959 = ~n4912 & n5958 ;
  assign n5960 = n5959 ^ n5521 ^ 1'b0 ;
  assign n5961 = ( n1197 & n1247 ) | ( n1197 & ~n3562 ) | ( n1247 & ~n3562 ) ;
  assign n5962 = n2463 | n5961 ;
  assign n5963 = ( n2362 & ~n4000 ) | ( n2362 & n5962 ) | ( ~n4000 & n5962 ) ;
  assign n5964 = n3826 ^ n1037 ^ 1'b0 ;
  assign n5965 = n2517 & ~n5964 ;
  assign n5966 = n5568 ^ n5354 ^ 1'b0 ;
  assign n5967 = n789 ^ n758 ^ n642 ;
  assign n5968 = n1730 | n4320 ;
  assign n5969 = n5968 ^ n892 ^ 1'b0 ;
  assign n5970 = x254 & ~n5969 ;
  assign n5971 = n5967 & ~n5970 ;
  assign n5972 = n338 & n3770 ;
  assign n5973 = ( ~n562 & n5224 ) | ( ~n562 & n5972 ) | ( n5224 & n5972 ) ;
  assign n5974 = n2681 ^ n1665 ^ 1'b0 ;
  assign n5975 = ~n2656 & n3761 ;
  assign n5976 = n5975 ^ n4742 ^ n4137 ;
  assign n5977 = n4867 ^ n3958 ^ n1266 ;
  assign n5978 = n5977 ^ n4470 ^ 1'b0 ;
  assign n5980 = n1842 ^ n1630 ^ 1'b0 ;
  assign n5979 = n1932 | n2941 ;
  assign n5981 = n5980 ^ n5979 ^ 1'b0 ;
  assign n5982 = n3122 ^ n2499 ^ n800 ;
  assign n5983 = x103 & ~n387 ;
  assign n5984 = n5982 & n5983 ;
  assign n5985 = ( n2073 & n4774 ) | ( n2073 & n5332 ) | ( n4774 & n5332 ) ;
  assign n5986 = n4462 ^ n600 ^ n449 ;
  assign n5987 = n5986 ^ n2454 ^ x237 ;
  assign n5988 = n1833 | n5987 ;
  assign n5989 = n1278 ^ x207 ^ 1'b0 ;
  assign n5990 = n3333 ^ n3094 ^ 1'b0 ;
  assign n5991 = n3770 | n5990 ;
  assign n5997 = n2768 ^ x244 ^ x224 ;
  assign n5992 = n1838 ^ n1590 ^ x227 ;
  assign n5993 = ( n347 & n1571 ) | ( n347 & n1590 ) | ( n1571 & n1590 ) ;
  assign n5994 = n5993 ^ n4787 ^ n3332 ;
  assign n5995 = n1075 & n5994 ;
  assign n5996 = n5992 & n5995 ;
  assign n5998 = n5997 ^ n5996 ^ 1'b0 ;
  assign n5999 = ~n5991 & n5998 ;
  assign n6001 = ~n1695 & n2404 ;
  assign n6000 = ~n1878 & n2989 ;
  assign n6002 = n6001 ^ n6000 ^ 1'b0 ;
  assign n6003 = n3097 & ~n6002 ;
  assign n6004 = n1863 ^ n1692 ^ 1'b0 ;
  assign n6005 = x243 & ~n6004 ;
  assign n6006 = n599 & ~n5246 ;
  assign n6007 = n2555 & n6006 ;
  assign n6008 = n3678 | n6007 ;
  assign n6009 = n6005 | n6008 ;
  assign n6010 = n4016 & n6009 ;
  assign n6011 = n6010 ^ n5383 ^ 1'b0 ;
  assign n6012 = n6011 ^ n5584 ^ n486 ;
  assign n6013 = ~n2132 & n2775 ;
  assign n6017 = x213 & n2294 ;
  assign n6018 = ~n853 & n6017 ;
  assign n6019 = x153 | n6018 ;
  assign n6014 = n1113 & n3270 ;
  assign n6015 = n3395 & n6014 ;
  assign n6016 = n2680 | n6015 ;
  assign n6020 = n6019 ^ n6016 ^ 1'b0 ;
  assign n6021 = n6013 & n6020 ;
  assign n6022 = n2751 & ~n3617 ;
  assign n6023 = ( n2709 & ~n5513 ) | ( n2709 & n6022 ) | ( ~n5513 & n6022 ) ;
  assign n6024 = n4774 & ~n6023 ;
  assign n6025 = ~n3912 & n6024 ;
  assign n6026 = n1877 | n2194 ;
  assign n6027 = n6026 ^ n5399 ^ 1'b0 ;
  assign n6028 = n6027 ^ n1687 ^ 1'b0 ;
  assign n6029 = ( n4242 & n5711 ) | ( n4242 & ~n6028 ) | ( n5711 & ~n6028 ) ;
  assign n6030 = n3540 & ~n6029 ;
  assign n6031 = x202 & n543 ;
  assign n6032 = n4836 & ~n5813 ;
  assign n6033 = ~n6031 & n6032 ;
  assign n6034 = n2399 & ~n3524 ;
  assign n6035 = n2017 ^ n693 ^ 1'b0 ;
  assign n6036 = x101 & n4281 ;
  assign n6037 = n5672 ^ n3034 ^ 1'b0 ;
  assign n6038 = n6036 & ~n6037 ;
  assign n6041 = n2271 ^ n2071 ^ 1'b0 ;
  assign n6039 = n1105 | n1526 ;
  assign n6040 = n423 & ~n6039 ;
  assign n6042 = n6041 ^ n6040 ^ 1'b0 ;
  assign n6043 = n4496 ^ n319 ^ 1'b0 ;
  assign n6044 = n3953 & ~n6043 ;
  assign n6052 = n1223 & n3148 ;
  assign n6053 = n6052 ^ n2608 ^ 1'b0 ;
  assign n6045 = n509 | n1000 ;
  assign n6046 = n743 | n6045 ;
  assign n6047 = n6046 ^ n447 ^ 1'b0 ;
  assign n6048 = x137 & n6047 ;
  assign n6049 = n6048 ^ n2372 ^ 1'b0 ;
  assign n6050 = n6049 ^ n5687 ^ 1'b0 ;
  assign n6051 = n4544 & n6050 ;
  assign n6054 = n6053 ^ n6051 ^ 1'b0 ;
  assign n6056 = n1498 & n4245 ;
  assign n6057 = n6056 ^ n3908 ^ 1'b0 ;
  assign n6055 = n4662 & ~n5155 ;
  assign n6058 = n6057 ^ n6055 ^ 1'b0 ;
  assign n6059 = x36 & n5676 ;
  assign n6060 = n6059 ^ n3271 ^ 1'b0 ;
  assign n6061 = ~n3002 & n3138 ;
  assign n6062 = n1806 | n3751 ;
  assign n6063 = n6062 ^ n2585 ^ 1'b0 ;
  assign n6064 = n4670 ^ n1943 ^ 1'b0 ;
  assign n6065 = n4881 ^ n2907 ^ 1'b0 ;
  assign n6066 = n743 | n6065 ;
  assign n6070 = n740 & ~n4743 ;
  assign n6071 = n5370 & n6070 ;
  assign n6067 = n4476 ^ n1707 ^ 1'b0 ;
  assign n6068 = n4016 & n6067 ;
  assign n6069 = n2165 & n6068 ;
  assign n6072 = n6071 ^ n6069 ^ 1'b0 ;
  assign n6073 = n1311 & n3305 ;
  assign n6074 = n6073 ^ n3399 ^ 1'b0 ;
  assign n6075 = n2093 ^ x252 ^ 1'b0 ;
  assign n6076 = n6075 ^ n3115 ^ 1'b0 ;
  assign n6077 = n2918 & ~n6076 ;
  assign n6078 = n317 | n2502 ;
  assign n6079 = x170 | n6078 ;
  assign n6080 = n1053 ^ n306 ^ 1'b0 ;
  assign n6081 = n3489 & ~n6080 ;
  assign n6082 = ( n4355 & ~n6079 ) | ( n4355 & n6081 ) | ( ~n6079 & n6081 ) ;
  assign n6083 = n6077 & n6082 ;
  assign n6084 = n6083 ^ n3293 ^ 1'b0 ;
  assign n6085 = ( n1795 & n2156 ) | ( n1795 & n2250 ) | ( n2156 & n2250 ) ;
  assign n6086 = x200 & ~n1005 ;
  assign n6087 = n6086 ^ n3557 ^ 1'b0 ;
  assign n6088 = n5150 & ~n6087 ;
  assign n6089 = ~n1160 & n4718 ;
  assign n6090 = n5757 | n6089 ;
  assign n6091 = n3439 | n6090 ;
  assign n6092 = ~n2080 & n3642 ;
  assign n6093 = n2275 ^ n1196 ^ 1'b0 ;
  assign n6094 = n6093 ^ n5641 ^ 1'b0 ;
  assign n6095 = n1518 & n6094 ;
  assign n6096 = n6095 ^ n2959 ^ 1'b0 ;
  assign n6097 = x89 ^ x12 ^ 1'b0 ;
  assign n6098 = ~n2732 & n6097 ;
  assign n6099 = x39 & n6098 ;
  assign n6100 = n6099 ^ n4703 ^ 1'b0 ;
  assign n6101 = n1833 & n6100 ;
  assign n6102 = n805 & ~n1370 ;
  assign n6103 = n1259 & n6102 ;
  assign n6104 = n1158 & ~n5226 ;
  assign n6105 = n6104 ^ n2423 ^ 1'b0 ;
  assign n6106 = n6105 ^ n924 ^ 1'b0 ;
  assign n6107 = n4913 & ~n6106 ;
  assign n6108 = n2130 ^ x178 ^ 1'b0 ;
  assign n6109 = n4505 ^ n2216 ^ 1'b0 ;
  assign n6110 = n6108 | n6109 ;
  assign n6111 = ~n5635 & n6110 ;
  assign n6112 = n6111 ^ n2982 ^ 1'b0 ;
  assign n6113 = n6112 ^ n2881 ^ 1'b0 ;
  assign n6114 = n6107 & n6113 ;
  assign n6115 = n4819 ^ n2929 ^ 1'b0 ;
  assign n6116 = ~n711 & n918 ;
  assign n6117 = n1404 & n6116 ;
  assign n6118 = n3942 & ~n6117 ;
  assign n6119 = n2158 & n6118 ;
  assign n6120 = n6119 ^ n3229 ^ 1'b0 ;
  assign n6121 = n6115 | n6120 ;
  assign n6122 = n3946 | n5410 ;
  assign n6123 = n947 & ~n1349 ;
  assign n6124 = n1582 & n2975 ;
  assign n6125 = x42 & n2701 ;
  assign n6126 = n365 & n6125 ;
  assign n6127 = ~n6124 & n6126 ;
  assign n6128 = n552 | n2302 ;
  assign n6129 = ~n2055 & n6128 ;
  assign n6130 = ~n1624 & n1677 ;
  assign n6131 = n6130 ^ n5336 ^ 1'b0 ;
  assign n6132 = ~n2493 & n4361 ;
  assign n6133 = n6132 ^ n2895 ^ 1'b0 ;
  assign n6134 = n3015 & ~n6133 ;
  assign n6135 = n729 | n4278 ;
  assign n6136 = n6135 ^ n2995 ^ 1'b0 ;
  assign n6137 = n5629 & ~n6136 ;
  assign n6138 = n3919 & n6137 ;
  assign n6139 = n6138 ^ n3659 ^ n429 ;
  assign n6140 = n1024 & ~n4746 ;
  assign n6141 = n5872 & ~n6140 ;
  assign n6144 = n960 & ~n3316 ;
  assign n6145 = n2036 & n6144 ;
  assign n6142 = n2525 | n5289 ;
  assign n6143 = ~n774 & n6142 ;
  assign n6146 = n6145 ^ n6143 ^ 1'b0 ;
  assign n6147 = n677 & n1070 ;
  assign n6148 = n6147 ^ n4139 ^ 1'b0 ;
  assign n6149 = n2462 | n6148 ;
  assign n6150 = n2532 ^ n1015 ^ n363 ;
  assign n6151 = n2057 ^ n472 ^ 1'b0 ;
  assign n6152 = ~n1481 & n1992 ;
  assign n6153 = n1600 & ~n3147 ;
  assign n6154 = n2504 | n6153 ;
  assign n6155 = n5610 | n6154 ;
  assign n6156 = n4580 | n6155 ;
  assign n6157 = n6152 | n6156 ;
  assign n6158 = n6151 | n6157 ;
  assign n6159 = ( ~x42 & n774 ) | ( ~x42 & n3783 ) | ( n774 & n3783 ) ;
  assign n6160 = n3554 ^ n2002 ^ 1'b0 ;
  assign n6161 = ~n6159 & n6160 ;
  assign n6162 = n1213 ^ n338 ^ 1'b0 ;
  assign n6163 = n1585 & ~n6162 ;
  assign n6164 = ~n5315 & n6163 ;
  assign n6165 = n2701 ^ x24 ^ 1'b0 ;
  assign n6166 = x58 & n6165 ;
  assign n6167 = n6166 ^ n4256 ^ n2277 ;
  assign n6168 = n3425 ^ n3338 ^ 1'b0 ;
  assign n6169 = n5697 | n6168 ;
  assign n6170 = ( n3958 & n4339 ) | ( n3958 & ~n5366 ) | ( n4339 & ~n5366 ) ;
  assign n6171 = n1547 & n1622 ;
  assign n6172 = ~n2605 & n6171 ;
  assign n6173 = n3704 ^ n1196 ^ 1'b0 ;
  assign n6174 = n2586 & n6173 ;
  assign n6175 = n5163 ^ n1821 ^ 1'b0 ;
  assign n6176 = n6174 & n6175 ;
  assign n6177 = n2744 ^ n668 ^ n383 ;
  assign n6178 = n3445 & ~n6177 ;
  assign n6179 = n6178 ^ n5050 ^ 1'b0 ;
  assign n6180 = n5010 & n5230 ;
  assign n6181 = n4100 ^ n2219 ^ 1'b0 ;
  assign n6182 = n1581 & ~n6181 ;
  assign n6183 = n3318 ^ n1062 ^ 1'b0 ;
  assign n6184 = n6011 & n6183 ;
  assign n6185 = n5124 ^ n432 ^ 1'b0 ;
  assign n6186 = n6185 ^ n3806 ^ n3687 ;
  assign n6187 = n5079 ^ n4779 ^ 1'b0 ;
  assign n6188 = n2711 | n6187 ;
  assign n6189 = n3862 | n6188 ;
  assign n6190 = x122 & n2684 ;
  assign n6191 = ~n3470 & n6190 ;
  assign n6194 = n4509 ^ n677 ^ 1'b0 ;
  assign n6192 = ( x156 & n1691 ) | ( x156 & n4604 ) | ( n1691 & n4604 ) ;
  assign n6193 = n6192 ^ n3229 ^ 1'b0 ;
  assign n6195 = n6194 ^ n6193 ^ 1'b0 ;
  assign n6196 = ~n6191 & n6195 ;
  assign n6197 = ~n5605 & n5997 ;
  assign n6198 = n6197 ^ n1101 ^ 1'b0 ;
  assign n6199 = ~n5347 & n6198 ;
  assign n6200 = n6199 ^ x90 ^ 1'b0 ;
  assign n6201 = n711 ^ n565 ^ 1'b0 ;
  assign n6202 = n1495 | n6201 ;
  assign n6203 = n6202 ^ n4450 ^ 1'b0 ;
  assign n6204 = n4626 ^ n3466 ^ n2986 ;
  assign n6205 = n4689 ^ n1782 ^ n1574 ;
  assign n6206 = n6205 ^ n4361 ^ n1232 ;
  assign n6207 = n5830 ^ n1808 ^ 1'b0 ;
  assign n6211 = n3586 | n5125 ;
  assign n6208 = n4558 | n4779 ;
  assign n6209 = n6208 ^ n283 ^ 1'b0 ;
  assign n6210 = n4656 & ~n6209 ;
  assign n6212 = n6211 ^ n6210 ^ 1'b0 ;
  assign n6213 = ( x135 & ~n4398 ) | ( x135 & n4565 ) | ( ~n4398 & n4565 ) ;
  assign n6214 = n4031 ^ x218 ^ 1'b0 ;
  assign n6215 = n1587 & n6214 ;
  assign n6216 = ~n2849 & n5443 ;
  assign n6217 = n2024 ^ n301 ^ 1'b0 ;
  assign n6218 = x135 & ~n6217 ;
  assign n6219 = n6218 ^ n1486 ^ 1'b0 ;
  assign n6220 = x97 & n6219 ;
  assign n6221 = x205 | n4091 ;
  assign n6222 = x172 & ~n304 ;
  assign n6223 = n6222 ^ n1418 ^ 1'b0 ;
  assign n6224 = n1374 & n6223 ;
  assign n6225 = n6224 ^ n536 ^ 1'b0 ;
  assign n6226 = n3970 ^ n1970 ^ 1'b0 ;
  assign n6227 = n6225 & n6226 ;
  assign n6228 = n2783 ^ n594 ^ 1'b0 ;
  assign n6229 = n3947 ^ n1842 ^ 1'b0 ;
  assign n6230 = n6228 & n6229 ;
  assign n6231 = n5246 ^ n729 ^ 1'b0 ;
  assign n6232 = ~n1120 & n6231 ;
  assign n6233 = n3170 | n6096 ;
  assign n6234 = n2935 | n6233 ;
  assign n6235 = n3096 ^ n671 ^ 1'b0 ;
  assign n6236 = n6235 ^ n3777 ^ n2276 ;
  assign n6237 = n6236 ^ n1213 ^ 1'b0 ;
  assign n6238 = n1798 & ~n6237 ;
  assign n6239 = n1164 & ~n1781 ;
  assign n6240 = n1616 & n6239 ;
  assign n6241 = ( x163 & ~n1776 ) | ( x163 & n6240 ) | ( ~n1776 & n6240 ) ;
  assign n6242 = n6241 ^ n2895 ^ 1'b0 ;
  assign n6250 = x11 & n704 ;
  assign n6243 = n480 | n4123 ;
  assign n6244 = n985 & ~n6243 ;
  assign n6245 = x104 & ~n6244 ;
  assign n6246 = ~n1129 & n6245 ;
  assign n6247 = ~n2951 & n3690 ;
  assign n6248 = n6247 ^ n841 ^ 1'b0 ;
  assign n6249 = ( n5029 & n6246 ) | ( n5029 & ~n6248 ) | ( n6246 & ~n6248 ) ;
  assign n6251 = n6250 ^ n6249 ^ n2064 ;
  assign n6252 = n484 & n6251 ;
  assign n6253 = n6252 ^ n4758 ^ 1'b0 ;
  assign n6254 = x19 & ~n2261 ;
  assign n6255 = n6253 & n6254 ;
  assign n6256 = n1026 | n4330 ;
  assign n6257 = n6256 ^ n3160 ^ 1'b0 ;
  assign n6258 = n5877 & n6128 ;
  assign n6259 = n3988 ^ n1254 ^ 1'b0 ;
  assign n6260 = n2615 ^ n2081 ^ 1'b0 ;
  assign n6261 = n6260 ^ n4229 ^ 1'b0 ;
  assign n6262 = n3783 & n6261 ;
  assign n6263 = ~n3671 & n6262 ;
  assign n6264 = n6263 ^ n5830 ^ 1'b0 ;
  assign n6265 = n944 & ~n2068 ;
  assign n6266 = x152 & ~n6265 ;
  assign n6267 = n6266 ^ n3439 ^ 1'b0 ;
  assign n6268 = n5185 ^ n456 ^ 1'b0 ;
  assign n6269 = n3056 ^ x197 ^ 1'b0 ;
  assign n6270 = n4719 & n6269 ;
  assign n6271 = n3048 ^ n989 ^ 1'b0 ;
  assign n6272 = n5657 ^ n1155 ^ 1'b0 ;
  assign n6273 = n1278 ^ n283 ^ 1'b0 ;
  assign n6274 = x44 & n616 ;
  assign n6275 = n6274 ^ n4383 ^ 1'b0 ;
  assign n6276 = n6273 & n6275 ;
  assign n6280 = n5232 ^ n1170 ^ 1'b0 ;
  assign n6281 = n1476 & n6280 ;
  assign n6277 = n444 | n5418 ;
  assign n6278 = n6277 ^ n2751 ^ 1'b0 ;
  assign n6279 = n6278 ^ n3427 ^ n1593 ;
  assign n6282 = n6281 ^ n6279 ^ n2925 ;
  assign n6283 = n6282 ^ n4247 ^ 1'b0 ;
  assign n6284 = n4363 & n6283 ;
  assign n6285 = n880 & ~n4624 ;
  assign n6286 = n2808 & ~n6285 ;
  assign n6287 = ~n1689 & n4728 ;
  assign n6288 = n4315 ^ n563 ^ 1'b0 ;
  assign n6289 = n3119 ^ x185 ^ 1'b0 ;
  assign n6290 = ~n3811 & n6289 ;
  assign n6291 = ( x80 & ~n4359 ) | ( x80 & n6290 ) | ( ~n4359 & n6290 ) ;
  assign n6292 = n2100 ^ n1582 ^ n1535 ;
  assign n6293 = n5735 & ~n6292 ;
  assign n6294 = n6293 ^ n1520 ^ 1'b0 ;
  assign n6295 = n2213 & ~n3951 ;
  assign n6296 = n2823 ^ n881 ^ x67 ;
  assign n6297 = n940 ^ n733 ^ 1'b0 ;
  assign n6298 = ( ~n1797 & n1851 ) | ( ~n1797 & n6297 ) | ( n1851 & n6297 ) ;
  assign n6299 = ( n833 & n6296 ) | ( n833 & ~n6298 ) | ( n6296 & ~n6298 ) ;
  assign n6300 = n2148 | n6299 ;
  assign n6301 = n2685 & n3170 ;
  assign n6302 = n6301 ^ n1234 ^ 1'b0 ;
  assign n6303 = n6302 ^ n4446 ^ n409 ;
  assign n6304 = n6303 ^ n2401 ^ 1'b0 ;
  assign n6305 = n3528 | n6304 ;
  assign n6306 = n5772 ^ n3901 ^ 1'b0 ;
  assign n6307 = ~n1823 & n6306 ;
  assign n6308 = n5137 ^ n4286 ^ 1'b0 ;
  assign n6309 = n3751 | n6308 ;
  assign n6310 = n6309 ^ n2051 ^ n1702 ;
  assign n6311 = n4876 ^ n1099 ^ 1'b0 ;
  assign n6312 = n6310 & n6311 ;
  assign n6313 = x101 & ~n3852 ;
  assign n6314 = n6262 ^ n5768 ^ n4413 ;
  assign n6315 = n2289 | n4761 ;
  assign n6316 = n4760 & ~n6315 ;
  assign n6317 = n6316 ^ n4544 ^ n1256 ;
  assign n6318 = n3328 & n6317 ;
  assign n6319 = n4261 ^ n2347 ^ 1'b0 ;
  assign n6321 = n2160 ^ n1658 ^ 1'b0 ;
  assign n6320 = x74 & ~n1037 ;
  assign n6322 = n6321 ^ n6320 ^ 1'b0 ;
  assign n6323 = ~n5025 & n6322 ;
  assign n6324 = n2684 & n6323 ;
  assign n6325 = n6324 ^ n3423 ^ 1'b0 ;
  assign n6326 = ~n798 & n4145 ;
  assign n6327 = n3670 & n6326 ;
  assign n6328 = n1140 & ~n5004 ;
  assign n6329 = ~n1767 & n6328 ;
  assign n6330 = n6329 ^ n4042 ^ n3009 ;
  assign n6331 = n646 & n3567 ;
  assign n6332 = n1197 ^ n474 ^ 1'b0 ;
  assign n6333 = x26 & ~n1113 ;
  assign n6334 = ~n3817 & n6333 ;
  assign n6335 = n4964 & ~n6334 ;
  assign n6336 = n6335 ^ n3889 ^ 1'b0 ;
  assign n6337 = n4986 & n4995 ;
  assign n6338 = n1179 | n4093 ;
  assign n6339 = n6338 ^ n1665 ^ 1'b0 ;
  assign n6340 = n6337 & ~n6339 ;
  assign n6341 = n4768 ^ n3316 ^ 1'b0 ;
  assign n6342 = n1000 | n1758 ;
  assign n6343 = ~n2571 & n6342 ;
  assign n6344 = n6343 ^ n2434 ^ 1'b0 ;
  assign n6345 = ( n2990 & n6341 ) | ( n2990 & n6344 ) | ( n6341 & n6344 ) ;
  assign n6346 = n6340 & ~n6345 ;
  assign n6347 = n3122 | n3216 ;
  assign n6348 = n6347 ^ n4894 ^ 1'b0 ;
  assign n6349 = ~n3383 & n3498 ;
  assign n6350 = n4340 & ~n6349 ;
  assign n6351 = x40 & n5398 ;
  assign n6352 = n1187 & ~n2340 ;
  assign n6353 = n6352 ^ n6093 ^ n5733 ;
  assign n6354 = n4661 ^ n3232 ^ n2895 ;
  assign n6355 = n6354 ^ n1021 ^ 1'b0 ;
  assign n6356 = ~n3201 & n6355 ;
  assign n6357 = n1111 & n6356 ;
  assign n6358 = n2812 ^ n2653 ^ 1'b0 ;
  assign n6359 = x67 & n6358 ;
  assign n6360 = ( n1427 & ~n4189 ) | ( n1427 & n5565 ) | ( ~n4189 & n5565 ) ;
  assign n6361 = n6360 ^ n6312 ^ 1'b0 ;
  assign n6362 = ( ~n3041 & n6359 ) | ( ~n3041 & n6361 ) | ( n6359 & n6361 ) ;
  assign n6363 = n3088 & n3598 ;
  assign n6364 = n4657 ^ n2040 ^ 1'b0 ;
  assign n6365 = n2802 | n6364 ;
  assign n6369 = n3089 ^ n1999 ^ 1'b0 ;
  assign n6366 = n2843 ^ n881 ^ 1'b0 ;
  assign n6367 = n1693 | n2524 ;
  assign n6368 = n6366 | n6367 ;
  assign n6370 = n6369 ^ n6368 ^ 1'b0 ;
  assign n6371 = ( x160 & ~n591 ) | ( x160 & n4610 ) | ( ~n591 & n4610 ) ;
  assign n6372 = n3786 ^ n2312 ^ 1'b0 ;
  assign n6373 = n5600 & n6372 ;
  assign n6374 = n526 & n783 ;
  assign n6375 = ~x124 & n6374 ;
  assign n6376 = n6375 ^ n2952 ^ 1'b0 ;
  assign n6377 = n6049 | n6376 ;
  assign n6378 = x22 & ~n4857 ;
  assign n6379 = n5184 & n6378 ;
  assign n6380 = n896 ^ n484 ^ 1'b0 ;
  assign n6381 = ~n1876 & n6380 ;
  assign n6382 = ~n1755 & n6381 ;
  assign n6383 = ( ~n2096 & n6119 ) | ( ~n2096 & n6382 ) | ( n6119 & n6382 ) ;
  assign n6384 = n4150 & ~n6000 ;
  assign n6385 = n357 | n1108 ;
  assign n6386 = n6385 ^ n3296 ^ n2513 ;
  assign n6387 = n1024 & ~n2350 ;
  assign n6388 = ~n6386 & n6387 ;
  assign n6389 = n3295 ^ n1256 ^ n358 ;
  assign n6390 = ~n5838 & n6389 ;
  assign n6396 = x96 & x198 ;
  assign n6397 = n1711 & n6396 ;
  assign n6391 = ~n446 & n1249 ;
  assign n6393 = n1528 ^ n397 ^ 1'b0 ;
  assign n6392 = n438 & n926 ;
  assign n6394 = n6393 ^ n6392 ^ 1'b0 ;
  assign n6395 = ~n6391 & n6394 ;
  assign n6398 = n6397 ^ n6395 ^ 1'b0 ;
  assign n6399 = n3242 & ~n3620 ;
  assign n6400 = n6399 ^ n5014 ^ 1'b0 ;
  assign n6401 = n2176 & ~n6375 ;
  assign n6402 = n6401 ^ n5038 ^ n756 ;
  assign n6403 = n1930 & ~n3598 ;
  assign n6404 = n5962 ^ n1033 ^ 1'b0 ;
  assign n6405 = n6403 | n6404 ;
  assign n6406 = n2274 ^ x81 ^ 1'b0 ;
  assign n6407 = x166 & n2344 ;
  assign n6408 = n1595 & n6407 ;
  assign n6409 = n4382 | n6408 ;
  assign n6410 = n1150 ^ n304 ^ 1'b0 ;
  assign n6411 = x160 & ~n6410 ;
  assign n6412 = ~n1938 & n6411 ;
  assign n6413 = x84 & n760 ;
  assign n6414 = ( ~n3671 & n3917 ) | ( ~n3671 & n6413 ) | ( n3917 & n6413 ) ;
  assign n6415 = n3067 ^ n1006 ^ 1'b0 ;
  assign n6416 = n1875 & n6415 ;
  assign n6417 = ~n2465 & n6416 ;
  assign n6418 = n6417 ^ n3793 ^ 1'b0 ;
  assign n6419 = n6414 & ~n6418 ;
  assign n6420 = n6412 & ~n6419 ;
  assign n6421 = n4435 ^ n1120 ^ 1'b0 ;
  assign n6422 = ( n1703 & n2313 ) | ( n1703 & n5887 ) | ( n2313 & n5887 ) ;
  assign n6423 = n6422 ^ n5744 ^ 1'b0 ;
  assign n6425 = n2522 ^ n2241 ^ 1'b0 ;
  assign n6424 = n1102 ^ n766 ^ 1'b0 ;
  assign n6426 = n6425 ^ n6424 ^ 1'b0 ;
  assign n6427 = ~n2002 & n6426 ;
  assign n6428 = n6427 ^ n2641 ^ 1'b0 ;
  assign n6429 = n3806 ^ n3084 ^ 1'b0 ;
  assign n6430 = ~n1571 & n1827 ;
  assign n6431 = n2735 ^ n1698 ^ 1'b0 ;
  assign n6432 = ~n2068 & n6431 ;
  assign n6433 = n6432 ^ n3932 ^ 1'b0 ;
  assign n6434 = n6430 & ~n6433 ;
  assign n6435 = ~n4220 & n6434 ;
  assign n6436 = n6435 ^ n3704 ^ 1'b0 ;
  assign n6437 = n4661 ^ n2191 ^ 1'b0 ;
  assign n6438 = n3001 | n6437 ;
  assign n6439 = n1773 & ~n5077 ;
  assign n6440 = ~n5722 & n6439 ;
  assign n6441 = n4157 | n6440 ;
  assign n6442 = n2618 | n6441 ;
  assign n6443 = ~n1214 & n1348 ;
  assign n6444 = n6443 ^ n288 ^ 1'b0 ;
  assign n6445 = n1264 & ~n2061 ;
  assign n6446 = n4305 ^ n471 ^ 1'b0 ;
  assign n6447 = ~n2610 & n6446 ;
  assign n6448 = n1000 & ~n6447 ;
  assign n6449 = x25 & ~n2434 ;
  assign n6450 = n6449 ^ n399 ^ 1'b0 ;
  assign n6451 = n353 & ~n2044 ;
  assign n6452 = ( n462 & n1608 ) | ( n462 & n6451 ) | ( n1608 & n6451 ) ;
  assign n6453 = n1433 & n6452 ;
  assign n6454 = n2690 ^ n1559 ^ 1'b0 ;
  assign n6455 = ~n2648 & n6454 ;
  assign n6456 = n1976 & ~n4739 ;
  assign n6460 = n3493 ^ n488 ^ 1'b0 ;
  assign n6461 = n6460 ^ n1453 ^ 1'b0 ;
  assign n6457 = ~n974 & n1496 ;
  assign n6458 = n3584 & n6457 ;
  assign n6459 = n6458 ^ n783 ^ 1'b0 ;
  assign n6462 = n6461 ^ n6459 ^ n1489 ;
  assign n6463 = x12 & ~n1090 ;
  assign n6464 = n6463 ^ n5652 ^ 1'b0 ;
  assign n6465 = n930 | n6414 ;
  assign n6466 = n5804 | n6465 ;
  assign n6467 = x110 & ~n5179 ;
  assign n6468 = n3710 & ~n3754 ;
  assign n6469 = ( n2896 & ~n4084 ) | ( n2896 & n6468 ) | ( ~n4084 & n6468 ) ;
  assign n6470 = n681 & n2133 ;
  assign n6471 = x6 & ~n6470 ;
  assign n6472 = ~n2692 & n6471 ;
  assign n6475 = n4471 ^ n393 ^ 1'b0 ;
  assign n6476 = n2720 & ~n6475 ;
  assign n6477 = n2407 | n5769 ;
  assign n6478 = n6476 | n6477 ;
  assign n6473 = n357 & ~n593 ;
  assign n6474 = n4300 & n6473 ;
  assign n6479 = n6478 ^ n6474 ^ 1'b0 ;
  assign n6480 = n5338 ^ n2392 ^ 1'b0 ;
  assign n6481 = n6479 & ~n6480 ;
  assign n6482 = n3472 & ~n6481 ;
  assign n6483 = n669 & n6482 ;
  assign n6484 = n2676 ^ n892 ^ 1'b0 ;
  assign n6485 = n6484 ^ n3269 ^ 1'b0 ;
  assign n6487 = n3922 ^ n805 ^ 1'b0 ;
  assign n6488 = n742 & ~n6487 ;
  assign n6486 = x37 & n3414 ;
  assign n6489 = n6488 ^ n6486 ^ 1'b0 ;
  assign n6490 = n2692 & ~n6489 ;
  assign n6491 = ~n6485 & n6490 ;
  assign n6492 = n2553 | n3429 ;
  assign n6493 = n6492 ^ n1213 ^ 1'b0 ;
  assign n6494 = ( ~n3445 & n3926 ) | ( ~n3445 & n5634 ) | ( n3926 & n5634 ) ;
  assign n6495 = n4289 ^ n3542 ^ 1'b0 ;
  assign n6496 = n2830 & n6495 ;
  assign n6497 = ~n2076 & n5653 ;
  assign n6498 = ~n6496 & n6497 ;
  assign n6499 = n261 | n5326 ;
  assign n6500 = n6499 ^ n3078 ^ 1'b0 ;
  assign n6501 = n1980 ^ n1605 ^ 1'b0 ;
  assign n6502 = ( n2214 & n4281 ) | ( n2214 & ~n6501 ) | ( n4281 & ~n6501 ) ;
  assign n6504 = n5991 ^ n4012 ^ 1'b0 ;
  assign n6503 = x38 & ~n4759 ;
  assign n6505 = n6504 ^ n6503 ^ 1'b0 ;
  assign n6506 = ~n6502 & n6505 ;
  assign n6507 = n3233 | n3281 ;
  assign n6510 = n1708 ^ n1388 ^ 1'b0 ;
  assign n6511 = ~n4556 & n6510 ;
  assign n6512 = n3958 & n6511 ;
  assign n6508 = n5343 ^ n3147 ^ 1'b0 ;
  assign n6509 = ( n939 & n5720 ) | ( n939 & ~n6508 ) | ( n5720 & ~n6508 ) ;
  assign n6513 = n6512 ^ n6509 ^ 1'b0 ;
  assign n6514 = n2708 | n5997 ;
  assign n6515 = n1768 ^ n922 ^ 1'b0 ;
  assign n6516 = ( ~n3222 & n5567 ) | ( ~n3222 & n6089 ) | ( n5567 & n6089 ) ;
  assign n6517 = n1358 & n5367 ;
  assign n6518 = n4306 & ~n6517 ;
  assign n6519 = ~n940 & n5629 ;
  assign n6520 = n1532 & n6519 ;
  assign n6521 = n2093 | n6520 ;
  assign n6522 = n6521 ^ n3878 ^ 1'b0 ;
  assign n6523 = ~n441 & n6522 ;
  assign n6524 = n6523 ^ n399 ^ 1'b0 ;
  assign n6525 = ~n4215 & n6524 ;
  assign n6526 = n4097 ^ n4037 ^ 1'b0 ;
  assign n6527 = n2241 ^ n1842 ^ 1'b0 ;
  assign n6528 = x52 & ~n6527 ;
  assign n6529 = n4926 | n6528 ;
  assign n6530 = n3126 & n6529 ;
  assign n6531 = n6530 ^ n1400 ^ 1'b0 ;
  assign n6532 = n6526 & n6531 ;
  assign n6533 = n6532 ^ n1610 ^ 1'b0 ;
  assign n6536 = n6080 ^ n3567 ^ 1'b0 ;
  assign n6537 = x99 | n6536 ;
  assign n6538 = n6537 ^ n744 ^ 1'b0 ;
  assign n6539 = n3643 & n6538 ;
  assign n6540 = ~n3694 & n6539 ;
  assign n6534 = n1113 & n4573 ;
  assign n6535 = n5468 & n6534 ;
  assign n6541 = n6540 ^ n6535 ^ 1'b0 ;
  assign n6542 = n1176 & ~n5687 ;
  assign n6543 = ( n1590 & n4056 ) | ( n1590 & n5315 ) | ( n4056 & n5315 ) ;
  assign n6545 = n931 & ~n2342 ;
  assign n6546 = n6545 ^ n1553 ^ 1'b0 ;
  assign n6544 = n3645 ^ n3362 ^ n1930 ;
  assign n6547 = n6546 ^ n6544 ^ 1'b0 ;
  assign n6548 = n2292 | n6547 ;
  assign n6549 = ~x22 & n405 ;
  assign n6550 = n6549 ^ n1716 ^ 1'b0 ;
  assign n6551 = n6484 | n6550 ;
  assign n6552 = n1776 | n6551 ;
  assign n6553 = n6552 ^ n5830 ^ 1'b0 ;
  assign n6554 = n6548 | n6553 ;
  assign n6555 = n6554 ^ n1253 ^ 1'b0 ;
  assign n6556 = ~n1302 & n1865 ;
  assign n6557 = x132 & n1955 ;
  assign n6558 = n4238 & n6557 ;
  assign n6559 = n5543 | n6558 ;
  assign n6560 = n926 & n1473 ;
  assign n6561 = ~n6559 & n6560 ;
  assign n6562 = n6561 ^ n2166 ^ 1'b0 ;
  assign n6563 = n2748 | n6562 ;
  assign n6564 = n5203 & ~n6563 ;
  assign n6565 = ~n6556 & n6564 ;
  assign n6566 = n4137 ^ n1707 ^ 1'b0 ;
  assign n6567 = n3344 & ~n6566 ;
  assign n6568 = n2735 ^ n2209 ^ 1'b0 ;
  assign n6569 = ~n3481 & n6568 ;
  assign n6570 = n704 & n2578 ;
  assign n6571 = ~n6569 & n6570 ;
  assign n6572 = n2921 & ~n6571 ;
  assign n6573 = ( x135 & n6054 ) | ( x135 & n6572 ) | ( n6054 & n6572 ) ;
  assign n6574 = n1832 & ~n2065 ;
  assign n6575 = ( n1053 & ~n2324 ) | ( n1053 & n4969 ) | ( ~n2324 & n4969 ) ;
  assign n6576 = x37 & ~n2504 ;
  assign n6577 = n1851 & n6576 ;
  assign n6578 = ( n970 & n1717 ) | ( n970 & n6577 ) | ( n1717 & n6577 ) ;
  assign n6583 = n445 ^ n261 ^ 1'b0 ;
  assign n6584 = n1223 & ~n6583 ;
  assign n6582 = n1572 | n1771 ;
  assign n6585 = n6584 ^ n6582 ^ 1'b0 ;
  assign n6581 = ~n3434 & n5476 ;
  assign n6586 = n6585 ^ n6581 ^ 1'b0 ;
  assign n6587 = n1823 ^ n1585 ^ 1'b0 ;
  assign n6588 = n6586 | n6587 ;
  assign n6579 = ( ~n1991 & n2156 ) | ( ~n1991 & n4126 ) | ( n2156 & n4126 ) ;
  assign n6580 = n3032 & n6579 ;
  assign n6589 = n6588 ^ n6580 ^ 1'b0 ;
  assign n6590 = n2653 ^ n683 ^ 1'b0 ;
  assign n6591 = n2959 & ~n6372 ;
  assign n6592 = ( n2274 & n5805 ) | ( n2274 & ~n5861 ) | ( n5805 & ~n5861 ) ;
  assign n6593 = n4004 ^ n3088 ^ x147 ;
  assign n6594 = ~n3376 & n6593 ;
  assign n6595 = n3864 & ~n6594 ;
  assign n6596 = n5231 ^ n2360 ^ 1'b0 ;
  assign n6597 = n2210 ^ n785 ^ 1'b0 ;
  assign n6603 = ~n480 & n1736 ;
  assign n6604 = n6603 ^ n1058 ^ 1'b0 ;
  assign n6601 = n3291 ^ n2580 ^ 1'b0 ;
  assign n6598 = x196 & ~n813 ;
  assign n6599 = n1648 & n6598 ;
  assign n6600 = n6599 ^ n1075 ^ 1'b0 ;
  assign n6602 = n6601 ^ n6600 ^ n307 ;
  assign n6605 = n6604 ^ n6602 ^ n306 ;
  assign n6606 = ( ~n947 & n1941 ) | ( ~n947 & n5759 ) | ( n1941 & n5759 ) ;
  assign n6607 = n4129 ^ n3081 ^ 1'b0 ;
  assign n6608 = n6604 ^ n1701 ^ n462 ;
  assign n6609 = n6608 ^ n3283 ^ 1'b0 ;
  assign n6610 = n6609 ^ n778 ^ 1'b0 ;
  assign n6611 = ~n1308 & n2525 ;
  assign n6612 = n3112 & n6611 ;
  assign n6613 = ~n4284 & n6612 ;
  assign n6614 = n4080 | n6613 ;
  assign n6615 = x15 | n6614 ;
  assign n6616 = n6408 ^ n317 ^ 1'b0 ;
  assign n6617 = n4608 & ~n6616 ;
  assign n6618 = ( n5652 & ~n6136 ) | ( n5652 & n6617 ) | ( ~n6136 & n6617 ) ;
  assign n6621 = x3 & ~n4964 ;
  assign n6620 = ~n545 & n2884 ;
  assign n6622 = n6621 ^ n6620 ^ 1'b0 ;
  assign n6619 = n2059 & ~n5095 ;
  assign n6623 = n6622 ^ n6619 ^ 1'b0 ;
  assign n6624 = ( n1431 & n2368 ) | ( n1431 & ~n3062 ) | ( n2368 & ~n3062 ) ;
  assign n6625 = n3254 & ~n6624 ;
  assign n6626 = n1448 & ~n4573 ;
  assign n6627 = n6626 ^ n1826 ^ 1'b0 ;
  assign n6628 = x160 | n1629 ;
  assign n6629 = x14 & n6628 ;
  assign n6630 = n6627 & n6629 ;
  assign n6631 = n6630 ^ n4281 ^ 1'b0 ;
  assign n6632 = n6625 | n6631 ;
  assign n6633 = x73 & ~n908 ;
  assign n6634 = n908 & n6633 ;
  assign n6635 = n2544 | n2941 ;
  assign n6636 = n6635 ^ n4808 ^ 1'b0 ;
  assign n6637 = n6636 ^ n3564 ^ 1'b0 ;
  assign n6638 = n1742 & n6637 ;
  assign n6639 = n6638 ^ n4978 ^ 1'b0 ;
  assign n6640 = ~n6634 & n6639 ;
  assign n6642 = n298 | n1475 ;
  assign n6643 = n2449 & ~n6642 ;
  assign n6644 = n2144 & n5804 ;
  assign n6645 = ( ~n663 & n6643 ) | ( ~n663 & n6644 ) | ( n6643 & n6644 ) ;
  assign n6641 = n2436 | n5404 ;
  assign n6646 = n6645 ^ n6641 ^ n5790 ;
  assign n6652 = n2522 ^ x167 ^ 1'b0 ;
  assign n6653 = ~n5693 & n6652 ;
  assign n6654 = n6653 ^ n2483 ^ n2481 ;
  assign n6647 = ~x111 & n3410 ;
  assign n6648 = n6647 ^ n2414 ^ 1'b0 ;
  assign n6649 = n3887 & ~n6648 ;
  assign n6650 = n6649 ^ n5980 ^ 1'b0 ;
  assign n6651 = x174 & n6650 ;
  assign n6655 = n6654 ^ n6651 ^ n5114 ;
  assign n6656 = n1517 ^ n1049 ^ n642 ;
  assign n6657 = ~n2973 & n6656 ;
  assign n6658 = ~n3095 & n6657 ;
  assign n6661 = ~x121 & n1978 ;
  assign n6662 = n6007 ^ x12 ^ 1'b0 ;
  assign n6663 = n572 | n6662 ;
  assign n6664 = n6661 | n6663 ;
  assign n6665 = n1107 | n6664 ;
  assign n6659 = x239 & n821 ;
  assign n6660 = n6659 ^ n2578 ^ 1'b0 ;
  assign n6666 = n6665 ^ n6660 ^ 1'b0 ;
  assign n6667 = n1685 | n6666 ;
  assign n6668 = n5621 | n6667 ;
  assign n6669 = n570 & n4480 ;
  assign n6670 = ( n1113 & ~n3551 ) | ( n1113 & n6669 ) | ( ~n3551 & n6669 ) ;
  assign n6671 = ( n818 & ~n1666 ) | ( n818 & n6670 ) | ( ~n1666 & n6670 ) ;
  assign n6672 = n6671 ^ n3469 ^ n1648 ;
  assign n6673 = n1961 & ~n2135 ;
  assign n6674 = n6279 | n6673 ;
  assign n6675 = n314 & n5893 ;
  assign n6676 = ~n6674 & n6675 ;
  assign n6677 = n4527 & ~n5849 ;
  assign n6678 = n2884 & ~n2907 ;
  assign n6679 = n6678 ^ n520 ^ 1'b0 ;
  assign n6680 = x175 & n1337 ;
  assign n6681 = ~n4080 & n6680 ;
  assign n6682 = ( n1170 & n6448 ) | ( n1170 & n6681 ) | ( n6448 & n6681 ) ;
  assign n6683 = n6682 ^ n3520 ^ 1'b0 ;
  assign n6684 = ( ~n1681 & n2133 ) | ( ~n1681 & n4993 ) | ( n2133 & n4993 ) ;
  assign n6685 = x17 & n2690 ;
  assign n6686 = n6685 ^ n2549 ^ 1'b0 ;
  assign n6687 = n6362 ^ n898 ^ 1'b0 ;
  assign n6688 = n5762 | n6687 ;
  assign n6692 = n436 & ~n4413 ;
  assign n6689 = n2020 & ~n2968 ;
  assign n6690 = n6689 ^ n639 ^ 1'b0 ;
  assign n6691 = ~n5989 & n6690 ;
  assign n6693 = n6692 ^ n6691 ^ 1'b0 ;
  assign n6695 = n1306 ^ x169 ^ 1'b0 ;
  assign n6696 = n1875 & ~n6695 ;
  assign n6694 = ~x247 & n4073 ;
  assign n6697 = n6696 ^ n6694 ^ n3804 ;
  assign n6698 = n6697 ^ n2949 ^ 1'b0 ;
  assign n6699 = x175 & ~n6698 ;
  assign n6700 = ~n3716 & n6699 ;
  assign n6701 = ~n3785 & n4704 ;
  assign n6702 = n6299 ^ n4153 ^ 1'b0 ;
  assign n6703 = n6701 & ~n6702 ;
  assign n6704 = ~n967 & n5453 ;
  assign n6705 = n629 & ~n1253 ;
  assign n6707 = ~n504 & n1690 ;
  assign n6708 = ~n1988 & n6707 ;
  assign n6706 = x95 & ~n3852 ;
  assign n6709 = n6708 ^ n6706 ^ 1'b0 ;
  assign n6710 = n6084 ^ n3019 ^ 1'b0 ;
  assign n6711 = n275 & ~n6710 ;
  assign n6712 = x163 & ~n2623 ;
  assign n6713 = n6712 ^ n3579 ^ 1'b0 ;
  assign n6714 = n3102 & n6713 ;
  assign n6715 = n1802 | n6714 ;
  assign n6716 = n2881 | n5634 ;
  assign n6717 = n6716 ^ n3245 ^ 1'b0 ;
  assign n6718 = n4600 & ~n4749 ;
  assign n6719 = ~n6717 & n6718 ;
  assign n6721 = n4661 | n4784 ;
  assign n6722 = n6721 ^ n3696 ^ n1233 ;
  assign n6723 = ( n1913 & ~n5540 ) | ( n1913 & n6722 ) | ( ~n5540 & n6722 ) ;
  assign n6720 = n2777 & n3180 ;
  assign n6724 = n6723 ^ n6720 ^ n2929 ;
  assign n6725 = n2630 | n4462 ;
  assign n6726 = n6711 & n6725 ;
  assign n6727 = ( n286 & n4245 ) | ( n286 & n4451 ) | ( n4245 & n4451 ) ;
  assign n6728 = ~n1285 & n1755 ;
  assign n6729 = ~n4057 & n6728 ;
  assign n6730 = n6729 ^ n2752 ^ 1'b0 ;
  assign n6731 = n3786 ^ n2253 ^ 1'b0 ;
  assign n6732 = n835 | n6731 ;
  assign n6733 = n2449 & ~n6732 ;
  assign n6734 = n6733 ^ n3633 ^ 1'b0 ;
  assign n6737 = n4494 ^ n2608 ^ 1'b0 ;
  assign n6735 = n1795 | n2860 ;
  assign n6736 = n6735 ^ n5140 ^ 1'b0 ;
  assign n6738 = n6737 ^ n6736 ^ 1'b0 ;
  assign n6739 = n4193 & n6738 ;
  assign n6740 = n4537 & n6198 ;
  assign n6741 = ~n1603 & n6740 ;
  assign n6742 = n6741 ^ n5089 ^ 1'b0 ;
  assign n6743 = n4242 & ~n6742 ;
  assign n6744 = x147 & n4996 ;
  assign n6745 = n6744 ^ n1874 ^ 1'b0 ;
  assign n6746 = n5052 & ~n6745 ;
  assign n6747 = n6746 ^ n6352 ^ 1'b0 ;
  assign n6748 = n3973 | n6571 ;
  assign n6749 = n5924 ^ n2232 ^ n2188 ;
  assign n6750 = x95 & ~n1033 ;
  assign n6751 = n6750 ^ n1967 ^ 1'b0 ;
  assign n6754 = ( ~x138 & n2020 ) | ( ~x138 & n3293 ) | ( n2020 & n3293 ) ;
  assign n6753 = n1913 & n2436 ;
  assign n6755 = n6754 ^ n6753 ^ 1'b0 ;
  assign n6756 = n3166 & n6755 ;
  assign n6752 = ~n886 & n4570 ;
  assign n6757 = n6756 ^ n6752 ^ 1'b0 ;
  assign n6758 = ( n2877 & n5498 ) | ( n2877 & ~n6757 ) | ( n5498 & ~n6757 ) ;
  assign n6759 = n3982 & n6758 ;
  assign n6760 = n6751 & n6759 ;
  assign n6761 = n2715 & n2943 ;
  assign n6762 = n6761 ^ n5818 ^ 1'b0 ;
  assign n6766 = n1826 & ~n6460 ;
  assign n6763 = n1840 ^ n1179 ^ 1'b0 ;
  assign n6764 = x176 & n6763 ;
  assign n6765 = ~n5671 & n6764 ;
  assign n6767 = n6766 ^ n6765 ^ 1'b0 ;
  assign n6768 = n3666 & n4934 ;
  assign n6769 = x39 & ~n6768 ;
  assign n6770 = n6767 & n6769 ;
  assign n6771 = n6553 ^ n3720 ^ n1213 ;
  assign n6772 = n5448 ^ n4573 ^ n3220 ;
  assign n6773 = n6166 ^ n5310 ^ 1'b0 ;
  assign n6774 = ( n471 & n1600 ) | ( n471 & ~n2849 ) | ( n1600 & ~n2849 ) ;
  assign n6775 = ~n365 & n6774 ;
  assign n6776 = n5825 ^ n1202 ^ n700 ;
  assign n6777 = n6775 | n6776 ;
  assign n6778 = ( ~n2536 & n4542 ) | ( ~n2536 & n6047 ) | ( n4542 & n6047 ) ;
  assign n6779 = n5306 ^ n1236 ^ x253 ;
  assign n6780 = n6778 | n6779 ;
  assign n6781 = n2901 ^ n723 ^ n320 ;
  assign n6782 = ~n2462 & n6781 ;
  assign n6783 = n6782 ^ n1631 ^ 1'b0 ;
  assign n6784 = n1255 ^ n492 ^ 1'b0 ;
  assign n6785 = ( ~n2697 & n3316 ) | ( ~n2697 & n6784 ) | ( n3316 & n6784 ) ;
  assign n6786 = n6785 ^ n5918 ^ 1'b0 ;
  assign n6787 = n6783 | n6786 ;
  assign n6788 = ~n1705 & n3108 ;
  assign n6789 = n1334 & n6788 ;
  assign n6790 = ~n3827 & n6789 ;
  assign n6792 = n6528 ^ n4494 ^ n634 ;
  assign n6791 = ~n3021 & n3310 ;
  assign n6793 = n6792 ^ n6791 ^ 1'b0 ;
  assign n6794 = n6793 ^ n5711 ^ 1'b0 ;
  assign n6795 = n5288 | n6794 ;
  assign n6796 = n1460 & n5915 ;
  assign n6797 = ~n5065 & n6796 ;
  assign n6798 = n2048 ^ x89 ^ 1'b0 ;
  assign n6799 = n1633 & n6798 ;
  assign n6800 = n1302 & n6799 ;
  assign n6801 = ( x111 & ~n1978 ) | ( x111 & n6800 ) | ( ~n1978 & n6800 ) ;
  assign n6802 = ~n1553 & n2563 ;
  assign n6803 = n6802 ^ n2132 ^ 1'b0 ;
  assign n6804 = ~n4278 & n6803 ;
  assign n6805 = n3232 ^ n797 ^ 1'b0 ;
  assign n6806 = n6805 ^ n2029 ^ 1'b0 ;
  assign n6807 = n6804 & n6806 ;
  assign n6808 = n6807 ^ n402 ^ 1'b0 ;
  assign n6809 = n2799 ^ n915 ^ 1'b0 ;
  assign n6810 = ~n4808 & n6809 ;
  assign n6814 = n2397 & n3215 ;
  assign n6811 = n1462 & n5877 ;
  assign n6812 = ~n3583 & n6811 ;
  assign n6813 = ~n3545 & n6812 ;
  assign n6815 = n6814 ^ n6813 ^ 1'b0 ;
  assign n6816 = n5479 ^ n3595 ^ n3538 ;
  assign n6817 = n4761 ^ n1122 ^ 1'b0 ;
  assign n6818 = n4349 | n6817 ;
  assign n6819 = n5729 ^ n1913 ^ 1'b0 ;
  assign n6820 = n3773 | n6819 ;
  assign n6821 = ( ~x19 & n1460 ) | ( ~x19 & n6114 ) | ( n1460 & n6114 ) ;
  assign n6822 = x107 | n6821 ;
  assign n6823 = n2100 & n3648 ;
  assign n6824 = n4689 & n6823 ;
  assign n6825 = ( n296 & ~n3917 ) | ( n296 & n5298 ) | ( ~n3917 & n5298 ) ;
  assign n6826 = n970 & n3116 ;
  assign n6827 = ~n4231 & n6826 ;
  assign n6828 = n6827 ^ n1468 ^ 1'b0 ;
  assign n6829 = x153 & ~n571 ;
  assign n6830 = ~n2221 & n6829 ;
  assign n6831 = n3929 ^ n2553 ^ 1'b0 ;
  assign n6832 = n1017 & n1096 ;
  assign n6833 = n2711 & n6832 ;
  assign n6834 = n4462 | n6833 ;
  assign n6835 = ( n1974 & n2066 ) | ( n1974 & n2649 ) | ( n2066 & n2649 ) ;
  assign n6836 = ~n856 & n946 ;
  assign n6837 = n6836 ^ n1987 ^ 1'b0 ;
  assign n6838 = ( n2998 & n5640 ) | ( n2998 & ~n6837 ) | ( n5640 & ~n6837 ) ;
  assign n6839 = n6835 | n6838 ;
  assign n6840 = n6839 ^ n961 ^ 1'b0 ;
  assign n6841 = ( ~n942 & n3438 ) | ( ~n942 & n3979 ) | ( n3438 & n3979 ) ;
  assign n6842 = ( ~n723 & n1019 ) | ( ~n723 & n1985 ) | ( n1019 & n1985 ) ;
  assign n6843 = n6022 ^ n4330 ^ 1'b0 ;
  assign n6844 = ~n6842 & n6843 ;
  assign n6845 = ~n2775 & n6844 ;
  assign n6846 = ~n5021 & n6845 ;
  assign n6847 = n694 | n3603 ;
  assign n6848 = n3047 & ~n6847 ;
  assign n6849 = n6848 ^ n5573 ^ 1'b0 ;
  assign n6850 = n2448 ^ n2278 ^ n2276 ;
  assign n6851 = n2306 & ~n3597 ;
  assign n6852 = ~n725 & n5364 ;
  assign n6853 = n1595 | n2286 ;
  assign n6854 = n3360 ^ n922 ^ x222 ;
  assign n6860 = ~n2387 & n4784 ;
  assign n6861 = n6860 ^ n2521 ^ 1'b0 ;
  assign n6862 = n3770 ^ n1504 ^ 1'b0 ;
  assign n6863 = n3417 & ~n6862 ;
  assign n6864 = n6863 ^ n599 ^ 1'b0 ;
  assign n6865 = ~n6861 & n6864 ;
  assign n6855 = ~n2212 & n2756 ;
  assign n6856 = n6855 ^ n1894 ^ 1'b0 ;
  assign n6857 = ~n6117 & n6856 ;
  assign n6858 = ~n4042 & n6857 ;
  assign n6859 = n6858 ^ n2466 ^ 1'b0 ;
  assign n6866 = n6865 ^ n6859 ^ 1'b0 ;
  assign n6867 = ( n4081 & ~n4587 ) | ( n4081 & n6442 ) | ( ~n4587 & n6442 ) ;
  assign n6868 = n5140 ^ n4170 ^ x78 ;
  assign n6869 = ~n3639 & n5025 ;
  assign n6870 = n2176 & n6476 ;
  assign n6871 = ~n1462 & n4718 ;
  assign n6872 = n5973 & ~n6871 ;
  assign n6873 = n6870 & n6872 ;
  assign n6874 = n371 ^ x103 ^ 1'b0 ;
  assign n6875 = n1228 ^ n354 ^ 1'b0 ;
  assign n6876 = ~n6874 & n6875 ;
  assign n6877 = n6876 ^ n5721 ^ 1'b0 ;
  assign n6879 = ~n1650 & n4602 ;
  assign n6880 = n6879 ^ n1125 ^ 1'b0 ;
  assign n6881 = n6880 ^ n5713 ^ 1'b0 ;
  assign n6878 = n570 & ~n1462 ;
  assign n6882 = n6881 ^ n6878 ^ 1'b0 ;
  assign n6883 = n905 & n2913 ;
  assign n6884 = n6883 ^ n1213 ^ 1'b0 ;
  assign n6885 = n6884 ^ n6140 ^ 1'b0 ;
  assign n6886 = n1808 ^ n496 ^ 1'b0 ;
  assign n6887 = n1427 & n6886 ;
  assign n6888 = n6415 ^ n2124 ^ n1807 ;
  assign n6889 = ~n6887 & n6888 ;
  assign n6890 = n911 ^ n283 ^ 1'b0 ;
  assign n6891 = n455 | n6890 ;
  assign n6892 = n972 ^ n596 ^ 1'b0 ;
  assign n6893 = n6891 | n6892 ;
  assign n6894 = n3216 & ~n6893 ;
  assign n6895 = n3253 ^ n2728 ^ n1572 ;
  assign n6896 = ~x219 & n6895 ;
  assign n6897 = n6896 ^ n5635 ^ 1'b0 ;
  assign n6898 = ~n3283 & n6897 ;
  assign n6899 = x170 | n2528 ;
  assign n6900 = n3010 & ~n6899 ;
  assign n6901 = n6900 ^ x31 ^ 1'b0 ;
  assign n6902 = n2644 | n5071 ;
  assign n6903 = n6902 ^ n3056 ^ 1'b0 ;
  assign n6910 = n1196 & n4959 ;
  assign n6909 = ( n3812 & n5326 ) | ( n3812 & ~n5521 ) | ( n5326 & ~n5521 ) ;
  assign n6907 = ( ~n3558 & n3783 ) | ( ~n3558 & n4216 ) | ( n3783 & n4216 ) ;
  assign n6905 = n1972 | n3696 ;
  assign n6906 = n5311 & ~n6905 ;
  assign n6904 = n6501 ^ n3225 ^ 1'b0 ;
  assign n6908 = n6907 ^ n6906 ^ n6904 ;
  assign n6911 = n6910 ^ n6909 ^ n6908 ;
  assign n6912 = ( n1117 & n2682 ) | ( n1117 & n4981 ) | ( n2682 & n4981 ) ;
  assign n6913 = n2406 | n6912 ;
  assign n6914 = n6913 ^ n6054 ^ 1'b0 ;
  assign n6915 = n6069 ^ n4182 ^ 1'b0 ;
  assign n6918 = n467 | n2422 ;
  assign n6919 = n5630 | n6918 ;
  assign n6916 = n1127 ^ x10 ^ 1'b0 ;
  assign n6917 = n4964 & ~n6916 ;
  assign n6920 = n6919 ^ n6917 ^ 1'b0 ;
  assign n6921 = n1327 ^ x65 ^ 1'b0 ;
  assign n6922 = ( n4007 & n6215 ) | ( n4007 & n6921 ) | ( n6215 & n6921 ) ;
  assign n6923 = n6922 ^ n2162 ^ 1'b0 ;
  assign n6925 = n4505 ^ n524 ^ 1'b0 ;
  assign n6926 = n1362 & ~n6925 ;
  assign n6924 = ~n1404 & n3209 ;
  assign n6927 = n6926 ^ n6924 ^ 1'b0 ;
  assign n6928 = x118 & n6051 ;
  assign n6929 = n6928 ^ n2231 ^ 1'b0 ;
  assign n6930 = n6929 ^ n3937 ^ n3145 ;
  assign n6931 = ( n3332 & n6927 ) | ( n3332 & n6930 ) | ( n6927 & n6930 ) ;
  assign n6932 = n2728 ^ n1404 ^ 1'b0 ;
  assign n6933 = n3074 & ~n6932 ;
  assign n6934 = n6933 ^ n2085 ^ 1'b0 ;
  assign n6935 = n6921 ^ n1005 ^ 1'b0 ;
  assign n6936 = n2153 & ~n6935 ;
  assign n6937 = n1665 ^ n315 ^ 1'b0 ;
  assign n6938 = ~n4039 & n6937 ;
  assign n6939 = n3884 | n6725 ;
  assign n6940 = n5550 | n6939 ;
  assign n6941 = x225 & n1366 ;
  assign n6942 = n6941 ^ n4644 ^ 1'b0 ;
  assign n6943 = n3536 | n6942 ;
  assign n6944 = ~n1423 & n4434 ;
  assign n6945 = ~n760 & n6944 ;
  assign n6946 = n2930 & n4905 ;
  assign n6947 = ~n6945 & n6946 ;
  assign n6948 = n4627 | n6947 ;
  assign n6949 = n6943 & ~n6948 ;
  assign n6950 = n2276 & n4002 ;
  assign n6951 = n3272 & n4938 ;
  assign n6952 = n6951 ^ n978 ^ 1'b0 ;
  assign n6953 = ( n1613 & ~n1980 ) | ( n1613 & n2543 ) | ( ~n1980 & n2543 ) ;
  assign n6954 = ~n2015 & n6953 ;
  assign n6955 = n6442 ^ n2437 ^ n2174 ;
  assign n6956 = n5690 ^ n1278 ^ x245 ;
  assign n6957 = ~n1916 & n3737 ;
  assign n6958 = ~n6232 & n6957 ;
  assign n6959 = n2778 & ~n4534 ;
  assign n6960 = n2101 & n6959 ;
  assign n6961 = n2838 ^ n1653 ^ 1'b0 ;
  assign n6962 = n6960 & n6961 ;
  assign n6964 = n345 | n1594 ;
  assign n6963 = n2421 & ~n5464 ;
  assign n6965 = n6964 ^ n6963 ^ 1'b0 ;
  assign n6966 = n1222 & n6965 ;
  assign n6967 = x186 & n2226 ;
  assign n6968 = n6967 ^ n2023 ^ 1'b0 ;
  assign n6969 = n3759 ^ x161 ^ 1'b0 ;
  assign n6973 = n2202 ^ n982 ^ 1'b0 ;
  assign n6974 = n6973 ^ n1490 ^ 1'b0 ;
  assign n6975 = n6638 & n6974 ;
  assign n6970 = n312 & n1798 ;
  assign n6971 = n6970 ^ n4368 ^ 1'b0 ;
  assign n6972 = n915 & ~n6971 ;
  assign n6976 = n6975 ^ n6972 ^ 1'b0 ;
  assign n6977 = n4715 ^ n3111 ^ 1'b0 ;
  assign n6978 = x159 & ~n3499 ;
  assign n6979 = ~n6977 & n6978 ;
  assign n6980 = x28 & ~n2303 ;
  assign n6981 = ( x158 & n3515 ) | ( x158 & n6980 ) | ( n3515 & n6980 ) ;
  assign n6982 = n6981 ^ n4618 ^ x181 ;
  assign n6983 = n5329 & n5464 ;
  assign n6984 = n6983 ^ n2463 ^ 1'b0 ;
  assign n6985 = ~n1055 & n3342 ;
  assign n6986 = n6167 ^ n4096 ^ n3764 ;
  assign n6987 = n6415 ^ n3806 ^ 1'b0 ;
  assign n6988 = n6103 ^ n1631 ^ 1'b0 ;
  assign n6992 = n6488 ^ n4454 ^ 1'b0 ;
  assign n6989 = n4960 | n6698 ;
  assign n6990 = n5449 | n6989 ;
  assign n6991 = n4969 & n6990 ;
  assign n6993 = n6992 ^ n6991 ^ 1'b0 ;
  assign n6994 = ( n2078 & ~n2216 ) | ( n2078 & n4438 ) | ( ~n2216 & n4438 ) ;
  assign n6995 = n1349 ^ x248 ^ 1'b0 ;
  assign n6996 = n3073 & n4588 ;
  assign n6997 = ~n6995 & n6996 ;
  assign n6998 = ( n3154 & ~n4358 ) | ( n3154 & n6997 ) | ( ~n4358 & n6997 ) ;
  assign n7002 = n2276 | n4995 ;
  assign n6999 = x102 & x217 ;
  assign n7000 = n6999 ^ n434 ^ 1'b0 ;
  assign n7001 = ( n1967 & ~n2871 ) | ( n1967 & n7000 ) | ( ~n2871 & n7000 ) ;
  assign n7003 = n7002 ^ n7001 ^ n2434 ;
  assign n7004 = n6690 ^ x132 ^ 1'b0 ;
  assign n7005 = n2851 ^ n1148 ^ 1'b0 ;
  assign n7006 = n3126 & ~n7005 ;
  assign n7007 = ~n7004 & n7006 ;
  assign n7008 = n557 & n4509 ;
  assign n7009 = x75 ^ x49 ^ 1'b0 ;
  assign n7010 = n1332 & n7009 ;
  assign n7011 = ~n3246 & n7010 ;
  assign n7012 = n1342 & n7011 ;
  assign n7013 = n7012 ^ n1021 ^ 1'b0 ;
  assign n7014 = x233 & n4326 ;
  assign n7015 = ( n1324 & ~n2702 ) | ( n1324 & n7014 ) | ( ~n2702 & n7014 ) ;
  assign n7016 = n4296 & ~n7015 ;
  assign n7017 = n2320 & n2676 ;
  assign n7018 = x2 & ~n2653 ;
  assign n7019 = ~n2206 & n7018 ;
  assign n7020 = n5515 ^ n604 ^ 1'b0 ;
  assign n7021 = n7020 ^ n6756 ^ n259 ;
  assign n7022 = x27 & ~n7021 ;
  assign n7023 = n3369 & n7022 ;
  assign n7024 = n733 & ~n1368 ;
  assign n7025 = n7024 ^ n5195 ^ 1'b0 ;
  assign n7026 = ~n7023 & n7025 ;
  assign n7027 = n4815 ^ n2481 ^ n1798 ;
  assign n7028 = n2414 ^ n481 ^ n407 ;
  assign n7029 = n1272 & ~n3094 ;
  assign n7030 = n7029 ^ n3270 ^ 1'b0 ;
  assign n7031 = n3249 & ~n7030 ;
  assign n7032 = x169 & n7031 ;
  assign n7033 = n7028 & n7032 ;
  assign n7034 = n1619 & n5684 ;
  assign n7035 = n7034 ^ n2975 ^ 1'b0 ;
  assign n7036 = x234 & n6197 ;
  assign n7037 = n1200 & n3907 ;
  assign n7038 = n7037 ^ n6641 ^ 1'b0 ;
  assign n7039 = ( n622 & n2322 ) | ( n622 & ~n3834 ) | ( n2322 & ~n3834 ) ;
  assign n7040 = n4980 ^ n4317 ^ n2998 ;
  assign n7041 = n2365 & ~n7040 ;
  assign n7042 = n4117 & ~n7041 ;
  assign n7043 = ~n5357 & n7042 ;
  assign n7044 = ~x178 & n265 ;
  assign n7045 = n7044 ^ n425 ^ 1'b0 ;
  assign n7046 = n4309 & ~n7045 ;
  assign n7047 = n6898 ^ n5142 ^ 1'b0 ;
  assign n7048 = n1592 & ~n3517 ;
  assign n7049 = n7048 ^ n4194 ^ 1'b0 ;
  assign n7053 = n1733 & ~n2823 ;
  assign n7052 = n326 & n1090 ;
  assign n7054 = n7053 ^ n7052 ^ n4917 ;
  assign n7050 = n3746 ^ n1561 ^ 1'b0 ;
  assign n7051 = n761 & ~n7050 ;
  assign n7055 = n7054 ^ n7051 ^ 1'b0 ;
  assign n7056 = n2183 ^ n1693 ^ n753 ;
  assign n7057 = n3335 & n7056 ;
  assign n7058 = ( x33 & n2183 ) | ( x33 & ~n7057 ) | ( n2183 & ~n7057 ) ;
  assign n7059 = n1156 ^ n718 ^ 1'b0 ;
  assign n7060 = n6656 & n7059 ;
  assign n7061 = n2910 | n6445 ;
  assign n7062 = n7060 | n7061 ;
  assign n7063 = ~n1763 & n2680 ;
  assign n7064 = ( n2699 & ~n5079 ) | ( n2699 & n7063 ) | ( ~n5079 & n7063 ) ;
  assign n7065 = n2122 & ~n4655 ;
  assign n7066 = n7065 ^ n1486 ^ 1'b0 ;
  assign n7067 = n3740 & n7066 ;
  assign n7068 = n7064 & ~n7067 ;
  assign n7069 = n5547 & n6337 ;
  assign n7070 = n7069 ^ n3913 ^ 1'b0 ;
  assign n7071 = n1332 & n6370 ;
  assign n7072 = ( x84 & n1932 ) | ( x84 & ~n6352 ) | ( n1932 & ~n6352 ) ;
  assign n7073 = n2300 ^ n512 ^ 1'b0 ;
  assign n7074 = n7073 ^ n4823 ^ n3926 ;
  assign n7076 = ~n1350 & n1558 ;
  assign n7077 = n6352 & n7076 ;
  assign n7075 = n5034 ^ n1762 ^ 1'b0 ;
  assign n7078 = n7077 ^ n7075 ^ n1237 ;
  assign n7079 = n3263 ^ n785 ^ 1'b0 ;
  assign n7080 = n3718 | n7079 ;
  assign n7081 = n1126 | n7080 ;
  assign n7082 = n3183 & n4731 ;
  assign n7083 = n7082 ^ n4721 ^ 1'b0 ;
  assign n7084 = n1958 & ~n2915 ;
  assign n7085 = n7084 ^ n581 ^ 1'b0 ;
  assign n7086 = ( n2605 & n2770 ) | ( n2605 & ~n7085 ) | ( n2770 & ~n7085 ) ;
  assign n7087 = ~n535 & n3202 ;
  assign n7088 = n2864 ^ n2340 ^ 1'b0 ;
  assign n7089 = ( x146 & n7087 ) | ( x146 & n7088 ) | ( n7087 & n7088 ) ;
  assign n7090 = n4644 & ~n5511 ;
  assign n7091 = x199 & ~n6140 ;
  assign n7093 = n1752 ^ n1737 ^ 1'b0 ;
  assign n7094 = n2378 | n4555 ;
  assign n7095 = n7094 ^ n2658 ^ 1'b0 ;
  assign n7096 = ~x76 & n1311 ;
  assign n7097 = n4761 ^ n1608 ^ 1'b0 ;
  assign n7098 = n7097 ^ n2457 ^ 1'b0 ;
  assign n7099 = n7096 | n7098 ;
  assign n7100 = n7095 & ~n7099 ;
  assign n7101 = ~n7093 & n7100 ;
  assign n7092 = x226 & n1767 ;
  assign n7102 = n7101 ^ n7092 ^ 1'b0 ;
  assign n7103 = n4611 ^ n4480 ^ 1'b0 ;
  assign n7104 = n1643 ^ n1501 ^ 1'b0 ;
  assign n7105 = ~n7103 & n7104 ;
  assign n7106 = ( n347 & ~n2675 ) | ( n347 & n4990 ) | ( ~n2675 & n4990 ) ;
  assign n7107 = n983 | n1015 ;
  assign n7108 = x244 & n7107 ;
  assign n7109 = ~n5575 & n7108 ;
  assign n7110 = ~n7106 & n7109 ;
  assign n7111 = n7110 ^ n6197 ^ 1'b0 ;
  assign n7112 = n463 & n7111 ;
  assign n7113 = n1766 | n7112 ;
  assign n7114 = ( x43 & n4286 ) | ( x43 & ~n6337 ) | ( n4286 & ~n6337 ) ;
  assign n7115 = n2081 ^ n1033 ^ 1'b0 ;
  assign n7116 = n7115 ^ n5930 ^ n1582 ;
  assign n7117 = ~n3757 & n7116 ;
  assign n7118 = n7117 ^ n6435 ^ 1'b0 ;
  assign n7119 = n5059 ^ n3198 ^ n1486 ;
  assign n7120 = n1369 & ~n4074 ;
  assign n7121 = ~n1404 & n7120 ;
  assign n7122 = ( n504 & n2096 ) | ( n504 & ~n7121 ) | ( n2096 & ~n7121 ) ;
  assign n7123 = n1203 | n4193 ;
  assign n7124 = n2527 ^ n1134 ^ 1'b0 ;
  assign n7125 = ~n2124 & n7124 ;
  assign n7126 = n7125 ^ n1764 ^ 1'b0 ;
  assign n7127 = n261 & ~n4034 ;
  assign n7128 = n6776 ^ n4463 ^ n1980 ;
  assign n7129 = ~n4413 & n7128 ;
  assign n7130 = n7129 ^ n4223 ^ 1'b0 ;
  assign n7131 = n445 & ~n6292 ;
  assign n7132 = n7131 ^ n1052 ^ 1'b0 ;
  assign n7133 = n5040 ^ n2262 ^ 1'b0 ;
  assign n7134 = x219 & ~n7133 ;
  assign n7135 = n2138 & n7134 ;
  assign n7136 = n5094 ^ x93 ^ 1'b0 ;
  assign n7137 = n1795 & ~n7136 ;
  assign n7143 = n4839 | n5540 ;
  assign n7138 = x143 & n6604 ;
  assign n7139 = n7138 ^ n2797 ^ 1'b0 ;
  assign n7140 = n4980 ^ n1510 ^ 1'b0 ;
  assign n7141 = n7139 | n7140 ;
  assign n7142 = n5695 | n7141 ;
  assign n7144 = n7143 ^ n7142 ^ 1'b0 ;
  assign n7145 = n4878 ^ n3687 ^ n3438 ;
  assign n7146 = n979 & ~n1512 ;
  assign n7147 = n1107 & ~n7146 ;
  assign n7148 = ~n2763 & n7147 ;
  assign n7149 = n7148 ^ n7041 ^ n6021 ;
  assign n7150 = x132 & ~n1319 ;
  assign n7151 = n7150 ^ n4689 ^ 1'b0 ;
  assign n7152 = n527 & ~n5151 ;
  assign n7153 = n7151 & ~n7152 ;
  assign n7154 = ~n6102 & n7153 ;
  assign n7155 = n3705 | n6071 ;
  assign n7156 = n4600 & n7155 ;
  assign n7157 = ( n2260 & n4280 ) | ( n2260 & n5603 ) | ( n4280 & n5603 ) ;
  assign n7158 = ~n6392 & n7157 ;
  assign n7159 = n7158 ^ n449 ^ 1'b0 ;
  assign n7160 = n5660 & n7159 ;
  assign n7161 = ~n506 & n3590 ;
  assign n7163 = n5594 ^ n4694 ^ 1'b0 ;
  assign n7164 = n2972 & n7163 ;
  assign n7162 = n2972 & ~n5233 ;
  assign n7165 = n7164 ^ n7162 ^ 1'b0 ;
  assign n7166 = n3695 & ~n7165 ;
  assign n7167 = ~n7161 & n7166 ;
  assign n7168 = n263 ^ x7 ^ 1'b0 ;
  assign n7169 = n6807 & ~n7168 ;
  assign n7170 = n434 ^ x111 ^ 1'b0 ;
  assign n7171 = ( n3198 & n6871 ) | ( n3198 & n7170 ) | ( n6871 & n7170 ) ;
  assign n7172 = n2210 & n3449 ;
  assign n7173 = ~n948 & n3466 ;
  assign n7174 = n7172 & n7173 ;
  assign n7175 = n3797 | n6690 ;
  assign n7176 = n7175 ^ n2261 ^ 1'b0 ;
  assign n7177 = n4268 & n7176 ;
  assign n7178 = x75 & n7177 ;
  assign n7179 = ~n915 & n5666 ;
  assign n7180 = n5308 & n7179 ;
  assign n7181 = n463 | n7180 ;
  assign n7182 = n7181 ^ x125 ^ 1'b0 ;
  assign n7183 = n3099 | n4340 ;
  assign n7184 = n7182 | n7183 ;
  assign n7185 = n256 & ~n3435 ;
  assign n7190 = ~n1873 & n3506 ;
  assign n7186 = ( n342 & ~n1916 ) | ( n342 & n3335 ) | ( ~n1916 & n3335 ) ;
  assign n7187 = ~n1858 & n7186 ;
  assign n7188 = ~n546 & n7187 ;
  assign n7189 = n942 | n7188 ;
  assign n7191 = n7190 ^ n7189 ^ 1'b0 ;
  assign n7192 = n2237 & ~n3903 ;
  assign n7193 = n1232 & n7192 ;
  assign n7194 = n7193 ^ n397 ^ 1'b0 ;
  assign n7195 = n7194 ^ n5102 ^ 1'b0 ;
  assign n7196 = ~x101 & n7195 ;
  assign n7197 = x113 & ~x178 ;
  assign n7198 = n7197 ^ n3447 ^ 1'b0 ;
  assign n7199 = n3039 | n7198 ;
  assign n7200 = n919 & n6197 ;
  assign n7201 = n1874 | n7200 ;
  assign n7202 = n7201 ^ n2357 ^ 1'b0 ;
  assign n7203 = n7199 & n7202 ;
  assign n7204 = n7203 ^ n3513 ^ n2839 ;
  assign n7205 = n502 | n3534 ;
  assign n7206 = n7205 ^ n4622 ^ 1'b0 ;
  assign n7207 = n2345 ^ n2156 ^ 1'b0 ;
  assign n7208 = n3733 & n7207 ;
  assign n7209 = n7206 & ~n7208 ;
  assign n7210 = n4400 ^ n1995 ^ 1'b0 ;
  assign n7211 = n7210 ^ n1671 ^ 1'b0 ;
  assign n7212 = n709 ^ n589 ^ 1'b0 ;
  assign n7213 = ~n2380 & n7212 ;
  assign n7214 = n4458 ^ n3354 ^ 1'b0 ;
  assign n7215 = n7214 ^ n3433 ^ 1'b0 ;
  assign n7216 = n7213 & ~n7215 ;
  assign n7217 = ~n458 & n3693 ;
  assign n7218 = n2033 ^ n560 ^ 1'b0 ;
  assign n7219 = n1502 & n7218 ;
  assign n7220 = n7219 ^ n3645 ^ 1'b0 ;
  assign n7221 = n3504 & ~n7220 ;
  assign n7222 = n547 & ~n2443 ;
  assign n7223 = n1546 | n7222 ;
  assign n7224 = n4776 & n7223 ;
  assign n7225 = ~n7221 & n7224 ;
  assign n7226 = ( x135 & ~n2311 ) | ( x135 & n6762 ) | ( ~n2311 & n6762 ) ;
  assign n7227 = ( n601 & ~n5389 ) | ( n601 & n7226 ) | ( ~n5389 & n7226 ) ;
  assign n7228 = n3596 & ~n4578 ;
  assign n7229 = ~n666 & n7228 ;
  assign n7230 = n4126 ^ n2603 ^ 1'b0 ;
  assign n7231 = ~x22 & n2249 ;
  assign n7232 = n7230 & n7231 ;
  assign n7233 = n7229 & n7232 ;
  assign n7234 = n3767 ^ n1600 ^ 1'b0 ;
  assign n7235 = x126 & ~n7234 ;
  assign n7236 = n1097 & n2726 ;
  assign n7237 = ~n489 & n7236 ;
  assign n7238 = n2318 & ~n7237 ;
  assign n7239 = n7238 ^ n1493 ^ 1'b0 ;
  assign n7240 = n7239 ^ x61 ^ 1'b0 ;
  assign n7241 = ~n5310 & n7240 ;
  assign n7243 = ~n533 & n3594 ;
  assign n7244 = n7243 ^ n5267 ^ 1'b0 ;
  assign n7242 = n4054 & n6600 ;
  assign n7245 = n7244 ^ n7242 ^ 1'b0 ;
  assign n7246 = n7245 ^ n5765 ^ n3490 ;
  assign n7247 = ( x85 & n1295 ) | ( x85 & ~n7066 ) | ( n1295 & ~n7066 ) ;
  assign n7251 = ( ~n2006 & n3555 ) | ( ~n2006 & n3901 ) | ( n3555 & n3901 ) ;
  assign n7249 = n3480 ^ n1798 ^ 1'b0 ;
  assign n7250 = ~n4468 & n7249 ;
  assign n7248 = n5386 ^ n1369 ^ 1'b0 ;
  assign n7252 = n7251 ^ n7250 ^ n7248 ;
  assign n7253 = n5471 ^ n3242 ^ 1'b0 ;
  assign n7254 = x140 | n7253 ;
  assign n7255 = n6577 ^ n3056 ^ n572 ;
  assign n7256 = n4024 | n7255 ;
  assign n7257 = n7254 | n7256 ;
  assign n7258 = n3899 & n6726 ;
  assign n7259 = n3352 ^ x133 ^ 1'b0 ;
  assign n7260 = n7152 ^ n5993 ^ n5323 ;
  assign n7261 = n7260 ^ x44 ^ 1'b0 ;
  assign n7262 = n7261 ^ n755 ^ 1'b0 ;
  assign n7263 = n4315 ^ n3403 ^ 1'b0 ;
  assign n7264 = ( n2799 & n4739 ) | ( n2799 & ~n5534 ) | ( n4739 & ~n5534 ) ;
  assign n7265 = n7146 | n7264 ;
  assign n7270 = n4154 & ~n5290 ;
  assign n7266 = n4867 & ~n7175 ;
  assign n7267 = n4827 & n7266 ;
  assign n7268 = n838 | n7267 ;
  assign n7269 = n7268 ^ n1358 ^ 1'b0 ;
  assign n7271 = n7270 ^ n7269 ^ n5790 ;
  assign n7272 = ~n781 & n1736 ;
  assign n7273 = n7272 ^ n6016 ^ 1'b0 ;
  assign n7274 = n7115 & n7273 ;
  assign n7275 = n2590 ^ n852 ^ 1'b0 ;
  assign n7276 = n1665 & n7275 ;
  assign n7277 = n1321 & n7276 ;
  assign n7278 = n1730 & n2257 ;
  assign n7279 = n1793 & n5010 ;
  assign n7280 = n747 & n7279 ;
  assign n7281 = ( n1196 & ~n2048 ) | ( n1196 & n7280 ) | ( ~n2048 & n7280 ) ;
  assign n7282 = n4703 | n5283 ;
  assign n7283 = n1946 & ~n6012 ;
  assign n7284 = ~n2794 & n5825 ;
  assign n7285 = n2794 & n7284 ;
  assign n7286 = n2216 & ~n3248 ;
  assign n7287 = n3248 & n7286 ;
  assign n7288 = n1760 & ~n7287 ;
  assign n7289 = ~n1760 & n7288 ;
  assign n7290 = n2144 & ~n7289 ;
  assign n7291 = ~n7285 & n7290 ;
  assign n7293 = n814 ^ n274 ^ 1'b0 ;
  assign n7292 = n3577 & ~n5127 ;
  assign n7294 = n7293 ^ n7292 ^ 1'b0 ;
  assign n7295 = n7294 ^ n1332 ^ 1'b0 ;
  assign n7296 = n4174 & n7295 ;
  assign n7297 = n2046 ^ n1742 ^ 1'b0 ;
  assign n7298 = n5984 | n7126 ;
  assign n7299 = n647 & n2057 ;
  assign n7300 = ~n896 & n7299 ;
  assign n7303 = ( x42 & ~n677 ) | ( x42 & n4440 ) | ( ~n677 & n4440 ) ;
  assign n7304 = n1233 & ~n7303 ;
  assign n7305 = n7304 ^ n902 ^ 1'b0 ;
  assign n7306 = n7305 ^ n1965 ^ 1'b0 ;
  assign n7301 = n2736 & n5859 ;
  assign n7302 = n6182 & ~n7301 ;
  assign n7307 = n7306 ^ n7302 ^ 1'b0 ;
  assign n7308 = n5773 ^ n2612 ^ 1'b0 ;
  assign n7309 = n543 & n6781 ;
  assign n7310 = ~n1236 & n7309 ;
  assign n7311 = ( n5538 & n6667 ) | ( n5538 & n7310 ) | ( n6667 & n7310 ) ;
  assign n7312 = n1830 & ~n7311 ;
  assign n7313 = ~n5672 & n7312 ;
  assign n7314 = n6808 ^ n2981 ^ 1'b0 ;
  assign n7315 = n2076 | n2318 ;
  assign n7316 = n690 & ~n1717 ;
  assign n7317 = n5153 ^ n2247 ^ 1'b0 ;
  assign n7318 = ( ~n5944 & n7316 ) | ( ~n5944 & n7317 ) | ( n7316 & n7317 ) ;
  assign n7319 = n3728 & ~n5687 ;
  assign n7320 = n7319 ^ n7244 ^ 1'b0 ;
  assign n7321 = ~n747 & n7320 ;
  assign n7324 = n4451 ^ n1101 ^ 1'b0 ;
  assign n7325 = n2358 & n7324 ;
  assign n7322 = n6375 ^ n883 ^ 1'b0 ;
  assign n7323 = n7322 ^ n6460 ^ x9 ;
  assign n7326 = n7325 ^ n7323 ^ n5264 ;
  assign n7327 = n7326 ^ n6579 ^ n2054 ;
  assign n7328 = n485 ^ x62 ^ 1'b0 ;
  assign n7329 = n931 & n7328 ;
  assign n7330 = n1763 & n7329 ;
  assign n7331 = n2161 & n7330 ;
  assign n7332 = ~n308 & n3547 ;
  assign n7333 = n694 & n7332 ;
  assign n7334 = ( n2696 & n3525 ) | ( n2696 & ~n7333 ) | ( n3525 & ~n7333 ) ;
  assign n7335 = n7334 ^ n2421 ^ 1'b0 ;
  assign n7336 = n2797 ^ n1158 ^ 1'b0 ;
  assign n7337 = ( ~n1253 & n3094 ) | ( ~n1253 & n5432 ) | ( n3094 & n5432 ) ;
  assign n7338 = n1360 & n1504 ;
  assign n7339 = n2881 & n7338 ;
  assign n7340 = x11 & n7339 ;
  assign n7341 = n7337 & n7340 ;
  assign n7342 = n519 ^ x150 ^ 1'b0 ;
  assign n7343 = x213 & n5003 ;
  assign n7344 = ~n7342 & n7343 ;
  assign n7345 = n1150 & ~n1346 ;
  assign n7346 = ~n7144 & n7345 ;
  assign n7347 = n3642 | n3662 ;
  assign n7348 = n867 & ~n7347 ;
  assign n7349 = ~n2984 & n3271 ;
  assign n7350 = ~n7348 & n7349 ;
  assign n7351 = n7350 ^ n4521 ^ 1'b0 ;
  assign n7352 = n5807 | n7351 ;
  assign n7355 = n3557 ^ n2299 ^ 1'b0 ;
  assign n7356 = ~n3984 & n7355 ;
  assign n7357 = n1429 ^ n972 ^ 1'b0 ;
  assign n7358 = ~n6152 & n7357 ;
  assign n7359 = ( n3088 & n7356 ) | ( n3088 & n7358 ) | ( n7356 & n7358 ) ;
  assign n7353 = n1212 & n5192 ;
  assign n7354 = n7353 ^ n5519 ^ 1'b0 ;
  assign n7360 = n7359 ^ n7354 ^ 1'b0 ;
  assign n7361 = n2397 ^ n259 ^ 1'b0 ;
  assign n7362 = ~n4029 & n7361 ;
  assign n7363 = n674 & ~n7362 ;
  assign n7364 = n1625 ^ n631 ^ 1'b0 ;
  assign n7365 = ~n6646 & n7364 ;
  assign n7366 = n4220 ^ n1732 ^ 1'b0 ;
  assign n7367 = n4259 & n7366 ;
  assign n7368 = ~n2412 & n7367 ;
  assign n7369 = n7368 ^ n3894 ^ 1'b0 ;
  assign n7370 = n5006 | n5294 ;
  assign n7371 = n358 & ~n842 ;
  assign n7372 = ~n4781 & n7371 ;
  assign n7373 = n2922 ^ n1842 ^ 1'b0 ;
  assign n7374 = n7372 | n7373 ;
  assign n7375 = n4264 | n7067 ;
  assign n7376 = n3973 & ~n7375 ;
  assign n7377 = ( ~n802 & n1577 ) | ( ~n802 & n5305 ) | ( n1577 & n5305 ) ;
  assign n7378 = ~x247 & n2285 ;
  assign n7379 = n5699 & n7378 ;
  assign n7380 = n7379 ^ n5567 ^ 1'b0 ;
  assign n7382 = n3651 ^ n1470 ^ n432 ;
  assign n7381 = n7010 ^ n575 ^ 1'b0 ;
  assign n7383 = n7382 ^ n7381 ^ n2973 ;
  assign n7384 = n7383 ^ n6960 ^ n5945 ;
  assign n7385 = n7384 ^ n5398 ^ 1'b0 ;
  assign n7389 = ~n5473 & n5769 ;
  assign n7386 = x29 & n2642 ;
  assign n7387 = n3055 & n7386 ;
  assign n7388 = n2915 | n7387 ;
  assign n7390 = n7389 ^ n7388 ^ 1'b0 ;
  assign n7391 = n4012 | n5261 ;
  assign n7392 = ( n3526 & ~n4196 ) | ( n3526 & n4808 ) | ( ~n4196 & n4808 ) ;
  assign n7393 = n918 & n7392 ;
  assign n7394 = ( ~n797 & n7261 ) | ( ~n797 & n7393 ) | ( n7261 & n7393 ) ;
  assign n7395 = ~n1026 & n1235 ;
  assign n7396 = n7395 ^ n3369 ^ 1'b0 ;
  assign n7397 = n4915 ^ n4272 ^ 1'b0 ;
  assign n7398 = x174 & n7397 ;
  assign n7399 = n7398 ^ n790 ^ 1'b0 ;
  assign n7400 = n5639 ^ n1430 ^ x117 ;
  assign n7401 = ~n947 & n1963 ;
  assign n7402 = n4218 ^ n2026 ^ 1'b0 ;
  assign n7403 = ( ~n2979 & n7401 ) | ( ~n2979 & n7402 ) | ( n7401 & n7402 ) ;
  assign n7404 = n1631 ^ n791 ^ 1'b0 ;
  assign n7405 = n7404 ^ n1489 ^ 1'b0 ;
  assign n7406 = n4652 ^ n3409 ^ 1'b0 ;
  assign n7407 = n3093 ^ n635 ^ 1'b0 ;
  assign n7408 = ( x26 & n7406 ) | ( x26 & n7407 ) | ( n7406 & n7407 ) ;
  assign n7409 = n2010 & ~n7408 ;
  assign n7410 = n2726 ^ n429 ^ 1'b0 ;
  assign n7411 = ~n1148 & n7410 ;
  assign n7412 = n1086 & n4966 ;
  assign n7413 = n880 & n7412 ;
  assign n7414 = n3821 | n7413 ;
  assign n7415 = n6956 | n7414 ;
  assign n7416 = n1206 & n3737 ;
  assign n7417 = ~n633 & n7416 ;
  assign n7418 = ( n3659 & n3908 ) | ( n3659 & n7417 ) | ( n3908 & n7417 ) ;
  assign n7419 = n984 & n1393 ;
  assign n7420 = ~n7418 & n7419 ;
  assign n7421 = ~n1037 & n4259 ;
  assign n7422 = n7421 ^ n1833 ^ 1'b0 ;
  assign n7423 = n2843 | n7422 ;
  assign n7424 = n6100 ^ n3727 ^ 1'b0 ;
  assign n7425 = n1808 | n7057 ;
  assign n7426 = n2111 | n7425 ;
  assign n7427 = n6322 ^ n2558 ^ 1'b0 ;
  assign n7428 = ~n5634 & n7427 ;
  assign n7429 = n6307 ^ n2158 ^ 1'b0 ;
  assign n7430 = n6121 ^ n3459 ^ 1'b0 ;
  assign n7431 = n1550 & n7430 ;
  assign n7432 = ~n1137 & n1919 ;
  assign n7433 = n7432 ^ n562 ^ 1'b0 ;
  assign n7434 = n7244 & n7433 ;
  assign n7435 = ~x130 & n7434 ;
  assign n7436 = n3369 & ~n7435 ;
  assign n7437 = n4890 ^ n2005 ^ 1'b0 ;
  assign n7438 = n4214 & ~n7437 ;
  assign n7439 = n7438 ^ n1982 ^ 1'b0 ;
  assign n7440 = n5986 ^ n2156 ^ 1'b0 ;
  assign n7443 = n4077 ^ n2291 ^ 1'b0 ;
  assign n7441 = n2006 & n4091 ;
  assign n7442 = n559 & n7441 ;
  assign n7444 = n7443 ^ n7442 ^ 1'b0 ;
  assign n7445 = ( n6459 & ~n7440 ) | ( n6459 & n7444 ) | ( ~n7440 & n7444 ) ;
  assign n7446 = n594 & ~n3666 ;
  assign n7447 = n5769 & n7446 ;
  assign n7448 = n7447 ^ n650 ^ 1'b0 ;
  assign n7449 = n1209 & ~n5616 ;
  assign n7450 = ~n486 & n7449 ;
  assign n7451 = ~n904 & n6079 ;
  assign n7452 = n7451 ^ n5970 ^ 1'b0 ;
  assign n7453 = n702 & n5721 ;
  assign n7454 = n4216 ^ n4174 ^ n569 ;
  assign n7455 = n7454 ^ n1023 ^ x88 ;
  assign n7456 = n1327 & n6406 ;
  assign n7457 = n7455 & n7456 ;
  assign n7458 = n2065 & n3579 ;
  assign n7459 = x230 & n4031 ;
  assign n7460 = ~n1184 & n7459 ;
  assign n7461 = n4278 ^ n3369 ^ 1'b0 ;
  assign n7462 = n7460 | n7461 ;
  assign n7463 = n7458 & ~n7462 ;
  assign n7464 = n7204 ^ n7053 ^ n4872 ;
  assign n7465 = n5363 ^ n2855 ^ 1'b0 ;
  assign n7466 = n2630 ^ n2292 ^ 1'b0 ;
  assign n7467 = n972 | n7466 ;
  assign n7468 = n7467 ^ n5541 ^ 1'b0 ;
  assign n7469 = n6003 ^ n5230 ^ n3504 ;
  assign n7470 = n6927 | n7469 ;
  assign n7471 = n7468 & ~n7470 ;
  assign n7472 = n1325 ^ n865 ^ 1'b0 ;
  assign n7473 = n1716 & n7472 ;
  assign n7474 = n2991 & n7473 ;
  assign n7475 = n4710 ^ n3756 ^ 1'b0 ;
  assign n7476 = ( ~n3271 & n7474 ) | ( ~n3271 & n7475 ) | ( n7474 & n7475 ) ;
  assign n7477 = n3718 ^ n663 ^ x239 ;
  assign n7478 = n7477 ^ n5569 ^ 1'b0 ;
  assign n7479 = ~n4123 & n7478 ;
  assign n7480 = n7479 ^ n4726 ^ 1'b0 ;
  assign n7481 = n873 & n4550 ;
  assign n7482 = n3958 ^ n1140 ^ 1'b0 ;
  assign n7483 = n7482 ^ n6834 ^ 1'b0 ;
  assign n7484 = n7481 | n7483 ;
  assign n7485 = ~n5519 & n7096 ;
  assign n7486 = x98 & ~n5038 ;
  assign n7487 = ~n3096 & n7486 ;
  assign n7488 = n7487 ^ n2286 ^ n2009 ;
  assign n7489 = n7488 ^ n6888 ^ n4187 ;
  assign n7491 = x76 & ~n3723 ;
  assign n7492 = ~n4249 & n7491 ;
  assign n7493 = n7492 ^ n6417 ^ 1'b0 ;
  assign n7494 = n2521 & n7493 ;
  assign n7495 = n3414 & n7494 ;
  assign n7496 = x119 ^ x35 ^ 1'b0 ;
  assign n7497 = ~n1308 & n7496 ;
  assign n7498 = n3551 & n7497 ;
  assign n7499 = ~n7495 & n7498 ;
  assign n7490 = n471 ^ n397 ^ 1'b0 ;
  assign n7500 = n7499 ^ n7490 ^ 1'b0 ;
  assign n7501 = ( ~n587 & n2125 ) | ( ~n587 & n2164 ) | ( n2125 & n2164 ) ;
  assign n7502 = n6842 | n7174 ;
  assign n7503 = n7502 ^ x124 ^ 1'b0 ;
  assign n7504 = x55 & n7503 ;
  assign n7505 = n7501 & n7504 ;
  assign n7506 = n4553 ^ x179 ^ 1'b0 ;
  assign n7507 = ~n623 & n7506 ;
  assign n7508 = n599 & n3021 ;
  assign n7509 = n7508 ^ n2749 ^ 1'b0 ;
  assign n7510 = n7509 ^ n1365 ^ 1'b0 ;
  assign n7511 = n7510 ^ n4852 ^ 1'b0 ;
  assign n7512 = n881 | n7511 ;
  assign n7513 = ~n824 & n1107 ;
  assign n7514 = n7513 ^ n2632 ^ 1'b0 ;
  assign n7515 = n2823 & n7514 ;
  assign n7516 = n5546 ^ n1761 ^ 1'b0 ;
  assign n7517 = n455 | n7516 ;
  assign n7518 = ( n5841 & n7515 ) | ( n5841 & ~n7517 ) | ( n7515 & ~n7517 ) ;
  assign n7519 = n2341 | n5887 ;
  assign n7520 = n7519 ^ n3239 ^ 1'b0 ;
  assign n7521 = n7520 ^ n4084 ^ n1978 ;
  assign n7522 = n3806 ^ x202 ^ 1'b0 ;
  assign n7523 = n7301 ^ n4647 ^ 1'b0 ;
  assign n7524 = n7523 ^ n1396 ^ 1'b0 ;
  assign n7525 = n6868 | n7524 ;
  assign n7526 = n7161 ^ n3842 ^ 1'b0 ;
  assign n7527 = n5540 | n7526 ;
  assign n7528 = n3647 ^ n473 ^ 1'b0 ;
  assign n7529 = n7487 | n7528 ;
  assign n7530 = ~n7527 & n7529 ;
  assign n7531 = n842 | n5019 ;
  assign n7532 = n401 | n1695 ;
  assign n7533 = ( n4236 & n7531 ) | ( n4236 & n7532 ) | ( n7531 & n7532 ) ;
  assign n7534 = n3680 & n7533 ;
  assign n7535 = ~x159 & n3043 ;
  assign n7536 = ~x81 & x142 ;
  assign n7537 = x22 & ~n7306 ;
  assign n7538 = ~n7536 & n7537 ;
  assign n7539 = n1343 | n4779 ;
  assign n7540 = n5588 | n7303 ;
  assign n7541 = n7539 | n7540 ;
  assign n7542 = n7541 ^ n5477 ^ 1'b0 ;
  assign n7543 = n4320 ^ x94 ^ 1'b0 ;
  assign n7544 = n7543 ^ n4072 ^ 1'b0 ;
  assign n7545 = n7544 ^ n5157 ^ 1'b0 ;
  assign n7546 = ~n335 & n7545 ;
  assign n7551 = x240 & n484 ;
  assign n7552 = n7551 ^ x4 ^ 1'b0 ;
  assign n7553 = n3949 | n7552 ;
  assign n7554 = n7553 ^ n4544 ^ 1'b0 ;
  assign n7547 = n1293 | n1677 ;
  assign n7548 = x143 & n7547 ;
  assign n7549 = n3048 & n7548 ;
  assign n7550 = n4479 | n7549 ;
  assign n7555 = n7554 ^ n7550 ^ 1'b0 ;
  assign n7556 = n2006 | n4015 ;
  assign n7557 = n7555 & ~n7556 ;
  assign n7558 = n6221 & n7557 ;
  assign n7559 = n2786 ^ n1467 ^ 1'b0 ;
  assign n7560 = n3587 & n7559 ;
  assign n7567 = n3666 ^ x240 ^ 1'b0 ;
  assign n7563 = ~n1019 & n6411 ;
  assign n7564 = ~n984 & n7563 ;
  assign n7561 = n1655 | n5070 ;
  assign n7562 = n555 | n7561 ;
  assign n7565 = n7564 ^ n7562 ^ n2895 ;
  assign n7566 = n570 & n7565 ;
  assign n7568 = n7567 ^ n7566 ^ 1'b0 ;
  assign n7569 = ( ~n1215 & n1295 ) | ( ~n1215 & n4435 ) | ( n1295 & n4435 ) ;
  assign n7570 = n6352 & n7569 ;
  assign n7571 = n1271 | n4925 ;
  assign n7572 = n5739 & ~n7571 ;
  assign n7573 = ~n2070 & n4058 ;
  assign n7574 = n7185 ^ n3897 ^ 1'b0 ;
  assign n7575 = n7573 & ~n7574 ;
  assign n7576 = n6800 | n7469 ;
  assign n7577 = n4661 ^ n1645 ^ n832 ;
  assign n7578 = ( x101 & n1876 ) | ( x101 & ~n7577 ) | ( n1876 & ~n7577 ) ;
  assign n7579 = n337 | n7578 ;
  assign n7580 = n383 | n7579 ;
  assign n7581 = ~n6641 & n7580 ;
  assign n7582 = n5725 ^ n3195 ^ 1'b0 ;
  assign n7583 = n1006 & n7582 ;
  assign n7584 = ~x222 & n3383 ;
  assign n7585 = n7584 ^ n7314 ^ 1'b0 ;
  assign n7600 = n3308 | n5341 ;
  assign n7597 = ~n942 & n1701 ;
  assign n7598 = n7597 ^ n5210 ^ n4620 ;
  assign n7586 = n5510 ^ n1451 ^ 1'b0 ;
  assign n7587 = n2335 & ~n7586 ;
  assign n7588 = ~n4483 & n7587 ;
  assign n7589 = n7588 ^ n1981 ^ 1'b0 ;
  assign n7590 = n539 & n1190 ;
  assign n7591 = n737 & n4574 ;
  assign n7592 = ~n4574 & n7591 ;
  assign n7593 = n7592 ^ n6045 ^ n2720 ;
  assign n7594 = n7590 & ~n7593 ;
  assign n7595 = ~n5040 & n7594 ;
  assign n7596 = n7589 | n7595 ;
  assign n7599 = n7598 ^ n7596 ^ 1'b0 ;
  assign n7601 = n7600 ^ n7599 ^ n1315 ;
  assign n7602 = n6172 ^ n4046 ^ 1'b0 ;
  assign n7603 = n5338 ^ n3678 ^ x164 ;
  assign n7604 = n7225 | n7603 ;
  assign n7607 = ( n872 & ~n3183 ) | ( n872 & n3817 ) | ( ~n3183 & n3817 ) ;
  assign n7605 = n5184 ^ n4507 ^ 1'b0 ;
  assign n7606 = ~n527 & n7605 ;
  assign n7608 = n7607 ^ n7606 ^ 1'b0 ;
  assign n7609 = n4626 | n7608 ;
  assign n7610 = n5527 ^ n265 ^ 1'b0 ;
  assign n7611 = n2243 & ~n7610 ;
  assign n7612 = ( ~n1872 & n3673 ) | ( ~n1872 & n4513 ) | ( n3673 & n4513 ) ;
  assign n7613 = n7612 ^ n4115 ^ n1033 ;
  assign n7614 = n7613 ^ n4710 ^ 1'b0 ;
  assign n7615 = n2315 & ~n7614 ;
  assign n7616 = n2816 & n7615 ;
  assign n7617 = n2259 & ~n7616 ;
  assign n7618 = ~n4713 & n7617 ;
  assign n7619 = ~n7611 & n7618 ;
  assign n7620 = n1653 | n7283 ;
  assign n7621 = n7620 ^ n1097 ^ 1'b0 ;
  assign n7622 = n7621 ^ n2519 ^ 1'b0 ;
  assign n7623 = n5289 ^ x183 ^ 1'b0 ;
  assign n7624 = n2649 | n7623 ;
  assign n7625 = x9 & ~n954 ;
  assign n7626 = n7624 & n7625 ;
  assign n7627 = n1091 | n7626 ;
  assign n7628 = n4435 ^ n438 ^ 1'b0 ;
  assign n7629 = x254 & n7628 ;
  assign n7630 = ( n478 & ~n833 ) | ( n478 & n7629 ) | ( ~n833 & n7629 ) ;
  assign n7631 = x7 & n412 ;
  assign n7632 = n7631 ^ n3747 ^ 1'b0 ;
  assign n7633 = n7632 ^ n647 ^ 1'b0 ;
  assign n7635 = n1376 ^ n946 ^ 1'b0 ;
  assign n7636 = n1991 & n7635 ;
  assign n7634 = n1630 | n2751 ;
  assign n7637 = n7636 ^ n7634 ^ 1'b0 ;
  assign n7642 = x78 & x189 ;
  assign n7643 = n7642 ^ n1407 ^ 1'b0 ;
  assign n7640 = x166 & ~n5613 ;
  assign n7641 = n7640 ^ n402 ^ 1'b0 ;
  assign n7638 = n2922 ^ n635 ^ 1'b0 ;
  assign n7639 = n887 & n7638 ;
  assign n7644 = n7643 ^ n7641 ^ n7639 ;
  assign n7645 = ( n2699 & ~n7637 ) | ( n2699 & n7644 ) | ( ~n7637 & n7644 ) ;
  assign n7646 = n5848 ^ n1263 ^ 1'b0 ;
  assign n7647 = n7646 ^ x150 ^ 1'b0 ;
  assign n7648 = n469 & n1926 ;
  assign n7649 = n7648 ^ n3911 ^ 1'b0 ;
  assign n7650 = n7649 ^ n803 ^ 1'b0 ;
  assign n7651 = n2101 ^ n1758 ^ n1509 ;
  assign n7652 = n3884 ^ x159 ^ 1'b0 ;
  assign n7653 = n7651 & ~n7652 ;
  assign n7654 = ~n5242 & n7653 ;
  assign n7655 = n459 | n7654 ;
  assign n7656 = n7655 ^ n580 ^ 1'b0 ;
  assign n7658 = n1006 & n5170 ;
  assign n7659 = n6147 & n7658 ;
  assign n7660 = n7659 ^ n6960 ^ 1'b0 ;
  assign n7657 = n2586 & ~n5013 ;
  assign n7661 = n7660 ^ n7657 ^ 1'b0 ;
  assign n7662 = x153 & ~n7661 ;
  assign n7663 = n7662 ^ n5021 ^ 1'b0 ;
  assign n7664 = n1098 & n5660 ;
  assign n7665 = n7329 ^ n2686 ^ n1785 ;
  assign n7666 = n3918 | n7665 ;
  assign n7667 = n7666 ^ n5835 ^ x201 ;
  assign n7668 = n3007 ^ n347 ^ 1'b0 ;
  assign n7669 = n7668 ^ n1347 ^ 1'b0 ;
  assign n7670 = ~n4023 & n7669 ;
  assign n7671 = n7670 ^ n4435 ^ 1'b0 ;
  assign n7672 = n4047 ^ n2392 ^ n1071 ;
  assign n7673 = n7672 ^ n865 ^ 1'b0 ;
  assign n7674 = n5338 ^ n5224 ^ n1788 ;
  assign n7675 = n7674 ^ n1081 ^ 1'b0 ;
  assign n7676 = n7675 ^ n5720 ^ 1'b0 ;
  assign n7677 = n7673 & ~n7676 ;
  assign n7678 = n4154 ^ n2719 ^ x164 ;
  assign n7679 = n7678 ^ n3986 ^ 1'b0 ;
  assign n7680 = ~n6405 & n7641 ;
  assign n7681 = ~n3639 & n6412 ;
  assign n7682 = n7681 ^ n7002 ^ 1'b0 ;
  assign n7683 = n4548 ^ n3552 ^ 1'b0 ;
  assign n7687 = n3534 ^ x133 ^ 1'b0 ;
  assign n7684 = n1519 & n2048 ;
  assign n7685 = n7684 ^ x112 ^ 1'b0 ;
  assign n7686 = n1797 | n7685 ;
  assign n7688 = n7687 ^ n7686 ^ 1'b0 ;
  assign n7689 = ~n789 & n3970 ;
  assign n7690 = ~n2276 & n7689 ;
  assign n7691 = ~n4287 & n7690 ;
  assign n7692 = n5934 & ~n7691 ;
  assign n7693 = n4995 & n7692 ;
  assign n7694 = n2305 | n7693 ;
  assign n7695 = n2958 | n3979 ;
  assign n7696 = ( n4909 & n7630 ) | ( n4909 & n7695 ) | ( n7630 & n7695 ) ;
  assign n7697 = n1170 | n2127 ;
  assign n7698 = n7697 ^ n5762 ^ 1'b0 ;
  assign n7699 = n5108 & ~n7698 ;
  assign n7700 = ~n4080 & n7699 ;
  assign n7701 = ~x122 & n832 ;
  assign n7702 = n939 & ~n3573 ;
  assign n7703 = n7702 ^ n1626 ^ 1'b0 ;
  assign n7704 = n7703 ^ n4703 ^ 1'b0 ;
  assign n7705 = n4281 & n7704 ;
  assign n7706 = n7705 ^ n849 ^ 1'b0 ;
  assign n7708 = n6015 ^ n5096 ^ 1'b0 ;
  assign n7707 = n3627 ^ n2877 ^ 1'b0 ;
  assign n7709 = n7708 ^ n7707 ^ n5667 ;
  assign n7710 = n2575 & n7709 ;
  assign n7711 = ~x153 & n3783 ;
  assign n7712 = n3061 & n4500 ;
  assign n7713 = ~n1470 & n7712 ;
  assign n7714 = n2785 ^ n1998 ^ 1'b0 ;
  assign n7715 = ( x49 & n315 ) | ( x49 & n1846 ) | ( n315 & n1846 ) ;
  assign n7716 = ~n3124 & n5725 ;
  assign n7717 = n3853 & ~n6458 ;
  assign n7718 = n7717 ^ n4719 ^ 1'b0 ;
  assign n7719 = n1953 & ~n5869 ;
  assign n7720 = n5963 ^ n2476 ^ 1'b0 ;
  assign n7721 = ~n1596 & n7720 ;
  assign n7722 = n755 & n7721 ;
  assign n7723 = n7722 ^ n3557 ^ 1'b0 ;
  assign n7725 = ~n1515 & n2309 ;
  assign n7726 = n3343 & n7725 ;
  assign n7724 = n3215 ^ n2642 ^ x182 ;
  assign n7727 = n7726 ^ n7724 ^ 1'b0 ;
  assign n7728 = n5216 ^ n2543 ^ 1'b0 ;
  assign n7729 = n4132 | n7728 ;
  assign n7730 = n2469 | n3761 ;
  assign n7731 = n7730 ^ n6964 ^ 1'b0 ;
  assign n7732 = n7731 ^ n7344 ^ n4998 ;
  assign n7734 = n2471 | n2598 ;
  assign n7733 = ~n2036 & n2922 ;
  assign n7735 = n7734 ^ n7733 ^ 1'b0 ;
  assign n7736 = n1344 & n7521 ;
  assign n7737 = n7736 ^ n5637 ^ 1'b0 ;
  assign n7738 = ~n512 & n7260 ;
  assign n7739 = n3600 & n7738 ;
  assign n7740 = n7612 ^ n7501 ^ 1'b0 ;
  assign n7741 = n2580 & ~n7740 ;
  assign n7744 = n6811 ^ n2561 ^ 1'b0 ;
  assign n7745 = n4947 | n7744 ;
  assign n7742 = n6756 ^ x208 ^ 1'b0 ;
  assign n7743 = ~n2547 & n7742 ;
  assign n7746 = n7745 ^ n7743 ^ 1'b0 ;
  assign n7747 = n3912 & ~n5077 ;
  assign n7748 = ~n2882 & n7747 ;
  assign n7749 = n7748 ^ n3395 ^ 1'b0 ;
  assign n7750 = n3135 ^ n1892 ^ 1'b0 ;
  assign n7751 = n2804 & n3102 ;
  assign n7752 = n5816 & n7751 ;
  assign n7753 = ( n3672 & ~n5175 ) | ( n3672 & n7752 ) | ( ~n5175 & n7752 ) ;
  assign n7754 = n3399 | n4211 ;
  assign n7755 = n2182 | n6244 ;
  assign n7756 = n6193 | n6203 ;
  assign n7757 = n7755 | n7756 ;
  assign n7758 = n7754 & ~n7757 ;
  assign n7760 = ( ~n1004 & n1657 ) | ( ~n1004 & n3737 ) | ( n1657 & n3737 ) ;
  assign n7759 = ~n6169 & n6964 ;
  assign n7761 = n7760 ^ n7759 ^ 1'b0 ;
  assign n7762 = n2390 | n2404 ;
  assign n7763 = n4563 | n7762 ;
  assign n7764 = x109 | n7763 ;
  assign n7765 = n5463 & n7764 ;
  assign n7766 = n2718 ^ n1598 ^ 1'b0 ;
  assign n7768 = n979 ^ n672 ^ 1'b0 ;
  assign n7769 = n7567 | n7768 ;
  assign n7767 = n432 & ~n1342 ;
  assign n7770 = n7769 ^ n7767 ^ 1'b0 ;
  assign n7771 = n6677 & n7770 ;
  assign n7772 = n6303 ^ x118 ^ 1'b0 ;
  assign n7773 = n1145 & n7772 ;
  assign n7774 = n7773 ^ n1378 ^ 1'b0 ;
  assign n7775 = n2488 & n7774 ;
  assign n7776 = n2389 & n7775 ;
  assign n7777 = n2686 & ~n4193 ;
  assign n7779 = n2707 ^ x59 ^ 1'b0 ;
  assign n7780 = ~n1712 & n7779 ;
  assign n7781 = n1127 | n7780 ;
  assign n7778 = x120 | n5361 ;
  assign n7782 = n7781 ^ n7778 ^ n6359 ;
  assign n7783 = n6792 | n7782 ;
  assign n7784 = n1084 | n7783 ;
  assign n7785 = n7784 ^ n854 ^ 1'b0 ;
  assign n7786 = ( ~x7 & n600 ) | ( ~x7 & n7785 ) | ( n600 & n7785 ) ;
  assign n7788 = ( n1343 & n2670 ) | ( n1343 & n3707 ) | ( n2670 & n3707 ) ;
  assign n7787 = n5603 ^ n2871 ^ n2219 ;
  assign n7789 = n7788 ^ n7787 ^ 1'b0 ;
  assign n7790 = ~n3513 & n7789 ;
  assign n7791 = n4823 & ~n7477 ;
  assign n7792 = n2539 | n4957 ;
  assign n7793 = x71 | n7792 ;
  assign n7794 = n7619 ^ n4302 ^ 1'b0 ;
  assign n7795 = ( n702 & n6379 ) | ( n702 & ~n7644 ) | ( n6379 & ~n7644 ) ;
  assign n7796 = ~x107 & n2966 ;
  assign n7797 = n7796 ^ n6451 ^ n2979 ;
  assign n7798 = n7797 ^ n7690 ^ 1'b0 ;
  assign n7803 = n6214 ^ x119 ^ 1'b0 ;
  assign n7804 = n5121 & ~n7803 ;
  assign n7800 = n1396 ^ n933 ^ 1'b0 ;
  assign n7801 = x181 & n7800 ;
  assign n7799 = n7157 ^ n2135 ^ n803 ;
  assign n7802 = n7801 ^ n7799 ^ n2131 ;
  assign n7805 = n7804 ^ n7802 ^ 1'b0 ;
  assign n7806 = n7805 ^ n5613 ^ n5054 ;
  assign n7807 = ~n706 & n5746 ;
  assign n7809 = n2207 & ~n2548 ;
  assign n7808 = n3911 & ~n4358 ;
  assign n7810 = n7809 ^ n7808 ^ 1'b0 ;
  assign n7811 = ~n2528 & n7810 ;
  assign n7812 = n5103 ^ n4010 ^ 1'b0 ;
  assign n7813 = ( n7807 & ~n7811 ) | ( n7807 & n7812 ) | ( ~n7811 & n7812 ) ;
  assign n7814 = ~n2856 & n7789 ;
  assign n7819 = x36 & n3423 ;
  assign n7820 = n369 & n7819 ;
  assign n7816 = n1297 & ~n1863 ;
  assign n7817 = ~n635 & n7816 ;
  assign n7818 = n2414 | n7817 ;
  assign n7821 = n7820 ^ n7818 ^ 1'b0 ;
  assign n7815 = n4649 | n5449 ;
  assign n7822 = n7821 ^ n7815 ^ 1'b0 ;
  assign n7823 = n2915 ^ n2537 ^ n1871 ;
  assign n7824 = x182 | n7823 ;
  assign n7825 = n3234 & n6386 ;
  assign n7826 = ~n7824 & n7825 ;
  assign n7827 = n3551 & n4509 ;
  assign n7828 = ~n6944 & n7827 ;
  assign n7829 = n7828 ^ n4998 ^ 1'b0 ;
  assign n7830 = ~n7826 & n7829 ;
  assign n7831 = n7830 ^ n6520 ^ n4994 ;
  assign n7843 = n3646 ^ n455 ^ 1'b0 ;
  assign n7834 = n6579 ^ n2250 ^ 1'b0 ;
  assign n7835 = n304 | n3886 ;
  assign n7836 = n7835 ^ x180 ^ 1'b0 ;
  assign n7837 = ~n476 & n7836 ;
  assign n7838 = ~n3259 & n7837 ;
  assign n7839 = n7838 ^ n2059 ^ 1'b0 ;
  assign n7840 = n1850 & ~n7839 ;
  assign n7841 = n7840 ^ n2951 ^ 1'b0 ;
  assign n7842 = ( n2172 & n7834 ) | ( n2172 & n7841 ) | ( n7834 & n7841 ) ;
  assign n7832 = n1088 & ~n1376 ;
  assign n7833 = n7832 ^ n624 ^ 1'b0 ;
  assign n7844 = n7843 ^ n7842 ^ n7833 ;
  assign n7845 = ~n3584 & n5729 ;
  assign n7846 = n7844 & n7845 ;
  assign n7847 = n1502 & ~n4535 ;
  assign n7848 = n7847 ^ n3233 ^ 1'b0 ;
  assign n7849 = x179 & ~n7848 ;
  assign n7850 = ~n2028 & n2737 ;
  assign n7851 = n7850 ^ n4021 ^ 1'b0 ;
  assign n7852 = x35 & n7851 ;
  assign n7853 = ( n535 & n7849 ) | ( n535 & n7852 ) | ( n7849 & n7852 ) ;
  assign n7854 = n4026 | n6895 ;
  assign n7855 = x213 & n1914 ;
  assign n7856 = n1212 & n7855 ;
  assign n7857 = n2537 ^ n1781 ^ n935 ;
  assign n7858 = n6488 | n7857 ;
  assign n7859 = ( ~n2597 & n7856 ) | ( ~n2597 & n7858 ) | ( n7856 & n7858 ) ;
  assign n7860 = n5684 & n7859 ;
  assign n7861 = n2748 ^ n1007 ^ 1'b0 ;
  assign n7862 = n7860 & n7861 ;
  assign n7863 = n7862 ^ n2864 ^ 1'b0 ;
  assign n7864 = ( ~n3297 & n6484 ) | ( ~n3297 & n7863 ) | ( n6484 & n7863 ) ;
  assign n7865 = ~n1865 & n5430 ;
  assign n7866 = ~n1130 & n7865 ;
  assign n7868 = x200 & n372 ;
  assign n7869 = n7868 ^ n441 ^ 1'b0 ;
  assign n7867 = n5157 ^ n806 ^ 1'b0 ;
  assign n7870 = n7869 ^ n7867 ^ 1'b0 ;
  assign n7871 = n4253 ^ n2261 ^ 1'b0 ;
  assign n7872 = n6389 ^ n5127 ^ 1'b0 ;
  assign n7873 = n7871 | n7872 ;
  assign n7874 = n392 & ~n3852 ;
  assign n7875 = n7874 ^ n7839 ^ 1'b0 ;
  assign n7876 = n7875 ^ n5880 ^ n1862 ;
  assign n7877 = ( ~x244 & n553 ) | ( ~x244 & n1350 ) | ( n553 & n1350 ) ;
  assign n7878 = n5550 & n7877 ;
  assign n7879 = n7878 ^ n835 ^ 1'b0 ;
  assign n7880 = n902 & n2636 ;
  assign n7881 = n5588 ^ n3365 ^ 1'b0 ;
  assign n7882 = n7881 ^ n3124 ^ 1'b0 ;
  assign n7883 = n7880 & ~n7882 ;
  assign n7884 = n4657 ^ n4124 ^ 1'b0 ;
  assign n7885 = ~n3489 & n7884 ;
  assign n7886 = n3388 & n7885 ;
  assign n7887 = n5713 ^ x188 ^ 1'b0 ;
  assign n7888 = n1630 & n2390 ;
  assign n7889 = n7888 ^ n329 ^ 1'b0 ;
  assign n7890 = ~n2463 & n7889 ;
  assign n7891 = ~n1321 & n5549 ;
  assign n7892 = ~n7890 & n7891 ;
  assign n7893 = n7892 ^ n5055 ^ 1'b0 ;
  assign n7894 = n732 & ~n7893 ;
  assign n7895 = n7894 ^ n2832 ^ n275 ;
  assign n7896 = n541 | n2155 ;
  assign n7897 = n4787 | n7896 ;
  assign n7898 = ~n4216 & n7897 ;
  assign n7899 = n7898 ^ n6725 ^ 1'b0 ;
  assign n7900 = n4259 | n6700 ;
  assign n7901 = n7900 ^ n4168 ^ 1'b0 ;
  assign n7902 = n7564 ^ n3438 ^ n2224 ;
  assign n7903 = n7902 ^ n7764 ^ n2800 ;
  assign n7904 = ~n4926 & n7073 ;
  assign n7905 = n7904 ^ n2730 ^ 1'b0 ;
  assign n7906 = n519 & n6988 ;
  assign n7907 = n758 ^ x156 ^ 1'b0 ;
  assign n7908 = n2344 & ~n7907 ;
  assign n7909 = n5824 ^ n1464 ^ 1'b0 ;
  assign n7910 = ( n634 & n7908 ) | ( n634 & n7909 ) | ( n7908 & n7909 ) ;
  assign n7911 = n5962 ^ n781 ^ 1'b0 ;
  assign n7912 = ~n7910 & n7911 ;
  assign n7913 = n1955 ^ n539 ^ 1'b0 ;
  assign n7914 = n1416 & ~n1882 ;
  assign n7915 = ( n1103 & ~n7913 ) | ( n1103 & n7914 ) | ( ~n7913 & n7914 ) ;
  assign n7916 = ~n752 & n4034 ;
  assign n7917 = n7916 ^ n374 ^ 1'b0 ;
  assign n7918 = ~n5806 & n7917 ;
  assign n7919 = n4860 ^ n3788 ^ 1'b0 ;
  assign n7920 = n1105 | n3499 ;
  assign n7921 = n7919 | n7920 ;
  assign n7922 = ( n569 & n3034 ) | ( n569 & n7122 ) | ( n3034 & n7122 ) ;
  assign n7923 = ( ~n802 & n2131 ) | ( ~n802 & n2765 ) | ( n2131 & n2765 ) ;
  assign n7924 = n7923 ^ n4313 ^ 1'b0 ;
  assign n7925 = n1645 | n3097 ;
  assign n7926 = n2394 ^ n2197 ^ 1'b0 ;
  assign n7927 = n3391 | n7926 ;
  assign n7928 = n7925 & ~n7927 ;
  assign n7929 = n4196 ^ n2005 ^ 1'b0 ;
  assign n7930 = ~n2337 & n7929 ;
  assign n7931 = ~n4945 & n7930 ;
  assign n7932 = n7931 ^ x126 ^ 1'b0 ;
  assign n7933 = n2697 & ~n3770 ;
  assign n7934 = n7317 & n7933 ;
  assign n7935 = n7934 ^ n7879 ^ n259 ;
  assign n7936 = n7674 ^ n4943 ^ 1'b0 ;
  assign n7937 = n1108 & n4036 ;
  assign n7938 = ~n4391 & n4587 ;
  assign n7939 = ~n7937 & n7938 ;
  assign n7940 = n7758 | n7939 ;
  assign n7941 = n2050 & n5772 ;
  assign n7942 = n1720 ^ n1102 ^ 1'b0 ;
  assign n7943 = n4287 ^ n3583 ^ 1'b0 ;
  assign n7944 = n7942 | n7943 ;
  assign n7945 = n4781 & ~n7294 ;
  assign n7946 = n7945 ^ n3296 ^ n2723 ;
  assign n7949 = n1411 | n3286 ;
  assign n7950 = n7949 ^ n4207 ^ 1'b0 ;
  assign n7951 = n5864 & ~n7950 ;
  assign n7952 = n7665 & n7951 ;
  assign n7947 = ~n411 & n2075 ;
  assign n7948 = n2575 | n7947 ;
  assign n7953 = n7952 ^ n7948 ^ 1'b0 ;
  assign n7954 = ( ~n6952 & n7946 ) | ( ~n6952 & n7953 ) | ( n7946 & n7953 ) ;
  assign n7955 = n3778 ^ n1808 ^ 1'b0 ;
  assign n7956 = n5575 ^ n2354 ^ 1'b0 ;
  assign n7957 = n7955 & ~n7956 ;
  assign n7958 = n4517 ^ x58 ^ 1'b0 ;
  assign n7959 = n410 & ~n1066 ;
  assign n7960 = n4440 & n7959 ;
  assign n7961 = n4150 | n7960 ;
  assign n7962 = n7961 ^ x109 ^ 1'b0 ;
  assign n7963 = n963 & n2956 ;
  assign n7964 = n1838 & n5331 ;
  assign n7965 = ~n1027 & n7964 ;
  assign n7966 = n2831 | n7965 ;
  assign n7967 = n5250 | n5519 ;
  assign n7968 = n7966 & ~n7967 ;
  assign n7969 = ( n6958 & ~n7963 ) | ( n6958 & n7968 ) | ( ~n7963 & n7968 ) ;
  assign n7970 = n4395 ^ n1134 ^ n537 ;
  assign n7971 = n7930 ^ n4483 ^ 1'b0 ;
  assign n7972 = ~n5169 & n6577 ;
  assign n7974 = n3038 ^ n2676 ^ n2226 ;
  assign n7973 = n1139 | n3842 ;
  assign n7975 = n7974 ^ n7973 ^ 1'b0 ;
  assign n7982 = n6091 ^ n2744 ^ n2326 ;
  assign n7976 = n1651 | n6253 ;
  assign n7978 = n5411 ^ n1726 ^ 1'b0 ;
  assign n7977 = ~n5599 & n6323 ;
  assign n7979 = n7978 ^ n7977 ^ 1'b0 ;
  assign n7980 = ~n7976 & n7979 ;
  assign n7981 = n1557 & n7980 ;
  assign n7983 = n7982 ^ n7981 ^ 1'b0 ;
  assign n7984 = n974 ^ n774 ^ 1'b0 ;
  assign n7985 = n7984 ^ n6215 ^ 1'b0 ;
  assign n7986 = n2942 & n7985 ;
  assign n7987 = n1164 | n1451 ;
  assign n7989 = n265 & ~n3002 ;
  assign n7990 = ~n3737 & n7989 ;
  assign n7991 = n1701 ^ n1657 ^ 1'b0 ;
  assign n7992 = n1870 & ~n7991 ;
  assign n7993 = n1732 & n3466 ;
  assign n7994 = ~n7992 & n7993 ;
  assign n7995 = n7994 ^ n4134 ^ x84 ;
  assign n7996 = n5914 | n7995 ;
  assign n7997 = n7990 & ~n7996 ;
  assign n7988 = n1691 ^ x14 ^ 1'b0 ;
  assign n7998 = n7997 ^ n7988 ^ 1'b0 ;
  assign n7999 = n7987 & n7998 ;
  assign n8000 = n1132 & n5970 ;
  assign n8001 = n1850 & n2057 ;
  assign n8002 = ( n2519 & n5843 ) | ( n2519 & n7063 ) | ( n5843 & n7063 ) ;
  assign n8003 = n4867 ^ x25 ^ 1'b0 ;
  assign n8004 = n8002 & ~n8003 ;
  assign n8005 = n8001 & n8004 ;
  assign n8006 = n5350 ^ n4575 ^ 1'b0 ;
  assign n8007 = n5661 | n8006 ;
  assign n8008 = n4038 & ~n8007 ;
  assign n8009 = n2951 & n8008 ;
  assign n8010 = n3566 ^ n2412 ^ 1'b0 ;
  assign n8011 = n2210 & n8010 ;
  assign n8012 = n5141 ^ n4902 ^ 1'b0 ;
  assign n8013 = n8011 & n8012 ;
  assign n8014 = n8013 ^ n305 ^ 1'b0 ;
  assign n8015 = n2212 | n5809 ;
  assign n8016 = n3800 | n8015 ;
  assign n8017 = n5043 & n8016 ;
  assign n8018 = n4137 & ~n7871 ;
  assign n8021 = n3304 ^ n1692 ^ 1'b0 ;
  assign n8022 = n1270 & ~n8021 ;
  assign n8019 = ( n2692 & n4422 ) | ( n2692 & ~n4889 ) | ( n4422 & ~n4889 ) ;
  assign n8020 = n8019 ^ n8007 ^ 1'b0 ;
  assign n8023 = n8022 ^ n8020 ^ 1'b0 ;
  assign n8024 = n648 & ~n8023 ;
  assign n8026 = n7974 ^ n7127 ^ n2869 ;
  assign n8025 = n5090 | n7250 ;
  assign n8027 = n8026 ^ n8025 ^ 1'b0 ;
  assign n8028 = n405 ^ n256 ^ 1'b0 ;
  assign n8029 = n3077 | n8028 ;
  assign n8030 = n8029 ^ n3613 ^ 1'b0 ;
  assign n8036 = n300 | n1646 ;
  assign n8037 = n572 & ~n8036 ;
  assign n8032 = n3617 ^ n1472 ^ x101 ;
  assign n8033 = x175 & n8032 ;
  assign n8034 = n2632 & ~n8033 ;
  assign n8031 = x163 & n6982 ;
  assign n8035 = n8034 ^ n8031 ^ 1'b0 ;
  assign n8038 = n8037 ^ n8035 ^ 1'b0 ;
  assign n8039 = ~n1376 & n4865 ;
  assign n8040 = ~n1524 & n4796 ;
  assign n8041 = n2076 & n6844 ;
  assign n8042 = x233 & n7404 ;
  assign n8043 = n3918 ^ x14 ^ 1'b0 ;
  assign n8044 = n4550 & n8043 ;
  assign n8045 = n1421 & ~n1804 ;
  assign n8046 = n6012 & n8045 ;
  assign n8047 = n2296 | n6692 ;
  assign n8048 = n5814 | n8047 ;
  assign n8049 = x182 & ~n4570 ;
  assign n8050 = n8049 ^ n4409 ^ 1'b0 ;
  assign n8051 = n1328 & n8050 ;
  assign n8052 = n8051 ^ n1823 ^ 1'b0 ;
  assign n8053 = ~n481 & n833 ;
  assign n8054 = n2350 & ~n8053 ;
  assign n8055 = n3881 ^ n2638 ^ 1'b0 ;
  assign n8056 = n4529 ^ n1377 ^ 1'b0 ;
  assign n8057 = ( n2374 & n4346 ) | ( n2374 & n8056 ) | ( n4346 & n8056 ) ;
  assign n8058 = ~n1304 & n8057 ;
  assign n8059 = n8055 | n8058 ;
  assign n8060 = n8059 ^ n4191 ^ 1'b0 ;
  assign n8061 = n5324 ^ n3779 ^ 1'b0 ;
  assign n8062 = n5057 | n8061 ;
  assign n8063 = n6450 & ~n8062 ;
  assign n8064 = n2696 & n8063 ;
  assign n8065 = ( n445 & n3297 ) | ( n445 & ~n6312 ) | ( n3297 & ~n6312 ) ;
  assign n8066 = n2216 & n8065 ;
  assign n8067 = n936 & n4984 ;
  assign n8068 = n6352 & n8067 ;
  assign n8069 = ~n1107 & n8068 ;
  assign n8070 = n8069 ^ n7584 ^ 1'b0 ;
  assign n8071 = n8066 & ~n8070 ;
  assign n8072 = n831 & ~n4349 ;
  assign n8073 = n8072 ^ n3747 ^ 1'b0 ;
  assign n8074 = n5922 & ~n8073 ;
  assign n8075 = n6299 & n8074 ;
  assign n8076 = n7003 | n8075 ;
  assign n8077 = n2864 & ~n3363 ;
  assign n8078 = n5522 ^ n1139 ^ 1'b0 ;
  assign n8079 = n8077 | n8078 ;
  assign n8080 = n5235 & ~n8079 ;
  assign n8081 = n5017 ^ n3251 ^ 1'b0 ;
  assign n8082 = n4676 | n6352 ;
  assign n8083 = n8082 ^ n5277 ^ 1'b0 ;
  assign n8084 = n8083 ^ n6345 ^ n4784 ;
  assign n8085 = x219 | n5720 ;
  assign n8086 = n3288 & n6976 ;
  assign n8087 = ~n4787 & n8086 ;
  assign n8088 = ( x205 & ~n1575 ) | ( x205 & n2954 ) | ( ~n1575 & n2954 ) ;
  assign n8089 = n5586 | n7756 ;
  assign n8090 = n7492 & ~n8089 ;
  assign n8091 = n1458 & ~n5411 ;
  assign n8092 = n2105 ^ x199 ^ 1'b0 ;
  assign n8093 = n459 & ~n8092 ;
  assign n8094 = n2214 & n8093 ;
  assign n8095 = n2091 ^ n610 ^ 1'b0 ;
  assign n8096 = ~x201 & n8095 ;
  assign n8097 = ~n940 & n8096 ;
  assign n8098 = ~n1164 & n8097 ;
  assign n8099 = n8094 | n8098 ;
  assign n8100 = n5617 | n8099 ;
  assign n8101 = n6297 ^ n5591 ^ n1082 ;
  assign n8102 = n8101 ^ n2838 ^ 1'b0 ;
  assign n8103 = ( n2800 & ~n3566 ) | ( n2800 & n8102 ) | ( ~n3566 & n8102 ) ;
  assign n8104 = n2770 | n4089 ;
  assign n8105 = n8104 ^ n6774 ^ 1'b0 ;
  assign n8106 = ~n8103 & n8105 ;
  assign n8107 = ~n734 & n8106 ;
  assign n8108 = n2777 & n4541 ;
  assign n8109 = n361 & n8108 ;
  assign n8110 = n8109 ^ n800 ^ 1'b0 ;
  assign n8111 = ~n764 & n8110 ;
  assign n8112 = n8111 ^ n5772 ^ 1'b0 ;
  assign n8113 = ( ~n3313 & n3924 ) | ( ~n3313 & n7707 ) | ( n3924 & n7707 ) ;
  assign n8114 = n8113 ^ n2966 ^ 1'b0 ;
  assign n8115 = n1281 | n6309 ;
  assign n8116 = n8115 ^ n5971 ^ 1'b0 ;
  assign n8117 = n5456 | n8116 ;
  assign n8118 = ~n1720 & n8117 ;
  assign n8119 = n3063 ^ x247 ^ 1'b0 ;
  assign n8120 = n8119 ^ n271 ^ 1'b0 ;
  assign n8121 = n283 | n4719 ;
  assign n8122 = n3078 ^ n2654 ^ 1'b0 ;
  assign n8123 = n3550 ^ n952 ^ 1'b0 ;
  assign n8124 = n2518 ^ n2247 ^ 1'b0 ;
  assign n8127 = n4896 ^ n3112 ^ 1'b0 ;
  assign n8128 = ~n2455 & n8127 ;
  assign n8125 = n2216 | n2571 ;
  assign n8126 = n8125 ^ n1413 ^ 1'b0 ;
  assign n8129 = n8128 ^ n8126 ^ 1'b0 ;
  assign n8130 = n2605 & ~n8129 ;
  assign n8131 = ( ~n1565 & n2076 ) | ( ~n1565 & n3705 ) | ( n2076 & n3705 ) ;
  assign n8132 = n2183 | n8131 ;
  assign n8133 = n6528 | n8132 ;
  assign n8134 = n2668 & ~n3242 ;
  assign n8135 = n4015 | n8134 ;
  assign n8136 = n5485 | n8135 ;
  assign n8137 = n8133 & n8136 ;
  assign n8138 = ~n4901 & n7609 ;
  assign n8139 = ~n2866 & n3933 ;
  assign n8140 = x109 & ~n1850 ;
  assign n8141 = ~n365 & n967 ;
  assign n8142 = n8141 ^ n1958 ^ 1'b0 ;
  assign n8143 = n6811 & ~n8142 ;
  assign n8144 = n8143 ^ n5054 ^ 1'b0 ;
  assign n8145 = n3438 ^ n2793 ^ 1'b0 ;
  assign n8146 = n8145 ^ n7752 ^ 1'b0 ;
  assign n8147 = n4729 ^ n3369 ^ 1'b0 ;
  assign n8148 = n8146 | n8147 ;
  assign n8149 = ~n3888 & n8148 ;
  assign n8151 = n4174 ^ n476 ^ 1'b0 ;
  assign n8150 = x136 & n7615 ;
  assign n8152 = n8151 ^ n8150 ^ 1'b0 ;
  assign n8153 = n8152 ^ n5145 ^ 1'b0 ;
  assign n8154 = n6572 ^ n1129 ^ n1113 ;
  assign n8155 = x17 & ~n5193 ;
  assign n8156 = n978 & n8155 ;
  assign n8157 = n8156 ^ n6646 ^ 1'b0 ;
  assign n8158 = n3773 & ~n8157 ;
  assign n8159 = n4010 ^ n1150 ^ 1'b0 ;
  assign n8160 = n8159 ^ n698 ^ 1'b0 ;
  assign n8161 = n3904 | n8160 ;
  assign n8162 = n2804 & n5228 ;
  assign n8163 = ~n2601 & n8162 ;
  assign n8164 = n988 ^ x199 ^ x94 ;
  assign n8165 = n5550 | n8164 ;
  assign n8170 = ~n2371 & n4764 ;
  assign n8166 = n718 | n6874 ;
  assign n8167 = n887 | n8166 ;
  assign n8168 = ~n4361 & n8167 ;
  assign n8169 = ~x37 & n8168 ;
  assign n8171 = n8170 ^ n8169 ^ 1'b0 ;
  assign n8172 = n2274 | n6625 ;
  assign n8173 = n5232 | n8172 ;
  assign n8174 = n2284 | n4524 ;
  assign n8175 = n8174 ^ n5431 ^ 1'b0 ;
  assign n8176 = n1524 & ~n8175 ;
  assign n8177 = x137 & n2240 ;
  assign n8178 = n8177 ^ n1024 ^ 1'b0 ;
  assign n8179 = ( x15 & n2148 ) | ( x15 & n6192 ) | ( n2148 & n6192 ) ;
  assign n8180 = n652 & n8179 ;
  assign n8181 = n8178 & n8180 ;
  assign n8182 = ~n444 & n3254 ;
  assign n8183 = n8182 ^ n5350 ^ 1'b0 ;
  assign n8184 = n8183 ^ n7817 ^ 1'b0 ;
  assign n8185 = n3548 & ~n8184 ;
  assign n8186 = n8185 ^ n4956 ^ 1'b0 ;
  assign n8187 = ~n8181 & n8186 ;
  assign n8188 = n1626 & ~n2698 ;
  assign n8189 = ~n8187 & n8188 ;
  assign n8190 = n8189 ^ n3113 ^ n1478 ;
  assign n8191 = n4383 & n7801 ;
  assign n8192 = n3121 ^ n677 ^ 1'b0 ;
  assign n8193 = n2746 & n8192 ;
  assign n8194 = ( n565 & n8191 ) | ( n565 & ~n8193 ) | ( n8191 & ~n8193 ) ;
  assign n8195 = x49 | n1011 ;
  assign n8196 = n7223 ^ n669 ^ 1'b0 ;
  assign n8197 = n6430 & ~n8196 ;
  assign n8198 = n4932 & n8197 ;
  assign n8201 = n4878 & ~n7329 ;
  assign n8199 = n908 ^ x19 ^ 1'b0 ;
  assign n8200 = n4652 & ~n8199 ;
  assign n8202 = n8201 ^ n8200 ^ n3239 ;
  assign n8203 = ( n1453 & ~n7421 ) | ( n1453 & n8202 ) | ( ~n7421 & n8202 ) ;
  assign n8215 = n3698 ^ n3472 ^ n982 ;
  assign n8212 = n2430 & n6628 ;
  assign n8213 = n8212 ^ n4735 ^ n345 ;
  assign n8214 = n8213 ^ n3913 ^ n939 ;
  assign n8204 = n3467 & ~n4569 ;
  assign n8205 = n8204 ^ n3651 ^ 1'b0 ;
  assign n8206 = n5071 | n5728 ;
  assign n8207 = n2097 & ~n8206 ;
  assign n8208 = n7037 & ~n8207 ;
  assign n8209 = ~x36 & n8208 ;
  assign n8210 = n1553 & ~n8209 ;
  assign n8211 = ~n8205 & n8210 ;
  assign n8216 = n8215 ^ n8214 ^ n8211 ;
  assign n8217 = x136 & ~n6330 ;
  assign n8218 = ( x228 & n3034 ) | ( x228 & n7923 ) | ( n3034 & n7923 ) ;
  assign n8219 = x36 | n645 ;
  assign n8220 = ~n6417 & n8207 ;
  assign n8221 = n4774 ^ n3014 ^ 1'b0 ;
  assign n8222 = ~n1561 & n8221 ;
  assign n8223 = ~n467 & n531 ;
  assign n8224 = n8223 ^ n1920 ^ 1'b0 ;
  assign n8225 = n1353 | n8224 ;
  assign n8226 = ( ~n395 & n8222 ) | ( ~n395 & n8225 ) | ( n8222 & n8225 ) ;
  assign n8227 = n8226 ^ n7667 ^ n3256 ;
  assign n8228 = ~n2707 & n4271 ;
  assign n8229 = n8228 ^ n5117 ^ 1'b0 ;
  assign n8230 = n4536 ^ n335 ^ 1'b0 ;
  assign n8231 = n8229 & ~n8230 ;
  assign n8232 = n2190 | n8231 ;
  assign n8233 = ~n1129 & n8232 ;
  assign n8234 = n1213 & n4289 ;
  assign n8235 = ~n974 & n4205 ;
  assign n8236 = n8235 ^ n2085 ^ x58 ;
  assign n8237 = n1220 & ~n8236 ;
  assign n8238 = n4434 & n8237 ;
  assign n8239 = n8238 ^ n1254 ^ 1'b0 ;
  assign n8240 = ~n1781 & n8239 ;
  assign n8241 = n8240 ^ n6852 ^ n2279 ;
  assign n8242 = ~n8234 & n8241 ;
  assign n8243 = n8242 ^ n4369 ^ 1'b0 ;
  assign n8244 = n2986 | n6541 ;
  assign n8245 = x52 & n6489 ;
  assign n8246 = n8245 ^ n6602 ^ n4542 ;
  assign n8249 = n7597 ^ n1550 ^ 1'b0 ;
  assign n8250 = n5877 & n8249 ;
  assign n8247 = ( ~n745 & n1036 ) | ( ~n745 & n1068 ) | ( n1036 & n1068 ) ;
  assign n8248 = ~n2900 & n8247 ;
  assign n8251 = n8250 ^ n8248 ^ 1'b0 ;
  assign n8252 = ( n369 & n2659 ) | ( n369 & ~n8156 ) | ( n2659 & ~n8156 ) ;
  assign n8253 = ( ~n692 & n2448 ) | ( ~n692 & n8252 ) | ( n2448 & n8252 ) ;
  assign n8255 = n2768 & ~n5077 ;
  assign n8256 = n8255 ^ n3652 ^ n579 ;
  assign n8254 = n4213 & ~n8034 ;
  assign n8257 = n8256 ^ n8254 ^ 1'b0 ;
  assign n8260 = ~n3288 & n4078 ;
  assign n8258 = n5914 ^ n2320 ^ 1'b0 ;
  assign n8259 = n3041 & n8258 ;
  assign n8261 = n8260 ^ n8259 ^ 1'b0 ;
  assign n8262 = n607 & n6390 ;
  assign n8263 = ~n5644 & n6814 ;
  assign n8264 = n8263 ^ n8236 ^ 1'b0 ;
  assign n8265 = n8264 ^ n4334 ^ 1'b0 ;
  assign n8266 = ~n2447 & n3472 ;
  assign n8267 = n5177 ^ n446 ^ 1'b0 ;
  assign n8268 = n614 | n8267 ;
  assign n8269 = n2592 | n8268 ;
  assign n8270 = n8266 & ~n8269 ;
  assign n8271 = n8118 & n8270 ;
  assign n8272 = x191 & ~x222 ;
  assign n8273 = ~n3128 & n8272 ;
  assign n8274 = n8273 ^ n768 ^ 1'b0 ;
  assign n8275 = n8274 ^ n312 ^ 1'b0 ;
  assign n8276 = n4521 ^ n1187 ^ 1'b0 ;
  assign n8280 = ~n4430 & n4774 ;
  assign n8281 = ~n6307 & n8280 ;
  assign n8277 = ( x115 & x196 ) | ( x115 & n681 ) | ( x196 & n681 ) ;
  assign n8278 = n8277 ^ n5043 ^ 1'b0 ;
  assign n8279 = n1328 & n8278 ;
  assign n8282 = n8281 ^ n8279 ^ 1'b0 ;
  assign n8283 = n5359 & n7644 ;
  assign n8284 = n5852 ^ n5639 ^ 1'b0 ;
  assign n8285 = n1486 & ~n1533 ;
  assign n8286 = n1762 & n8285 ;
  assign n8287 = n514 & ~n8286 ;
  assign n8288 = n3513 ^ n1108 ^ 1'b0 ;
  assign n8289 = n8288 ^ n2166 ^ 1'b0 ;
  assign n8290 = ~n5445 & n8289 ;
  assign n8291 = ( n3405 & ~n5110 ) | ( n3405 & n8290 ) | ( ~n5110 & n8290 ) ;
  assign n8292 = n2113 | n2794 ;
  assign n8293 = n8291 | n8292 ;
  assign n8294 = n7008 ^ n5449 ^ 1'b0 ;
  assign n8295 = n2260 & n4887 ;
  assign n8296 = ~n1063 & n4853 ;
  assign n8297 = n1584 & n8296 ;
  assign n8298 = ~n8295 & n8297 ;
  assign n8299 = ( n3915 & n4338 ) | ( n3915 & n6064 ) | ( n4338 & n6064 ) ;
  assign n8300 = n7023 ^ n5138 ^ n3765 ;
  assign n8301 = n2332 & ~n8300 ;
  assign n8302 = n2169 & n5402 ;
  assign n8303 = n853 & n6114 ;
  assign n8306 = n5807 ^ n3150 ^ n2953 ;
  assign n8304 = n1700 & ~n4780 ;
  assign n8305 = n8304 ^ n1817 ^ 1'b0 ;
  assign n8307 = n8306 ^ n8305 ^ 1'b0 ;
  assign n8309 = n3682 ^ n2759 ^ 1'b0 ;
  assign n8308 = n319 & ~n2955 ;
  assign n8310 = n8309 ^ n8308 ^ 1'b0 ;
  assign n8311 = n3225 & ~n8310 ;
  assign n8312 = ( n1992 & n6031 ) | ( n1992 & ~n6579 ) | ( n6031 & ~n6579 ) ;
  assign n8313 = n8312 ^ n3386 ^ 1'b0 ;
  assign n8314 = n5159 | n8313 ;
  assign n8315 = n8037 ^ n1989 ^ 1'b0 ;
  assign n8316 = ( n984 & ~n5650 ) | ( n984 & n8315 ) | ( ~n5650 & n8315 ) ;
  assign n8317 = n1496 & n2053 ;
  assign n8318 = n8317 ^ n3536 ^ 1'b0 ;
  assign n8319 = n8318 ^ n3826 ^ n552 ;
  assign n8320 = n2195 ^ n1273 ^ 1'b0 ;
  assign n8321 = n1677 ^ n1162 ^ 1'b0 ;
  assign n8322 = ~n1168 & n3763 ;
  assign n8323 = n8322 ^ n7833 ^ 1'b0 ;
  assign n8324 = n677 & n838 ;
  assign n8325 = n3926 ^ n1450 ^ n1281 ;
  assign n8326 = n8117 ^ n7028 ^ 1'b0 ;
  assign n8327 = n1835 & n8326 ;
  assign n8328 = n4533 & ~n5600 ;
  assign n8329 = n8328 ^ n302 ^ 1'b0 ;
  assign n8330 = n2852 ^ x65 ^ 1'b0 ;
  assign n8331 = ~n258 & n4174 ;
  assign n8332 = n8331 ^ n758 ^ 1'b0 ;
  assign n8333 = x26 & n8332 ;
  assign n8334 = n8333 ^ n326 ^ 1'b0 ;
  assign n8335 = n8334 ^ n4964 ^ 1'b0 ;
  assign n8336 = n8330 & n8335 ;
  assign n8337 = ~n1418 & n6645 ;
  assign n8338 = ~n650 & n8337 ;
  assign n8339 = n8338 ^ n3059 ^ 1'b0 ;
  assign n8340 = ( n3402 & n3785 ) | ( n3402 & ~n4719 ) | ( n3785 & ~n4719 ) ;
  assign n8341 = n881 | n2329 ;
  assign n8342 = n3282 & ~n8341 ;
  assign n8343 = n8342 ^ n2953 ^ n2600 ;
  assign n8344 = ( ~x39 & n2106 ) | ( ~x39 & n4636 ) | ( n2106 & n4636 ) ;
  assign n8345 = ~n8343 & n8344 ;
  assign n8346 = x177 | n8144 ;
  assign n8347 = n1239 & ~n5716 ;
  assign n8348 = n8347 ^ x239 ^ 1'b0 ;
  assign n8349 = n2203 & ~n8348 ;
  assign n8350 = n8349 ^ n6321 ^ 1'b0 ;
  assign n8351 = n7577 ^ n6202 ^ 1'b0 ;
  assign n8352 = ( n4655 & n6717 ) | ( n4655 & ~n8351 ) | ( n6717 & ~n8351 ) ;
  assign n8353 = x153 & n4191 ;
  assign n8354 = ~n6798 & n8353 ;
  assign n8355 = n709 & ~n8354 ;
  assign n8356 = n8355 ^ n1172 ^ 1'b0 ;
  assign n8357 = ~n4817 & n8356 ;
  assign n8358 = ~n4284 & n8357 ;
  assign n8359 = ~n650 & n1733 ;
  assign n8360 = n8359 ^ n7172 ^ 1'b0 ;
  assign n8361 = ~n721 & n3088 ;
  assign n8362 = ~n8360 & n8361 ;
  assign n8363 = n6605 & n7462 ;
  assign n8364 = n2460 & ~n8363 ;
  assign n8366 = n7127 ^ n6119 ^ n5939 ;
  assign n8365 = n883 & n5810 ;
  assign n8367 = n8366 ^ n8365 ^ 1'b0 ;
  assign n8368 = ( n5510 & n5972 ) | ( n5510 & ~n8145 ) | ( n5972 & ~n8145 ) ;
  assign n8369 = n2755 & n8368 ;
  assign n8370 = n6682 ^ n5398 ^ x188 ;
  assign n8371 = ~n4840 & n8370 ;
  assign n8372 = ~x112 & n8371 ;
  assign n8373 = n2841 & ~n5411 ;
  assign n8374 = ~n1310 & n8373 ;
  assign n8375 = n956 | n8374 ;
  assign n8376 = n8372 | n8375 ;
  assign n8377 = ~n1472 & n5752 ;
  assign n8378 = n993 & n3448 ;
  assign n8380 = n5672 ^ n1592 ^ 1'b0 ;
  assign n8381 = n5188 | n8380 ;
  assign n8379 = ~n1364 & n2648 ;
  assign n8382 = n8381 ^ n8379 ^ 1'b0 ;
  assign n8383 = n3212 | n4356 ;
  assign n8384 = ( n3274 & n6302 ) | ( n3274 & n8383 ) | ( n6302 & n8383 ) ;
  assign n8385 = n1156 | n2174 ;
  assign n8386 = n6973 | n8385 ;
  assign n8387 = ~n6561 & n8386 ;
  assign n8388 = n5117 ^ n3604 ^ 1'b0 ;
  assign n8389 = n8388 ^ n6708 ^ n790 ;
  assign n8390 = n7672 & ~n8389 ;
  assign n8391 = ( n417 & n5576 ) | ( n417 & n6264 ) | ( n5576 & n6264 ) ;
  assign n8392 = n6285 ^ n2617 ^ 1'b0 ;
  assign n8393 = n7969 | n8392 ;
  assign n8394 = n6236 ^ n4224 ^ 1'b0 ;
  assign n8395 = ( n1358 & n4827 ) | ( n1358 & n8394 ) | ( n4827 & n8394 ) ;
  assign n8397 = n2166 ^ n1655 ^ 1'b0 ;
  assign n8398 = n6884 & ~n8397 ;
  assign n8396 = n1955 & ~n4701 ;
  assign n8399 = n8398 ^ n8396 ^ 1'b0 ;
  assign n8401 = ~n4298 & n6394 ;
  assign n8402 = n8401 ^ n7330 ^ 1'b0 ;
  assign n8400 = n4542 & ~n6737 ;
  assign n8403 = n8402 ^ n8400 ^ 1'b0 ;
  assign n8404 = n3650 ^ x159 ^ 1'b0 ;
  assign n8405 = n1201 | n8404 ;
  assign n8406 = ~n2610 & n4548 ;
  assign n8407 = n8405 & ~n8406 ;
  assign n8408 = n8403 | n8407 ;
  assign n8409 = n5426 ^ n960 ^ 1'b0 ;
  assign n8410 = n5350 & n5967 ;
  assign n8411 = n6895 & ~n8410 ;
  assign n8412 = ~n2182 & n3787 ;
  assign n8413 = ~n5115 & n8412 ;
  assign n8414 = n2249 & ~n8413 ;
  assign n8415 = n8414 ^ n1189 ^ 1'b0 ;
  assign n8416 = n1880 & ~n8415 ;
  assign n8417 = ~n5019 & n8416 ;
  assign n8418 = n2707 & ~n8417 ;
  assign n8419 = ~n3638 & n8418 ;
  assign n8420 = n2547 ^ n946 ^ 1'b0 ;
  assign n8421 = n3111 & ~n4936 ;
  assign n8422 = n4231 & n8421 ;
  assign n8423 = n8422 ^ x143 ^ 1'b0 ;
  assign n8424 = n1442 & ~n5762 ;
  assign n8425 = ~n1077 & n4137 ;
  assign n8426 = ~n1304 & n5315 ;
  assign n8427 = ~n8425 & n8426 ;
  assign n8428 = n8427 ^ n7229 ^ n5404 ;
  assign n8429 = ~n402 & n599 ;
  assign n8430 = ~n1675 & n8429 ;
  assign n8431 = n6665 & ~n8430 ;
  assign n8432 = n8431 ^ n3723 ^ 1'b0 ;
  assign n8433 = n4168 ^ n3275 ^ 1'b0 ;
  assign n8434 = n2151 & ~n3929 ;
  assign n8435 = n8434 ^ n1508 ^ 1'b0 ;
  assign n8436 = n3711 | n5122 ;
  assign n8437 = n8436 ^ n8049 ^ 1'b0 ;
  assign n8438 = ( ~n397 & n937 ) | ( ~n397 & n5246 ) | ( n937 & n5246 ) ;
  assign n8439 = n2768 | n8438 ;
  assign n8440 = n5663 | n8439 ;
  assign n8441 = x244 & n5043 ;
  assign n8442 = n8440 & n8441 ;
  assign n8443 = ~n5522 & n8442 ;
  assign n8444 = n5036 & ~n8443 ;
  assign n8445 = n8437 & n8444 ;
  assign n8447 = n6534 ^ n6198 ^ n498 ;
  assign n8448 = n1919 & ~n3714 ;
  assign n8449 = ~n8447 & n8448 ;
  assign n8446 = n7976 ^ n7650 ^ 1'b0 ;
  assign n8450 = n8449 ^ n8446 ^ 1'b0 ;
  assign n8451 = n7849 ^ n6976 ^ 1'b0 ;
  assign n8452 = x138 & ~n4903 ;
  assign n8453 = n8452 ^ n1369 ^ 1'b0 ;
  assign n8454 = n3244 & ~n8453 ;
  assign n8455 = n8454 ^ n3451 ^ 1'b0 ;
  assign n8456 = n8455 ^ n7354 ^ 1'b0 ;
  assign n8457 = n4222 & n8456 ;
  assign n8458 = n7316 ^ n6614 ^ 1'b0 ;
  assign n8459 = n1152 | n8458 ;
  assign n8460 = n410 & n1234 ;
  assign n8461 = n2730 & n8460 ;
  assign n8462 = n2142 & ~n8461 ;
  assign n8463 = n8459 & n8462 ;
  assign n8464 = n8308 ^ n6644 ^ 1'b0 ;
  assign n8465 = n5586 | n8464 ;
  assign n8466 = n7492 | n8465 ;
  assign n8467 = n8466 ^ x247 ^ 1'b0 ;
  assign n8468 = n2667 | n8467 ;
  assign n8469 = ~n2051 & n8432 ;
  assign n8470 = n8469 ^ n7918 ^ 1'b0 ;
  assign n8471 = n3791 ^ x10 ^ 1'b0 ;
  assign n8472 = n2204 ^ n1917 ^ 1'b0 ;
  assign n8473 = n1932 & ~n8472 ;
  assign n8474 = n8473 ^ n485 ^ 1'b0 ;
  assign n8475 = x112 & x185 ;
  assign n8476 = n6833 & n8475 ;
  assign n8477 = ( n259 & n8474 ) | ( n259 & ~n8476 ) | ( n8474 & ~n8476 ) ;
  assign n8478 = n8471 & ~n8477 ;
  assign n8479 = n3938 ^ n806 ^ 1'b0 ;
  assign n8480 = n411 & n8479 ;
  assign n8481 = ~n4977 & n8480 ;
  assign n8482 = ~n822 & n5501 ;
  assign n8483 = x98 & ~n3212 ;
  assign n8484 = n8483 ^ x166 ^ 1'b0 ;
  assign n8485 = n6814 ^ n2223 ^ 1'b0 ;
  assign n8486 = n2975 & n5457 ;
  assign n8487 = ~n8485 & n8486 ;
  assign n8488 = ( n4312 & n8484 ) | ( n4312 & ~n8487 ) | ( n8484 & ~n8487 ) ;
  assign n8489 = n6049 ^ n2521 ^ 1'b0 ;
  assign n8490 = n8488 | n8489 ;
  assign n8491 = ( n2138 & n2442 ) | ( n2138 & ~n3775 ) | ( n2442 & ~n3775 ) ;
  assign n8492 = n2155 | n8491 ;
  assign n8493 = n8490 & ~n8492 ;
  assign n8494 = n2490 & ~n7540 ;
  assign n8495 = n886 & n4222 ;
  assign n8496 = n1084 & n8495 ;
  assign n8497 = n3926 ^ n1895 ^ 1'b0 ;
  assign n8499 = n1067 ^ n831 ^ 1'b0 ;
  assign n8500 = n8178 | n8499 ;
  assign n8498 = n2584 & ~n3070 ;
  assign n8501 = n8500 ^ n8498 ^ 1'b0 ;
  assign n8502 = n3113 ^ n1250 ^ 1'b0 ;
  assign n8503 = n5680 | n8502 ;
  assign n8504 = n8503 ^ n5934 ^ 1'b0 ;
  assign n8505 = n7482 & ~n8504 ;
  assign n8506 = n5067 ^ n3338 ^ 1'b0 ;
  assign n8507 = n1124 | n8506 ;
  assign n8508 = n5376 | n8507 ;
  assign n8509 = n7088 | n8508 ;
  assign n8510 = n7823 ^ n2571 ^ 1'b0 ;
  assign n8511 = n6556 ^ n4201 ^ n2935 ;
  assign n8512 = n3721 & ~n8511 ;
  assign n8513 = n8512 ^ n7376 ^ 1'b0 ;
  assign n8514 = n858 & ~n3201 ;
  assign n8515 = ~n2368 & n8514 ;
  assign n8516 = n5687 | n8515 ;
  assign n8517 = n8516 ^ n8302 ^ 1'b0 ;
  assign n8520 = n7809 ^ n7012 ^ 1'b0 ;
  assign n8518 = n1255 & n2421 ;
  assign n8519 = ~n3045 & n8518 ;
  assign n8521 = n8520 ^ n8519 ^ 1'b0 ;
  assign n8522 = n7515 ^ n4560 ^ n1811 ;
  assign n8523 = n4481 | n8522 ;
  assign n8524 = ( ~x216 & n6914 ) | ( ~x216 & n8523 ) | ( n6914 & n8523 ) ;
  assign n8525 = n4417 | n6124 ;
  assign n8526 = n8525 ^ n3672 ^ 1'b0 ;
  assign n8527 = x15 & n4722 ;
  assign n8528 = n8527 ^ n2359 ^ 1'b0 ;
  assign n8529 = n317 & ~n824 ;
  assign n8530 = n8529 ^ n3959 ^ n1807 ;
  assign n8531 = n8530 ^ n405 ^ 1'b0 ;
  assign n8532 = n3995 | n8531 ;
  assign n8534 = n1444 | n3431 ;
  assign n8535 = n3051 & ~n8534 ;
  assign n8536 = n4469 | n8535 ;
  assign n8537 = n8536 ^ n933 ^ 1'b0 ;
  assign n8538 = n8537 ^ n5162 ^ n3000 ;
  assign n8539 = n8538 ^ n527 ^ 1'b0 ;
  assign n8533 = n3926 & ~n4752 ;
  assign n8540 = n8539 ^ n8533 ^ 1'b0 ;
  assign n8541 = n4526 & ~n8540 ;
  assign n8542 = ( ~n966 & n8532 ) | ( ~n966 & n8541 ) | ( n8532 & n8541 ) ;
  assign n8543 = ( n332 & n377 ) | ( n332 & ~n1153 ) | ( n377 & ~n1153 ) ;
  assign n8544 = x238 | n8543 ;
  assign n8545 = n8544 ^ n1144 ^ 1'b0 ;
  assign n8546 = ~n1801 & n8545 ;
  assign n8547 = n5045 & n8546 ;
  assign n8548 = n4205 & ~n8547 ;
  assign n8549 = n2713 ^ n836 ^ 1'b0 ;
  assign n8550 = n8549 ^ n5412 ^ 1'b0 ;
  assign n8553 = x110 & n610 ;
  assign n8554 = ~x123 & n8553 ;
  assign n8551 = n1922 & n3495 ;
  assign n8552 = ~n7337 & n8551 ;
  assign n8555 = n8554 ^ n8552 ^ 1'b0 ;
  assign n8556 = ( n2495 & n6771 ) | ( n2495 & n8555 ) | ( n6771 & n8555 ) ;
  assign n8557 = n6202 & n8556 ;
  assign n8558 = n2395 & ~n5305 ;
  assign n8559 = ~n7139 & n7617 ;
  assign n8560 = n8559 ^ n7251 ^ 1'b0 ;
  assign n8561 = n2523 & n4768 ;
  assign n8562 = ~n4036 & n8561 ;
  assign n8563 = x164 & n411 ;
  assign n8564 = n8563 ^ n2147 ^ 1'b0 ;
  assign n8565 = n433 | n8564 ;
  assign n8566 = ~n2162 & n8565 ;
  assign n8567 = n8562 & n8566 ;
  assign n8568 = n5618 & ~n6122 ;
  assign n8569 = ~n610 & n8568 ;
  assign n8570 = n8569 ^ n6385 ^ 1'b0 ;
  assign n8571 = n6412 ^ n979 ^ 1'b0 ;
  assign n8572 = n1750 & ~n8571 ;
  assign n8573 = ~n1489 & n3714 ;
  assign n8574 = n8572 & n8573 ;
  assign n8575 = n8539 & n8574 ;
  assign n8576 = n2402 ^ n1085 ^ 1'b0 ;
  assign n8577 = n6875 & n8576 ;
  assign n8578 = n6185 ^ n5828 ^ n5411 ;
  assign n8579 = n6185 ^ n4590 ^ 1'b0 ;
  assign n8580 = n8579 ^ n5954 ^ 1'b0 ;
  assign n8581 = n7621 & ~n8580 ;
  assign n8582 = n3627 ^ n686 ^ 1'b0 ;
  assign n8583 = n6122 | n8582 ;
  assign n8584 = n5804 ^ n736 ^ 1'b0 ;
  assign n8585 = ~n3477 & n4693 ;
  assign n8586 = ( n3831 & n4658 ) | ( n3831 & ~n6393 ) | ( n4658 & ~n6393 ) ;
  assign n8587 = n6544 & n8586 ;
  assign n8588 = ~n405 & n5326 ;
  assign n8589 = n2706 ^ n880 ^ n793 ;
  assign n8590 = n6420 ^ n5289 ^ n4624 ;
  assign n8591 = n8589 | n8590 ;
  assign n8592 = n8588 & ~n8591 ;
  assign n8593 = n5131 ^ n4615 ^ 1'b0 ;
  assign n8594 = n3128 & n8593 ;
  assign n8599 = n3744 ^ n742 ^ 1'b0 ;
  assign n8596 = n6528 ^ n288 ^ 1'b0 ;
  assign n8597 = n768 | n8596 ;
  assign n8595 = ~n3972 & n5490 ;
  assign n8598 = n8597 ^ n8595 ^ 1'b0 ;
  assign n8600 = n8599 ^ n8598 ^ 1'b0 ;
  assign n8601 = n8594 & n8600 ;
  assign n8602 = n8601 ^ n8065 ^ x235 ;
  assign n8603 = ( n4342 & n4376 ) | ( n4342 & n8512 ) | ( n4376 & n8512 ) ;
  assign n8604 = n1063 | n8603 ;
  assign n8605 = n8077 & ~n8604 ;
  assign n8606 = n7172 ^ n4651 ^ 1'b0 ;
  assign n8607 = x115 & n3129 ;
  assign n8608 = n8607 ^ n6665 ^ 1'b0 ;
  assign n8609 = n4784 & ~n8608 ;
  assign n8610 = n8606 & n8609 ;
  assign n8611 = n1707 ^ n616 ^ 1'b0 ;
  assign n8612 = ~n872 & n8611 ;
  assign n8613 = n6182 & ~n8612 ;
  assign n8614 = n8613 ^ n3721 ^ 1'b0 ;
  assign n8617 = n2694 ^ x47 ^ 1'b0 ;
  assign n8618 = n4891 & ~n8617 ;
  assign n8615 = n7916 ^ n3122 ^ 1'b0 ;
  assign n8616 = n2350 | n8615 ;
  assign n8619 = n8618 ^ n8616 ^ 1'b0 ;
  assign n8620 = n5903 & ~n8619 ;
  assign n8621 = ( x161 & n8449 ) | ( x161 & n8620 ) | ( n8449 & n8620 ) ;
  assign n8622 = n8237 ^ n1838 ^ 1'b0 ;
  assign n8623 = n8622 ^ n7338 ^ n921 ;
  assign n8624 = ~n856 & n5210 ;
  assign n8625 = n8624 ^ n4380 ^ 1'b0 ;
  assign n8626 = ~n1724 & n4153 ;
  assign n8627 = ~n1639 & n8626 ;
  assign n8628 = n2465 ^ n311 ^ 1'b0 ;
  assign n8629 = ~n1106 & n8628 ;
  assign n8630 = n8629 ^ n7066 ^ 1'b0 ;
  assign n8631 = n8627 | n8630 ;
  assign n8632 = n8625 & ~n8631 ;
  assign n8633 = ~n3308 & n6973 ;
  assign n8634 = n8632 & n8633 ;
  assign n8635 = x211 & n8634 ;
  assign n8636 = n4200 & ~n4622 ;
  assign n8637 = n557 | n5968 ;
  assign n8638 = n2118 ^ n906 ^ 1'b0 ;
  assign n8639 = n2959 & n8638 ;
  assign n8640 = n607 & n2010 ;
  assign n8641 = n8640 ^ n2847 ^ 1'b0 ;
  assign n8642 = x167 & ~n8641 ;
  assign n8643 = ~n3273 & n8086 ;
  assign n8644 = x54 & ~n2445 ;
  assign n8645 = n8644 ^ n1548 ^ 1'b0 ;
  assign n8646 = n1288 & n8645 ;
  assign n8647 = n8646 ^ n1705 ^ 1'b0 ;
  assign n8648 = n1648 & n8647 ;
  assign n8649 = n3738 & ~n4241 ;
  assign n8650 = n5028 & ~n8649 ;
  assign n8651 = n8648 & n8650 ;
  assign n8652 = n2781 | n8090 ;
  assign n8653 = n8652 ^ x229 ^ 1'b0 ;
  assign n8654 = ( n1360 & ~n2046 ) | ( n1360 & n3466 ) | ( ~n2046 & n3466 ) ;
  assign n8655 = n1663 & ~n8654 ;
  assign n8656 = n3757 & ~n7745 ;
  assign n8657 = n8656 ^ n985 ^ 1'b0 ;
  assign n8658 = n1785 & n7010 ;
  assign n8659 = n8658 ^ n4846 ^ 1'b0 ;
  assign n8660 = ~n2162 & n3716 ;
  assign n8661 = n8660 ^ n1559 ^ 1'b0 ;
  assign n8662 = n8661 ^ n3282 ^ n1555 ;
  assign n8663 = n7569 & ~n8662 ;
  assign n8664 = ~n3707 & n8663 ;
  assign n8665 = ~n4676 & n5918 ;
  assign n8666 = n7960 ^ n5966 ^ 1'b0 ;
  assign n8667 = n8665 & ~n8666 ;
  assign n8668 = n6049 | n8667 ;
  assign n8669 = n8668 ^ n7364 ^ 1'b0 ;
  assign n8670 = n6015 ^ n4335 ^ 1'b0 ;
  assign n8671 = n3984 | n8670 ;
  assign n8672 = n1119 | n8671 ;
  assign n8673 = n7703 & n8672 ;
  assign n8674 = ~n2752 & n8673 ;
  assign n8675 = n2569 & ~n3572 ;
  assign n8676 = n6249 ^ n1816 ^ 1'b0 ;
  assign n8677 = n8675 & n8676 ;
  assign n8678 = n5581 ^ x253 ^ 1'b0 ;
  assign n8679 = n3196 & ~n4334 ;
  assign n8680 = ~n3487 & n8679 ;
  assign n8682 = n8547 ^ n647 ^ 1'b0 ;
  assign n8683 = ~n5728 & n8682 ;
  assign n8681 = n3259 & n5714 ;
  assign n8684 = n8683 ^ n8681 ^ n8526 ;
  assign n8685 = n2846 ^ n2320 ^ 1'b0 ;
  assign n8686 = n7300 | n8685 ;
  assign n8687 = n1868 & n2558 ;
  assign n8688 = ~n2390 & n8687 ;
  assign n8689 = n2858 ^ n2345 ^ n719 ;
  assign n8690 = n8689 ^ n6142 ^ x15 ;
  assign n8691 = n8688 & ~n8690 ;
  assign n8692 = ~n3413 & n7137 ;
  assign n8693 = n1633 & n3410 ;
  assign n8694 = ~n4694 & n8693 ;
  assign n8695 = n2276 | n3003 ;
  assign n8696 = n4703 & ~n8695 ;
  assign n8697 = ~n5778 & n8271 ;
  assign n8698 = n1536 | n6309 ;
  assign n8699 = n8698 ^ n1944 ^ 1'b0 ;
  assign n8700 = n6775 & n7668 ;
  assign n8701 = n8700 ^ n2108 ^ 1'b0 ;
  assign n8702 = ~x7 & n2856 ;
  assign n8703 = ~n8701 & n8702 ;
  assign n8704 = ~n3874 & n8703 ;
  assign n8705 = n3723 & ~n8073 ;
  assign n8706 = ~n5116 & n5804 ;
  assign n8707 = ~n3939 & n8706 ;
  assign n8708 = n288 & ~n8707 ;
  assign n8709 = n7527 ^ n5417 ^ 1'b0 ;
  assign n8711 = n1889 & n4027 ;
  assign n8710 = n536 & ~n3847 ;
  assign n8712 = n8711 ^ n8710 ^ 1'b0 ;
  assign n8714 = x17 & ~n8313 ;
  assign n8715 = n8714 ^ n1823 ^ 1'b0 ;
  assign n8713 = n5833 | n6268 ;
  assign n8716 = n8715 ^ n8713 ^ 1'b0 ;
  assign n8717 = n7107 ^ n4835 ^ n1680 ;
  assign n8718 = n6136 | n8717 ;
  assign n8719 = n6161 | n8718 ;
  assign n8720 = n8719 ^ x247 ^ 1'b0 ;
  assign n8721 = n5016 ^ n4436 ^ 1'b0 ;
  assign n8722 = ( n747 & n1021 ) | ( n747 & n8721 ) | ( n1021 & n8721 ) ;
  assign n8723 = n2227 ^ n1188 ^ x190 ;
  assign n8724 = n1031 | n2438 ;
  assign n8725 = n8724 ^ x210 ^ 1'b0 ;
  assign n8726 = ( n4409 & n8723 ) | ( n4409 & n8725 ) | ( n8723 & n8725 ) ;
  assign n8727 = ~n4042 & n8726 ;
  assign n8728 = ~n8722 & n8727 ;
  assign n8729 = ( n6087 & n7685 ) | ( n6087 & n8728 ) | ( n7685 & n8728 ) ;
  assign n8734 = n6211 ^ x63 ^ 1'b0 ;
  assign n8733 = n3709 | n5375 ;
  assign n8735 = n8734 ^ n8733 ^ 1'b0 ;
  assign n8736 = n8735 ^ n2965 ^ 1'b0 ;
  assign n8737 = ~n3894 & n8736 ;
  assign n8730 = ~n2076 & n4595 ;
  assign n8731 = n8730 ^ n2444 ^ 1'b0 ;
  assign n8732 = n5874 | n8731 ;
  assign n8738 = n8737 ^ n8732 ^ 1'b0 ;
  assign n8739 = n8729 & n8738 ;
  assign n8740 = ( ~n1769 & n3467 ) | ( ~n1769 & n3640 ) | ( n3467 & n3640 ) ;
  assign n8741 = n538 & ~n6352 ;
  assign n8742 = n8741 ^ n7616 ^ 1'b0 ;
  assign n8743 = n3145 ^ n2903 ^ 1'b0 ;
  assign n8744 = n4135 & ~n8743 ;
  assign n8745 = n8742 & n8744 ;
  assign n8746 = ~n8740 & n8745 ;
  assign n8747 = n1033 ^ x88 ^ 1'b0 ;
  assign n8748 = n8747 ^ n3140 ^ 1'b0 ;
  assign n8749 = n6296 | n8748 ;
  assign n8750 = n2827 & ~n8749 ;
  assign n8751 = n8750 ^ n896 ^ 1'b0 ;
  assign n8752 = n8751 ^ n7077 ^ n3583 ;
  assign n8753 = x15 & ~n6820 ;
  assign n8754 = n8753 ^ n4721 ^ 1'b0 ;
  assign n8755 = n2703 ^ n1451 ^ x182 ;
  assign n8758 = n599 & ~n3232 ;
  assign n8759 = n8758 ^ n5811 ^ 1'b0 ;
  assign n8756 = n2500 ^ n358 ^ 1'b0 ;
  assign n8757 = ~n650 & n8756 ;
  assign n8760 = n8759 ^ n8757 ^ 1'b0 ;
  assign n8761 = n8760 ^ x220 ^ 1'b0 ;
  assign n8762 = n8755 & ~n8761 ;
  assign n8763 = ( n471 & n1152 ) | ( n471 & n1581 ) | ( n1152 & n1581 ) ;
  assign n8764 = n869 & n2024 ;
  assign n8765 = n8764 ^ n2893 ^ 1'b0 ;
  assign n8766 = n8765 ^ n2418 ^ 1'b0 ;
  assign n8767 = ~n8763 & n8766 ;
  assign n8768 = n8767 ^ n7607 ^ 1'b0 ;
  assign n8769 = n4257 & n8768 ;
  assign n8770 = n4493 & ~n5663 ;
  assign n8771 = n1275 | n5667 ;
  assign n8772 = n8770 & ~n8771 ;
  assign n8773 = n3410 ^ n1304 ^ 1'b0 ;
  assign n8774 = n8773 ^ n8216 ^ 1'b0 ;
  assign n8775 = ( ~n3821 & n7654 ) | ( ~n3821 & n8774 ) | ( n7654 & n8774 ) ;
  assign n8776 = n3915 ^ n2939 ^ n2184 ;
  assign n8777 = ( ~n677 & n843 ) | ( ~n677 & n2543 ) | ( n843 & n2543 ) ;
  assign n8778 = n8777 ^ n6417 ^ n3664 ;
  assign n8779 = n8778 ^ n3725 ^ 1'b0 ;
  assign n8780 = ( n6548 & n8776 ) | ( n6548 & ~n8779 ) | ( n8776 & ~n8779 ) ;
  assign n8781 = n319 | n5479 ;
  assign n8782 = ( n3118 & n8632 ) | ( n3118 & ~n8781 ) | ( n8632 & ~n8781 ) ;
  assign n8784 = n4175 ^ n1540 ^ 1'b0 ;
  assign n8785 = n1665 & ~n8784 ;
  assign n8783 = n3738 & ~n8413 ;
  assign n8786 = n8785 ^ n8783 ^ 1'b0 ;
  assign n8787 = ~n6259 & n8786 ;
  assign n8788 = n4060 ^ n894 ^ 1'b0 ;
  assign n8789 = n485 & n8788 ;
  assign n8790 = n6101 & n8789 ;
  assign n8791 = ( x121 & ~n3382 ) | ( x121 & n4351 ) | ( ~n3382 & n4351 ) ;
  assign n8792 = n6176 & n6841 ;
  assign n8793 = ~n8791 & n8792 ;
  assign n8794 = n1088 & n5306 ;
  assign n8795 = ~n2522 & n8794 ;
  assign n8796 = n8795 ^ n4584 ^ 1'b0 ;
  assign n8797 = ~n405 & n8796 ;
  assign n8798 = n8797 ^ n5338 ^ 1'b0 ;
  assign n8799 = ~n4880 & n8798 ;
  assign n8800 = n1809 & ~n2247 ;
  assign n8801 = ~n3523 & n6714 ;
  assign n8802 = ~n8800 & n8801 ;
  assign n8803 = ( x111 & n3232 ) | ( x111 & ~n3615 ) | ( n3232 & ~n3615 ) ;
  assign n8804 = n8803 ^ n6715 ^ 1'b0 ;
  assign n8805 = n4535 & ~n8804 ;
  assign n8806 = n3324 | n5433 ;
  assign n8807 = n4820 & ~n8806 ;
  assign n8808 = n7439 ^ n5840 ^ 1'b0 ;
  assign n8809 = n5920 ^ n1999 ^ n838 ;
  assign n8810 = n8809 ^ n7778 ^ n3183 ;
  assign n8811 = n8810 ^ n636 ^ 1'b0 ;
  assign n8812 = ~n1390 & n2335 ;
  assign n8813 = n8812 ^ n480 ^ 1'b0 ;
  assign n8814 = ~n948 & n2260 ;
  assign n8815 = n8814 ^ n3832 ^ 1'b0 ;
  assign n8816 = n8815 ^ n5882 ^ 1'b0 ;
  assign n8817 = n8813 & ~n8816 ;
  assign n8818 = n6074 ^ n3829 ^ 1'b0 ;
  assign n8819 = ~n5698 & n8818 ;
  assign n8820 = n5541 ^ n4114 ^ n3879 ;
  assign n8821 = n2768 ^ n2224 ^ 1'b0 ;
  assign n8822 = ~n5410 & n8821 ;
  assign n8823 = n8822 ^ x82 ^ 1'b0 ;
  assign n8824 = n8823 ^ n2213 ^ 1'b0 ;
  assign n8825 = n7068 & n7847 ;
  assign n8826 = n7001 ^ n5149 ^ 1'b0 ;
  assign n8827 = n488 & ~n4912 ;
  assign n8828 = n2155 & n8827 ;
  assign n8830 = n1589 ^ n446 ^ x245 ;
  assign n8829 = n1564 & ~n1724 ;
  assign n8831 = n8830 ^ n8829 ^ n3021 ;
  assign n8832 = ~n8828 & n8831 ;
  assign n8833 = ~n6926 & n8832 ;
  assign n8834 = x169 & ~n8833 ;
  assign n8835 = n7910 ^ n5396 ^ n1947 ;
  assign n8836 = n8835 ^ n8421 ^ 1'b0 ;
  assign n8837 = x96 & ~n867 ;
  assign n8838 = n8837 ^ n5334 ^ 1'b0 ;
  assign n8839 = n2854 & ~n8838 ;
  assign n8840 = n6152 ^ n636 ^ 1'b0 ;
  assign n8841 = n2749 & ~n8840 ;
  assign n8842 = n8841 ^ n1780 ^ x10 ;
  assign n8843 = n8842 ^ x254 ^ 1'b0 ;
  assign n8844 = n2947 | n8843 ;
  assign n8845 = ( x113 & ~n1423 ) | ( x113 & n5635 ) | ( ~n1423 & n5635 ) ;
  assign n8846 = n3239 ^ n3138 ^ 1'b0 ;
  assign n8847 = n4775 ^ n1724 ^ 1'b0 ;
  assign n8848 = ( n8664 & ~n8846 ) | ( n8664 & n8847 ) | ( ~n8846 & n8847 ) ;
  assign n8849 = n629 & ~n2712 ;
  assign n8850 = ~n4758 & n8849 ;
  assign n8851 = n2454 & n8850 ;
  assign n8852 = n5532 & ~n5801 ;
  assign n8853 = n2455 | n8852 ;
  assign n8854 = n8853 ^ n8328 ^ 1'b0 ;
  assign n8855 = n8851 | n8854 ;
  assign n8856 = n2968 & ~n4890 ;
  assign n8857 = n5383 ^ n1877 ^ 1'b0 ;
  assign n8858 = ~n3425 & n8857 ;
  assign n8859 = n1650 & ~n1780 ;
  assign n8860 = n8858 & ~n8859 ;
  assign n8861 = n8860 ^ n8101 ^ 1'b0 ;
  assign n8862 = ( ~n2495 & n6669 ) | ( ~n2495 & n8861 ) | ( n6669 & n8861 ) ;
  assign n8863 = n5538 & n5879 ;
  assign n8864 = n8863 ^ n6967 ^ 1'b0 ;
  assign n8865 = n8864 ^ n3375 ^ 1'b0 ;
  assign n8867 = n610 ^ n347 ^ 1'b0 ;
  assign n8868 = x43 & ~n312 ;
  assign n8869 = ~x43 & n8868 ;
  assign n8870 = n1261 | n8869 ;
  assign n8871 = n1261 & ~n8870 ;
  assign n8872 = n8867 & ~n8871 ;
  assign n8873 = ~n8867 & n8872 ;
  assign n8874 = n835 | n8873 ;
  assign n8875 = n8873 & ~n8874 ;
  assign n8876 = n8875 ^ n3095 ^ 1'b0 ;
  assign n8866 = n4518 ^ n2681 ^ x79 ;
  assign n8877 = n8876 ^ n8866 ^ n6866 ;
  assign n8878 = n1601 | n3021 ;
  assign n8879 = n8878 ^ n8648 ^ 1'b0 ;
  assign n8880 = n5367 & ~n8879 ;
  assign n8881 = n3126 & n8834 ;
  assign n8882 = n8881 ^ n3395 ^ 1'b0 ;
  assign n8883 = n4758 & n4806 ;
  assign n8884 = n8883 ^ n1111 ^ 1'b0 ;
  assign n8885 = n2269 & n3068 ;
  assign n8886 = n8885 ^ n2887 ^ 1'b0 ;
  assign n8887 = n8886 ^ n5748 ^ n972 ;
  assign n8888 = n8887 ^ n5223 ^ n1495 ;
  assign n8889 = n6737 ^ n4406 ^ n2907 ;
  assign n8890 = n4072 ^ n706 ^ 1'b0 ;
  assign n8891 = n6267 | n8890 ;
  assign n8892 = n8891 ^ n3429 ^ 1'b0 ;
  assign n8893 = n4980 & n8515 ;
  assign n8894 = ( n481 & ~n4183 ) | ( n481 & n8893 ) | ( ~n4183 & n8893 ) ;
  assign n8895 = n681 & n7495 ;
  assign n8899 = n3502 ^ n1943 ^ n877 ;
  assign n8900 = n3770 | n8899 ;
  assign n8896 = n1767 & n1780 ;
  assign n8897 = ~n1584 & n8896 ;
  assign n8898 = n8897 ^ n5361 ^ 1'b0 ;
  assign n8901 = n8900 ^ n8898 ^ n6458 ;
  assign n8902 = ( n1594 & n2739 ) | ( n1594 & ~n3845 ) | ( n2739 & ~n3845 ) ;
  assign n8903 = n8902 ^ n1837 ^ 1'b0 ;
  assign n8904 = n4821 ^ x63 ^ 1'b0 ;
  assign n8905 = n6246 | n8904 ;
  assign n8906 = ( ~n7499 & n8374 ) | ( ~n7499 & n8905 ) | ( n8374 & n8905 ) ;
  assign n8907 = ~n2329 & n3213 ;
  assign n8908 = ~n1660 & n8907 ;
  assign n8909 = n4917 ^ n4545 ^ 1'b0 ;
  assign n8910 = n8908 | n8909 ;
  assign n8911 = n869 & n8910 ;
  assign n8913 = n5305 ^ n4736 ^ n4322 ;
  assign n8912 = n6458 ^ n5172 ^ 1'b0 ;
  assign n8914 = n8913 ^ n8912 ^ n6425 ;
  assign n8915 = n6360 ^ n1230 ^ 1'b0 ;
  assign n8916 = n8915 ^ n898 ^ 1'b0 ;
  assign n8917 = n3533 & ~n8916 ;
  assign n8918 = n8917 ^ n5851 ^ 1'b0 ;
  assign n8919 = n655 | n8918 ;
  assign n8920 = n601 ^ n288 ^ 1'b0 ;
  assign n8921 = n8919 | n8920 ;
  assign n8922 = n8167 & ~n8921 ;
  assign n8923 = n8922 ^ x235 ^ 1'b0 ;
  assign n8924 = x178 | n3641 ;
  assign n8925 = ~n4072 & n8924 ;
  assign n8926 = n8925 ^ n2775 ^ 1'b0 ;
  assign n8927 = ~n3552 & n8926 ;
  assign n8928 = n2352 & n6585 ;
  assign n8929 = ~n8236 & n8928 ;
  assign n8930 = n1685 | n1911 ;
  assign n8931 = n8930 ^ x245 ^ 1'b0 ;
  assign n8932 = n1261 | n8375 ;
  assign n8933 = n995 ^ n773 ^ 1'b0 ;
  assign n8934 = n8933 ^ n4041 ^ n3275 ;
  assign n8935 = x83 & n8934 ;
  assign n8936 = ~n6003 & n8935 ;
  assign n8937 = n4872 | n6260 ;
  assign n8938 = n8937 ^ n2168 ^ 1'b0 ;
  assign n8939 = n8938 ^ n2795 ^ 1'b0 ;
  assign n8940 = ~n8305 & n8939 ;
  assign n8941 = n5977 ^ n2008 ^ 1'b0 ;
  assign n8942 = n7226 ^ n5216 ^ n2234 ;
  assign n8943 = n7313 & n8942 ;
  assign n8944 = n8943 ^ n5313 ^ 1'b0 ;
  assign n8945 = n1462 ^ n1026 ^ 1'b0 ;
  assign n8946 = ( n1106 & n4812 ) | ( n1106 & n5421 ) | ( n4812 & n5421 ) ;
  assign n8947 = ( n3888 & n4160 ) | ( n3888 & n6344 ) | ( n4160 & n6344 ) ;
  assign n8948 = ( ~n271 & n8946 ) | ( ~n271 & n8947 ) | ( n8946 & n8947 ) ;
  assign n8949 = n5930 ^ n3085 ^ n1518 ;
  assign n8950 = n8949 ^ n7488 ^ 1'b0 ;
  assign n8951 = n1378 | n8950 ;
  assign n8955 = n2941 | n4520 ;
  assign n8952 = n5092 & n5339 ;
  assign n8953 = ~n1585 & n8952 ;
  assign n8954 = n8826 & ~n8953 ;
  assign n8956 = n8955 ^ n8954 ^ 1'b0 ;
  assign n8957 = ( x22 & n872 ) | ( x22 & n2706 ) | ( n872 & n2706 ) ;
  assign n8958 = n6402 | n8957 ;
  assign n8959 = n2635 | n8958 ;
  assign n8960 = n6223 ^ n3024 ^ 1'b0 ;
  assign n8961 = n5613 & ~n8960 ;
  assign n8962 = n3445 & n7418 ;
  assign n8963 = x73 & n8962 ;
  assign n8964 = n4432 ^ n1140 ^ 1'b0 ;
  assign n8965 = n8964 ^ n6866 ^ n1311 ;
  assign n8966 = n2248 | n8712 ;
  assign n8969 = ~n1515 & n2638 ;
  assign n8970 = n3617 ^ n1947 ^ 1'b0 ;
  assign n8971 = ~n8969 & n8970 ;
  assign n8972 = ( n558 & n838 ) | ( n558 & ~n8971 ) | ( n838 & ~n8971 ) ;
  assign n8967 = n5014 ^ n1877 ^ 1'b0 ;
  assign n8968 = n5834 | n8967 ;
  assign n8973 = n8972 ^ n8968 ^ 1'b0 ;
  assign n8974 = n3378 & n8973 ;
  assign n8975 = n847 & ~n1546 ;
  assign n8976 = ~n2437 & n8975 ;
  assign n8977 = n8976 ^ n7832 ^ n5460 ;
  assign n8978 = n5471 ^ n4820 ^ n937 ;
  assign n8979 = x183 ^ x74 ^ 1'b0 ;
  assign n8980 = ~n1313 & n8979 ;
  assign n8981 = n5973 & n8980 ;
  assign n8982 = n8981 ^ n6565 ^ 1'b0 ;
  assign n8983 = n7690 ^ n1540 ^ 1'b0 ;
  assign n8984 = n3088 & ~n8983 ;
  assign n8985 = n4826 & n8984 ;
  assign n8986 = n8985 ^ n1692 ^ n922 ;
  assign n8987 = n8982 & n8986 ;
  assign n8988 = n8978 & n8987 ;
  assign n8989 = n8134 ^ n686 ^ 1'b0 ;
  assign n8990 = ( n3759 & n8590 ) | ( n3759 & ~n8989 ) | ( n8590 & ~n8989 ) ;
  assign n8991 = n5099 ^ n2547 ^ 1'b0 ;
  assign n8992 = n5954 | n8991 ;
  assign n8993 = n8992 ^ n412 ^ 1'b0 ;
  assign n8994 = ~n2447 & n8622 ;
  assign n8995 = n1976 & n6504 ;
  assign n8996 = n5243 ^ n3435 ^ 1'b0 ;
  assign n8997 = ( ~n1148 & n6001 ) | ( ~n1148 & n6842 ) | ( n6001 & n6842 ) ;
  assign n8998 = n8996 & ~n8997 ;
  assign n8999 = n3294 ^ n924 ^ 1'b0 ;
  assign n9000 = ~n1788 & n8999 ;
  assign n9001 = n5647 & n9000 ;
  assign n9002 = n8030 ^ n5247 ^ 1'b0 ;
  assign n9007 = n3548 & n8545 ;
  assign n9008 = ~n3116 & n9007 ;
  assign n9003 = x89 | n2597 ;
  assign n9004 = n436 | n9003 ;
  assign n9005 = n2550 & ~n9004 ;
  assign n9006 = n9005 ^ n3126 ^ n2877 ;
  assign n9009 = n9008 ^ n9006 ^ 1'b0 ;
  assign n9010 = n547 & n1860 ;
  assign n9011 = n9010 ^ n963 ^ 1'b0 ;
  assign n9012 = ~n2179 & n9011 ;
  assign n9013 = n8548 | n9012 ;
  assign n9014 = n9009 & ~n9013 ;
  assign n9015 = n8893 ^ n4701 ^ n3727 ;
  assign n9016 = n281 & ~n6071 ;
  assign n9017 = n9016 ^ x15 ^ 1'b0 ;
  assign n9018 = ~n1200 & n2806 ;
  assign n9019 = n9018 ^ n6882 ^ 1'b0 ;
  assign n9020 = n9017 & ~n9019 ;
  assign n9021 = n3136 ^ n1678 ^ 1'b0 ;
  assign n9022 = n704 ^ x247 ^ 1'b0 ;
  assign n9023 = ~n3958 & n9022 ;
  assign n9024 = ( n5098 & n9021 ) | ( n5098 & ~n9023 ) | ( n9021 & ~n9023 ) ;
  assign n9025 = n1063 ^ n527 ^ 1'b0 ;
  assign n9026 = n5629 ^ n1150 ^ 1'b0 ;
  assign n9027 = n9025 | n9026 ;
  assign n9028 = ( n4406 & n6338 ) | ( n4406 & ~n8773 ) | ( n6338 & ~n8773 ) ;
  assign n9029 = n3404 | n4960 ;
  assign n9030 = n9028 & n9029 ;
  assign n9031 = n1625 | n5473 ;
  assign n9032 = n6824 & ~n9031 ;
  assign n9033 = n9032 ^ n3421 ^ 1'b0 ;
  assign n9034 = n4455 & ~n5428 ;
  assign n9035 = ~n7070 & n8961 ;
  assign n9037 = n744 & ~n3675 ;
  assign n9038 = ~n5357 & n9037 ;
  assign n9039 = n9038 ^ n4031 ^ n1205 ;
  assign n9036 = n6140 ^ n4852 ^ 1'b0 ;
  assign n9040 = n9039 ^ n9036 ^ 1'b0 ;
  assign n9041 = ~n3348 & n5584 ;
  assign n9042 = ~n5282 & n9041 ;
  assign n9043 = n519 ^ n380 ^ 1'b0 ;
  assign n9044 = ~n9042 & n9043 ;
  assign n9045 = n4033 ^ n2322 ^ 1'b0 ;
  assign n9046 = n9045 ^ n1323 ^ 1'b0 ;
  assign n9047 = n2287 & n9046 ;
  assign n9048 = n4909 & ~n7887 ;
  assign n9049 = n3526 & n5791 ;
  assign n9050 = n8927 & n9049 ;
  assign n9051 = n4241 & n9050 ;
  assign n9052 = ~n2585 & n5341 ;
  assign n9053 = n4714 | n8547 ;
  assign n9054 = n1717 & ~n9053 ;
  assign n9055 = n616 | n2502 ;
  assign n9056 = n407 | n9055 ;
  assign n9057 = n2099 ^ n2008 ^ 1'b0 ;
  assign n9058 = n2014 & n5023 ;
  assign n9059 = ( x8 & ~n3588 ) | ( x8 & n8250 ) | ( ~n3588 & n8250 ) ;
  assign n9060 = n5837 ^ n3652 ^ n357 ;
  assign n9061 = ~n2431 & n9060 ;
  assign n9062 = n9061 ^ n4020 ^ 1'b0 ;
  assign n9063 = ~n4909 & n5020 ;
  assign n9064 = n9063 ^ n1980 ^ 1'b0 ;
  assign n9065 = ~n2250 & n7399 ;
  assign n9066 = n3098 | n7305 ;
  assign n9067 = n5744 ^ n2869 ^ n2656 ;
  assign n9068 = n9021 | n9067 ;
  assign n9069 = n9068 ^ n3688 ^ 1'b0 ;
  assign n9070 = n6937 ^ n5172 ^ 1'b0 ;
  assign n9071 = n1129 & n2882 ;
  assign n9072 = n9071 ^ n5888 ^ 1'b0 ;
  assign n9073 = n6228 ^ n2010 ^ 1'b0 ;
  assign n9074 = ~n3233 & n9073 ;
  assign n9075 = ( ~n1665 & n9072 ) | ( ~n1665 & n9074 ) | ( n9072 & n9074 ) ;
  assign n9076 = n840 | n981 ;
  assign n9077 = n9076 ^ n5968 ^ 1'b0 ;
  assign n9078 = n9077 ^ n2188 ^ 1'b0 ;
  assign n9079 = ( ~n2172 & n3746 ) | ( ~n2172 & n9078 ) | ( n3746 & n9078 ) ;
  assign n9080 = ~n3534 & n9079 ;
  assign n9081 = n8354 & n9080 ;
  assign n9082 = n3051 ^ n1517 ^ 1'b0 ;
  assign n9083 = ~n2467 & n9082 ;
  assign n9084 = n4808 ^ n3265 ^ n1641 ;
  assign n9085 = n2276 & n4236 ;
  assign n9086 = n9085 ^ n2240 ^ 1'b0 ;
  assign n9087 = ( x191 & ~n9084 ) | ( x191 & n9086 ) | ( ~n9084 & n9086 ) ;
  assign n9088 = n429 & ~n7310 ;
  assign n9089 = n5025 | n6128 ;
  assign n9090 = n9089 ^ n7674 ^ 1'b0 ;
  assign n9091 = ( n5302 & n9088 ) | ( n5302 & n9090 ) | ( n9088 & n9090 ) ;
  assign n9092 = ~n7828 & n9091 ;
  assign n9093 = n9092 ^ n4048 ^ 1'b0 ;
  assign n9094 = ( n2203 & n2296 ) | ( n2203 & n9093 ) | ( n2296 & n9093 ) ;
  assign n9095 = n7869 ^ n7261 ^ 1'b0 ;
  assign n9096 = n6758 & n9095 ;
  assign n9102 = ( n332 & ~n8629 ) | ( n332 & n8867 ) | ( ~n8629 & n8867 ) ;
  assign n9103 = n5736 | n9102 ;
  assign n9097 = n1489 ^ n387 ^ 1'b0 ;
  assign n9098 = n3548 & n5985 ;
  assign n9099 = n9097 & n9098 ;
  assign n9100 = n9099 ^ n4535 ^ 1'b0 ;
  assign n9101 = n1788 | n9100 ;
  assign n9104 = n9103 ^ n9101 ^ n2957 ;
  assign n9105 = ~n4719 & n5836 ;
  assign n9107 = n3403 ^ n3281 ^ 1'b0 ;
  assign n9108 = x221 & ~n9107 ;
  assign n9106 = n2539 & ~n2728 ;
  assign n9109 = n9108 ^ n9106 ^ 1'b0 ;
  assign n9110 = ~n7529 & n9109 ;
  assign n9111 = n1176 ^ n488 ^ 1'b0 ;
  assign n9112 = n3698 | n6377 ;
  assign n9116 = n679 & ~n3642 ;
  assign n9117 = n3814 & n9116 ;
  assign n9114 = n3492 ^ n1285 ^ 1'b0 ;
  assign n9115 = ~n3201 & n9114 ;
  assign n9118 = n9117 ^ n9115 ^ 1'b0 ;
  assign n9113 = n8334 ^ n3586 ^ 1'b0 ;
  assign n9119 = n9118 ^ n9113 ^ 1'b0 ;
  assign n9120 = n6342 ^ n5055 ^ 1'b0 ;
  assign n9121 = n4180 & ~n9120 ;
  assign n9125 = ~n1548 & n2023 ;
  assign n9126 = ~n3430 & n9125 ;
  assign n9122 = n5315 & ~n6117 ;
  assign n9123 = n6889 & n9122 ;
  assign n9124 = n5562 & ~n9123 ;
  assign n9127 = n9126 ^ n9124 ^ 1'b0 ;
  assign n9128 = n1679 ^ n1675 ^ 1'b0 ;
  assign n9129 = n6352 & ~n9128 ;
  assign n9130 = ~n9127 & n9129 ;
  assign n9131 = n6309 ^ n856 ^ 1'b0 ;
  assign n9132 = n4842 & ~n9131 ;
  assign n9133 = n4698 ^ n3256 ^ 1'b0 ;
  assign n9134 = ( n3296 & n7984 ) | ( n3296 & n9133 ) | ( n7984 & n9133 ) ;
  assign n9135 = n8616 ^ n2537 ^ 1'b0 ;
  assign n9136 = ~n3711 & n9135 ;
  assign n9137 = n9136 ^ n6751 ^ 1'b0 ;
  assign n9138 = n1850 & ~n2943 ;
  assign n9139 = ~n1250 & n9138 ;
  assign n9140 = n9139 ^ n3601 ^ 1'b0 ;
  assign n9141 = n3095 | n9140 ;
  assign n9142 = x101 & n5562 ;
  assign n9143 = n1066 & n9142 ;
  assign n9144 = n5185 & ~n9143 ;
  assign n9145 = x36 & ~n8151 ;
  assign n9146 = n9145 ^ n4286 ^ 1'b0 ;
  assign n9147 = n7024 ^ n2501 ^ 1'b0 ;
  assign n9148 = n4648 & ~n9147 ;
  assign n9149 = n3839 ^ n833 ^ 1'b0 ;
  assign n9150 = n3749 | n9149 ;
  assign n9151 = ( n5159 & n9148 ) | ( n5159 & n9150 ) | ( n9148 & n9150 ) ;
  assign n9152 = n1190 & ~n8501 ;
  assign n9153 = n1389 ^ x213 ^ 1'b0 ;
  assign n9154 = x71 | n3009 ;
  assign n9155 = n5130 ^ n332 ^ 1'b0 ;
  assign n9156 = n3652 | n4339 ;
  assign n9157 = n2473 ^ n271 ^ 1'b0 ;
  assign n9158 = n9157 ^ n7161 ^ 1'b0 ;
  assign n9159 = ~n3769 & n9158 ;
  assign n9160 = n353 & n9159 ;
  assign n9161 = n8032 & n9160 ;
  assign n9162 = n2166 & n5758 ;
  assign n9163 = n2292 & n9162 ;
  assign n9164 = ~n9161 & n9163 ;
  assign n9165 = n8543 ^ n2560 ^ x18 ;
  assign n9166 = n513 & ~n2171 ;
  assign n9167 = ~n6871 & n9166 ;
  assign n9168 = n9167 ^ n545 ^ 1'b0 ;
  assign n9169 = n9165 & ~n9168 ;
  assign n9170 = n3495 | n8164 ;
  assign n9171 = ~n4620 & n7338 ;
  assign n9172 = ~n5296 & n9171 ;
  assign n9173 = n298 & ~n3001 ;
  assign n9174 = ~n6694 & n9173 ;
  assign n9175 = ( ~n981 & n1498 ) | ( ~n981 & n2096 ) | ( n1498 & n2096 ) ;
  assign n9176 = n5079 & ~n9175 ;
  assign n9177 = n9176 ^ n8016 ^ 1'b0 ;
  assign n9178 = n8618 ^ n2539 ^ 1'b0 ;
  assign n9179 = n3150 | n9178 ;
  assign n9181 = n549 & ~n7172 ;
  assign n9182 = n9181 ^ n5460 ^ 1'b0 ;
  assign n9183 = ~n6138 & n9182 ;
  assign n9180 = ~n1108 & n1991 ;
  assign n9184 = n9183 ^ n9180 ^ 1'b0 ;
  assign n9185 = n9179 & ~n9184 ;
  assign n9186 = ~n9177 & n9185 ;
  assign n9187 = ~n6352 & n9186 ;
  assign n9188 = n2416 & n4195 ;
  assign n9189 = n5851 ^ n3515 ^ 1'b0 ;
  assign n9190 = n4549 & n9189 ;
  assign n9191 = n9190 ^ n5215 ^ 1'b0 ;
  assign n9192 = ~n2411 & n9191 ;
  assign n9193 = n9188 & n9192 ;
  assign n9194 = n9193 ^ x83 ^ 1'b0 ;
  assign n9195 = ( n2995 & n3624 ) | ( n2995 & n8231 ) | ( n3624 & n8231 ) ;
  assign n9196 = n7076 ^ n1619 ^ 1'b0 ;
  assign n9197 = n4868 ^ n1138 ^ 1'b0 ;
  assign n9198 = n759 & n9197 ;
  assign n9199 = n3132 ^ n543 ^ 1'b0 ;
  assign n9200 = n2492 ^ n1164 ^ 1'b0 ;
  assign n9201 = ~n2547 & n9200 ;
  assign n9202 = n9199 & n9201 ;
  assign n9203 = n9202 ^ n8024 ^ 1'b0 ;
  assign n9204 = ( n9196 & ~n9198 ) | ( n9196 & n9203 ) | ( ~n9198 & n9203 ) ;
  assign n9205 = ( ~x205 & n3466 ) | ( ~x205 & n4662 ) | ( n3466 & n4662 ) ;
  assign n9206 = n4205 | n4824 ;
  assign n9207 = n791 & ~n5264 ;
  assign n9208 = ( ~n2681 & n9206 ) | ( ~n2681 & n9207 ) | ( n9206 & n9207 ) ;
  assign n9209 = n9205 | n9208 ;
  assign n9210 = ~n1023 & n3095 ;
  assign n9211 = n9210 ^ n2224 ^ 1'b0 ;
  assign n9212 = n9211 ^ n6980 ^ 1'b0 ;
  assign n9213 = n7145 ^ n2549 ^ 1'b0 ;
  assign n9214 = n1098 & ~n8562 ;
  assign n9215 = n8223 ^ n4049 ^ n791 ;
  assign n9216 = n7112 ^ n5536 ^ 1'b0 ;
  assign n9217 = n9215 & n9216 ;
  assign n9218 = n1528 & n8645 ;
  assign n9219 = n9218 ^ n2626 ^ 1'b0 ;
  assign n9220 = n1066 & n7201 ;
  assign n9221 = n5976 ^ n1044 ^ 1'b0 ;
  assign n9229 = n2697 & ~n6616 ;
  assign n9230 = n9229 ^ n4812 ^ 1'b0 ;
  assign n9222 = n1017 ^ n347 ^ x172 ;
  assign n9223 = n9222 ^ n1691 ^ 1'b0 ;
  assign n9224 = n1874 & ~n9223 ;
  assign n9225 = x162 & ~n4701 ;
  assign n9226 = ~n3450 & n9225 ;
  assign n9227 = ( ~n2495 & n9224 ) | ( ~n2495 & n9226 ) | ( n9224 & n9226 ) ;
  assign n9228 = ~n6597 & n9227 ;
  assign n9231 = n9230 ^ n9228 ^ 1'b0 ;
  assign n9232 = ( ~n9220 & n9221 ) | ( ~n9220 & n9231 ) | ( n9221 & n9231 ) ;
  assign n9233 = ( n3176 & ~n6196 ) | ( n3176 & n9232 ) | ( ~n6196 & n9232 ) ;
  assign n9234 = n972 | n1421 ;
  assign n9235 = n1688 & ~n2463 ;
  assign n9236 = ~n1380 & n9235 ;
  assign n9237 = n3898 & n9236 ;
  assign n9238 = n727 | n9237 ;
  assign n9239 = n4591 | n9238 ;
  assign n9240 = n2558 & n7088 ;
  assign n9241 = n9240 ^ n1068 ^ 1'b0 ;
  assign n9242 = n7135 | n9241 ;
  assign n9243 = n4004 & n4748 ;
  assign n9244 = n2983 & n9243 ;
  assign n9245 = n9244 ^ n1671 ^ 1'b0 ;
  assign n9246 = n6389 ^ n449 ^ 1'b0 ;
  assign n9247 = n9032 ^ n4097 ^ n2116 ;
  assign n9248 = n2065 | n9247 ;
  assign n9249 = n9246 & ~n9248 ;
  assign n9250 = n4776 & n6914 ;
  assign n9251 = n9250 ^ n2991 ^ 1'b0 ;
  assign n9252 = n4881 ^ n1346 ^ 1'b0 ;
  assign n9253 = n5274 ^ n928 ^ 1'b0 ;
  assign n9254 = n3002 | n4440 ;
  assign n9255 = n9254 ^ x128 ^ 1'b0 ;
  assign n9256 = ~n6025 & n9255 ;
  assign n9257 = n9253 & n9256 ;
  assign n9259 = n749 & ~n4216 ;
  assign n9258 = n5887 ^ n5592 ^ n4342 ;
  assign n9260 = n9259 ^ n9258 ^ n2563 ;
  assign n9261 = n2342 | n9260 ;
  assign n9267 = n417 | n1741 ;
  assign n9262 = n6205 ^ n1266 ^ 1'b0 ;
  assign n9263 = n1048 & ~n9262 ;
  assign n9264 = n4701 ^ n1739 ^ 1'b0 ;
  assign n9265 = n2924 & n9264 ;
  assign n9266 = ~n9263 & n9265 ;
  assign n9268 = n9267 ^ n9266 ^ 1'b0 ;
  assign n9269 = ( n1308 & n2613 ) | ( n1308 & ~n9268 ) | ( n2613 & ~n9268 ) ;
  assign n9270 = n4041 | n7024 ;
  assign n9271 = n1129 & ~n9270 ;
  assign n9272 = n9271 ^ n729 ^ 1'b0 ;
  assign n9273 = n2436 & n9272 ;
  assign n9274 = n9273 ^ n2723 ^ n1213 ;
  assign n9275 = ( x254 & n2005 ) | ( x254 & n3121 ) | ( n2005 & n3121 ) ;
  assign n9276 = ( n1155 & n2336 ) | ( n1155 & ~n9275 ) | ( n2336 & ~n9275 ) ;
  assign n9277 = n9276 ^ n3371 ^ 1'b0 ;
  assign n9278 = n8143 & n9277 ;
  assign n9279 = n3424 ^ n3055 ^ x8 ;
  assign n9280 = n9279 ^ n1356 ^ x60 ;
  assign n9281 = x217 & ~n9280 ;
  assign n9282 = n9281 ^ n3164 ^ n2913 ;
  assign n9283 = n1530 | n4243 ;
  assign n9284 = n9283 ^ n3363 ^ 1'b0 ;
  assign n9285 = n1442 | n9284 ;
  assign n9286 = n9285 ^ n570 ^ 1'b0 ;
  assign n9287 = n9286 ^ n3648 ^ n2017 ;
  assign n9288 = n2824 | n5680 ;
  assign n9289 = n9288 ^ n3842 ^ 1'b0 ;
  assign n9290 = ( n3249 & ~n5443 ) | ( n3249 & n9289 ) | ( ~n5443 & n9289 ) ;
  assign n9291 = ~n8803 & n9290 ;
  assign n9292 = n9291 ^ n3326 ^ 1'b0 ;
  assign n9293 = n3465 & ~n4770 ;
  assign n9294 = ~n2338 & n6098 ;
  assign n9295 = n9294 ^ n3907 ^ 1'b0 ;
  assign n9296 = n9295 ^ n7679 ^ n6776 ;
  assign n9297 = n6838 & ~n8517 ;
  assign n9298 = n3710 ^ n2668 ^ 1'b0 ;
  assign n9299 = ( n2702 & n2728 ) | ( n2702 & n9298 ) | ( n2728 & n9298 ) ;
  assign n9300 = n9299 ^ n4927 ^ 1'b0 ;
  assign n9304 = ~n1481 & n1850 ;
  assign n9301 = n2769 | n4172 ;
  assign n9302 = n9301 ^ n1594 ^ 1'b0 ;
  assign n9303 = n2138 | n9302 ;
  assign n9305 = n9304 ^ n9303 ^ 1'b0 ;
  assign n9306 = ~n1564 & n6696 ;
  assign n9307 = n9306 ^ n5339 ^ 1'b0 ;
  assign n9308 = n9209 ^ n559 ^ 1'b0 ;
  assign n9309 = ~n9307 & n9308 ;
  assign n9310 = n358 & n1570 ;
  assign n9311 = ~n677 & n9310 ;
  assign n9312 = n3203 & ~n9311 ;
  assign n9313 = ~x97 & n9312 ;
  assign n9314 = n1689 ^ x74 ^ x67 ;
  assign n9315 = n817 & ~n5094 ;
  assign n9316 = n9314 & n9315 ;
  assign n9317 = ~n1697 & n9316 ;
  assign n9318 = n9317 ^ n8632 ^ 1'b0 ;
  assign n9319 = n3521 | n7995 ;
  assign n9320 = n3009 ^ n467 ^ 1'b0 ;
  assign n9321 = n5618 & ~n9320 ;
  assign n9322 = ~n7760 & n9321 ;
  assign n9323 = n3145 & ~n9322 ;
  assign n9324 = n9319 & n9323 ;
  assign n9325 = ~n6461 & n7000 ;
  assign n9326 = ~n1928 & n9325 ;
  assign n9327 = n9326 ^ n8421 ^ n6851 ;
  assign n9328 = ~n4917 & n6590 ;
  assign n9329 = ~x67 & n9328 ;
  assign n9331 = x5 & ~n4970 ;
  assign n9332 = n9331 ^ n4945 ^ 1'b0 ;
  assign n9330 = n2294 & n7577 ;
  assign n9333 = n9332 ^ n9330 ^ 1'b0 ;
  assign n9339 = n1527 ^ x34 ^ 1'b0 ;
  assign n9334 = n2181 & n7539 ;
  assign n9335 = x109 & ~n9334 ;
  assign n9336 = n9335 ^ n6375 ^ 1'b0 ;
  assign n9337 = n1404 | n9336 ;
  assign n9338 = n9337 ^ n3741 ^ 1'b0 ;
  assign n9340 = n9339 ^ n9338 ^ 1'b0 ;
  assign n9342 = n536 & ~n2019 ;
  assign n9343 = n681 | n9342 ;
  assign n9341 = x217 | n3920 ;
  assign n9344 = n9343 ^ n9341 ^ 1'b0 ;
  assign n9345 = ~n7527 & n9344 ;
  assign n9346 = ~n4895 & n6077 ;
  assign n9347 = n9035 | n9346 ;
  assign n9348 = ~n1201 & n8367 ;
  assign n9349 = ~n1793 & n9348 ;
  assign n9350 = ( x111 & ~n2959 ) | ( x111 & n4990 ) | ( ~n2959 & n4990 ) ;
  assign n9351 = ~n7406 & n9350 ;
  assign n9352 = ( ~n1232 & n2038 ) | ( ~n1232 & n3523 ) | ( n2038 & n3523 ) ;
  assign n9353 = n6681 & ~n9352 ;
  assign n9354 = n7580 & ~n9353 ;
  assign n9355 = n9354 ^ n5976 ^ 1'b0 ;
  assign n9356 = ( n8082 & n9351 ) | ( n8082 & ~n9355 ) | ( n9351 & ~n9355 ) ;
  assign n9357 = n1370 | n7549 ;
  assign n9358 = n9357 ^ n527 ^ 1'b0 ;
  assign n9359 = n9358 ^ n4913 ^ 1'b0 ;
  assign n9360 = ~n535 & n5504 ;
  assign n9361 = n9360 ^ n8139 ^ 1'b0 ;
  assign n9362 = n3212 & n3976 ;
  assign n9363 = ( x105 & n5669 ) | ( x105 & n7245 ) | ( n5669 & n7245 ) ;
  assign n9364 = n4077 ^ n1862 ^ n1253 ;
  assign n9365 = n9364 ^ x227 ^ 1'b0 ;
  assign n9366 = n3647 & n9365 ;
  assign n9367 = ( ~n2452 & n3175 ) | ( ~n2452 & n4244 ) | ( n3175 & n4244 ) ;
  assign n9368 = n3597 & n5141 ;
  assign n9369 = n9368 ^ n1360 ^ 1'b0 ;
  assign n9370 = x12 & n3733 ;
  assign n9371 = n2892 & n9370 ;
  assign n9372 = n7005 ^ n4580 ^ 1'b0 ;
  assign n9373 = ~n9371 & n9372 ;
  assign n9374 = n7378 ^ n5592 ^ n1233 ;
  assign n9377 = n872 | n4571 ;
  assign n9378 = n2517 & ~n9377 ;
  assign n9379 = n9378 ^ n2057 ^ 1'b0 ;
  assign n9375 = n4977 ^ n3672 ^ 1'b0 ;
  assign n9376 = n6591 & ~n9375 ;
  assign n9380 = n9379 ^ n9376 ^ 1'b0 ;
  assign n9381 = n9374 | n9380 ;
  assign n9382 = n6674 & ~n9364 ;
  assign n9383 = n9382 ^ n2174 ^ 1'b0 ;
  assign n9384 = n6951 ^ n5610 ^ 1'b0 ;
  assign n9385 = ~n9383 & n9384 ;
  assign n9386 = n3901 | n7925 ;
  assign n9387 = n9386 ^ n5415 ^ 1'b0 ;
  assign n9388 = x84 | n1604 ;
  assign n9389 = n3259 ^ n547 ^ 1'b0 ;
  assign n9390 = n9388 & n9389 ;
  assign n9391 = ~n7152 & n9390 ;
  assign n9392 = n9391 ^ n3781 ^ 1'b0 ;
  assign n9393 = n2087 & ~n9392 ;
  assign n9394 = ~n3454 & n9393 ;
  assign n9395 = n9150 ^ x53 ^ 1'b0 ;
  assign n9396 = n4338 & ~n9395 ;
  assign n9397 = n6236 & n9396 ;
  assign n9398 = ~n5853 & n9397 ;
  assign n9399 = n9398 ^ n6260 ^ n1004 ;
  assign n9400 = n6854 | n9399 ;
  assign n9401 = n9400 ^ n7598 ^ 1'b0 ;
  assign n9402 = n263 & ~n8989 ;
  assign n9403 = n3558 ^ n2715 ^ 1'b0 ;
  assign n9404 = n1340 & ~n9403 ;
  assign n9406 = ( n519 & n7001 ) | ( n519 & n9028 ) | ( n7001 & n9028 ) ;
  assign n9405 = ~n3842 & n8647 ;
  assign n9407 = n9406 ^ n9405 ^ 1'b0 ;
  assign n9408 = n1347 ^ x206 ^ 1'b0 ;
  assign n9409 = ( x228 & ~n9407 ) | ( x228 & n9408 ) | ( ~n9407 & n9408 ) ;
  assign n9410 = n1344 & ~n2900 ;
  assign n9411 = n9410 ^ n1021 ^ 1'b0 ;
  assign n9412 = n9411 ^ n2416 ^ 1'b0 ;
  assign n9413 = n921 & ~n9412 ;
  assign n9414 = n2441 | n8313 ;
  assign n9415 = n9414 ^ n6638 ^ 1'b0 ;
  assign n9416 = n9415 ^ n3716 ^ n2195 ;
  assign n9417 = n9413 & n9416 ;
  assign n9418 = ~n1716 & n9417 ;
  assign n9419 = ~n2081 & n4536 ;
  assign n9420 = n9419 ^ n7530 ^ 1'b0 ;
  assign n9421 = n6642 ^ n674 ^ 1'b0 ;
  assign n9422 = n451 & n5048 ;
  assign n9423 = n3961 ^ n3231 ^ n2135 ;
  assign n9424 = n292 | n3960 ;
  assign n9425 = n9424 ^ n7107 ^ 1'b0 ;
  assign n9426 = n9425 ^ n981 ^ 1'b0 ;
  assign n9427 = ~n4287 & n9426 ;
  assign n9428 = x187 & ~n6174 ;
  assign n9429 = n1055 & ~n9428 ;
  assign n9430 = ~n1701 & n5859 ;
  assign n9431 = n966 | n9430 ;
  assign n9434 = ~n1605 & n4901 ;
  assign n9435 = ~n3659 & n9434 ;
  assign n9433 = n2701 & n7476 ;
  assign n9436 = n9435 ^ n9433 ^ 1'b0 ;
  assign n9432 = n5719 ^ n4699 ^ n1645 ;
  assign n9437 = n9436 ^ n9432 ^ 1'b0 ;
  assign n9438 = ~n1208 & n3688 ;
  assign n9439 = n2785 | n9438 ;
  assign n9440 = n9439 ^ x122 ^ 1'b0 ;
  assign n9441 = n1138 & n8826 ;
  assign n9442 = n9441 ^ n2609 ^ 1'b0 ;
  assign n9443 = n7925 ^ n795 ^ 1'b0 ;
  assign n9444 = ~n4852 & n9443 ;
  assign n9445 = ~n4302 & n8931 ;
  assign n9446 = ~n2194 & n2317 ;
  assign n9447 = n9446 ^ n6305 ^ 1'b0 ;
  assign n9448 = ( n2713 & ~n4699 ) | ( n2713 & n5305 ) | ( ~n4699 & n5305 ) ;
  assign n9449 = n3001 ^ x33 ^ 1'b0 ;
  assign n9450 = n7488 | n9449 ;
  assign n9451 = ~n536 & n1418 ;
  assign n9452 = x118 & ~n5805 ;
  assign n9453 = n9452 ^ n8449 ^ 1'b0 ;
  assign n9454 = ~n5289 & n9453 ;
  assign n9455 = n9451 & n9454 ;
  assign n9456 = n7734 ^ n4769 ^ n1194 ;
  assign n9457 = n6995 ^ n6391 ^ 1'b0 ;
  assign n9458 = n5898 ^ n3547 ^ 1'b0 ;
  assign n9459 = n2993 & ~n9458 ;
  assign n9460 = n9459 ^ n9078 ^ 1'b0 ;
  assign n9461 = n3104 | n9460 ;
  assign n9462 = ( ~n438 & n9457 ) | ( ~n438 & n9461 ) | ( n9457 & n9461 ) ;
  assign n9463 = n9462 ^ n9331 ^ n7627 ;
  assign n9464 = n3225 & n9463 ;
  assign n9465 = n9464 ^ n6723 ^ 1'b0 ;
  assign n9468 = n338 & n2823 ;
  assign n9469 = n2601 | n9468 ;
  assign n9470 = n1488 | n9469 ;
  assign n9466 = n1767 & n2093 ;
  assign n9467 = ( n4896 & n5599 ) | ( n4896 & ~n9466 ) | ( n5599 & ~n9466 ) ;
  assign n9471 = n9470 ^ n9467 ^ n1850 ;
  assign n9474 = n2684 ^ n376 ^ 1'b0 ;
  assign n9475 = n5944 | n9474 ;
  assign n9472 = n2240 & ~n2352 ;
  assign n9473 = n4846 | n9472 ;
  assign n9476 = n9475 ^ n9473 ^ 1'b0 ;
  assign n9477 = ( n259 & n739 ) | ( n259 & ~n2984 ) | ( n739 & ~n2984 ) ;
  assign n9478 = n7950 ^ n1070 ^ 1'b0 ;
  assign n9479 = n3811 | n9478 ;
  assign n9480 = n7514 ^ n983 ^ n677 ;
  assign n9481 = ~n9479 & n9480 ;
  assign n9482 = ~n9477 & n9481 ;
  assign n9483 = n478 & ~n9482 ;
  assign n9484 = n3332 & ~n5023 ;
  assign n9485 = n5184 | n9484 ;
  assign n9486 = n9483 & ~n9485 ;
  assign n9487 = n9486 ^ n4797 ^ 1'b0 ;
  assign n9488 = n8980 & ~n9487 ;
  assign n9489 = n3475 | n3860 ;
  assign n9490 = n4123 & n5853 ;
  assign n9491 = n7342 ^ n2160 ^ 1'b0 ;
  assign n9492 = n8886 & ~n9491 ;
  assign n9493 = n7595 & n9492 ;
  assign n9494 = n9493 ^ n8651 ^ n1809 ;
  assign n9495 = n9490 | n9494 ;
  assign n9496 = n9489 | n9495 ;
  assign n9497 = n7976 ^ n3915 ^ n2291 ;
  assign n9499 = n1483 & n2066 ;
  assign n9500 = ~n1793 & n9499 ;
  assign n9501 = ( n3354 & n5811 ) | ( n3354 & n9500 ) | ( n5811 & n9500 ) ;
  assign n9502 = n3981 & ~n9501 ;
  assign n9498 = n6813 ^ n1228 ^ 1'b0 ;
  assign n9503 = n9502 ^ n9498 ^ 1'b0 ;
  assign n9504 = n3731 | n9503 ;
  assign n9505 = x122 & ~n5506 ;
  assign n9506 = n9505 ^ n7966 ^ 1'b0 ;
  assign n9507 = n4764 ^ n3728 ^ 1'b0 ;
  assign n9508 = n9506 & n9507 ;
  assign n9509 = ~n3806 & n9508 ;
  assign n9510 = ~n6621 & n9509 ;
  assign n9511 = n2841 & ~n4210 ;
  assign n9512 = ~n5483 & n9511 ;
  assign n9513 = n1590 & ~n9512 ;
  assign n9514 = ( n6912 & n8810 ) | ( n6912 & n9513 ) | ( n8810 & n9513 ) ;
  assign n9515 = n7210 & ~n9214 ;
  assign n9516 = n4966 & ~n6354 ;
  assign n9517 = n9516 ^ n8318 ^ 1'b0 ;
  assign n9518 = n3646 ^ n980 ^ n265 ;
  assign n9519 = n1861 & ~n2365 ;
  assign n9520 = n5677 & n9519 ;
  assign n9521 = n9520 ^ n4269 ^ 1'b0 ;
  assign n9522 = n9521 ^ n3281 ^ 1'b0 ;
  assign n9523 = n351 | n9522 ;
  assign n9524 = n9518 | n9523 ;
  assign n9526 = n2586 ^ n527 ^ n395 ;
  assign n9525 = n6214 ^ n3051 ^ x232 ;
  assign n9527 = n9526 ^ n9525 ^ 1'b0 ;
  assign n9528 = n4382 & n7581 ;
  assign n9529 = n4819 ^ n4097 ^ n2363 ;
  assign n9530 = n5661 ^ x235 ^ 1'b0 ;
  assign n9531 = ( n3584 & n3664 ) | ( n3584 & n9530 ) | ( n3664 & n9530 ) ;
  assign n9532 = n4002 | n9531 ;
  assign n9533 = n1869 & ~n4460 ;
  assign n9534 = n9533 ^ n4175 ^ 1'b0 ;
  assign n9535 = ( n548 & n1932 ) | ( n548 & n9534 ) | ( n1932 & n9534 ) ;
  assign n9536 = n1053 & n4878 ;
  assign n9537 = n9536 ^ n4943 ^ 1'b0 ;
  assign n9538 = ( n2431 & ~n5895 ) | ( n2431 & n9537 ) | ( ~n5895 & n9537 ) ;
  assign n9539 = n7138 ^ n5657 ^ n776 ;
  assign n9540 = n1807 & n9539 ;
  assign n9541 = n9540 ^ n1442 ^ 1'b0 ;
  assign n9542 = n5170 ^ n4146 ^ 1'b0 ;
  assign n9543 = n9542 ^ n3885 ^ 1'b0 ;
  assign n9544 = n326 & n9543 ;
  assign n9545 = n805 & ~n2910 ;
  assign n9546 = n9544 & ~n9545 ;
  assign n9547 = n3542 | n5467 ;
  assign n9548 = n1803 & ~n9547 ;
  assign n9549 = n9548 ^ x91 ^ 1'b0 ;
  assign n9550 = x191 & ~n9549 ;
  assign n9551 = x246 | n3558 ;
  assign n9552 = n3126 & ~n9551 ;
  assign n9553 = n9552 ^ n9381 ^ n8866 ;
  assign n9554 = n806 | n1343 ;
  assign n9555 = n9554 ^ n3600 ^ n3551 ;
  assign n9556 = n6667 ^ n5178 ^ 1'b0 ;
  assign n9557 = n3642 & ~n9556 ;
  assign n9558 = n9557 ^ n9456 ^ 1'b0 ;
  assign n9559 = ~x3 & n9558 ;
  assign n9560 = n2015 ^ x241 ^ 1'b0 ;
  assign n9561 = n8491 | n9560 ;
  assign n9562 = n9561 ^ n4150 ^ n2581 ;
  assign n9563 = n984 & n9562 ;
  assign n9564 = n3882 & n9563 ;
  assign n9565 = ~n822 & n5380 ;
  assign n9566 = ~n2203 & n9565 ;
  assign n9567 = x226 & n9566 ;
  assign n9568 = ~n3244 & n6534 ;
  assign n9569 = n1550 ^ n490 ^ 1'b0 ;
  assign n9570 = ~n1475 & n1752 ;
  assign n9571 = n9438 & n9570 ;
  assign n9572 = n5081 | n9571 ;
  assign n9573 = n636 & ~n9572 ;
  assign n9574 = ~n2678 & n9573 ;
  assign n9575 = n9574 ^ n5778 ^ 1'b0 ;
  assign n9576 = x86 ^ x15 ^ 1'b0 ;
  assign n9577 = n6760 | n9576 ;
  assign n9578 = n1056 & n4194 ;
  assign n9579 = n6047 ^ n5075 ^ 1'b0 ;
  assign n9580 = n9579 ^ n307 ^ 1'b0 ;
  assign n9581 = n9578 | n9580 ;
  assign n9582 = ( n2910 & n5462 ) | ( n2910 & n8616 ) | ( n5462 & n8616 ) ;
  assign n9583 = n1795 & ~n9582 ;
  assign n9584 = x61 & n3273 ;
  assign n9585 = ~n5053 & n9584 ;
  assign n9586 = n298 | n1281 ;
  assign n9587 = x59 & ~n9586 ;
  assign n9588 = ~n3193 & n9587 ;
  assign n9589 = n5208 ^ n3924 ^ 1'b0 ;
  assign n9590 = n9589 ^ x251 ^ 1'b0 ;
  assign n9591 = n5085 | n9590 ;
  assign n9592 = n9591 ^ n2692 ^ n932 ;
  assign n9593 = n7219 & n8887 ;
  assign n9594 = n9593 ^ n4050 ^ 1'b0 ;
  assign n9595 = n9594 ^ n3514 ^ 1'b0 ;
  assign n9597 = n647 | n694 ;
  assign n9598 = n9597 ^ x67 ^ 1'b0 ;
  assign n9596 = n7073 & n7793 ;
  assign n9599 = n9598 ^ n9596 ^ 1'b0 ;
  assign n9600 = ~n2463 & n5391 ;
  assign n9601 = n9600 ^ n6783 ^ n5629 ;
  assign n9602 = n721 | n9101 ;
  assign n9603 = n9602 ^ n8318 ^ 1'b0 ;
  assign n9604 = n5326 ^ n3316 ^ 1'b0 ;
  assign n9605 = x128 & n9604 ;
  assign n9606 = n4278 ^ n2661 ^ 1'b0 ;
  assign n9607 = ( n2503 & ~n4375 ) | ( n2503 & n9606 ) | ( ~n4375 & n9606 ) ;
  assign n9608 = n9607 ^ n4585 ^ 1'b0 ;
  assign n9609 = n8995 & ~n9608 ;
  assign n9610 = n9609 ^ n2688 ^ 1'b0 ;
  assign n9611 = n7776 ^ n1351 ^ n271 ;
  assign n9612 = x182 & ~n1212 ;
  assign n9613 = n6788 & ~n9612 ;
  assign n9614 = n5914 ^ n2882 ^ n1807 ;
  assign n9615 = ( n1179 & n2480 ) | ( n1179 & n9614 ) | ( n2480 & n9614 ) ;
  assign n9616 = n9448 & ~n9615 ;
  assign n9617 = ~n4057 & n4081 ;
  assign n9618 = ~n7678 & n9617 ;
  assign n9619 = n9618 ^ n6561 ^ 1'b0 ;
  assign n9620 = n6859 ^ n2899 ^ 1'b0 ;
  assign n9621 = n6030 & ~n9620 ;
  assign n9622 = n7997 & n9621 ;
  assign n9623 = n2549 ^ n626 ^ 1'b0 ;
  assign n9624 = n6681 ^ n5059 ^ 1'b0 ;
  assign n9625 = n2294 & n9624 ;
  assign n9626 = n8277 ^ n4194 ^ 1'b0 ;
  assign n9627 = n9625 & ~n9626 ;
  assign n9628 = n6955 & n9627 ;
  assign n9629 = ~n8350 & n9628 ;
  assign n9630 = n4918 & ~n5366 ;
  assign n9631 = n9630 ^ n5542 ^ 1'b0 ;
  assign n9632 = n9631 ^ n7666 ^ n2158 ;
  assign n9633 = n1801 & ~n9632 ;
  assign n9634 = n9633 ^ n1097 ^ 1'b0 ;
  assign n9635 = n596 & n995 ;
  assign n9636 = ~n6413 & n9635 ;
  assign n9637 = n3051 ^ n1900 ^ 1'b0 ;
  assign n9638 = n2847 & n9637 ;
  assign n9639 = n9638 ^ n3176 ^ n3127 ;
  assign n9640 = n1902 | n9639 ;
  assign n9641 = x144 & n443 ;
  assign n9642 = n9640 & n9641 ;
  assign n9643 = n1451 | n9642 ;
  assign n9644 = n9643 ^ n5049 ^ 1'b0 ;
  assign n9645 = n6985 | n9644 ;
  assign n9646 = ~n2281 & n7101 ;
  assign n9651 = n637 | n3705 ;
  assign n9652 = ( ~n4000 & n7577 ) | ( ~n4000 & n9651 ) | ( n7577 & n9651 ) ;
  assign n9648 = n745 ^ x62 ^ 1'b0 ;
  assign n9647 = n1732 & ~n3888 ;
  assign n9649 = n9648 ^ n9647 ^ 1'b0 ;
  assign n9650 = ~n4517 & n9649 ;
  assign n9653 = n9652 ^ n9650 ^ 1'b0 ;
  assign n9654 = n7318 ^ x37 ^ 1'b0 ;
  assign n9655 = ~n9653 & n9654 ;
  assign n9656 = ~x42 & n1509 ;
  assign n9657 = n5643 ^ n5311 ^ 1'b0 ;
  assign n9658 = n9656 & ~n9657 ;
  assign n9659 = n5235 ^ n4652 ^ 1'b0 ;
  assign n9660 = n9658 & ~n9659 ;
  assign n9661 = n9660 ^ n7778 ^ n6875 ;
  assign n9662 = ~x241 & n8744 ;
  assign n9663 = ~n821 & n9662 ;
  assign n9664 = n702 ^ n495 ^ 1'b0 ;
  assign n9665 = ~n3246 & n9664 ;
  assign n9666 = n2347 & n2963 ;
  assign n9667 = n9666 ^ n2444 ^ 1'b0 ;
  assign n9668 = n9667 ^ n7338 ^ n6414 ;
  assign n9669 = n9668 ^ n9500 ^ 1'b0 ;
  assign n9670 = ~n7381 & n9669 ;
  assign n9672 = ( n2031 & n6425 ) | ( n2031 & ~n9436 ) | ( n6425 & ~n9436 ) ;
  assign n9671 = n5673 ^ n1213 ^ 1'b0 ;
  assign n9673 = n9672 ^ n9671 ^ 1'b0 ;
  assign n9674 = n9119 | n9673 ;
  assign n9675 = n4084 & n8466 ;
  assign n9676 = ( ~n770 & n4209 ) | ( ~n770 & n4584 ) | ( n4209 & n4584 ) ;
  assign n9677 = n9676 ^ n860 ^ 1'b0 ;
  assign n9678 = n5131 | n9677 ;
  assign n9679 = n2882 & n3835 ;
  assign n9680 = n9679 ^ n8666 ^ 1'b0 ;
  assign n9681 = n2366 & ~n4216 ;
  assign n9682 = n2246 & n9681 ;
  assign n9683 = n2553 & ~n7613 ;
  assign n9684 = n9682 & n9683 ;
  assign n9685 = n9680 & ~n9684 ;
  assign n9686 = n9678 & n9685 ;
  assign n9687 = n8308 ^ n3436 ^ 1'b0 ;
  assign n9688 = n9687 ^ n399 ^ 1'b0 ;
  assign n9689 = ( n557 & ~n4034 ) | ( n557 & n9688 ) | ( ~n4034 & n9688 ) ;
  assign n9690 = n3953 ^ n3729 ^ 1'b0 ;
  assign n9691 = n2574 & n9690 ;
  assign n9692 = n9691 ^ n3301 ^ n402 ;
  assign n9693 = n4169 ^ n3493 ^ n3222 ;
  assign n9694 = n9693 ^ n6614 ^ n2544 ;
  assign n9695 = n2808 & ~n7685 ;
  assign n9696 = ~n781 & n1577 ;
  assign n9697 = n9696 ^ n1037 ^ 1'b0 ;
  assign n9698 = ~n9695 & n9697 ;
  assign n9699 = n9698 ^ n1091 ^ 1'b0 ;
  assign n9700 = n9699 ^ n6621 ^ n4853 ;
  assign n9701 = n5760 & n9090 ;
  assign n9702 = n3395 | n4582 ;
  assign n9703 = n7936 | n9702 ;
  assign n9704 = n9703 ^ n3362 ^ 1'b0 ;
  assign n9705 = n5131 ^ n3220 ^ 1'b0 ;
  assign n9706 = n2241 & n9705 ;
  assign n9707 = n4284 & ~n5294 ;
  assign n9708 = n9706 & n9707 ;
  assign n9709 = ~n3804 & n9699 ;
  assign n9710 = n1574 & ~n2597 ;
  assign n9711 = ( n5203 & ~n5647 ) | ( n5203 & n9710 ) | ( ~n5647 & n9710 ) ;
  assign n9712 = ~n9709 & n9711 ;
  assign n9713 = n9712 ^ n4776 ^ 1'b0 ;
  assign n9714 = n9713 ^ n7001 ^ 1'b0 ;
  assign n9715 = n9249 ^ n8507 ^ n388 ;
  assign n9716 = n365 & n4282 ;
  assign n9721 = n2922 ^ n1861 ^ 1'b0 ;
  assign n9722 = n1177 & n9721 ;
  assign n9723 = n9722 ^ n1605 ^ 1'b0 ;
  assign n9724 = n395 & ~n9723 ;
  assign n9717 = n1451 | n2284 ;
  assign n9718 = n9717 ^ n2264 ^ 1'b0 ;
  assign n9719 = n9718 ^ n6413 ^ 1'b0 ;
  assign n9720 = n559 & n9719 ;
  assign n9725 = n9724 ^ n9720 ^ n1027 ;
  assign n9726 = ~n9716 & n9725 ;
  assign n9727 = n6617 ^ n1079 ^ 1'b0 ;
  assign n9728 = n9199 ^ n6262 ^ 1'b0 ;
  assign n9729 = ~n367 & n9728 ;
  assign n9730 = n8525 ^ n4806 ^ n2561 ;
  assign n9731 = x132 | n2826 ;
  assign n9732 = n9730 & n9731 ;
  assign n9733 = ~n9729 & n9732 ;
  assign n9734 = n6388 ^ n1392 ^ 1'b0 ;
  assign n9735 = n4119 | n9734 ;
  assign n9736 = n9733 | n9735 ;
  assign n9737 = n9736 ^ n3917 ^ 1'b0 ;
  assign n9738 = n7161 ^ n4557 ^ 1'b0 ;
  assign n9739 = n4832 ^ n1657 ^ 1'b0 ;
  assign n9740 = ~n4466 & n9739 ;
  assign n9741 = n8782 & n9740 ;
  assign n9742 = n9741 ^ n9208 ^ 1'b0 ;
  assign n9743 = n6579 ^ n2694 ^ 1'b0 ;
  assign n9744 = n9743 ^ n987 ^ 1'b0 ;
  assign n9745 = n2523 | n9744 ;
  assign n9746 = ( n514 & n2991 ) | ( n514 & ~n8776 ) | ( n2991 & ~n8776 ) ;
  assign n9747 = n9746 ^ n1489 ^ 1'b0 ;
  assign n9748 = n6901 ^ n5804 ^ n3536 ;
  assign n9750 = ~n4191 & n5649 ;
  assign n9749 = n2907 | n4057 ;
  assign n9751 = n9750 ^ n9749 ^ 1'b0 ;
  assign n9752 = x106 & ~n4157 ;
  assign n9753 = n2368 & n4945 ;
  assign n9754 = n286 | n9753 ;
  assign n9755 = n9754 ^ n7674 ^ 1'b0 ;
  assign n9756 = x14 & ~n3910 ;
  assign n9757 = n1863 & n9756 ;
  assign n9758 = n707 & n5751 ;
  assign n9759 = ~n6604 & n9758 ;
  assign n9760 = n2182 | n9759 ;
  assign n9761 = n9757 & ~n9760 ;
  assign n9762 = n3979 ^ n3895 ^ 1'b0 ;
  assign n9763 = n7876 | n9762 ;
  assign n9764 = n3577 | n5473 ;
  assign n9765 = n9764 ^ n5637 ^ 1'b0 ;
  assign n9766 = n2640 | n5404 ;
  assign n9767 = n9766 ^ n4083 ^ 1'b0 ;
  assign n9768 = n9767 ^ x172 ^ 1'b0 ;
  assign n9769 = n2390 ^ n1396 ^ x199 ;
  assign n9770 = n7109 ^ n4787 ^ 1'b0 ;
  assign n9771 = n9769 & ~n9770 ;
  assign n9772 = n9771 ^ n3698 ^ 1'b0 ;
  assign n9773 = ( n3209 & ~n3394 ) | ( n3209 & n4272 ) | ( ~n3394 & n4272 ) ;
  assign n9774 = ( ~n6053 & n7426 ) | ( ~n6053 & n9773 ) | ( n7426 & n9773 ) ;
  assign n9775 = n5765 ^ n3712 ^ 1'b0 ;
  assign n9776 = n9775 ^ n2603 ^ n395 ;
  assign n9777 = ( ~n2883 & n3515 ) | ( ~n2883 & n9776 ) | ( n3515 & n9776 ) ;
  assign n9778 = n3517 & n9777 ;
  assign n9779 = n3150 | n9778 ;
  assign n9780 = n4077 ^ n3244 ^ n2630 ;
  assign n9781 = n9780 ^ x44 ^ 1'b0 ;
  assign n9782 = n6501 & n9781 ;
  assign n9783 = n8774 ^ n8163 ^ 1'b0 ;
  assign n9784 = n1938 ^ n1097 ^ 1'b0 ;
  assign n9785 = ( n7200 & n8447 ) | ( n7200 & ~n9784 ) | ( n8447 & ~n9784 ) ;
  assign n9786 = n6429 ^ n1155 ^ 1'b0 ;
  assign n9787 = n5193 | n8286 ;
  assign n9788 = n9786 | n9787 ;
  assign n9791 = n7992 ^ n1491 ^ 1'b0 ;
  assign n9789 = n4670 & n8824 ;
  assign n9790 = n7783 & n9789 ;
  assign n9792 = n9791 ^ n9790 ^ n5976 ;
  assign n9793 = n7557 ^ n5187 ^ 1'b0 ;
  assign n9794 = ~n5142 & n5232 ;
  assign n9795 = n9794 ^ n3333 ^ 1'b0 ;
  assign n9796 = ~n365 & n4344 ;
  assign n9797 = n9796 ^ n3740 ^ 1'b0 ;
  assign n9798 = n2726 & n3845 ;
  assign n9799 = n9798 ^ n6223 ^ 1'b0 ;
  assign n9800 = n4638 & ~n9799 ;
  assign n9801 = ~n9490 & n9800 ;
  assign n9802 = ~n5008 & n9801 ;
  assign n9803 = n9428 ^ n439 ^ 1'b0 ;
  assign n9804 = ~n9802 & n9803 ;
  assign n9805 = n9334 ^ n4186 ^ 1'b0 ;
  assign n9806 = n5521 ^ n1264 ^ 1'b0 ;
  assign n9807 = ~n9805 & n9806 ;
  assign n9809 = n6386 ^ n2129 ^ 1'b0 ;
  assign n9810 = n4148 | n9809 ;
  assign n9808 = n3205 & ~n6299 ;
  assign n9811 = n9810 ^ n9808 ^ n681 ;
  assign n9816 = x57 & ~n3689 ;
  assign n9812 = n1822 ^ n1466 ^ 1'b0 ;
  assign n9813 = n3551 & ~n9812 ;
  assign n9814 = n9813 ^ n3495 ^ 1'b0 ;
  assign n9815 = n2153 & ~n9814 ;
  assign n9817 = n9816 ^ n9815 ^ 1'b0 ;
  assign n9818 = n1233 | n5997 ;
  assign n9819 = n2574 | n9818 ;
  assign n9820 = n9819 ^ n2055 ^ x112 ;
  assign n9825 = x109 & x244 ;
  assign n9826 = n9825 ^ x61 ^ 1'b0 ;
  assign n9827 = n1450 | n8093 ;
  assign n9828 = n9827 ^ n6694 ^ 1'b0 ;
  assign n9829 = n9828 ^ n3316 ^ 1'b0 ;
  assign n9830 = ~n9826 & n9829 ;
  assign n9821 = n5565 ^ n4019 ^ 1'b0 ;
  assign n9822 = ~n5716 & n9821 ;
  assign n9823 = n2519 & n3453 ;
  assign n9824 = ~n9822 & n9823 ;
  assign n9831 = n9830 ^ n9824 ^ 1'b0 ;
  assign n9832 = n7578 ^ n535 ^ 1'b0 ;
  assign n9833 = ~n2888 & n3126 ;
  assign n9834 = n4026 | n9833 ;
  assign n9835 = n9832 & ~n9834 ;
  assign n9836 = n7884 ^ n2199 ^ 1'b0 ;
  assign n9837 = x243 & ~n1595 ;
  assign n9838 = n9837 ^ n2184 ^ 1'b0 ;
  assign n9839 = n6124 | n9838 ;
  assign n9840 = n3592 & ~n9839 ;
  assign n9841 = n3746 ^ n2497 ^ 1'b0 ;
  assign n9842 = n9840 | n9841 ;
  assign n9843 = n5331 & ~n8007 ;
  assign n9844 = ( ~n337 & n7365 ) | ( ~n337 & n7860 ) | ( n7365 & n7860 ) ;
  assign n9845 = ~n502 & n9844 ;
  assign n9846 = n1069 & n9845 ;
  assign n9847 = n5769 ^ n2838 ^ 1'b0 ;
  assign n9848 = ~n6262 & n6921 ;
  assign n9849 = n6988 ^ n6774 ^ 1'b0 ;
  assign n9850 = n7653 ^ n4371 ^ 1'b0 ;
  assign n9851 = n3939 & ~n9850 ;
  assign n9852 = n7785 & n9851 ;
  assign n9853 = n9852 ^ n1701 ^ 1'b0 ;
  assign n9854 = n2191 | n8688 ;
  assign n9855 = n3350 | n9854 ;
  assign n9856 = n9855 ^ n5790 ^ 1'b0 ;
  assign n9857 = n363 | n1913 ;
  assign n9858 = n3944 & n9857 ;
  assign n9859 = n4404 | n9858 ;
  assign n9860 = n9859 ^ n5828 ^ 1'b0 ;
  assign n9861 = n9860 ^ n2543 ^ n1500 ;
  assign n9862 = ~x127 & n9861 ;
  assign n9863 = n9856 & n9862 ;
  assign n9864 = n2970 & ~n4068 ;
  assign n9865 = n9864 ^ n4235 ^ 1'b0 ;
  assign n9866 = n9865 ^ x187 ^ 1'b0 ;
  assign n9867 = n803 & n9866 ;
  assign n9868 = n3625 | n9867 ;
  assign n9869 = n9868 ^ n7768 ^ 1'b0 ;
  assign n9870 = n1000 & n5645 ;
  assign n9871 = n9870 ^ n3443 ^ 1'b0 ;
  assign n9872 = ( ~n3320 & n3915 ) | ( ~n3320 & n5898 ) | ( n3915 & n5898 ) ;
  assign n9873 = n9872 ^ n9290 ^ 1'b0 ;
  assign n9874 = x129 & n1678 ;
  assign n9875 = x210 & ~n6064 ;
  assign n9876 = n9874 & n9875 ;
  assign n9877 = n9873 & n9876 ;
  assign n9878 = ~n5640 & n6982 ;
  assign n9879 = ~n6920 & n9878 ;
  assign n9880 = n3060 ^ n2365 ^ x172 ;
  assign n9881 = n2153 ^ n1024 ^ 1'b0 ;
  assign n9882 = n2241 & ~n8000 ;
  assign n9883 = n2542 ^ n2017 ^ 1'b0 ;
  assign n9884 = n9883 ^ n9374 ^ 1'b0 ;
  assign n9890 = n4723 ^ n637 ^ 1'b0 ;
  assign n9887 = ~n4832 & n6198 ;
  assign n9888 = n9887 ^ n1113 ^ 1'b0 ;
  assign n9889 = n2489 & n9888 ;
  assign n9891 = n9890 ^ n9889 ^ n3723 ;
  assign n9885 = n4500 ^ n3853 ^ 1'b0 ;
  assign n9886 = n5893 & ~n9885 ;
  assign n9892 = n9891 ^ n9886 ^ 1'b0 ;
  assign n9893 = n6531 & n9892 ;
  assign n9894 = n9893 ^ n3198 ^ 1'b0 ;
  assign n9895 = n1524 & n7937 ;
  assign n9898 = n1073 | n8539 ;
  assign n9899 = n9898 ^ n9222 ^ 1'b0 ;
  assign n9896 = n3340 ^ n604 ^ 1'b0 ;
  assign n9897 = ~n4957 & n9896 ;
  assign n9900 = n9899 ^ n9897 ^ n4002 ;
  assign n9901 = n2796 | n8771 ;
  assign n9902 = n4986 & n7709 ;
  assign n9903 = n7810 & ~n9902 ;
  assign n9904 = ~n2885 & n5575 ;
  assign n9905 = ( n1955 & ~n2748 ) | ( n1955 & n3077 ) | ( ~n2748 & n3077 ) ;
  assign n9906 = x77 & ~n2028 ;
  assign n9907 = n9906 ^ n3008 ^ 1'b0 ;
  assign n9908 = n9905 & n9907 ;
  assign n9909 = n1458 | n3859 ;
  assign n9913 = n1406 & n1646 ;
  assign n9914 = n9913 ^ n7569 ^ 1'b0 ;
  assign n9915 = n5115 ^ n3089 ^ 1'b0 ;
  assign n9916 = n9914 | n9915 ;
  assign n9910 = n8179 ^ n322 ^ 1'b0 ;
  assign n9911 = n694 | n9910 ;
  assign n9912 = n9911 ^ n8501 ^ 1'b0 ;
  assign n9917 = n9916 ^ n9912 ^ n4831 ;
  assign n9918 = n5361 ^ n1722 ^ 1'b0 ;
  assign n9919 = ( ~n2988 & n8884 ) | ( ~n2988 & n9918 ) | ( n8884 & n9918 ) ;
  assign n9920 = n1728 & ~n4209 ;
  assign n9921 = n9556 ^ n8133 ^ n7497 ;
  assign n9922 = n299 & n1317 ;
  assign n9923 = n9921 & n9922 ;
  assign n9925 = n7330 ^ n7087 ^ n3055 ;
  assign n9926 = n1823 | n9925 ;
  assign n9927 = n6296 & ~n9926 ;
  assign n9924 = x229 & n4145 ;
  assign n9928 = n9927 ^ n9924 ^ 1'b0 ;
  assign n9929 = ~n1287 & n2066 ;
  assign n9930 = n616 & n9929 ;
  assign n9931 = x98 & ~n9930 ;
  assign n9932 = ~n9928 & n9931 ;
  assign n9933 = n1567 ^ n911 ^ x46 ;
  assign n9934 = n9933 ^ n8231 ^ 1'b0 ;
  assign n9935 = n5110 & n5783 ;
  assign n9936 = n5528 & n9935 ;
  assign n9937 = n9411 & n9936 ;
  assign n9938 = ~n543 & n6543 ;
  assign n9939 = x234 & ~n9545 ;
  assign n9940 = n4657 ^ x220 ^ 1'b0 ;
  assign n9941 = n1827 & ~n9940 ;
  assign n9942 = n9941 ^ n7965 ^ n269 ;
  assign n9943 = n9942 ^ n4638 ^ 1'b0 ;
  assign n9944 = ~n2174 & n9943 ;
  assign n9945 = n2459 & ~n3246 ;
  assign n9946 = ( ~n3686 & n6349 ) | ( ~n3686 & n9945 ) | ( n6349 & n9945 ) ;
  assign n9947 = ~n2986 & n4144 ;
  assign n9948 = ~n4694 & n9947 ;
  assign n9949 = n3570 | n6381 ;
  assign n9950 = n6608 ^ n3325 ^ n2752 ;
  assign n9951 = n9950 ^ n3103 ^ 1'b0 ;
  assign n9952 = n5791 & ~n9951 ;
  assign n9953 = ( n3839 & ~n6420 ) | ( n3839 & n9952 ) | ( ~n6420 & n9952 ) ;
  assign n9954 = n4636 ^ n1929 ^ 1'b0 ;
  assign n9955 = n1965 & n9954 ;
  assign n9956 = n9955 ^ n4729 ^ n1887 ;
  assign n9957 = n3466 & n9143 ;
  assign n9958 = n3554 & ~n9957 ;
  assign n9959 = n4083 & n9958 ;
  assign n9960 = ( ~n5187 & n7753 ) | ( ~n5187 & n9959 ) | ( n7753 & n9959 ) ;
  assign n9961 = n2124 | n3132 ;
  assign n9962 = n2484 ^ n1840 ^ 1'b0 ;
  assign n9963 = ~n4759 & n9962 ;
  assign n9964 = n9963 ^ n6460 ^ 1'b0 ;
  assign n9965 = n9964 ^ n552 ^ 1'b0 ;
  assign n9966 = ( n2050 & n9961 ) | ( n2050 & ~n9965 ) | ( n9961 & ~n9965 ) ;
  assign n9967 = ~n4688 & n9207 ;
  assign n9968 = n9967 ^ n8105 ^ 1'b0 ;
  assign n9969 = ~n8394 & n8627 ;
  assign n9970 = n8589 | n9969 ;
  assign n9971 = n9968 & ~n9970 ;
  assign n9974 = n6282 ^ n4552 ^ 1'b0 ;
  assign n9975 = n4939 & n9974 ;
  assign n9972 = n1265 & n2996 ;
  assign n9973 = ~n4748 & n9972 ;
  assign n9976 = n9975 ^ n9973 ^ 1'b0 ;
  assign n9977 = n9976 ^ n1166 ^ 1'b0 ;
  assign n9978 = n9977 ^ n1255 ^ 1'b0 ;
  assign n9979 = ( ~n3163 & n5495 ) | ( ~n3163 & n6668 ) | ( n5495 & n6668 ) ;
  assign n9980 = n773 & n9979 ;
  assign n9981 = ~n9978 & n9980 ;
  assign n9982 = n3779 & ~n7515 ;
  assign n9983 = n7852 & ~n9982 ;
  assign n9984 = n2615 & n6567 ;
  assign n9985 = n9984 ^ n1041 ^ 1'b0 ;
  assign n9986 = n8537 ^ n5365 ^ n2232 ;
  assign n9987 = n7253 ^ n1150 ^ n1034 ;
  assign n9988 = ~n9255 & n9987 ;
  assign n9989 = ( ~n4703 & n9986 ) | ( ~n4703 & n9988 ) | ( n9986 & n9988 ) ;
  assign n9990 = n3734 & ~n3995 ;
  assign n9991 = n9990 ^ n4284 ^ 1'b0 ;
  assign n9992 = n2939 ^ n1633 ^ n1148 ;
  assign n9993 = n886 & n1170 ;
  assign n9994 = n4631 & ~n9993 ;
  assign n9995 = ~n9992 & n9994 ;
  assign n9998 = n2795 ^ n1495 ^ 1'b0 ;
  assign n9996 = x32 & ~n6197 ;
  assign n9997 = n9996 ^ n1289 ^ 1'b0 ;
  assign n9999 = n9998 ^ n9997 ^ 1'b0 ;
  assign n10000 = n5497 ^ n3202 ^ 1'b0 ;
  assign n10001 = ~n2246 & n10000 ;
  assign n10002 = n2284 & n9989 ;
  assign n10003 = n867 | n1021 ;
  assign n10004 = n10003 ^ n7093 ^ n547 ;
  assign n10005 = ~n6438 & n10004 ;
  assign n10006 = ~n3061 & n10005 ;
  assign n10012 = n7653 ^ n3164 ^ 1'b0 ;
  assign n10007 = n2617 ^ n640 ^ 1'b0 ;
  assign n10008 = n1677 & n10007 ;
  assign n10009 = n10008 ^ n263 ^ 1'b0 ;
  assign n10010 = n7769 | n10009 ;
  assign n10011 = n10010 ^ n2578 ^ n858 ;
  assign n10013 = n10012 ^ n10011 ^ n4410 ;
  assign n10014 = n5325 ^ n4626 ^ 1'b0 ;
  assign n10015 = n2425 & ~n3051 ;
  assign n10016 = ( x10 & ~n10014 ) | ( x10 & n10015 ) | ( ~n10014 & n10015 ) ;
  assign n10017 = n2548 & ~n6899 ;
  assign n10018 = n1856 | n4981 ;
  assign n10019 = n1645 & ~n10018 ;
  assign n10020 = n7607 ^ n5647 ^ n331 ;
  assign n10021 = n1991 & n10020 ;
  assign n10022 = n10021 ^ n7064 ^ 1'b0 ;
  assign n10023 = n10019 | n10022 ;
  assign n10024 = n387 | n3626 ;
  assign n10025 = n10024 ^ n732 ^ 1'b0 ;
  assign n10026 = n2605 & n10025 ;
  assign n10027 = ( n2365 & n4806 ) | ( n2365 & n8844 ) | ( n4806 & n8844 ) ;
  assign n10028 = ~n2656 & n5151 ;
  assign n10029 = n8213 ^ n6856 ^ 1'b0 ;
  assign n10030 = n8519 & n10029 ;
  assign n10031 = n1760 & n8899 ;
  assign n10032 = ~n443 & n10031 ;
  assign n10033 = n10032 ^ n4076 ^ 1'b0 ;
  assign n10034 = n317 | n3709 ;
  assign n10035 = n10034 ^ n7186 ^ 1'b0 ;
  assign n10036 = n10035 ^ n2246 ^ 1'b0 ;
  assign n10037 = n8837 ^ n2628 ^ 1'b0 ;
  assign n10038 = n6617 | n10037 ;
  assign n10039 = n10038 ^ n6822 ^ 1'b0 ;
  assign n10040 = ~n10036 & n10039 ;
  assign n10041 = n2336 & ~n2783 ;
  assign n10042 = n10041 ^ n787 ^ 1'b0 ;
  assign n10043 = ~n974 & n10042 ;
  assign n10049 = n3401 ^ n2428 ^ 1'b0 ;
  assign n10048 = n1932 & n5412 ;
  assign n10050 = n10049 ^ n10048 ^ 1'b0 ;
  assign n10044 = n2856 ^ n1173 ^ 1'b0 ;
  assign n10045 = n8037 | n10044 ;
  assign n10046 = ~n5366 & n7363 ;
  assign n10047 = n10045 | n10046 ;
  assign n10051 = n10050 ^ n10047 ^ 1'b0 ;
  assign n10052 = n6264 ^ n3821 ^ n1982 ;
  assign n10053 = n9456 ^ n5656 ^ 1'b0 ;
  assign n10054 = ( n6597 & n10052 ) | ( n6597 & n10053 ) | ( n10052 & n10053 ) ;
  assign n10055 = ~n6384 & n10054 ;
  assign n10056 = n5343 ^ x250 ^ 1'b0 ;
  assign n10057 = ( x188 & n10055 ) | ( x188 & n10056 ) | ( n10055 & n10056 ) ;
  assign n10058 = n2347 | n2516 ;
  assign n10059 = n1920 & ~n10058 ;
  assign n10063 = ( ~x11 & n6338 ) | ( ~x11 & n6429 ) | ( n6338 & n6429 ) ;
  assign n10060 = n2009 & ~n4132 ;
  assign n10061 = n10060 ^ n314 ^ 1'b0 ;
  assign n10062 = ~n2653 & n10061 ;
  assign n10064 = n10063 ^ n10062 ^ 1'b0 ;
  assign n10065 = n3642 & ~n4760 ;
  assign n10066 = n10065 ^ n3310 ^ 1'b0 ;
  assign n10069 = x175 & n2621 ;
  assign n10070 = n10069 ^ n2838 ^ 1'b0 ;
  assign n10067 = n2823 ^ n1323 ^ 1'b0 ;
  assign n10068 = n6851 | n10067 ;
  assign n10071 = n10070 ^ n10068 ^ 1'b0 ;
  assign n10072 = n10071 ^ n9280 ^ 1'b0 ;
  assign n10075 = n3959 ^ n3501 ^ 1'b0 ;
  assign n10076 = n6967 | n10075 ;
  assign n10077 = n10076 ^ n8190 ^ n620 ;
  assign n10073 = n2844 ^ n1712 ^ 1'b0 ;
  assign n10074 = ~n6373 & n10073 ;
  assign n10078 = n10077 ^ n10074 ^ 1'b0 ;
  assign n10079 = n5038 ^ n686 ^ 1'b0 ;
  assign n10080 = n928 | n8515 ;
  assign n10081 = n2269 | n10080 ;
  assign n10082 = n10081 ^ n3430 ^ 1'b0 ;
  assign n10083 = n9906 & n10082 ;
  assign n10084 = n10083 ^ n8251 ^ 1'b0 ;
  assign n10085 = ~n10079 & n10084 ;
  assign n10086 = n4145 ^ n2974 ^ 1'b0 ;
  assign n10087 = n2093 | n10086 ;
  assign n10088 = n10087 ^ n2797 ^ n1574 ;
  assign n10090 = n1515 | n8437 ;
  assign n10089 = n1766 & n2598 ;
  assign n10091 = n10090 ^ n10089 ^ n4707 ;
  assign n10093 = n1202 | n5513 ;
  assign n10092 = ~n4057 & n8828 ;
  assign n10094 = n10093 ^ n10092 ^ n6653 ;
  assign n10095 = n7261 ^ x90 ^ 1'b0 ;
  assign n10096 = n1225 | n9666 ;
  assign n10097 = n906 | n10096 ;
  assign n10101 = n1666 & ~n2563 ;
  assign n10102 = ~n3551 & n10101 ;
  assign n10103 = n6338 & n10102 ;
  assign n10098 = n2210 & ~n8220 ;
  assign n10099 = n10098 ^ n10008 ^ 1'b0 ;
  assign n10100 = n2890 & ~n10099 ;
  assign n10104 = n10103 ^ n10100 ^ 1'b0 ;
  assign n10105 = n10104 ^ n883 ^ 1'b0 ;
  assign n10106 = n10097 & n10105 ;
  assign n10107 = ~n381 & n3915 ;
  assign n10108 = n6064 & n10107 ;
  assign n10109 = n3301 & n4114 ;
  assign n10110 = n6268 | n10109 ;
  assign n10111 = n10110 ^ n4001 ^ 1'b0 ;
  assign n10112 = n10111 ^ n4868 ^ 1'b0 ;
  assign n10119 = n1979 ^ x109 ^ 1'b0 ;
  assign n10120 = n1393 & ~n10119 ;
  assign n10121 = n2714 ^ n1324 ^ 1'b0 ;
  assign n10122 = n10120 & n10121 ;
  assign n10116 = n967 & n4999 ;
  assign n10117 = ~n2831 & n4896 ;
  assign n10118 = n10116 & n10117 ;
  assign n10113 = n3063 ^ n1310 ^ 1'b0 ;
  assign n10114 = n360 & ~n10113 ;
  assign n10115 = n10114 ^ n1601 ^ 1'b0 ;
  assign n10123 = n10122 ^ n10118 ^ n10115 ;
  assign n10125 = n6424 ^ n906 ^ 1'b0 ;
  assign n10126 = n10125 ^ n5549 ^ 1'b0 ;
  assign n10124 = n2441 | n7331 ;
  assign n10127 = n10126 ^ n10124 ^ 1'b0 ;
  assign n10128 = n8884 ^ n1489 ^ n1166 ;
  assign n10129 = ( ~n2372 & n5124 ) | ( ~n2372 & n10128 ) | ( n5124 & n10128 ) ;
  assign n10130 = ~x107 & n4338 ;
  assign n10131 = n6723 & n10130 ;
  assign n10132 = n10129 & ~n10131 ;
  assign n10133 = ~n599 & n7443 ;
  assign n10134 = n3413 ^ n3362 ^ n1579 ;
  assign n10135 = ~n1203 & n10134 ;
  assign n10136 = n4921 ^ n4907 ^ 1'b0 ;
  assign n10137 = n1547 & n10136 ;
  assign n10138 = n5396 & ~n10137 ;
  assign n10139 = n6337 & ~n9684 ;
  assign n10140 = n10139 ^ n4766 ^ 1'b0 ;
  assign n10141 = n2122 ^ n1930 ^ 1'b0 ;
  assign n10142 = n10141 ^ n5095 ^ 1'b0 ;
  assign n10143 = n10052 ^ n6346 ^ 1'b0 ;
  assign n10144 = ( n1260 & n9652 ) | ( n1260 & n10143 ) | ( n9652 & n10143 ) ;
  assign n10145 = n10144 ^ n6375 ^ 1'b0 ;
  assign n10146 = n3102 ^ n2108 ^ n548 ;
  assign n10147 = n10146 ^ n2738 ^ 1'b0 ;
  assign n10148 = n1809 & n10147 ;
  assign n10149 = n9791 ^ n3834 ^ x167 ;
  assign n10150 = n10149 ^ n5923 ^ 1'b0 ;
  assign n10151 = ( x170 & n1701 ) | ( x170 & ~n7824 ) | ( n1701 & ~n7824 ) ;
  assign n10153 = ( ~x99 & n4709 ) | ( ~x99 & n4766 ) | ( n4709 & n4766 ) ;
  assign n10152 = x181 & ~n2739 ;
  assign n10154 = n10153 ^ n10152 ^ 1'b0 ;
  assign n10155 = n706 | n10154 ;
  assign n10156 = n10151 & ~n10155 ;
  assign n10157 = n10156 ^ n3550 ^ 1'b0 ;
  assign n10158 = n10150 & ~n10157 ;
  assign n10159 = ~n1085 & n1212 ;
  assign n10160 = n1678 & ~n10159 ;
  assign n10161 = n552 | n4184 ;
  assign n10162 = n10160 | n10161 ;
  assign n10163 = n1437 | n3904 ;
  assign n10164 = n10163 ^ n4970 ^ 1'b0 ;
  assign n10165 = n10162 & n10164 ;
  assign n10166 = n10165 ^ n2455 ^ 1'b0 ;
  assign n10167 = x209 & ~n10166 ;
  assign n10168 = ( n2294 & n4867 ) | ( n2294 & n9237 ) | ( n4867 & n9237 ) ;
  assign n10169 = ( n7847 & ~n9416 ) | ( n7847 & n10168 ) | ( ~n9416 & n10168 ) ;
  assign n10170 = n984 | n1360 ;
  assign n10171 = ~n5164 & n6770 ;
  assign n10172 = ~n2577 & n10171 ;
  assign n10173 = n7384 ^ n6068 ^ 1'b0 ;
  assign n10174 = ( n1026 & n4881 ) | ( n1026 & n10173 ) | ( n4881 & n10173 ) ;
  assign n10175 = ~n1907 & n2640 ;
  assign n10176 = x123 | n541 ;
  assign n10177 = n10176 ^ n1156 ^ 1'b0 ;
  assign n10178 = ~n1401 & n10177 ;
  assign n10179 = n5006 & ~n6692 ;
  assign n10180 = x197 & n981 ;
  assign n10181 = n10180 ^ n500 ^ 1'b0 ;
  assign n10182 = n10181 ^ n1296 ^ 1'b0 ;
  assign n10183 = n1296 & n2653 ;
  assign n10184 = n10183 ^ n3434 ^ 1'b0 ;
  assign n10185 = ~n10182 & n10184 ;
  assign n10189 = n3893 & n6601 ;
  assign n10186 = n2935 ^ n1196 ^ 1'b0 ;
  assign n10187 = ( n2160 & n9411 ) | ( n2160 & n10186 ) | ( n9411 & n10186 ) ;
  assign n10188 = n10187 ^ n5750 ^ 1'b0 ;
  assign n10190 = n10189 ^ n10188 ^ 1'b0 ;
  assign n10191 = n7492 | n10190 ;
  assign n10192 = n1766 & ~n10191 ;
  assign n10193 = n5538 ^ n1494 ^ 1'b0 ;
  assign n10194 = n1499 & n5726 ;
  assign n10195 = n1210 | n7267 ;
  assign n10196 = n10194 | n10195 ;
  assign n10197 = x253 & n1046 ;
  assign n10198 = n10197 ^ n7748 ^ 1'b0 ;
  assign n10199 = n9146 & n10198 ;
  assign n10200 = n1355 & n10199 ;
  assign n10203 = ~n875 & n1396 ;
  assign n10202 = x161 & ~n552 ;
  assign n10204 = n10203 ^ n10202 ^ 1'b0 ;
  assign n10205 = n10204 ^ n4047 ^ 1'b0 ;
  assign n10201 = ( n474 & n2402 ) | ( n474 & n4455 ) | ( n2402 & n4455 ) ;
  assign n10206 = n10205 ^ n10201 ^ 1'b0 ;
  assign n10207 = n10206 ^ n8643 ^ 1'b0 ;
  assign n10208 = ~n5963 & n7385 ;
  assign n10209 = ~n6290 & n10208 ;
  assign n10210 = n5922 & ~n7333 ;
  assign n10211 = ~n7386 & n10210 ;
  assign n10212 = n10211 ^ n4010 ^ 1'b0 ;
  assign n10213 = ~n3640 & n4417 ;
  assign n10214 = n8682 ^ n8356 ^ 1'b0 ;
  assign n10215 = n9336 ^ n1265 ^ n1007 ;
  assign n10216 = ( n520 & n706 ) | ( n520 & n875 ) | ( n706 & n875 ) ;
  assign n10217 = n10216 ^ n6460 ^ n4469 ;
  assign n10226 = x137 & ~n5522 ;
  assign n10221 = n395 & ~n583 ;
  assign n10220 = n459 & n981 ;
  assign n10222 = n10221 ^ n10220 ^ 1'b0 ;
  assign n10223 = ( n2797 & ~n3419 ) | ( n2797 & n10222 ) | ( ~n3419 & n10222 ) ;
  assign n10224 = n10223 ^ n3265 ^ 1'b0 ;
  assign n10225 = n9722 & n10224 ;
  assign n10227 = n10226 ^ n10225 ^ 1'b0 ;
  assign n10218 = n5398 ^ n4184 ^ 1'b0 ;
  assign n10219 = n4196 & n10218 ;
  assign n10228 = n10227 ^ n10219 ^ 1'b0 ;
  assign n10229 = n3501 ^ n1760 ^ 1'b0 ;
  assign n10230 = ~n5468 & n10229 ;
  assign n10231 = ~n7743 & n10230 ;
  assign n10232 = ~n2810 & n9636 ;
  assign n10233 = n4243 ^ n1272 ^ 1'b0 ;
  assign n10234 = n10233 ^ n9273 ^ 1'b0 ;
  assign n10235 = n1943 | n9630 ;
  assign n10236 = n10235 ^ n737 ^ 1'b0 ;
  assign n10237 = ~n2749 & n6623 ;
  assign n10238 = n10237 ^ n5098 ^ 1'b0 ;
  assign n10239 = n10236 & n10238 ;
  assign n10240 = n5113 ^ n1270 ^ 1'b0 ;
  assign n10241 = n2630 | n10240 ;
  assign n10242 = ~n4074 & n9559 ;
  assign n10243 = ~n10120 & n10242 ;
  assign n10244 = ~n2276 & n8936 ;
  assign n10245 = n9856 ^ n9575 ^ n1980 ;
  assign n10246 = x194 | n8905 ;
  assign n10247 = ~n4527 & n10246 ;
  assign n10248 = ~n988 & n10247 ;
  assign n10249 = ~n495 & n5807 ;
  assign n10250 = n7454 & n10249 ;
  assign n10251 = n269 & ~n10250 ;
  assign n10252 = n10251 ^ n4284 ^ 1'b0 ;
  assign n10253 = n3144 & ~n3615 ;
  assign n10254 = n8225 | n9137 ;
  assign n10255 = n10254 ^ n9374 ^ 1'b0 ;
  assign n10257 = n6833 ^ n2905 ^ 1'b0 ;
  assign n10256 = n3239 & ~n3518 ;
  assign n10258 = n10257 ^ n10256 ^ 1'b0 ;
  assign n10259 = n428 | n620 ;
  assign n10260 = n6166 | n10259 ;
  assign n10261 = n9271 & n10260 ;
  assign n10262 = n1096 & ~n3859 ;
  assign n10263 = n1297 & n2970 ;
  assign n10264 = n10263 ^ n3688 ^ 1'b0 ;
  assign n10265 = ~n5396 & n10264 ;
  assign n10268 = n369 | n3624 ;
  assign n10266 = n2131 | n4066 ;
  assign n10267 = n8332 | n10266 ;
  assign n10269 = n10268 ^ n10267 ^ 1'b0 ;
  assign n10270 = n10265 | n10269 ;
  assign n10272 = n8625 ^ n7386 ^ n686 ;
  assign n10271 = n565 & ~n7116 ;
  assign n10273 = n10272 ^ n10271 ^ n5124 ;
  assign n10274 = n2799 ^ n1296 ^ 1'b0 ;
  assign n10275 = n9561 ^ n5858 ^ n496 ;
  assign n10276 = n10275 ^ n5131 ^ 1'b0 ;
  assign n10277 = ( n8618 & n10274 ) | ( n8618 & ~n10276 ) | ( n10274 & ~n10276 ) ;
  assign n10278 = ~n1681 & n6674 ;
  assign n10279 = n1278 & n10278 ;
  assign n10280 = n4148 ^ n3911 ^ 1'b0 ;
  assign n10281 = n482 | n10280 ;
  assign n10282 = n10281 ^ x160 ^ 1'b0 ;
  assign n10283 = n3729 ^ x87 ^ 1'b0 ;
  assign n10284 = ~n1191 & n10283 ;
  assign n10285 = n5684 & ~n10284 ;
  assign n10286 = n6351 ^ n1486 ^ 1'b0 ;
  assign n10287 = n6540 | n10286 ;
  assign n10288 = n10287 ^ n6136 ^ 1'b0 ;
  assign n10289 = n2699 & ~n4260 ;
  assign n10290 = n9049 & n10289 ;
  assign n10291 = ~x33 & n10290 ;
  assign n10292 = n5624 ^ n4220 ^ 1'b0 ;
  assign n10293 = n6741 | n10292 ;
  assign n10294 = n6847 ^ n2502 ^ 1'b0 ;
  assign n10295 = n3413 | n10294 ;
  assign n10296 = ( n886 & n3307 ) | ( n886 & ~n8134 ) | ( n3307 & ~n8134 ) ;
  assign n10297 = n10295 | n10296 ;
  assign n10298 = n8393 & ~n10297 ;
  assign n10300 = n347 & ~n1180 ;
  assign n10301 = ~n1312 & n10300 ;
  assign n10302 = n10301 ^ n3850 ^ 1'b0 ;
  assign n10299 = n1369 & ~n7977 ;
  assign n10303 = n10302 ^ n10299 ^ 1'b0 ;
  assign n10304 = n4812 ^ n1571 ^ 1'b0 ;
  assign n10305 = n5684 & ~n10304 ;
  assign n10306 = n10305 ^ n1000 ^ 1'b0 ;
  assign n10311 = ( x130 & n2430 ) | ( x130 & ~n4124 ) | ( n2430 & ~n4124 ) ;
  assign n10312 = ~n9076 & n10311 ;
  assign n10313 = n10312 ^ n9777 ^ n2246 ;
  assign n10314 = n7599 & ~n10313 ;
  assign n10307 = n1021 & n7653 ;
  assign n10308 = n10307 ^ n883 ^ 1'b0 ;
  assign n10309 = n10308 ^ n5417 ^ n3577 ;
  assign n10310 = ~n3003 & n10309 ;
  assign n10315 = n10314 ^ n10310 ^ n2359 ;
  assign n10316 = n1605 ^ x21 ^ 1'b0 ;
  assign n10317 = n10316 ^ n4556 ^ n896 ;
  assign n10318 = n2271 & n4124 ;
  assign n10319 = n10318 ^ n3158 ^ 1'b0 ;
  assign n10320 = n10319 ^ n5146 ^ 1'b0 ;
  assign n10321 = n10317 & n10320 ;
  assign n10322 = ( ~n518 & n6940 ) | ( ~n518 & n7901 ) | ( n6940 & n7901 ) ;
  assign n10323 = n5391 & ~n5468 ;
  assign n10325 = n1470 ^ n1129 ^ 1'b0 ;
  assign n10324 = n6604 ^ n5193 ^ 1'b0 ;
  assign n10326 = n10325 ^ n10324 ^ n2371 ;
  assign n10327 = n10326 ^ n4396 ^ 1'b0 ;
  assign n10328 = n7945 ^ n1886 ^ 1'b0 ;
  assign n10329 = n449 & ~n10328 ;
  assign n10330 = n10329 ^ n9866 ^ 1'b0 ;
  assign n10331 = n8001 | n10330 ;
  assign n10332 = n3357 ^ n2239 ^ x103 ;
  assign n10333 = ( n8121 & n9881 ) | ( n8121 & ~n10332 ) | ( n9881 & ~n10332 ) ;
  assign n10336 = n8245 ^ n2002 ^ 1'b0 ;
  assign n10337 = x54 & n10336 ;
  assign n10338 = ~n1348 & n10337 ;
  assign n10334 = n4355 ^ n4267 ^ 1'b0 ;
  assign n10335 = ~n4925 & n10334 ;
  assign n10339 = n10338 ^ n10335 ^ 1'b0 ;
  assign n10340 = n4355 ^ x39 ^ 1'b0 ;
  assign n10341 = ~n10339 & n10340 ;
  assign n10342 = n2075 & ~n3958 ;
  assign n10343 = n10342 ^ n4402 ^ 1'b0 ;
  assign n10344 = n8598 ^ n8051 ^ n2285 ;
  assign n10345 = n2082 ^ n1798 ^ 1'b0 ;
  assign n10346 = n2936 & n10345 ;
  assign n10347 = ~n8515 & n10346 ;
  assign n10348 = ~n5805 & n10347 ;
  assign n10349 = ( n1060 & n6912 ) | ( n1060 & ~n10348 ) | ( n6912 & ~n10348 ) ;
  assign n10350 = n3251 ^ n2052 ^ 1'b0 ;
  assign n10351 = n2140 & n10350 ;
  assign n10352 = ~n4087 & n10351 ;
  assign n10353 = n2414 | n10352 ;
  assign n10354 = n10353 ^ n8957 ^ 1'b0 ;
  assign n10355 = n1313 & ~n8413 ;
  assign n10356 = n10355 ^ n9034 ^ 1'b0 ;
  assign n10357 = n6625 ^ n5006 ^ 1'b0 ;
  assign n10358 = n3296 | n3312 ;
  assign n10359 = n10357 & ~n10358 ;
  assign n10360 = n358 | n6089 ;
  assign n10361 = n10360 ^ n6625 ^ 1'b0 ;
  assign n10364 = n1500 ^ n607 ^ 1'b0 ;
  assign n10362 = ~n1512 & n7570 ;
  assign n10363 = n1520 & n10362 ;
  assign n10365 = n10364 ^ n10363 ^ 1'b0 ;
  assign n10366 = n8605 ^ n1865 ^ 1'b0 ;
  assign n10367 = n6018 ^ n4361 ^ 1'b0 ;
  assign n10368 = n903 & n10367 ;
  assign n10369 = n10368 ^ n372 ^ 1'b0 ;
  assign n10370 = n1629 | n3920 ;
  assign n10371 = n10370 ^ n10204 ^ 1'b0 ;
  assign n10372 = n10371 ^ n1023 ^ 1'b0 ;
  assign n10373 = ~n5013 & n10372 ;
  assign n10374 = n10369 & n10373 ;
  assign n10375 = n3596 | n7799 ;
  assign n10378 = n4462 | n7984 ;
  assign n10376 = ~n5188 & n5513 ;
  assign n10377 = n10376 ^ n9640 ^ 1'b0 ;
  assign n10379 = n10378 ^ n10377 ^ 1'b0 ;
  assign n10380 = ( n762 & ~n3391 ) | ( n762 & n6768 ) | ( ~n3391 & n6768 ) ;
  assign n10381 = n1620 & n5653 ;
  assign n10382 = ~n3776 & n10381 ;
  assign n10383 = n1730 & n10382 ;
  assign n10384 = n3982 & ~n5361 ;
  assign n10385 = n10384 ^ n5489 ^ 1'b0 ;
  assign n10386 = n10385 ^ n4077 ^ 1'b0 ;
  assign n10387 = n9752 ^ n8316 ^ n2332 ;
  assign n10388 = n8236 ^ n7911 ^ 1'b0 ;
  assign n10389 = n8634 & n10388 ;
  assign n10390 = n913 & n8255 ;
  assign n10391 = ~n1091 & n10390 ;
  assign n10392 = n2455 | n10204 ;
  assign n10393 = n10392 ^ n6736 ^ 1'b0 ;
  assign n10394 = n7519 ^ n1107 ^ 1'b0 ;
  assign n10395 = ~n4364 & n10379 ;
  assign n10396 = ( n4616 & ~n6423 ) | ( n4616 & n7847 ) | ( ~n6423 & n7847 ) ;
  assign n10397 = n806 & n3365 ;
  assign n10398 = n7064 | n9067 ;
  assign n10399 = ~n963 & n7358 ;
  assign n10400 = n10399 ^ n4342 ^ 1'b0 ;
  assign n10401 = n2378 ^ x186 ^ 1'b0 ;
  assign n10402 = n10400 & ~n10401 ;
  assign n10403 = n5499 | n6713 ;
  assign n10404 = n10403 ^ n7605 ^ 1'b0 ;
  assign n10405 = n2642 ^ n2282 ^ n1785 ;
  assign n10406 = n10405 ^ n2046 ^ x174 ;
  assign n10407 = n10406 ^ n3062 ^ 1'b0 ;
  assign n10408 = n7897 & n10407 ;
  assign n10410 = ~n1372 & n6223 ;
  assign n10411 = ~n7093 & n10410 ;
  assign n10412 = ~n8081 & n10411 ;
  assign n10409 = n2668 & n4722 ;
  assign n10413 = n10412 ^ n10409 ^ 1'b0 ;
  assign n10414 = n4284 & ~n9804 ;
  assign n10415 = n5918 & ~n8605 ;
  assign n10416 = ~n7735 & n10415 ;
  assign n10417 = n2634 ^ n1369 ^ 1'b0 ;
  assign n10418 = n7781 ^ n677 ^ 1'b0 ;
  assign n10419 = x73 & ~n10418 ;
  assign n10420 = n8728 | n10419 ;
  assign n10421 = n5529 ^ n5465 ^ 1'b0 ;
  assign n10422 = n10421 ^ n950 ^ 1'b0 ;
  assign n10424 = n4405 ^ n4046 ^ 1'b0 ;
  assign n10423 = n7405 ^ n6720 ^ n3693 ;
  assign n10425 = n10424 ^ n10423 ^ n3254 ;
  assign n10428 = n2913 & ~n8113 ;
  assign n10426 = n2231 ^ n379 ^ 1'b0 ;
  assign n10427 = ~n1106 & n10426 ;
  assign n10429 = n10428 ^ n10427 ^ 1'b0 ;
  assign n10430 = n6096 ^ n2638 ^ 1'b0 ;
  assign n10431 = ~n10429 & n10430 ;
  assign n10432 = n4284 | n7666 ;
  assign n10433 = n1616 | n3135 ;
  assign n10434 = n10432 | n10433 ;
  assign n10435 = n1295 & ~n9805 ;
  assign n10436 = ~n10434 & n10435 ;
  assign n10437 = x145 & ~n7973 ;
  assign n10438 = n3680 & n10437 ;
  assign n10439 = n706 & ~n10438 ;
  assign n10440 = n5701 ^ n1773 ^ 1'b0 ;
  assign n10450 = ~n861 & n1376 ;
  assign n10451 = n8841 & n10233 ;
  assign n10452 = ( n8768 & n10450 ) | ( n8768 & ~n10451 ) | ( n10450 & ~n10451 ) ;
  assign n10446 = n3147 ^ x158 ^ 1'b0 ;
  assign n10447 = n333 | n10446 ;
  assign n10441 = n4286 ^ n2327 ^ n530 ;
  assign n10442 = n3693 & n10441 ;
  assign n10443 = n10442 ^ n2501 ^ 1'b0 ;
  assign n10444 = n10443 ^ n2610 ^ 1'b0 ;
  assign n10445 = n10444 ^ n7567 ^ 1'b0 ;
  assign n10448 = n10447 ^ n10445 ^ n8685 ;
  assign n10449 = n897 & n10448 ;
  assign n10453 = n10452 ^ n10449 ^ 1'b0 ;
  assign n10454 = n283 | n4606 ;
  assign n10455 = ( n1200 & n5864 ) | ( n1200 & ~n10454 ) | ( n5864 & ~n10454 ) ;
  assign n10456 = ~n6189 & n9151 ;
  assign n10457 = ~n10455 & n10456 ;
  assign n10458 = n2587 ^ n1929 ^ 1'b0 ;
  assign n10459 = n2673 | n10458 ;
  assign n10460 = n8893 & n10459 ;
  assign n10461 = n2483 | n10460 ;
  assign n10462 = n10461 ^ n6286 ^ 1'b0 ;
  assign n10463 = n2685 & ~n5744 ;
  assign n10464 = n1353 & n10463 ;
  assign n10465 = n6709 & ~n10464 ;
  assign n10466 = n6501 & n10465 ;
  assign n10467 = n9054 ^ n5677 ^ 1'b0 ;
  assign n10468 = n3504 & n10467 ;
  assign n10469 = n4290 ^ x21 ^ 1'b0 ;
  assign n10470 = n8728 | n10469 ;
  assign n10471 = n3084 & ~n10470 ;
  assign n10472 = n6507 | n10471 ;
  assign n10473 = n3088 & n10472 ;
  assign n10474 = n8417 ^ n6793 ^ n1567 ;
  assign n10475 = n1838 & n5729 ;
  assign n10476 = n2077 | n4514 ;
  assign n10477 = n10475 | n10476 ;
  assign n10478 = n10477 ^ n1312 ^ 1'b0 ;
  assign n10479 = n4303 | n10478 ;
  assign n10480 = n5418 ^ n4718 ^ n974 ;
  assign n10481 = n7880 & ~n10480 ;
  assign n10482 = n1433 & n9735 ;
  assign n10483 = ~n10481 & n10482 ;
  assign n10484 = n1296 & n2925 ;
  assign n10485 = n2178 & n6213 ;
  assign n10486 = ~n10484 & n10485 ;
  assign n10487 = n10436 ^ n3690 ^ 1'b0 ;
  assign n10488 = n4412 | n10487 ;
  assign n10489 = n841 & ~n8057 ;
  assign n10490 = n10489 ^ n1601 ^ 1'b0 ;
  assign n10491 = n6302 & ~n10490 ;
  assign n10492 = n1232 & ~n5705 ;
  assign n10493 = ~n2973 & n4398 ;
  assign n10494 = ~n2384 & n10493 ;
  assign n10495 = ( ~n3558 & n5391 ) | ( ~n3558 & n7577 ) | ( n5391 & n7577 ) ;
  assign n10496 = ~n3630 & n10495 ;
  assign n10497 = ~n6975 & n10496 ;
  assign n10498 = n4230 & ~n8968 ;
  assign n10499 = n4644 & n10498 ;
  assign n10500 = n2201 & ~n2549 ;
  assign n10501 = ~n2654 & n10500 ;
  assign n10502 = ( n5227 & n9472 ) | ( n5227 & ~n10501 ) | ( n9472 & ~n10501 ) ;
  assign n10503 = n3253 ^ n579 ^ 1'b0 ;
  assign n10504 = n7002 ^ n2763 ^ 1'b0 ;
  assign n10505 = n10503 & ~n10504 ;
  assign n10506 = ~n3430 & n10505 ;
  assign n10507 = n10205 ^ n3800 ^ 1'b0 ;
  assign n10508 = ~n10506 & n10507 ;
  assign n10509 = n1460 & n6528 ;
  assign n10510 = n911 ^ n783 ^ 1'b0 ;
  assign n10511 = n5135 ^ n4712 ^ 1'b0 ;
  assign n10512 = n10510 & ~n10511 ;
  assign n10513 = n10512 ^ x133 ^ 1'b0 ;
  assign n10514 = n10509 | n10513 ;
  assign n10515 = n2186 | n7110 ;
  assign n10516 = n9527 ^ n8862 ^ 1'b0 ;
  assign n10517 = ( ~n2014 & n5703 ) | ( ~n2014 & n6461 ) | ( n5703 & n6461 ) ;
  assign n10518 = n10517 ^ n1252 ^ x158 ;
  assign n10519 = n1708 | n3628 ;
  assign n10520 = n5497 & ~n10519 ;
  assign n10521 = n4547 & n10520 ;
  assign n10524 = n3239 & n6223 ;
  assign n10525 = ~n1504 & n10524 ;
  assign n10523 = n2995 | n3680 ;
  assign n10526 = n10525 ^ n10523 ^ 1'b0 ;
  assign n10522 = n10284 ^ n8866 ^ n7830 ;
  assign n10527 = n10526 ^ n10522 ^ n2488 ;
  assign n10528 = n5430 & n10527 ;
  assign n10529 = n10528 ^ n5373 ^ 1'b0 ;
  assign n10530 = n3920 ^ n1486 ^ 1'b0 ;
  assign n10531 = n845 & n3023 ;
  assign n10532 = n10531 ^ n2924 ^ 1'b0 ;
  assign n10533 = n10530 | n10532 ;
  assign n10534 = n5034 ^ n1450 ^ x113 ;
  assign n10535 = n3278 & n3620 ;
  assign n10536 = n3881 ^ n505 ^ 1'b0 ;
  assign n10537 = n10535 & ~n10536 ;
  assign n10538 = n4588 & ~n10537 ;
  assign n10539 = n10538 ^ n2337 ^ 1'b0 ;
  assign n10540 = n10534 | n10539 ;
  assign n10541 = x209 | n10540 ;
  assign n10542 = ~n4096 & n10541 ;
  assign n10543 = ~n3647 & n10542 ;
  assign n10544 = n6494 | n10543 ;
  assign n10545 = n10533 & ~n10544 ;
  assign n10546 = n4351 | n9011 ;
  assign n10547 = n10546 ^ n6985 ^ 1'b0 ;
  assign n10548 = n903 ^ n436 ^ 1'b0 ;
  assign n10549 = n5145 & n9962 ;
  assign n10550 = n10549 ^ n1298 ^ 1'b0 ;
  assign n10551 = n6825 ^ n3620 ^ 1'b0 ;
  assign n10552 = ~n817 & n10551 ;
  assign n10553 = ( x58 & ~n1340 ) | ( x58 & n7844 ) | ( ~n1340 & n7844 ) ;
  assign n10554 = n5289 | n8768 ;
  assign n10555 = n7354 | n10554 ;
  assign n10556 = n1124 & ~n3584 ;
  assign n10557 = n4105 & n10556 ;
  assign n10558 = n5770 | n10557 ;
  assign n10559 = n1052 | n7782 ;
  assign n10560 = n6098 | n10559 ;
  assign n10561 = n4855 & ~n5984 ;
  assign n10562 = ~n8755 & n10561 ;
  assign n10563 = x115 & ~n5885 ;
  assign n10564 = n5276 & n10563 ;
  assign n10565 = n10564 ^ n2741 ^ 1'b0 ;
  assign n10566 = n7200 & ~n10565 ;
  assign n10567 = ( x153 & ~n3525 ) | ( x153 & n10566 ) | ( ~n3525 & n10566 ) ;
  assign n10568 = n7026 & ~n10567 ;
  assign n10569 = n1963 | n3383 ;
  assign n10570 = ~n9840 & n10569 ;
  assign n10571 = ~n7677 & n10570 ;
  assign n10572 = ( ~n2161 & n5304 ) | ( ~n2161 & n10571 ) | ( n5304 & n10571 ) ;
  assign n10573 = n6302 & n10572 ;
  assign n10574 = n1543 ^ n429 ^ 1'b0 ;
  assign n10575 = ( x231 & n399 ) | ( x231 & ~n10574 ) | ( n399 & ~n10574 ) ;
  assign n10576 = n6919 ^ n4110 ^ 1'b0 ;
  assign n10577 = ( n3394 & n3998 ) | ( n3394 & n10576 ) | ( n3998 & n10576 ) ;
  assign n10578 = n10577 ^ n9990 ^ 1'b0 ;
  assign n10579 = n1707 ^ n357 ^ 1'b0 ;
  assign n10580 = ~n3413 & n10579 ;
  assign n10581 = n10083 ^ n978 ^ 1'b0 ;
  assign n10582 = n3834 | n10581 ;
  assign n10583 = n5687 ^ x17 ^ 1'b0 ;
  assign n10584 = n3741 | n10583 ;
  assign n10587 = n328 | n4034 ;
  assign n10588 = n10587 ^ n9857 ^ 1'b0 ;
  assign n10585 = n6303 ^ n4394 ^ n4114 ;
  assign n10586 = n2686 & n10585 ;
  assign n10589 = n10588 ^ n10586 ^ n6129 ;
  assign n10590 = n3376 ^ n793 ^ n711 ;
  assign n10591 = n6734 ^ n1058 ^ 1'b0 ;
  assign n10592 = n10590 & n10591 ;
  assign n10593 = n9939 ^ n9498 ^ 1'b0 ;
  assign n10594 = n3376 ^ x81 ^ 1'b0 ;
  assign n10595 = ( n2394 & n6807 ) | ( n2394 & ~n10594 ) | ( n6807 & ~n10594 ) ;
  assign n10599 = ~n1951 & n3185 ;
  assign n10600 = n1313 & n10599 ;
  assign n10601 = ~n3904 & n10600 ;
  assign n10602 = n10601 ^ n1776 ^ 1'b0 ;
  assign n10596 = n4246 & n4422 ;
  assign n10597 = ~n277 & n5882 ;
  assign n10598 = ~n10596 & n10597 ;
  assign n10603 = n10602 ^ n10598 ^ n1720 ;
  assign n10605 = n6079 ^ n5071 ^ 1'b0 ;
  assign n10604 = n6228 & n8130 ;
  assign n10606 = n10605 ^ n10604 ^ 1'b0 ;
  assign n10607 = n1612 & n4797 ;
  assign n10608 = ~n2272 & n4109 ;
  assign n10609 = ~n3506 & n10608 ;
  assign n10610 = n2993 & n3382 ;
  assign n10611 = n7514 & n10610 ;
  assign n10612 = n1443 | n7943 ;
  assign n10614 = x67 & ~n6476 ;
  assign n10613 = n3737 & n6609 ;
  assign n10615 = n10614 ^ n10613 ^ 1'b0 ;
  assign n10616 = n713 | n10615 ;
  assign n10617 = n10612 | n10616 ;
  assign n10618 = n785 | n5464 ;
  assign n10619 = ~n6741 & n10618 ;
  assign n10620 = ~n1214 & n10619 ;
  assign n10621 = n275 & n8551 ;
  assign n10622 = n2921 | n9840 ;
  assign n10623 = n1622 | n10622 ;
  assign n10624 = n6874 ^ n2947 ^ 1'b0 ;
  assign n10625 = n7408 ^ n7101 ^ 1'b0 ;
  assign n10626 = ~n10624 & n10625 ;
  assign n10627 = n5840 | n10626 ;
  assign n10628 = n1052 & ~n2739 ;
  assign n10629 = n7675 ^ n1073 ^ 1'b0 ;
  assign n10630 = ~n7406 & n10158 ;
  assign n10631 = n8807 & n10630 ;
  assign n10632 = ( n10628 & n10629 ) | ( n10628 & ~n10631 ) | ( n10629 & ~n10631 ) ;
  assign n10633 = n2955 & ~n3897 ;
  assign n10634 = n6209 & ~n10633 ;
  assign n10635 = ~n2998 & n10160 ;
  assign n10636 = n10635 ^ n7322 ^ 1'b0 ;
  assign n10637 = n7833 & ~n10636 ;
  assign n10638 = x172 & ~n4021 ;
  assign n10639 = n10638 ^ n4812 ^ 1'b0 ;
  assign n10640 = x54 | n2623 ;
  assign n10641 = ~n5224 & n10640 ;
  assign n10642 = ~x7 & n10641 ;
  assign n10643 = n10639 | n10642 ;
  assign n10644 = ~n7182 & n10643 ;
  assign n10645 = n5719 ^ n591 ^ 1'b0 ;
  assign n10646 = ~n9965 & n10645 ;
  assign n10647 = n3742 & n5339 ;
  assign n10648 = x187 & ~n514 ;
  assign n10649 = ( n3872 & n9793 ) | ( n3872 & n10648 ) | ( n9793 & n10648 ) ;
  assign n10650 = n2584 ^ n1206 ^ 1'b0 ;
  assign n10651 = n4426 | n10650 ;
  assign n10656 = x8 & ~n2858 ;
  assign n10657 = n1254 & n10656 ;
  assign n10652 = n2333 & ~n5347 ;
  assign n10653 = n10652 ^ n650 ^ 1'b0 ;
  assign n10654 = n7404 ^ x167 ^ 1'b0 ;
  assign n10655 = n10653 & ~n10654 ;
  assign n10658 = n10657 ^ n10655 ^ 1'b0 ;
  assign n10659 = n6589 & ~n10658 ;
  assign n10660 = ~n5760 & n10659 ;
  assign n10661 = n2851 ^ n2197 ^ 1'b0 ;
  assign n10662 = n6473 & ~n10661 ;
  assign n10663 = n10662 ^ n9268 ^ 1'b0 ;
  assign n10664 = n9968 | n10663 ;
  assign n10665 = x90 & ~n7271 ;
  assign n10666 = ~n1916 & n10665 ;
  assign n10667 = n10666 ^ n559 ^ 1'b0 ;
  assign n10668 = n5266 | n7780 ;
  assign n10669 = n10668 ^ n9710 ^ 1'b0 ;
  assign n10672 = n1225 & ~n1878 ;
  assign n10673 = n10672 ^ n4469 ^ 1'b0 ;
  assign n10670 = n5963 | n9329 ;
  assign n10671 = n3279 | n10670 ;
  assign n10674 = n10673 ^ n10671 ^ 1'b0 ;
  assign n10675 = n860 & n10674 ;
  assign n10676 = ~n3891 & n10675 ;
  assign n10677 = ~n7130 & n10676 ;
  assign n10678 = ~n2858 & n6904 ;
  assign n10679 = n2575 & n10678 ;
  assign n10680 = n7229 ^ n5547 ^ n4246 ;
  assign n10682 = ( ~n545 & n3374 ) | ( ~n545 & n7105 ) | ( n3374 & n7105 ) ;
  assign n10681 = n1715 | n3538 ;
  assign n10683 = n10682 ^ n10681 ^ 1'b0 ;
  assign n10684 = n9056 ^ n6722 ^ n2345 ;
  assign n10685 = ~n6049 & n8247 ;
  assign n10686 = n269 | n2214 ;
  assign n10691 = n3523 ^ n1059 ^ n725 ;
  assign n10687 = ~n399 & n1091 ;
  assign n10688 = n2286 & n10687 ;
  assign n10689 = n10688 ^ n4494 ^ n3273 ;
  assign n10690 = n10689 ^ n7645 ^ 1'b0 ;
  assign n10692 = n10691 ^ n10690 ^ 1'b0 ;
  assign n10693 = n6517 ^ n5348 ^ 1'b0 ;
  assign n10694 = ~n4655 & n10693 ;
  assign n10695 = ~n8039 & n10694 ;
  assign n10696 = n10695 ^ n7664 ^ 1'b0 ;
  assign n10697 = ( n671 & n4344 ) | ( n671 & n6265 ) | ( n4344 & n6265 ) ;
  assign n10698 = n4765 & ~n5411 ;
  assign n10699 = n7995 & n10698 ;
  assign n10700 = n2467 | n10699 ;
  assign n10701 = n2902 | n10700 ;
  assign n10702 = n9018 & n10701 ;
  assign n10703 = n732 & ~n1228 ;
  assign n10704 = n1228 & n10703 ;
  assign n10705 = n2518 & ~n10704 ;
  assign n10706 = ( x103 & ~n5356 ) | ( x103 & n10705 ) | ( ~n5356 & n10705 ) ;
  assign n10707 = n9778 ^ n1809 ^ 1'b0 ;
  assign n10708 = x81 & n1782 ;
  assign n10709 = n10708 ^ n1764 ^ 1'b0 ;
  assign n10710 = n10707 | n10709 ;
  assign n10711 = n10710 ^ n6874 ^ 1'b0 ;
  assign n10712 = ~n840 & n1323 ;
  assign n10713 = n3632 & ~n6177 ;
  assign n10714 = n10712 & n10713 ;
  assign n10715 = n1346 & n10714 ;
  assign n10716 = n2223 ^ n947 ^ 1'b0 ;
  assign n10717 = n10716 ^ n3019 ^ 1'b0 ;
  assign n10718 = n8813 & ~n10717 ;
  assign n10720 = ~n3658 & n6141 ;
  assign n10719 = n2955 | n7457 ;
  assign n10721 = n10720 ^ n10719 ^ 1'b0 ;
  assign n10722 = ~n2156 & n6774 ;
  assign n10723 = n7087 & n10722 ;
  assign n10724 = n10723 ^ n8765 ^ n1595 ;
  assign n10725 = n5588 ^ n1063 ^ 1'b0 ;
  assign n10726 = n10724 & n10725 ;
  assign n10727 = ~n8447 & n10726 ;
  assign n10728 = ( ~n4445 & n4891 ) | ( ~n4445 & n10727 ) | ( n4891 & n10727 ) ;
  assign n10729 = n903 & ~n1064 ;
  assign n10730 = ~n903 & n10729 ;
  assign n10731 = n5067 | n10730 ;
  assign n10732 = n10728 & ~n10731 ;
  assign n10733 = n3035 & ~n9451 ;
  assign n10735 = ~n4743 & n5166 ;
  assign n10736 = n2719 & n10735 ;
  assign n10734 = ~n1515 & n5354 ;
  assign n10737 = n10736 ^ n10734 ^ 1'b0 ;
  assign n10740 = n1881 ^ n1009 ^ 1'b0 ;
  assign n10741 = ~n1772 & n10740 ;
  assign n10738 = n9857 ^ n3779 ^ x141 ;
  assign n10739 = n535 | n10738 ;
  assign n10742 = n10741 ^ n10739 ^ 1'b0 ;
  assign n10743 = n6312 & ~n10742 ;
  assign n10744 = ( ~n918 & n1764 ) | ( ~n918 & n3664 ) | ( n1764 & n3664 ) ;
  assign n10745 = n8823 ^ n5487 ^ n2118 ;
  assign n10746 = n9350 ^ n7962 ^ n1746 ;
  assign n10747 = n6074 ^ n2277 ^ 1'b0 ;
  assign n10748 = ( n1086 & n2393 ) | ( n1086 & n3335 ) | ( n2393 & n3335 ) ;
  assign n10749 = ~n5778 & n10748 ;
  assign n10750 = n10749 ^ n5776 ^ 1'b0 ;
  assign n10752 = ~n1943 & n2743 ;
  assign n10751 = n9230 ^ n3958 ^ x129 ;
  assign n10753 = n10752 ^ n10751 ^ n2448 ;
  assign n10754 = n2376 | n10037 ;
  assign n10755 = n10754 ^ n8255 ^ 1'b0 ;
  assign n10756 = n1298 & ~n1526 ;
  assign n10757 = n10756 ^ n1437 ^ 1'b0 ;
  assign n10758 = n10757 ^ x165 ^ 1'b0 ;
  assign n10759 = n9339 | n10758 ;
  assign n10760 = n6798 ^ n4718 ^ 1'b0 ;
  assign n10761 = ~n2089 & n10760 ;
  assign n10762 = ~n1024 & n2842 ;
  assign n10763 = n10762 ^ n1832 ^ 1'b0 ;
  assign n10764 = n3374 ^ n1667 ^ 1'b0 ;
  assign n10765 = n1946 | n5540 ;
  assign n10766 = n5489 & ~n10765 ;
  assign n10767 = n10766 ^ n6937 ^ n3895 ;
  assign n10768 = n3879 & ~n10767 ;
  assign n10769 = n2995 ^ n1620 ^ 1'b0 ;
  assign n10770 = n2267 | n10769 ;
  assign n10771 = n10770 ^ n5884 ^ 1'b0 ;
  assign n10772 = n10771 ^ n8947 ^ 1'b0 ;
  assign n10773 = ~n10768 & n10772 ;
  assign n10774 = ~n10764 & n10773 ;
  assign n10775 = n6085 ^ n6018 ^ 1'b0 ;
  assign n10776 = n10775 ^ n4172 ^ 1'b0 ;
  assign n10777 = x202 | n2146 ;
  assign n10778 = n10777 ^ n772 ^ 1'b0 ;
  assign n10779 = ~n341 & n579 ;
  assign n10780 = n7210 ^ n749 ^ 1'b0 ;
  assign n10781 = ( n7748 & n7847 ) | ( n7748 & ~n10780 ) | ( n7847 & ~n10780 ) ;
  assign n10782 = ( ~n5775 & n8477 ) | ( ~n5775 & n10781 ) | ( n8477 & n10781 ) ;
  assign n10783 = ~n10779 & n10782 ;
  assign n10784 = n1190 & ~n1464 ;
  assign n10785 = n10784 ^ n3283 ^ 1'b0 ;
  assign n10786 = n5875 | n10785 ;
  assign n10787 = n7313 & n9207 ;
  assign n10791 = n9259 ^ n1378 ^ 1'b0 ;
  assign n10788 = n1558 ^ n719 ^ 1'b0 ;
  assign n10789 = n3831 & n7312 ;
  assign n10790 = ~n10788 & n10789 ;
  assign n10792 = n10791 ^ n10790 ^ 1'b0 ;
  assign n10793 = n1919 & ~n10792 ;
  assign n10801 = n4286 ^ n4196 ^ 1'b0 ;
  assign n10802 = n7316 ^ n397 ^ 1'b0 ;
  assign n10803 = n10801 | n10802 ;
  assign n10804 = ~n4056 & n10803 ;
  assign n10794 = ( n995 & n1455 ) | ( n995 & n2552 ) | ( n1455 & n2552 ) ;
  assign n10795 = n2131 ^ n1271 ^ 1'b0 ;
  assign n10796 = n10794 & n10795 ;
  assign n10797 = ~n3343 & n10796 ;
  assign n10798 = n10797 ^ n5731 ^ 1'b0 ;
  assign n10799 = n9403 ^ n9255 ^ 1'b0 ;
  assign n10800 = n10798 & n10799 ;
  assign n10805 = n10804 ^ n10800 ^ 1'b0 ;
  assign n10806 = n605 | n10805 ;
  assign n10807 = ~n2955 & n9394 ;
  assign n10808 = n10807 ^ n1278 ^ 1'b0 ;
  assign n10809 = n9090 ^ x248 ^ 1'b0 ;
  assign n10810 = n1063 | n10809 ;
  assign n10811 = n10810 ^ n4552 ^ 1'b0 ;
  assign n10812 = n3245 | n10811 ;
  assign n10813 = n873 | n6117 ;
  assign n10814 = n10813 ^ n8662 ^ 1'b0 ;
  assign n10815 = ~n5295 & n10814 ;
  assign n10816 = ( n725 & n2814 ) | ( n725 & ~n5484 ) | ( n2814 & ~n5484 ) ;
  assign n10817 = n7474 ^ n1563 ^ 1'b0 ;
  assign n10818 = n4898 & ~n10817 ;
  assign n10819 = n10818 ^ n2797 ^ 1'b0 ;
  assign n10820 = n10816 & n10819 ;
  assign n10824 = ( x115 & n1767 ) | ( x115 & ~n6394 ) | ( n1767 & ~n6394 ) ;
  assign n10825 = ( n319 & n4552 ) | ( n319 & ~n10824 ) | ( n4552 & ~n10824 ) ;
  assign n10822 = n762 & n3111 ;
  assign n10823 = n5134 & n10822 ;
  assign n10826 = n10825 ^ n10823 ^ 1'b0 ;
  assign n10821 = n5684 & ~n10203 ;
  assign n10827 = n10826 ^ n10821 ^ 1'b0 ;
  assign n10828 = n4828 ^ n543 ^ 1'b0 ;
  assign n10832 = n6922 ^ n2648 ^ 1'b0 ;
  assign n10829 = n4732 ^ n4560 ^ n3152 ;
  assign n10830 = ( n778 & n6811 ) | ( n778 & n10829 ) | ( n6811 & n10829 ) ;
  assign n10831 = n9844 & n10830 ;
  assign n10833 = n10832 ^ n10831 ^ 1'b0 ;
  assign n10834 = n1324 ^ n478 ^ 1'b0 ;
  assign n10835 = n3096 & ~n10834 ;
  assign n10836 = n4232 ^ n2173 ^ 1'b0 ;
  assign n10837 = n3477 & ~n10836 ;
  assign n10838 = n10837 ^ n2479 ^ 1'b0 ;
  assign n10839 = n10835 & n10838 ;
  assign n10840 = ( n4848 & n5471 ) | ( n4848 & ~n8771 ) | ( n5471 & ~n8771 ) ;
  assign n10841 = n5061 | n10840 ;
  assign n10842 = n10841 ^ n1862 ^ 1'b0 ;
  assign n10843 = n4839 & n7930 ;
  assign n10844 = n7928 & n10843 ;
  assign n10845 = n9813 ^ n1170 ^ 1'b0 ;
  assign n10846 = n6842 ^ n863 ^ 1'b0 ;
  assign n10847 = n5929 & n7336 ;
  assign n10848 = ~n1546 & n10847 ;
  assign n10849 = n1223 & ~n5694 ;
  assign n10850 = ~n3545 & n10849 ;
  assign n10851 = n2259 ^ n488 ^ 1'b0 ;
  assign n10852 = n2523 ^ x235 ^ 1'b0 ;
  assign n10853 = n10851 | n10852 ;
  assign n10854 = n5193 | n7161 ;
  assign n10855 = n10854 ^ n8603 ^ 1'b0 ;
  assign n10856 = n5129 ^ n1046 ^ 1'b0 ;
  assign n10858 = n5217 ^ n4104 ^ 1'b0 ;
  assign n10859 = x90 & ~n10858 ;
  assign n10860 = n6887 & n10859 ;
  assign n10861 = n10860 ^ n7752 ^ 1'b0 ;
  assign n10862 = n2775 & ~n10861 ;
  assign n10857 = n1033 & n3545 ;
  assign n10863 = n10862 ^ n10857 ^ 1'b0 ;
  assign n10864 = n6232 & n10863 ;
  assign n10865 = n8345 ^ n7954 ^ 1'b0 ;
  assign n10867 = ( ~n1437 & n2213 ) | ( ~n1437 & n3908 ) | ( n2213 & n3908 ) ;
  assign n10866 = n909 & ~n4205 ;
  assign n10868 = n10867 ^ n10866 ^ 1'b0 ;
  assign n10869 = n8915 ^ n3904 ^ 1'b0 ;
  assign n10870 = n10868 | n10869 ;
  assign n10871 = ~n681 & n5675 ;
  assign n10872 = n10871 ^ n8001 ^ 1'b0 ;
  assign n10873 = n10872 ^ n907 ^ 1'b0 ;
  assign n10874 = n4985 & n10421 ;
  assign n10885 = ( n1467 & n1832 ) | ( n1467 & ~n4892 ) | ( n1832 & ~n4892 ) ;
  assign n10884 = ( n606 & n5577 ) | ( n606 & n6234 ) | ( n5577 & n6234 ) ;
  assign n10886 = n10885 ^ n10884 ^ n7014 ;
  assign n10887 = n631 ^ n522 ^ 1'b0 ;
  assign n10888 = ~n1712 & n10887 ;
  assign n10889 = n2766 & n10888 ;
  assign n10890 = ~n10886 & n10889 ;
  assign n10878 = n3376 & ~n4613 ;
  assign n10879 = ~n7362 & n10878 ;
  assign n10880 = n6574 & ~n10879 ;
  assign n10877 = n5022 | n7917 ;
  assign n10875 = n2900 & n4520 ;
  assign n10876 = ~n3195 & n10875 ;
  assign n10881 = n10880 ^ n10877 ^ n10876 ;
  assign n10882 = n6432 ^ n5596 ^ 1'b0 ;
  assign n10883 = ~n10881 & n10882 ;
  assign n10891 = n10890 ^ n10883 ^ 1'b0 ;
  assign n10892 = n4638 ^ n2445 ^ 1'b0 ;
  assign n10893 = n6871 | n10892 ;
  assign n10894 = n10893 ^ n9342 ^ 1'b0 ;
  assign n10895 = n9026 & n10894 ;
  assign n10896 = n5895 & ~n8623 ;
  assign n10897 = n3170 | n6349 ;
  assign n10898 = n4191 & n10897 ;
  assign n10899 = n4450 ^ n3566 ^ 1'b0 ;
  assign n10900 = n4249 & n10899 ;
  assign n10901 = n1930 & ~n10815 ;
  assign n10907 = n1874 & n6035 ;
  assign n10902 = n1979 | n7237 ;
  assign n10903 = ~n2015 & n2481 ;
  assign n10904 = n10903 ^ n1989 ^ 1'b0 ;
  assign n10905 = ~n7400 & n10904 ;
  assign n10906 = ( n4638 & n10902 ) | ( n4638 & ~n10905 ) | ( n10902 & ~n10905 ) ;
  assign n10908 = n10907 ^ n10906 ^ n5922 ;
  assign n10909 = ~n5162 & n8696 ;
  assign n10910 = x18 & n3716 ;
  assign n10911 = ~n3447 & n10910 ;
  assign n10912 = n985 | n3490 ;
  assign n10913 = n10911 & ~n10912 ;
  assign n10914 = n10913 ^ n1760 ^ 1'b0 ;
  assign n10915 = n3306 | n10914 ;
  assign n10916 = n4326 & ~n10915 ;
  assign n10917 = n10916 ^ n4999 ^ 1'b0 ;
  assign n10919 = n5967 ^ n5338 ^ n3088 ;
  assign n10918 = n269 & n10448 ;
  assign n10920 = n10919 ^ n10918 ^ 1'b0 ;
  assign n10921 = n8691 ^ n547 ^ 1'b0 ;
  assign n10927 = ~n480 & n9614 ;
  assign n10928 = n3798 & n10927 ;
  assign n10923 = n4410 | n4549 ;
  assign n10922 = n463 | n4573 ;
  assign n10924 = n10923 ^ n10922 ^ 1'b0 ;
  assign n10925 = n5352 | n10924 ;
  assign n10926 = n5621 & ~n10925 ;
  assign n10929 = n10928 ^ n10926 ^ 1'b0 ;
  assign n10930 = n9577 & ~n10929 ;
  assign n10931 = n2380 ^ n1186 ^ 1'b0 ;
  assign n10932 = ~n648 & n10931 ;
  assign n10933 = n6762 ^ n4816 ^ 1'b0 ;
  assign n10934 = n10932 & ~n10933 ;
  assign n10935 = n5565 ^ n3958 ^ n2814 ;
  assign n10936 = ~n6588 & n10935 ;
  assign n10937 = n10936 ^ n4558 ^ 1'b0 ;
  assign n10938 = ~n755 & n10937 ;
  assign n10939 = n4616 & n10938 ;
  assign n10940 = n369 & n1681 ;
  assign n10941 = ( n795 & ~n2134 ) | ( n795 & n3239 ) | ( ~n2134 & n3239 ) ;
  assign n10942 = n4016 & n10941 ;
  assign n10943 = ~n10940 & n10942 ;
  assign n10944 = x36 | n10566 ;
  assign n10945 = n9307 ^ n4394 ^ 1'b0 ;
  assign n10946 = ~n2989 & n10945 ;
  assign n10947 = n1669 ^ n1261 ^ 1'b0 ;
  assign n10948 = ( n3686 & n7460 ) | ( n3686 & ~n10947 ) | ( n7460 & ~n10947 ) ;
  assign n10949 = n10948 ^ x65 ^ 1'b0 ;
  assign n10950 = n8672 ^ n7946 ^ n7149 ;
  assign n10951 = n5785 & n10950 ;
  assign n10956 = n1622 & n2393 ;
  assign n10952 = n1879 & ~n2266 ;
  assign n10953 = n10480 & n10952 ;
  assign n10954 = n10953 ^ n10438 ^ 1'b0 ;
  assign n10955 = n1486 & n10954 ;
  assign n10957 = n10956 ^ n10955 ^ 1'b0 ;
  assign n10958 = n9920 | n10957 ;
  assign n10959 = n9072 ^ n2896 ^ 1'b0 ;
  assign n10960 = n5102 | n10959 ;
  assign n10961 = n5330 ^ n5084 ^ 1'b0 ;
  assign n10962 = n10550 & ~n10961 ;
  assign n10963 = n4545 | n5621 ;
  assign n10964 = ~n5172 & n10963 ;
  assign n10965 = n10964 ^ n7645 ^ 1'b0 ;
  assign n10966 = n10965 ^ n7101 ^ n3790 ;
  assign n10967 = n2457 ^ n1998 ^ 1'b0 ;
  assign n10968 = n10966 | n10967 ;
  assign n10969 = n1327 & n2278 ;
  assign n10970 = n10969 ^ n7149 ^ 1'b0 ;
  assign n10971 = n9740 ^ n6605 ^ 1'b0 ;
  assign n10972 = n3434 | n4429 ;
  assign n10973 = n10972 ^ n3088 ^ 1'b0 ;
  assign n10974 = n7381 ^ n4099 ^ 1'b0 ;
  assign n10975 = ~n10973 & n10974 ;
  assign n10976 = n2255 | n10454 ;
  assign n10977 = n538 ^ x161 ^ 1'b0 ;
  assign n10978 = n10977 ^ n8913 ^ 1'b0 ;
  assign n10979 = ~n7836 & n8645 ;
  assign n10981 = n5825 ^ n3843 ^ 1'b0 ;
  assign n10982 = n6366 & n10981 ;
  assign n10980 = n877 | n9011 ;
  assign n10983 = n10982 ^ n10980 ^ 1'b0 ;
  assign n10984 = n7074 & ~n10983 ;
  assign n10985 = n10320 ^ n1270 ^ 1'b0 ;
  assign n10990 = ( n3088 & n3419 ) | ( n3088 & n4331 ) | ( n3419 & n4331 ) ;
  assign n10988 = n4616 ^ n2879 ^ 1'b0 ;
  assign n10989 = ~n3029 & n10988 ;
  assign n10986 = n7105 ^ n6494 ^ 1'b0 ;
  assign n10987 = n4232 | n10986 ;
  assign n10991 = n10990 ^ n10989 ^ n10987 ;
  assign n10992 = n2778 ^ n1102 ^ n1027 ;
  assign n10993 = n673 & ~n1254 ;
  assign n10994 = n10993 ^ n535 ^ 1'b0 ;
  assign n10995 = ( n3877 & n10992 ) | ( n3877 & n10994 ) | ( n10992 & n10994 ) ;
  assign n10996 = n4389 ^ n2230 ^ n570 ;
  assign n10997 = n10996 ^ n7027 ^ n2785 ;
  assign n10998 = n10997 ^ n942 ^ 1'b0 ;
  assign n10999 = n1055 | n10998 ;
  assign n11000 = n7581 & n9068 ;
  assign n11002 = ~n787 & n4370 ;
  assign n11001 = x65 & ~n3144 ;
  assign n11003 = n11002 ^ n11001 ^ 1'b0 ;
  assign n11004 = x77 & n11003 ;
  assign n11005 = n11000 & n11004 ;
  assign n11006 = n11005 ^ n4271 ^ 1'b0 ;
  assign n11007 = n869 & n8603 ;
  assign n11008 = n11007 ^ n4696 ^ 1'b0 ;
  assign n11009 = n592 & ~n1129 ;
  assign n11010 = n11009 ^ n8007 ^ 1'b0 ;
  assign n11011 = n6573 ^ n1817 ^ 1'b0 ;
  assign n11012 = n4750 & n9961 ;
  assign n11013 = n3785 | n5961 ;
  assign n11014 = n10818 ^ n8516 ^ n1733 ;
  assign n11015 = ( ~n335 & n6555 ) | ( ~n335 & n11014 ) | ( n6555 & n11014 ) ;
  assign n11016 = n10029 ^ n560 ^ 1'b0 ;
  assign n11017 = n9026 & n11016 ;
  assign n11019 = n5772 ^ n2743 ^ 1'b0 ;
  assign n11020 = n3732 ^ n2818 ^ 1'b0 ;
  assign n11021 = ~n11019 & n11020 ;
  assign n11018 = n1289 & n8560 ;
  assign n11022 = n11021 ^ n11018 ^ 1'b0 ;
  assign n11023 = n894 & n5610 ;
  assign n11024 = n2226 & n11023 ;
  assign n11025 = n7682 ^ n4397 ^ 1'b0 ;
  assign n11026 = ~n11024 & n11025 ;
  assign n11027 = x43 & ~n4264 ;
  assign n11028 = n374 & n11027 ;
  assign n11029 = n447 & n474 ;
  assign n11030 = n11029 ^ x144 ^ 1'b0 ;
  assign n11031 = n2598 ^ x209 ^ 1'b0 ;
  assign n11032 = ( n5884 & n11030 ) | ( n5884 & ~n11031 ) | ( n11030 & ~n11031 ) ;
  assign n11033 = ( n1142 & n4520 ) | ( n1142 & n9241 ) | ( n4520 & n9241 ) ;
  assign n11034 = n11033 ^ n3692 ^ 1'b0 ;
  assign n11035 = n6926 & ~n11034 ;
  assign n11036 = ~n9542 & n11035 ;
  assign n11037 = n11036 ^ n3267 ^ 1'b0 ;
  assign n11041 = x84 & n1200 ;
  assign n11039 = ~n2713 & n5968 ;
  assign n11038 = n1144 | n5732 ;
  assign n11040 = n11039 ^ n11038 ^ 1'b0 ;
  assign n11042 = n11041 ^ n11040 ^ 1'b0 ;
  assign n11043 = n2824 ^ n1093 ^ 1'b0 ;
  assign n11044 = n2684 & n8867 ;
  assign n11045 = n11043 & n11044 ;
  assign n11046 = n5025 | n5108 ;
  assign n11047 = n3269 & ~n11046 ;
  assign n11050 = n674 ^ x241 ^ 1'b0 ;
  assign n11051 = n10445 ^ n690 ^ 1'b0 ;
  assign n11052 = n11050 | n11051 ;
  assign n11048 = n7316 ^ n3786 ^ 1'b0 ;
  assign n11049 = n3554 & ~n11048 ;
  assign n11053 = n11052 ^ n11049 ^ 1'b0 ;
  assign n11054 = n8659 ^ n2346 ^ 1'b0 ;
  assign n11055 = n2243 & n11054 ;
  assign n11056 = n11055 ^ n1831 ^ n1295 ;
  assign n11057 = n11056 ^ n6044 ^ 1'b0 ;
  assign n11058 = n9152 & ~n11057 ;
  assign n11059 = n9150 ^ n2158 ^ 1'b0 ;
  assign n11060 = n9044 & n11059 ;
  assign n11061 = ( n880 & n7508 ) | ( n880 & ~n11060 ) | ( n7508 & ~n11060 ) ;
  assign n11062 = n7443 ^ n3342 ^ 1'b0 ;
  assign n11063 = n11062 ^ n7314 ^ n3088 ;
  assign n11064 = n7035 ^ n3420 ^ 1'b0 ;
  assign n11065 = n11064 ^ n6969 ^ 1'b0 ;
  assign n11066 = n3427 ^ n1495 ^ 1'b0 ;
  assign n11067 = n8038 ^ n5917 ^ 1'b0 ;
  assign n11068 = ~n2653 & n11067 ;
  assign n11069 = n11068 ^ n10701 ^ 1'b0 ;
  assign n11070 = ~n4052 & n10724 ;
  assign n11071 = ~n3318 & n5215 ;
  assign n11072 = n11071 ^ n10203 ^ 1'b0 ;
  assign n11073 = ~n607 & n4063 ;
  assign n11074 = ~n11072 & n11073 ;
  assign n11075 = n8343 | n8887 ;
  assign n11076 = n455 | n11075 ;
  assign n11077 = ( n1823 & n6509 ) | ( n1823 & ~n6655 ) | ( n6509 & ~n6655 ) ;
  assign n11078 = n10633 ^ n2317 ^ 1'b0 ;
  assign n11079 = n411 & ~n11078 ;
  assign n11080 = n11079 ^ n7135 ^ 1'b0 ;
  assign n11081 = n11080 ^ n9366 ^ 1'b0 ;
  assign n11082 = ~n10925 & n11081 ;
  assign n11083 = n9769 ^ n3898 ^ n1872 ;
  assign n11084 = ~n3642 & n10854 ;
  assign n11085 = n4884 & n11084 ;
  assign n11086 = n4108 & n10256 ;
  assign n11087 = n2816 & n4565 ;
  assign n11088 = n2361 & n9577 ;
  assign n11089 = n2450 ^ n593 ^ 1'b0 ;
  assign n11090 = n6611 & ~n11089 ;
  assign n11091 = n8564 ^ n2327 ^ n1440 ;
  assign n11092 = ~n821 & n5663 ;
  assign n11093 = n1148 ^ x201 ^ 1'b0 ;
  assign n11094 = n11093 ^ n1813 ^ 1'b0 ;
  assign n11095 = ~n4132 & n11094 ;
  assign n11096 = ~n6472 & n11095 ;
  assign n11097 = n11092 & n11096 ;
  assign n11098 = ~n2395 & n7876 ;
  assign n11099 = n2839 ^ n685 ^ 1'b0 ;
  assign n11100 = ~n11030 & n11099 ;
  assign n11101 = n3163 | n11100 ;
  assign n11102 = n926 | n1254 ;
  assign n11103 = ~n2418 & n11102 ;
  assign n11104 = n3158 & ~n3979 ;
  assign n11105 = n11104 ^ n3516 ^ 1'b0 ;
  assign n11106 = ~n11103 & n11105 ;
  assign n11107 = ~n4962 & n11106 ;
  assign n11108 = n11107 ^ n1201 ^ 1'b0 ;
  assign n11109 = n4812 & ~n6484 ;
  assign n11110 = n2299 & n10114 ;
  assign n11111 = n1957 & n11110 ;
  assign n11112 = n11111 ^ x228 ^ 1'b0 ;
  assign n11113 = n11109 | n11112 ;
  assign n11114 = ~n1358 & n2692 ;
  assign n11115 = n2470 & ~n11114 ;
  assign n11118 = ~n4867 & n8815 ;
  assign n11119 = n11118 ^ n5912 ^ 1'b0 ;
  assign n11116 = x152 & ~n6493 ;
  assign n11117 = ~n6731 & n11116 ;
  assign n11120 = n11119 ^ n11117 ^ 1'b0 ;
  assign n11121 = ~n2178 & n11120 ;
  assign n11122 = n7263 ^ n6400 ^ n6018 ;
  assign n11123 = n974 | n5667 ;
  assign n11124 = n1471 | n6899 ;
  assign n11125 = n8232 | n8476 ;
  assign n11126 = n8071 & n11125 ;
  assign n11127 = ~n11124 & n11126 ;
  assign n11128 = ~n5348 & n9871 ;
  assign n11129 = n8661 & n11128 ;
  assign n11130 = n1928 & n4901 ;
  assign n11131 = ~x159 & n11130 ;
  assign n11132 = n5061 | n11131 ;
  assign n11133 = n11132 ^ n3939 ^ 1'b0 ;
  assign n11134 = n2811 ^ n610 ^ 1'b0 ;
  assign n11135 = n11134 ^ n11070 ^ 1'b0 ;
  assign n11136 = ~n4263 & n11046 ;
  assign n11140 = n10837 ^ n10749 ^ n5395 ;
  assign n11137 = n6777 & n7850 ;
  assign n11138 = ~n8038 & n11137 ;
  assign n11139 = n357 | n11138 ;
  assign n11141 = n11140 ^ n11139 ^ 1'b0 ;
  assign n11142 = n3617 & ~n5832 ;
  assign n11143 = ( x15 & n7063 ) | ( x15 & n11142 ) | ( n7063 & n11142 ) ;
  assign n11144 = n8011 | n11143 ;
  assign n11145 = n4446 ^ n2597 ^ 1'b0 ;
  assign n11146 = n4716 & ~n11145 ;
  assign n11147 = n11144 & ~n11146 ;
  assign n11148 = n5084 & ~n9334 ;
  assign n11149 = n11148 ^ n9520 ^ 1'b0 ;
  assign n11150 = n8002 & n11149 ;
  assign n11151 = ~n9694 & n11150 ;
  assign n11152 = n3032 & n6373 ;
  assign n11153 = ~n3073 & n4885 ;
  assign n11158 = n1121 & ~n3111 ;
  assign n11159 = n4662 & n9731 ;
  assign n11160 = ~n11158 & n11159 ;
  assign n11154 = n4513 ^ n2575 ^ 1'b0 ;
  assign n11155 = n6375 | n11154 ;
  assign n11156 = n11155 ^ n1877 ^ 1'b0 ;
  assign n11157 = ~n2628 & n11156 ;
  assign n11161 = n11160 ^ n11157 ^ n2768 ;
  assign n11162 = x142 & ~n6502 ;
  assign n11163 = ~n3244 & n11162 ;
  assign n11164 = n1232 ^ n998 ^ 1'b0 ;
  assign n11165 = n1951 ^ n1906 ^ 1'b0 ;
  assign n11167 = n9562 ^ n2524 ^ 1'b0 ;
  assign n11166 = n1938 | n6248 ;
  assign n11168 = n11167 ^ n11166 ^ 1'b0 ;
  assign n11169 = n332 & ~n8535 ;
  assign n11170 = n1453 & ~n3723 ;
  assign n11171 = n11170 ^ n6941 ^ 1'b0 ;
  assign n11172 = n3485 & ~n9076 ;
  assign n11173 = n11172 ^ n10884 ^ 1'b0 ;
  assign n11174 = n11173 ^ n6287 ^ 1'b0 ;
  assign n11175 = n3216 & n8933 ;
  assign n11185 = x176 & n6332 ;
  assign n11186 = n11185 ^ n2450 ^ 1'b0 ;
  assign n11180 = n842 & ~n9666 ;
  assign n11181 = n3040 & n11180 ;
  assign n11182 = n9500 & ~n11181 ;
  assign n11183 = n11182 ^ n4428 ^ 1'b0 ;
  assign n11176 = n4927 & ~n9026 ;
  assign n11177 = ~n8148 & n11176 ;
  assign n11178 = ~n5503 & n11177 ;
  assign n11179 = n480 | n11178 ;
  assign n11184 = n11183 ^ n11179 ^ 1'b0 ;
  assign n11187 = n11186 ^ n11184 ^ 1'b0 ;
  assign n11188 = ( n732 & n2234 ) | ( n732 & ~n4473 ) | ( n2234 & ~n4473 ) ;
  assign n11189 = n5219 | n11188 ;
  assign n11190 = n11189 ^ n2692 ^ 1'b0 ;
  assign n11191 = n489 & n3712 ;
  assign n11192 = n11075 ^ n4648 ^ 1'b0 ;
  assign n11193 = n11191 | n11192 ;
  assign n11194 = n11193 ^ n905 ^ 1'b0 ;
  assign n11195 = ~n711 & n6084 ;
  assign n11196 = n11195 ^ n7354 ^ 1'b0 ;
  assign n11197 = n5912 & ~n10628 ;
  assign n11198 = n7690 & n11197 ;
  assign n11199 = n9927 ^ n7344 ^ 1'b0 ;
  assign n11200 = ~n480 & n11199 ;
  assign n11201 = n882 & n3821 ;
  assign n11202 = ( x229 & n2433 ) | ( x229 & n11201 ) | ( n2433 & n11201 ) ;
  assign n11203 = n7020 ^ n5922 ^ 1'b0 ;
  assign n11204 = ( n6708 & ~n10457 ) | ( n6708 & n11203 ) | ( ~n10457 & n11203 ) ;
  assign n11205 = ~n653 & n1701 ;
  assign n11206 = n11205 ^ n1102 ^ 1'b0 ;
  assign n11207 = n5725 | n11206 ;
  assign n11208 = n6597 & ~n11207 ;
  assign n11209 = n1038 ^ x178 ^ 1'b0 ;
  assign n11210 = n2026 | n11209 ;
  assign n11211 = n3451 | n11210 ;
  assign n11212 = n11211 ^ n2253 ^ 1'b0 ;
  assign n11213 = ( ~n869 & n8328 ) | ( ~n869 & n11212 ) | ( n8328 & n11212 ) ;
  assign n11214 = n7010 & ~n10962 ;
  assign n11215 = n11214 ^ n3955 ^ 1'b0 ;
  assign n11216 = ( n4021 & ~n6354 ) | ( n4021 & n6676 ) | ( ~n6354 & n6676 ) ;
  assign n11217 = n6907 ^ n6780 ^ 1'b0 ;
  assign n11218 = n5502 & ~n11217 ;
  assign n11219 = n7654 & n11218 ;
  assign n11220 = n11219 ^ n6736 ^ 1'b0 ;
  assign n11221 = ~n11216 & n11220 ;
  assign n11222 = n5768 ^ n3716 ^ n2430 ;
  assign n11223 = ( n5190 & ~n10268 ) | ( n5190 & n11222 ) | ( ~n10268 & n11222 ) ;
  assign n11224 = n1871 ^ n1214 ^ 1'b0 ;
  assign n11225 = ~n948 & n11224 ;
  assign n11226 = n11225 ^ n9500 ^ n905 ;
  assign n11227 = ~n5070 & n11226 ;
  assign n11228 = ( n7239 & n10312 ) | ( n7239 & ~n11227 ) | ( n10312 & ~n11227 ) ;
  assign n11229 = n2723 & ~n11228 ;
  assign n11230 = n11223 & n11229 ;
  assign n11231 = n11230 ^ n4903 ^ n3806 ;
  assign n11234 = ~n813 & n4065 ;
  assign n11232 = n5449 ^ n2228 ^ 1'b0 ;
  assign n11233 = n2380 & n11232 ;
  assign n11235 = n11234 ^ n11233 ^ 1'b0 ;
  assign n11236 = n10886 ^ n3106 ^ n1233 ;
  assign n11237 = n6401 & n7564 ;
  assign n11238 = n2910 ^ n1597 ^ 1'b0 ;
  assign n11239 = n11237 & ~n11238 ;
  assign n11240 = n273 | n2320 ;
  assign n11241 = n11240 ^ n2169 ^ 1'b0 ;
  assign n11242 = n11241 ^ n3641 ^ 1'b0 ;
  assign n11243 = ~n6667 & n11242 ;
  assign n11244 = n11243 ^ n3924 ^ 1'b0 ;
  assign n11245 = ~n9611 & n11244 ;
  assign n11246 = ~n11239 & n11245 ;
  assign n11248 = n8702 ^ n5892 ^ 1'b0 ;
  assign n11247 = x254 & n7958 ;
  assign n11249 = n11248 ^ n11247 ^ 1'b0 ;
  assign n11250 = n6792 ^ n5051 ^ 1'b0 ;
  assign n11251 = n6405 | n11250 ;
  assign n11252 = n11251 ^ n10306 ^ 1'b0 ;
  assign n11253 = n3392 & n3396 ;
  assign n11254 = ~n3392 & n11253 ;
  assign n11255 = n11254 ^ n5772 ^ 1'b0 ;
  assign n11256 = ~n6553 & n11255 ;
  assign n11260 = x30 & ~n6140 ;
  assign n11261 = n11260 ^ n811 ^ 1'b0 ;
  assign n11262 = n2546 & n11261 ;
  assign n11263 = n298 | n4895 ;
  assign n11264 = n11262 & n11263 ;
  assign n11265 = n11264 ^ x176 ^ 1'b0 ;
  assign n11257 = n478 | n8037 ;
  assign n11258 = n11257 ^ n2471 ^ 1'b0 ;
  assign n11259 = ~n9961 & n11258 ;
  assign n11266 = n11265 ^ n11259 ^ 1'b0 ;
  assign n11267 = n6049 | n10453 ;
  assign n11268 = n10999 ^ n1705 ^ 1'b0 ;
  assign n11269 = ( n567 & ~n645 ) | ( n567 & n8893 ) | ( ~n645 & n8893 ) ;
  assign n11270 = ~n1346 & n9902 ;
  assign n11271 = n6131 & n11270 ;
  assign n11272 = n3557 | n10447 ;
  assign n11273 = ~n4831 & n7307 ;
  assign n11274 = n4446 ^ n363 ^ 1'b0 ;
  assign n11275 = ~n11273 & n11274 ;
  assign n11276 = x91 & n1736 ;
  assign n11277 = n9459 & n11242 ;
  assign n11278 = n11277 ^ n4268 ^ 1'b0 ;
  assign n11279 = n2291 & ~n11278 ;
  assign n11280 = n9531 & n11279 ;
  assign n11281 = ~n4218 & n7371 ;
  assign n11282 = n1382 | n7810 ;
  assign n11283 = n11282 ^ n5643 ^ 1'b0 ;
  assign n11284 = n11281 & ~n11283 ;
  assign n11285 = ~n1510 & n1880 ;
  assign n11286 = ( ~n3958 & n5762 ) | ( ~n3958 & n11285 ) | ( n5762 & n11285 ) ;
  assign n11287 = n4867 ^ n3304 ^ 1'b0 ;
  assign n11288 = ~n6686 & n11287 ;
  assign n11289 = ~n2206 & n11288 ;
  assign n11290 = n4135 | n8098 ;
  assign n11291 = n10102 ^ n6447 ^ n2826 ;
  assign n11292 = n3068 & ~n11291 ;
  assign n11293 = n8126 | n9215 ;
  assign n11294 = n11293 ^ x221 ^ 1'b0 ;
  assign n11295 = n8237 & n11294 ;
  assign n11296 = ~n4583 & n8351 ;
  assign n11297 = n11296 ^ n2212 ^ 1'b0 ;
  assign n11298 = n11297 ^ n8229 ^ n2082 ;
  assign n11299 = n11298 ^ n388 ^ 1'b0 ;
  assign n11300 = n1053 & ~n11299 ;
  assign n11301 = n6887 & n9986 ;
  assign n11302 = n11301 ^ n3555 ^ 1'b0 ;
  assign n11303 = n4626 ^ x239 ^ 1'b0 ;
  assign n11304 = n9038 ^ n3790 ^ 1'b0 ;
  assign n11305 = n6871 ^ n6316 ^ 1'b0 ;
  assign n11306 = n2521 | n11305 ;
  assign n11307 = n4853 ^ n1319 ^ 1'b0 ;
  assign n11308 = n9099 | n11307 ;
  assign n11312 = ( x16 & n456 ) | ( x16 & n2895 ) | ( n456 & n2895 ) ;
  assign n11309 = n5107 | n8543 ;
  assign n11310 = n6363 & ~n11309 ;
  assign n11311 = n5053 & ~n11310 ;
  assign n11313 = n11312 ^ n11311 ^ 1'b0 ;
  assign n11314 = n5575 ^ n3660 ^ 1'b0 ;
  assign n11315 = n4508 | n4984 ;
  assign n11316 = x137 | n11315 ;
  assign n11317 = n11314 & ~n11316 ;
  assign n11318 = n11317 ^ n5264 ^ 1'b0 ;
  assign n11319 = n9157 & n11318 ;
  assign n11320 = n875 | n5155 ;
  assign n11321 = n1739 | n11320 ;
  assign n11322 = ( n3251 & n5100 ) | ( n3251 & n11321 ) | ( n5100 & n11321 ) ;
  assign n11323 = n3126 & ~n11322 ;
  assign n11324 = ~n11319 & n11323 ;
  assign n11325 = x124 & ~n3850 ;
  assign n11326 = n11325 ^ n5380 ^ 1'b0 ;
  assign n11327 = n7455 ^ n6035 ^ 1'b0 ;
  assign n11328 = ~n11326 & n11327 ;
  assign n11329 = n1622 & ~n10842 ;
  assign n11330 = ~n11328 & n11329 ;
  assign n11331 = n3413 & n9952 ;
  assign n11332 = n11331 ^ n6798 ^ 1'b0 ;
  assign n11333 = n681 & n4193 ;
  assign n11334 = n11333 ^ n2649 ^ 1'b0 ;
  assign n11335 = ~n833 & n11334 ;
  assign n11336 = n10160 ^ n2430 ^ 1'b0 ;
  assign n11337 = ~n3318 & n4894 ;
  assign n11338 = n11337 ^ n7188 ^ n7093 ;
  assign n11339 = n3597 ^ n591 ^ 1'b0 ;
  assign n11340 = ~n1663 & n3417 ;
  assign n11341 = ~n10329 & n11340 ;
  assign n11344 = n1547 & n3521 ;
  assign n11345 = n1762 & ~n11344 ;
  assign n11342 = ( n1685 & n1690 ) | ( n1685 & n8458 ) | ( n1690 & n8458 ) ;
  assign n11343 = n3160 | n11342 ;
  assign n11346 = n11345 ^ n11343 ^ 1'b0 ;
  assign n11347 = n2336 ^ n875 ^ 1'b0 ;
  assign n11348 = n4373 | n11347 ;
  assign n11349 = ( n4789 & n8113 ) | ( n4789 & ~n9493 ) | ( n8113 & ~n9493 ) ;
  assign n11350 = ( n2632 & n7796 ) | ( n2632 & n11349 ) | ( n7796 & n11349 ) ;
  assign n11351 = ( n790 & ~n2228 ) | ( n790 & n2979 ) | ( ~n2228 & n2979 ) ;
  assign n11352 = n2232 | n2907 ;
  assign n11353 = n11352 ^ n4338 ^ 1'b0 ;
  assign n11354 = n11353 ^ n6829 ^ 1'b0 ;
  assign n11355 = n1478 & n11354 ;
  assign n11356 = n4209 | n7145 ;
  assign n11357 = n1119 | n11356 ;
  assign n11358 = n7812 & ~n9084 ;
  assign n11359 = ~n11357 & n11358 ;
  assign n11360 = ~n1351 & n3467 ;
  assign n11361 = n5151 ^ n4561 ^ n2380 ;
  assign n11362 = n5232 & n11361 ;
  assign n11363 = n11362 ^ n677 ^ 1'b0 ;
  assign n11364 = n7546 ^ n841 ^ 1'b0 ;
  assign n11365 = ~n11363 & n11364 ;
  assign n11366 = n972 ^ x9 ^ 1'b0 ;
  assign n11367 = n9735 | n11366 ;
  assign n11368 = n877 ^ n798 ^ 1'b0 ;
  assign n11369 = ( n474 & ~n3473 ) | ( n474 & n4417 ) | ( ~n3473 & n4417 ) ;
  assign n11370 = ~n9720 & n11369 ;
  assign n11371 = n3903 ^ n616 ^ 1'b0 ;
  assign n11372 = n5958 & n11371 ;
  assign n11374 = n4001 ^ n1208 ^ n481 ;
  assign n11376 = n304 | n2800 ;
  assign n11375 = n5432 | n7664 ;
  assign n11377 = n11376 ^ n11375 ^ 1'b0 ;
  assign n11378 = n8903 & n11377 ;
  assign n11379 = ~n11374 & n11378 ;
  assign n11373 = n1763 | n10790 ;
  assign n11380 = n11379 ^ n11373 ^ 1'b0 ;
  assign n11381 = n2271 & n2539 ;
  assign n11382 = n11381 ^ n4012 ^ 1'b0 ;
  assign n11383 = n2357 | n11382 ;
  assign n11384 = ~n8899 & n11383 ;
  assign n11385 = ~n8281 & n11384 ;
  assign n11393 = n4189 ^ n2641 ^ n1683 ;
  assign n11389 = n4455 ^ n3832 ^ n3257 ;
  assign n11386 = n3281 & ~n7010 ;
  assign n11387 = n2129 | n4467 ;
  assign n11388 = n11386 | n11387 ;
  assign n11390 = n11389 ^ n11388 ^ 1'b0 ;
  assign n11391 = n9479 | n11390 ;
  assign n11392 = n11282 & ~n11391 ;
  assign n11394 = n11393 ^ n11392 ^ 1'b0 ;
  assign n11398 = ~n3048 & n10948 ;
  assign n11399 = n519 & n3695 ;
  assign n11400 = n11398 & n11399 ;
  assign n11396 = n1777 & ~n2008 ;
  assign n11397 = n7934 | n11396 ;
  assign n11401 = n11400 ^ n11397 ^ 1'b0 ;
  assign n11395 = n3533 & n8066 ;
  assign n11402 = n11401 ^ n11395 ^ 1'b0 ;
  assign n11403 = n1249 & ~n2553 ;
  assign n11404 = n11403 ^ n7858 ^ 1'b0 ;
  assign n11405 = n10106 ^ n5182 ^ n4905 ;
  assign n11406 = n5381 ^ x138 ^ 1'b0 ;
  assign n11407 = n2149 & ~n3251 ;
  assign n11408 = n11407 ^ n1302 ^ 1'b0 ;
  assign n11409 = n11408 ^ n3993 ^ 1'b0 ;
  assign n11410 = n1013 & ~n11409 ;
  assign n11411 = n1369 & n6005 ;
  assign n11412 = n2346 & n11411 ;
  assign n11413 = n616 & n11412 ;
  assign n11414 = n8053 ^ n7719 ^ n5853 ;
  assign n11415 = ( n3893 & ~n10424 ) | ( n3893 & n11414 ) | ( ~n10424 & n11414 ) ;
  assign n11416 = n3376 | n5786 ;
  assign n11417 = ~n9435 & n11416 ;
  assign n11418 = ( ~n395 & n4114 ) | ( ~n395 & n11417 ) | ( n4114 & n11417 ) ;
  assign n11419 = n698 & n11418 ;
  assign n11421 = n936 ^ n557 ^ 1'b0 ;
  assign n11420 = n3806 ^ n3517 ^ 1'b0 ;
  assign n11422 = n11421 ^ n11420 ^ 1'b0 ;
  assign n11427 = x8 | n1304 ;
  assign n11424 = n1701 | n3675 ;
  assign n11425 = n6352 | n11424 ;
  assign n11423 = n2300 & ~n2378 ;
  assign n11426 = n11425 ^ n11423 ^ 1'b0 ;
  assign n11428 = n11427 ^ n11426 ^ 1'b0 ;
  assign n11429 = ~n2194 & n6153 ;
  assign n11430 = n7573 ^ n4296 ^ 1'b0 ;
  assign n11431 = n5825 & n11430 ;
  assign n11435 = ~x74 & n10935 ;
  assign n11432 = n5519 ^ n5090 ^ 1'b0 ;
  assign n11433 = n608 & ~n11432 ;
  assign n11434 = ~n2656 & n11433 ;
  assign n11436 = n11435 ^ n11434 ^ n9295 ;
  assign n11437 = n1440 & n11436 ;
  assign n11438 = ~n11431 & n11437 ;
  assign n11439 = n623 | n7647 ;
  assign n11440 = n11439 ^ n7777 ^ 1'b0 ;
  assign n11441 = n4296 & ~n5431 ;
  assign n11442 = ~n2777 & n11441 ;
  assign n11443 = n2831 | n10915 ;
  assign n11444 = ( n8756 & n11442 ) | ( n8756 & n11443 ) | ( n11442 & n11443 ) ;
  assign n11445 = n7834 & ~n9431 ;
  assign n11446 = n11445 ^ n9710 ^ 1'b0 ;
  assign n11447 = x199 & n818 ;
  assign n11448 = ~n10775 & n11447 ;
  assign n11451 = n1533 | n9561 ;
  assign n11452 = n11451 ^ n3259 ^ 1'b0 ;
  assign n11453 = ( n6440 & n10822 ) | ( n6440 & ~n11452 ) | ( n10822 & ~n11452 ) ;
  assign n11449 = ~x58 & n1919 ;
  assign n11450 = n6777 & n11449 ;
  assign n11454 = n11453 ^ n11450 ^ 1'b0 ;
  assign n11455 = n7867 ^ n3487 ^ 1'b0 ;
  assign n11457 = n895 & ~n1232 ;
  assign n11456 = n672 & n3010 ;
  assign n11458 = n11457 ^ n11456 ^ 1'b0 ;
  assign n11459 = n8673 & ~n11458 ;
  assign n11460 = x243 & ~n2266 ;
  assign n11461 = n11460 ^ n6531 ^ 1'b0 ;
  assign n11462 = n2997 | n11461 ;
  assign n11463 = n2761 | n11462 ;
  assign n11464 = n7405 | n11463 ;
  assign n11465 = n10088 ^ n5396 ^ x230 ;
  assign n11466 = ( n3109 & n3135 ) | ( n3109 & n3448 ) | ( n3135 & n3448 ) ;
  assign n11467 = n11466 ^ n10891 ^ n1466 ;
  assign n11468 = n1727 & n6967 ;
  assign n11469 = ~x251 & n7860 ;
  assign n11470 = n3978 & n11469 ;
  assign n11471 = n5812 & n11470 ;
  assign n11472 = n2638 ^ n2322 ^ 1'b0 ;
  assign n11473 = ~n4749 & n9375 ;
  assign n11474 = ~n11472 & n11473 ;
  assign n11475 = n11474 ^ n3325 ^ 1'b0 ;
  assign n11476 = n11475 ^ n10863 ^ 1'b0 ;
  assign n11477 = n3352 & ~n11476 ;
  assign n11478 = n11367 ^ n1308 ^ 1'b0 ;
  assign n11479 = n10464 ^ n7146 ^ 1'b0 ;
  assign n11480 = ~n7953 & n9697 ;
  assign n11481 = n11479 & ~n11480 ;
  assign n11482 = n11481 ^ n6461 ^ 1'b0 ;
  assign n11483 = ( n1381 & ~n6686 ) | ( n1381 & n6910 ) | ( ~n6686 & n6910 ) ;
  assign n11484 = ~n1777 & n6001 ;
  assign n11485 = ( x76 & ~n2359 ) | ( x76 & n8908 ) | ( ~n2359 & n8908 ) ;
  assign n11486 = ~n7339 & n8533 ;
  assign n11487 = n11485 | n11486 ;
  assign n11488 = n11487 ^ n5514 ^ 1'b0 ;
  assign n11489 = n8690 ^ n4232 ^ 1'b0 ;
  assign n11490 = n11489 ^ n7046 ^ n745 ;
  assign n11492 = n1353 | n3740 ;
  assign n11493 = n4833 | n11492 ;
  assign n11491 = n7073 & n7836 ;
  assign n11494 = n11493 ^ n11491 ^ 1'b0 ;
  assign n11495 = n11494 ^ n7599 ^ 1'b0 ;
  assign n11496 = n8800 & ~n11495 ;
  assign n11498 = n1900 ^ n1192 ^ 1'b0 ;
  assign n11497 = n2048 & ~n5844 ;
  assign n11499 = n11498 ^ n11497 ^ 1'b0 ;
  assign n11500 = x155 & ~n8543 ;
  assign n11501 = n8543 & n11500 ;
  assign n11502 = ~n1306 & n10185 ;
  assign n11503 = n1354 & n11502 ;
  assign n11504 = x183 & ~n1506 ;
  assign n11505 = n9483 & ~n11504 ;
  assign n11506 = n4824 | n11092 ;
  assign n11507 = n11506 ^ n5909 ^ 1'b0 ;
  assign n11508 = ( n358 & ~n5699 ) | ( n358 & n11507 ) | ( ~n5699 & n11507 ) ;
  assign n11509 = n1209 & n1693 ;
  assign n11510 = n4776 & n6216 ;
  assign n11511 = n8313 & n11510 ;
  assign n11512 = n4715 & n11511 ;
  assign n11513 = n2844 & ~n11512 ;
  assign n11514 = n11513 ^ n2430 ^ 1'b0 ;
  assign n11515 = n11509 | n11514 ;
  assign n11516 = n1144 & ~n7174 ;
  assign n11517 = n5666 & ~n11516 ;
  assign n11518 = n531 | n11517 ;
  assign n11519 = n10001 ^ n1360 ^ 1'b0 ;
  assign n11520 = n3632 | n6136 ;
  assign n11521 = n11520 ^ n519 ^ 1'b0 ;
  assign n11522 = n11521 ^ n8629 ^ x115 ;
  assign n11523 = n5163 ^ x86 ^ 1'b0 ;
  assign n11524 = n4741 ^ n3566 ^ 1'b0 ;
  assign n11525 = n11524 ^ n6402 ^ 1'b0 ;
  assign n11526 = n11523 & n11525 ;
  assign n11527 = n8659 & n11526 ;
  assign n11528 = n11527 ^ n8101 ^ 1'b0 ;
  assign n11529 = n7706 ^ n5754 ^ 1'b0 ;
  assign n11530 = n1824 | n11529 ;
  assign n11531 = n9011 ^ n643 ^ 1'b0 ;
  assign n11532 = n11531 ^ n8077 ^ n3712 ;
  assign n11533 = n5770 & ~n11532 ;
  assign n11534 = n10679 & n11533 ;
  assign n11535 = n6708 | n9432 ;
  assign n11536 = n639 & ~n11535 ;
  assign n11537 = n11536 ^ n2603 ^ 1'b0 ;
  assign n11538 = n1538 | n11537 ;
  assign n11539 = ~n6045 & n11538 ;
  assign n11540 = n9029 & n11539 ;
  assign n11541 = ( n1813 & n5976 ) | ( n1813 & ~n11540 ) | ( n5976 & ~n11540 ) ;
  assign n11542 = n1590 ^ x158 ^ 1'b0 ;
  assign n11543 = ~n2965 & n11542 ;
  assign n11544 = n8339 & n11543 ;
  assign n11545 = n2162 & n11544 ;
  assign n11549 = n1392 & n3360 ;
  assign n11550 = n11549 ^ n8437 ^ 1'b0 ;
  assign n11546 = n2968 | n6274 ;
  assign n11547 = n4818 | n11546 ;
  assign n11548 = ~n8388 & n11547 ;
  assign n11551 = n11550 ^ n11548 ^ 1'b0 ;
  assign n11552 = ~n2148 & n11551 ;
  assign n11553 = ( n3056 & n3369 ) | ( n3056 & ~n8273 ) | ( n3369 & ~n8273 ) ;
  assign n11554 = n5759 & n6908 ;
  assign n11555 = n4195 ^ n2168 ^ 1'b0 ;
  assign n11556 = ( ~n5522 & n6589 ) | ( ~n5522 & n10973 ) | ( n6589 & n10973 ) ;
  assign n11557 = ~n6121 & n11556 ;
  assign n11558 = n11555 & n11557 ;
  assign n11559 = n2966 | n6288 ;
  assign n11560 = ( n7085 & ~n7199 ) | ( n7085 & n11559 ) | ( ~n7199 & n11559 ) ;
  assign n11561 = n1706 & ~n7253 ;
  assign n11563 = n994 & ~n10777 ;
  assign n11562 = n5084 & ~n7790 ;
  assign n11564 = n11563 ^ n11562 ^ 1'b0 ;
  assign n11565 = n6976 & ~n10179 ;
  assign n11566 = n1073 & ~n7866 ;
  assign n11567 = ( x5 & ~x115 ) | ( x5 & n5725 ) | ( ~x115 & n5725 ) ;
  assign n11568 = n5116 ^ n2808 ^ 1'b0 ;
  assign n11569 = ~n4579 & n11568 ;
  assign n11570 = n8227 & n10279 ;
  assign n11571 = n2080 | n3702 ;
  assign n11572 = ~n6773 & n10225 ;
  assign n11573 = ~n7937 & n11572 ;
  assign n11574 = n9786 | n11573 ;
  assign n11575 = n4433 ^ n332 ^ 1'b0 ;
  assign n11576 = n1271 | n11575 ;
  assign n11577 = n11576 ^ n5052 ^ 1'b0 ;
  assign n11578 = n1200 & ~n9682 ;
  assign n11579 = ~n11577 & n11578 ;
  assign n11580 = n7860 ^ n5772 ^ n4454 ;
  assign n11581 = ( n610 & n2490 ) | ( n610 & ~n11580 ) | ( n2490 & ~n11580 ) ;
  assign n11582 = n10477 & n11581 ;
  assign n11583 = ~n6936 & n11582 ;
  assign n11584 = n2291 ^ n610 ^ 1'b0 ;
  assign n11585 = ~x44 & n11584 ;
  assign n11586 = ~n2681 & n4047 ;
  assign n11587 = ~n2272 & n11586 ;
  assign n11588 = ~n10664 & n11587 ;
  assign n11589 = n530 & ~n9430 ;
  assign n11590 = n11589 ^ n980 ^ 1'b0 ;
  assign n11591 = n1021 & ~n11590 ;
  assign n11592 = n4749 | n4890 ;
  assign n11593 = n11592 ^ n2401 ^ 1'b0 ;
  assign n11594 = n10205 & ~n11593 ;
  assign n11595 = n7726 ^ n5321 ^ 1'b0 ;
  assign n11596 = ~n4840 & n11595 ;
  assign n11597 = n11596 ^ n6577 ^ 1'b0 ;
  assign n11598 = n3073 & n7048 ;
  assign n11599 = n536 & n11598 ;
  assign n11600 = n11599 ^ n4777 ^ 1'b0 ;
  assign n11601 = n3456 & n11600 ;
  assign n11602 = n3438 & n11601 ;
  assign n11603 = ~n7321 & n11602 ;
  assign n11604 = n11603 ^ n7842 ^ 1'b0 ;
  assign n11605 = ~x114 & n635 ;
  assign n11606 = n11605 ^ n10611 ^ 1'b0 ;
  assign n11607 = n745 | n11606 ;
  assign n11613 = n3392 & ~n4607 ;
  assign n11614 = n11613 ^ n2821 ^ 1'b0 ;
  assign n11615 = ~n4355 & n11614 ;
  assign n11608 = ~n1228 & n10332 ;
  assign n11609 = n10019 ^ n8893 ^ 1'b0 ;
  assign n11610 = n2382 | n11609 ;
  assign n11611 = ( n4359 & n9722 ) | ( n4359 & n11610 ) | ( n9722 & n11610 ) ;
  assign n11612 = ~n11608 & n11611 ;
  assign n11616 = n11615 ^ n11612 ^ 1'b0 ;
  assign n11617 = n5558 ^ n4611 ^ 1'b0 ;
  assign n11618 = ~n1147 & n11617 ;
  assign n11619 = n11258 ^ n6309 ^ 1'b0 ;
  assign n11620 = x61 & n11619 ;
  assign n11621 = n11620 ^ n2253 ^ 1'b0 ;
  assign n11622 = n6617 ^ n952 ^ 1'b0 ;
  assign n11623 = ~n11621 & n11622 ;
  assign n11624 = n11623 ^ n719 ^ 1'b0 ;
  assign n11625 = n744 & ~n6444 ;
  assign n11626 = ~n2897 & n11625 ;
  assign n11627 = n10315 ^ n6366 ^ 1'b0 ;
  assign n11628 = n11088 & n11627 ;
  assign n11629 = n6484 ^ n1829 ^ 1'b0 ;
  assign n11630 = n2541 & ~n11629 ;
  assign n11631 = ( n690 & n2812 ) | ( n690 & n11630 ) | ( n2812 & n11630 ) ;
  assign n11632 = n3554 & n7220 ;
  assign n11633 = ~n11631 & n11632 ;
  assign n11634 = n6202 ^ n3601 ^ 1'b0 ;
  assign n11635 = n11634 ^ n7755 ^ 1'b0 ;
  assign n11636 = x105 & n11420 ;
  assign n11637 = n1989 | n7048 ;
  assign n11638 = n8013 | n11637 ;
  assign n11639 = n6811 & n11638 ;
  assign n11640 = n7188 & n11639 ;
  assign n11641 = ~n822 & n1858 ;
  assign n11642 = n11641 ^ n8723 ^ 1'b0 ;
  assign n11643 = ~n11640 & n11642 ;
  assign n11644 = ~n3369 & n11643 ;
  assign n11645 = ~n2687 & n11644 ;
  assign n11646 = n3791 ^ n926 ^ 1'b0 ;
  assign n11647 = n1744 & ~n11646 ;
  assign n11648 = n1697 | n5194 ;
  assign n11649 = n281 | n11648 ;
  assign n11650 = n3806 ^ n3668 ^ 1'b0 ;
  assign n11651 = n2401 | n11650 ;
  assign n11652 = n1900 | n11651 ;
  assign n11653 = n11652 ^ x229 ^ 1'b0 ;
  assign n11654 = n11649 & n11653 ;
  assign n11655 = n11654 ^ n4597 ^ 1'b0 ;
  assign n11656 = ( ~n4681 & n5669 ) | ( ~n4681 & n11073 ) | ( n5669 & n11073 ) ;
  assign n11657 = ~n1227 & n11656 ;
  assign n11658 = ( x198 & n5305 ) | ( x198 & ~n5632 ) | ( n5305 & ~n5632 ) ;
  assign n11659 = n3142 & ~n11658 ;
  assign n11660 = n4220 & n11659 ;
  assign n11661 = ( n519 & n1976 ) | ( n519 & ~n5765 ) | ( n1976 & ~n5765 ) ;
  assign n11662 = n5939 ^ n5079 ^ 1'b0 ;
  assign n11663 = n11547 & n11662 ;
  assign n11664 = ~n6536 & n11663 ;
  assign n11665 = ~n11661 & n11664 ;
  assign n11667 = ( n3051 & n7617 ) | ( n3051 & n7697 ) | ( n7617 & n7697 ) ;
  assign n11666 = ~n4752 & n10040 ;
  assign n11668 = n11667 ^ n11666 ^ 1'b0 ;
  assign n11669 = n2991 & ~n8239 ;
  assign n11670 = n11669 ^ n4093 ^ 1'b0 ;
  assign n11671 = n11670 ^ n5153 ^ 1'b0 ;
  assign n11672 = ~n7828 & n11671 ;
  assign n11673 = n4366 & n11672 ;
  assign n11674 = n11673 ^ n853 ^ 1'b0 ;
  assign n11675 = ~n1520 & n5303 ;
  assign n11676 = n11675 ^ n4986 ^ 1'b0 ;
  assign n11677 = n6907 & n11676 ;
  assign n11678 = n11677 ^ n4038 ^ n3777 ;
  assign n11679 = n10293 ^ n9791 ^ 1'b0 ;
  assign n11680 = x253 & ~n3059 ;
  assign n11681 = ~n10947 & n11680 ;
  assign n11682 = n11681 ^ n9704 ^ 1'b0 ;
  assign n11683 = n5129 & ~n11682 ;
  assign n11687 = ~n1808 & n3460 ;
  assign n11688 = n11687 ^ n851 ^ 1'b0 ;
  assign n11689 = n11688 ^ n6424 ^ n2469 ;
  assign n11685 = n3554 ^ n557 ^ 1'b0 ;
  assign n11686 = n9374 & ~n11685 ;
  assign n11684 = n2358 & ~n2549 ;
  assign n11690 = n11689 ^ n11686 ^ n11684 ;
  assign n11691 = n3245 ^ n1048 ^ 1'b0 ;
  assign n11692 = n7543 & n11691 ;
  assign n11693 = n6577 ^ n3919 ^ 1'b0 ;
  assign n11694 = ~n721 & n11693 ;
  assign n11695 = n6002 | n11694 ;
  assign n11696 = n789 & ~n11695 ;
  assign n11697 = n11696 ^ n6360 ^ 1'b0 ;
  assign n11698 = n11692 & ~n11697 ;
  assign n11699 = n11587 ^ n10999 ^ n451 ;
  assign n11710 = ~n1532 & n5122 ;
  assign n11708 = n5011 ^ n4526 ^ 1'b0 ;
  assign n11709 = ~n1719 & n11708 ;
  assign n11711 = n11710 ^ n11709 ^ 1'b0 ;
  assign n11712 = n11711 ^ n1001 ^ 1'b0 ;
  assign n11700 = n1151 & n3144 ;
  assign n11701 = ~n1780 & n11700 ;
  assign n11702 = n11701 ^ n906 ^ 1'b0 ;
  assign n11703 = n4132 | n11702 ;
  assign n11704 = n369 & ~n11703 ;
  assign n11705 = ~n5049 & n11704 ;
  assign n11706 = n2161 & ~n11705 ;
  assign n11707 = ~n11444 & n11706 ;
  assign n11713 = n11712 ^ n11707 ^ 1'b0 ;
  assign n11714 = n2100 & ~n7706 ;
  assign n11715 = n11714 ^ n8287 ^ 1'b0 ;
  assign n11716 = ~n5016 & n11715 ;
  assign n11717 = n5805 & ~n9752 ;
  assign n11720 = ~n1139 & n3172 ;
  assign n11718 = ( ~n3754 & n8567 ) | ( ~n3754 & n10877 ) | ( n8567 & n10877 ) ;
  assign n11719 = n5464 & n11718 ;
  assign n11721 = n11720 ^ n11719 ^ n7609 ;
  assign n11722 = n2430 ^ n1476 ^ 1'b0 ;
  assign n11723 = n11722 ^ n10093 ^ 1'b0 ;
  assign n11724 = n9362 & ~n11723 ;
  assign n11725 = ~n7200 & n7411 ;
  assign n11726 = ~n1895 & n6604 ;
  assign n11727 = n2839 ^ n2019 ^ 1'b0 ;
  assign n11728 = ~n11726 & n11727 ;
  assign n11729 = n11728 ^ n9619 ^ 1'b0 ;
  assign n11730 = ( ~n7490 & n7866 ) | ( ~n7490 & n11729 ) | ( n7866 & n11729 ) ;
  assign n11734 = n6891 | n7994 ;
  assign n11731 = n3195 | n3625 ;
  assign n11732 = n11731 ^ n6663 ^ 1'b0 ;
  assign n11733 = n10050 & ~n11732 ;
  assign n11735 = n11734 ^ n11733 ^ 1'b0 ;
  assign n11736 = n3269 | n11735 ;
  assign n11737 = n4762 & ~n11736 ;
  assign n11738 = n8202 ^ n7118 ^ x48 ;
  assign n11739 = n11738 ^ n455 ^ 1'b0 ;
  assign n11740 = n1437 | n11739 ;
  assign n11741 = n7797 & ~n11740 ;
  assign n11742 = n6463 ^ n2166 ^ 1'b0 ;
  assign n11743 = n1701 ^ n486 ^ 1'b0 ;
  assign n11744 = n11312 ^ n8790 ^ 1'b0 ;
  assign n11745 = n11743 & ~n11744 ;
  assign n11746 = ( ~n9281 & n11742 ) | ( ~n9281 & n11745 ) | ( n11742 & n11745 ) ;
  assign n11747 = n607 & ~n2075 ;
  assign n11748 = n3759 | n10526 ;
  assign n11749 = n824 & ~n11748 ;
  assign n11750 = ( x151 & ~n11225 ) | ( x151 & n11749 ) | ( ~n11225 & n11749 ) ;
  assign n11751 = n8974 ^ n8901 ^ 1'b0 ;
  assign n11752 = ~n8635 & n9456 ;
  assign n11753 = x88 & ~n6895 ;
  assign n11754 = n9607 ^ n7899 ^ 1'b0 ;
  assign n11755 = n5670 ^ n3534 ^ 1'b0 ;
  assign n11756 = ( ~n2255 & n9743 ) | ( ~n2255 & n11755 ) | ( n9743 & n11755 ) ;
  assign n11757 = n11756 ^ n4389 ^ 1'b0 ;
  assign n11758 = n6386 & ~n11757 ;
  assign n11759 = n7941 | n11758 ;
  assign n11760 = ~n5004 & n5135 ;
  assign n11761 = ~n4284 & n11760 ;
  assign n11762 = ~n2497 & n9185 ;
  assign n11763 = n11761 & n11762 ;
  assign n11764 = ( n7396 & n11759 ) | ( n7396 & ~n11763 ) | ( n11759 & ~n11763 ) ;
  assign n11765 = n7768 ^ n4766 ^ 1'b0 ;
  assign n11766 = ~n2412 & n11677 ;
  assign n11767 = n11766 ^ n560 ^ 1'b0 ;
  assign n11768 = n11765 | n11767 ;
  assign n11769 = n11768 ^ n8996 ^ 1'b0 ;
  assign n11770 = ( x83 & ~n1115 ) | ( x83 & n11769 ) | ( ~n1115 & n11769 ) ;
  assign n11771 = n10937 ^ n7748 ^ 1'b0 ;
  assign n11772 = n4268 ^ n1464 ^ 1'b0 ;
  assign n11773 = n565 & n2954 ;
  assign n11774 = n11772 & ~n11773 ;
  assign n11775 = ~n9913 & n11774 ;
  assign n11776 = ~n10196 & n11775 ;
  assign n11777 = n7817 ^ n6290 ^ 1'b0 ;
  assign n11778 = n9960 ^ n2873 ^ 1'b0 ;
  assign n11779 = n6756 & n10341 ;
  assign n11780 = n11779 ^ n11413 ^ 1'b0 ;
  assign n11781 = ~n2914 & n7301 ;
  assign n11782 = n1148 | n1488 ;
  assign n11783 = n3376 | n11782 ;
  assign n11787 = n5780 ^ n376 ^ 1'b0 ;
  assign n11788 = n4571 & ~n11787 ;
  assign n11784 = n2684 & ~n10121 ;
  assign n11785 = ~n374 & n11784 ;
  assign n11786 = n11785 ^ n1095 ^ 1'b0 ;
  assign n11789 = n11788 ^ n11786 ^ 1'b0 ;
  assign n11790 = n2711 | n11789 ;
  assign n11791 = ~n2663 & n11790 ;
  assign n11792 = n661 | n3241 ;
  assign n11793 = n1629 | n11792 ;
  assign n11794 = n11791 | n11793 ;
  assign n11795 = n11794 ^ n7106 ^ n2489 ;
  assign n11796 = ( n11374 & n11783 ) | ( n11374 & ~n11795 ) | ( n11783 & ~n11795 ) ;
  assign n11797 = x178 & n2534 ;
  assign n11798 = ~n9979 & n11797 ;
  assign n11799 = n3935 & ~n11798 ;
  assign n11800 = n7185 & ~n9911 ;
  assign n11802 = n4533 ^ n4452 ^ n3584 ;
  assign n11801 = n1833 | n6409 ;
  assign n11803 = n11802 ^ n11801 ^ 1'b0 ;
  assign n11804 = n11800 | n11803 ;
  assign n11805 = n3557 & n9425 ;
  assign n11806 = n2137 ^ n2080 ^ 1'b0 ;
  assign n11807 = n11805 | n11806 ;
  assign n11808 = n793 | n11807 ;
  assign n11809 = n11808 ^ n7497 ^ n5569 ;
  assign n11810 = n1097 & ~n8223 ;
  assign n11811 = n474 & ~n11810 ;
  assign n11812 = ~n4931 & n11811 ;
  assign n11813 = ( ~n2781 & n3084 ) | ( ~n2781 & n8245 ) | ( n3084 & n8245 ) ;
  assign n11814 = n8765 ^ n7305 ^ 1'b0 ;
  assign n11815 = ~n2460 & n11814 ;
  assign n11816 = n1203 & ~n1949 ;
  assign n11817 = n11816 ^ n11792 ^ 1'b0 ;
  assign n11818 = n2553 & n9477 ;
  assign n11819 = n8278 | n11818 ;
  assign n11820 = n10582 ^ n3157 ^ 1'b0 ;
  assign n11821 = n7795 | n11820 ;
  assign n11822 = n6393 | n6681 ;
  assign n11823 = n6775 & ~n11822 ;
  assign n11824 = n11377 ^ n3096 ^ 1'b0 ;
  assign n11825 = n11824 ^ n5895 ^ n5182 ;
  assign n11826 = n3695 & ~n9866 ;
  assign n11827 = n11825 & n11826 ;
  assign n11828 = n2063 & ~n11265 ;
  assign n11829 = n438 & n11828 ;
  assign n11830 = n5848 ^ n1766 ^ 1'b0 ;
  assign n11831 = n9304 ^ n1437 ^ 1'b0 ;
  assign n11832 = n10726 ^ n4271 ^ 1'b0 ;
  assign n11833 = ~n2293 & n11832 ;
  assign n11834 = ( n11804 & n11831 ) | ( n11804 & n11833 ) | ( n11831 & n11833 ) ;
  assign n11837 = n379 & ~n9913 ;
  assign n11835 = n1637 & ~n2392 ;
  assign n11836 = n11835 ^ n2674 ^ 1'b0 ;
  assign n11838 = n11837 ^ n11836 ^ 1'b0 ;
  assign n11839 = n2588 ^ n1764 ^ 1'b0 ;
  assign n11840 = n11838 | n11839 ;
  assign n11841 = ~n8052 & n11840 ;
  assign n11842 = ~n2704 & n3332 ;
  assign n11843 = n11842 ^ n8236 ^ 1'b0 ;
  assign n11844 = ~n3877 & n11843 ;
  assign n11845 = n7683 ^ n845 ^ 1'b0 ;
  assign n11846 = n1840 & n10223 ;
  assign n11847 = n5138 ^ n3518 ^ n1875 ;
  assign n11848 = n6352 & ~n11847 ;
  assign n11849 = n4440 ^ n1175 ^ n1145 ;
  assign n11850 = n7982 | n11849 ;
  assign n11851 = n5837 ^ n5817 ^ 1'b0 ;
  assign n11852 = n7088 & n11851 ;
  assign n11853 = n11850 & n11852 ;
  assign n11854 = n1279 & ~n3891 ;
  assign n11855 = n2581 | n11499 ;
  assign n11856 = n2419 | n8616 ;
  assign n11857 = n11856 ^ n6882 ^ 1'b0 ;
  assign n11858 = n6663 | n11857 ;
  assign n11859 = n776 & n1886 ;
  assign n11860 = n11859 ^ n10451 ^ 1'b0 ;
  assign n11861 = ~n5330 & n11860 ;
  assign n11862 = n9807 ^ n3993 ^ 1'b0 ;
  assign n11863 = n11861 & ~n11862 ;
  assign n11864 = x226 & ~n1200 ;
  assign n11865 = n4884 ^ n2751 ^ n1750 ;
  assign n11866 = n11865 ^ n3647 ^ 1'b0 ;
  assign n11867 = n11866 ^ n3920 ^ 1'b0 ;
  assign n11868 = n5115 ^ n4281 ^ 1'b0 ;
  assign n11869 = ~n2070 & n11868 ;
  assign n11870 = ( n11864 & ~n11867 ) | ( n11864 & n11869 ) | ( ~n11867 & n11869 ) ;
  assign n11871 = ~n1648 & n2654 ;
  assign n11872 = n1232 & n11871 ;
  assign n11873 = n2826 | n11872 ;
  assign n11874 = n9952 & n11873 ;
  assign n11875 = ( n9589 & n9857 ) | ( n9589 & n11874 ) | ( n9857 & n11874 ) ;
  assign n11876 = n3985 | n11875 ;
  assign n11877 = n4781 & ~n5133 ;
  assign n11878 = n11877 ^ n7063 ^ 1'b0 ;
  assign n11879 = ~n2674 & n11878 ;
  assign n11885 = n2627 | n5325 ;
  assign n11886 = n11885 ^ n7360 ^ 1'b0 ;
  assign n11880 = n9311 ^ n6536 ^ 1'b0 ;
  assign n11881 = n11734 ^ n1255 ^ 1'b0 ;
  assign n11882 = ~n8562 & n11881 ;
  assign n11883 = ~n11880 & n11882 ;
  assign n11884 = n11883 ^ n9366 ^ 1'b0 ;
  assign n11887 = n11886 ^ n11884 ^ 1'b0 ;
  assign n11888 = n6700 & ~n11887 ;
  assign n11889 = n627 & ~n3985 ;
  assign n11890 = n10329 ^ n9331 ^ 1'b0 ;
  assign n11891 = n1336 & n11890 ;
  assign n11892 = n7910 & n11891 ;
  assign n11893 = n11892 ^ n10420 ^ 1'b0 ;
  assign n11894 = n2746 & n4571 ;
  assign n11895 = ~n6198 & n11894 ;
  assign n11896 = n1538 | n2946 ;
  assign n11897 = n1212 & ~n11896 ;
  assign n11898 = ~n11895 & n11897 ;
  assign n11899 = n11406 ^ n7764 ^ 1'b0 ;
  assign n11900 = ~n8735 & n11899 ;
  assign n11901 = n8945 ^ n5042 ^ 1'b0 ;
  assign n11902 = n8659 | n10745 ;
  assign n11903 = n1553 & n3940 ;
  assign n11904 = ( x178 & n2219 ) | ( x178 & n11903 ) | ( n2219 & n11903 ) ;
  assign n11905 = n11904 ^ n5398 ^ n2285 ;
  assign n11906 = n9005 ^ n1404 ^ n413 ;
  assign n11907 = n2502 | n5538 ;
  assign n11908 = n11906 & ~n11907 ;
  assign n11909 = n2543 & ~n3530 ;
  assign n11910 = n3627 & n11909 ;
  assign n11911 = n7836 & ~n11910 ;
  assign n11912 = n2711 & n11911 ;
  assign n11915 = n10205 ^ n2257 ^ 1'b0 ;
  assign n11913 = n8955 ^ n6079 ^ n681 ;
  assign n11914 = n11913 ^ n8772 ^ n4576 ;
  assign n11916 = n11915 ^ n11914 ^ 1'b0 ;
  assign n11917 = ~n11912 & n11916 ;
  assign n11918 = n10978 ^ n8810 ^ 1'b0 ;
  assign n11919 = n2180 | n3723 ;
  assign n11920 = n11919 ^ n3136 ^ 1'b0 ;
  assign n11921 = n11920 ^ n967 ^ 1'b0 ;
  assign n11922 = n9451 ^ n1300 ^ 1'b0 ;
  assign n11923 = n8810 | n11922 ;
  assign n11924 = n11923 ^ n8938 ^ 1'b0 ;
  assign n11927 = n5898 ^ n2168 ^ 1'b0 ;
  assign n11925 = n2234 | n5074 ;
  assign n11926 = n3050 & ~n11925 ;
  assign n11928 = n11927 ^ n11926 ^ 1'b0 ;
  assign n11929 = n11615 ^ n867 ^ 1'b0 ;
  assign n11930 = n6278 & n9108 ;
  assign n11931 = ( ~n1453 & n8815 ) | ( ~n1453 & n11930 ) | ( n8815 & n11930 ) ;
  assign n11932 = n1451 & n11931 ;
  assign n11933 = ( ~x24 & n2264 ) | ( ~x24 & n11932 ) | ( n2264 & n11932 ) ;
  assign n11934 = n7925 ^ n2120 ^ 1'b0 ;
  assign n11935 = n1622 & n1862 ;
  assign n11936 = n2906 & ~n11935 ;
  assign n11937 = n1132 & n11936 ;
  assign n11938 = n1897 & n7836 ;
  assign n11939 = n9156 | n11938 ;
  assign n11940 = n4526 & ~n4716 ;
  assign n11941 = ( n645 & n7210 ) | ( n645 & ~n11940 ) | ( n7210 & ~n11940 ) ;
  assign n11942 = n2827 | n11941 ;
  assign n11943 = n6321 ^ n5850 ^ n1502 ;
  assign n11944 = n2801 & n4271 ;
  assign n11945 = ~n11943 & n11944 ;
  assign n11946 = n5124 & ~n11945 ;
  assign n11947 = n11946 ^ n8980 ^ 1'b0 ;
  assign n11948 = n10436 | n11947 ;
  assign n11949 = n9062 ^ n8218 ^ n2395 ;
  assign n11951 = n620 ^ n600 ^ 1'b0 ;
  assign n11950 = n4334 ^ n1550 ^ 1'b0 ;
  assign n11952 = n11951 ^ n11950 ^ 1'b0 ;
  assign n11953 = n9502 & n11952 ;
  assign n11954 = n5140 ^ n2541 ^ n1215 ;
  assign n11955 = ~n2262 & n11954 ;
  assign n11956 = x134 & ~n3860 ;
  assign n11957 = n488 | n6964 ;
  assign n11958 = n7939 & ~n11957 ;
  assign n11959 = n11958 ^ n3903 ^ 1'b0 ;
  assign n11960 = n9655 ^ n2168 ^ n2141 ;
  assign n11961 = n7382 ^ n2965 ^ 1'b0 ;
  assign n11962 = n4652 & ~n7549 ;
  assign n11963 = n11961 & n11962 ;
  assign n11966 = n3325 ^ n1231 ^ 1'b0 ;
  assign n11964 = n5119 & n11906 ;
  assign n11965 = n3413 & n11964 ;
  assign n11967 = n11966 ^ n11965 ^ n5329 ;
  assign n11968 = n11967 ^ n9390 ^ n1528 ;
  assign n11969 = ( n3765 & n4284 ) | ( n3765 & n5624 ) | ( n4284 & n5624 ) ;
  assign n11970 = ~n9529 & n10551 ;
  assign n11971 = n7172 & n11970 ;
  assign n11972 = ( n963 & n11969 ) | ( n963 & n11971 ) | ( n11969 & n11971 ) ;
  assign n11973 = n8026 ^ n1792 ^ 1'b0 ;
  assign n11974 = ~n1604 & n2601 ;
  assign n11975 = n2913 & ~n5179 ;
  assign n11976 = n11975 ^ n4454 ^ 1'b0 ;
  assign n11977 = n1495 & ~n11976 ;
  assign n11978 = n2871 & n6447 ;
  assign n11979 = n11978 ^ n3770 ^ 1'b0 ;
  assign n11980 = ~n3388 & n11979 ;
  assign n11981 = n8416 & n11980 ;
  assign n11982 = n1231 & ~n6153 ;
  assign n11983 = n11982 ^ n6646 ^ 1'b0 ;
  assign n11985 = n1130 & n7031 ;
  assign n11986 = n492 & n11985 ;
  assign n11984 = ( x56 & n1636 ) | ( x56 & n2103 ) | ( n1636 & n2103 ) ;
  assign n11987 = n11986 ^ n11984 ^ 1'b0 ;
  assign n11988 = n7668 & n11987 ;
  assign n11989 = n6903 ^ n2434 ^ 1'b0 ;
  assign n11990 = n9104 & n11686 ;
  assign n11991 = n3685 ^ n1228 ^ 1'b0 ;
  assign n11994 = n987 & ~n3725 ;
  assign n11995 = n11994 ^ n2282 ^ 1'b0 ;
  assign n11992 = n3937 ^ n392 ^ 1'b0 ;
  assign n11993 = n3047 & ~n11992 ;
  assign n11996 = n11995 ^ n11993 ^ 1'b0 ;
  assign n11997 = n5141 & ~n11996 ;
  assign n11998 = n8501 ^ n7675 ^ 1'b0 ;
  assign n11999 = n5439 ^ n5064 ^ 1'b0 ;
  assign n12005 = n1707 | n6508 ;
  assign n12006 = n12005 ^ n411 ^ 1'b0 ;
  assign n12000 = n1044 & ~n2068 ;
  assign n12001 = n12000 ^ n2588 ^ 1'b0 ;
  assign n12002 = ~n349 & n3499 ;
  assign n12003 = n12001 & ~n12002 ;
  assign n12004 = n12003 ^ n1442 ^ 1'b0 ;
  assign n12007 = n12006 ^ n12004 ^ 1'b0 ;
  assign n12008 = n7052 ^ n5334 ^ 1'b0 ;
  assign n12009 = n2344 ^ n645 ^ 1'b0 ;
  assign n12010 = n826 & n1737 ;
  assign n12011 = ~n3345 & n12010 ;
  assign n12012 = n8860 ^ n2029 ^ 1'b0 ;
  assign n12013 = ( n12009 & n12011 ) | ( n12009 & n12012 ) | ( n12011 & n12012 ) ;
  assign n12014 = n5225 ^ x230 ^ 1'b0 ;
  assign n12015 = n3297 & ~n12014 ;
  assign n12016 = n4846 | n12015 ;
  assign n12017 = n12016 ^ n11112 ^ 1'b0 ;
  assign n12018 = n5988 | n12017 ;
  assign n12019 = n2380 ^ x207 ^ 1'b0 ;
  assign n12020 = n1026 ^ x77 ^ 1'b0 ;
  assign n12021 = n1887 & n12020 ;
  assign n12022 = n1559 & n12021 ;
  assign n12023 = n12022 ^ n3728 ^ 1'b0 ;
  assign n12024 = ( n2224 & n4579 ) | ( n2224 & ~n12023 ) | ( n4579 & ~n12023 ) ;
  assign n12025 = n9725 | n12024 ;
  assign n12026 = n2325 & n6081 ;
  assign n12027 = n12026 ^ n5415 ^ 1'b0 ;
  assign n12028 = n8976 ^ n3034 ^ 1'b0 ;
  assign n12029 = n7597 & ~n12028 ;
  assign n12030 = n4134 | n4976 ;
  assign n12031 = n12030 ^ n5331 ^ 1'b0 ;
  assign n12032 = n783 & n12031 ;
  assign n12033 = ~n7369 & n12032 ;
  assign n12034 = ~n2190 & n4917 ;
  assign n12035 = n11308 & n12034 ;
  assign n12036 = n11518 ^ n2291 ^ 1'b0 ;
  assign n12037 = n1129 & n12036 ;
  assign n12038 = ~n5478 & n5645 ;
  assign n12039 = n2648 | n12038 ;
  assign n12040 = n11954 ^ n1681 ^ 1'b0 ;
  assign n12041 = n1726 | n12040 ;
  assign n12042 = n4039 ^ n1004 ^ 1'b0 ;
  assign n12043 = ~n10447 & n12042 ;
  assign n12044 = n12041 & n12043 ;
  assign n12045 = n10455 ^ n6945 ^ 1'b0 ;
  assign n12046 = n3659 | n4775 ;
  assign n12047 = n12046 ^ n6327 ^ 1'b0 ;
  assign n12048 = n6736 & ~n12047 ;
  assign n12049 = ~n3843 & n8478 ;
  assign n12050 = n11465 & ~n12049 ;
  assign n12051 = ~n3263 & n12050 ;
  assign n12052 = n793 ^ n306 ^ 1'b0 ;
  assign n12053 = n4368 | n12052 ;
  assign n12054 = n3843 ^ n1462 ^ 1'b0 ;
  assign n12055 = n3091 & ~n12054 ;
  assign n12056 = n3256 | n8503 ;
  assign n12057 = n12056 ^ n354 ^ 1'b0 ;
  assign n12058 = ( ~n9033 & n12055 ) | ( ~n9033 & n12057 ) | ( n12055 & n12057 ) ;
  assign n12059 = n11301 | n11873 ;
  assign n12060 = n11163 & n12059 ;
  assign n12061 = ( n2102 & n2806 ) | ( n2102 & ~n6146 ) | ( n2806 & ~n6146 ) ;
  assign n12062 = n3438 ^ n2890 ^ 1'b0 ;
  assign n12063 = ~n3380 & n8370 ;
  assign n12064 = n11429 & n12063 ;
  assign n12065 = ( x247 & n12062 ) | ( x247 & n12064 ) | ( n12062 & n12064 ) ;
  assign n12069 = n2882 & ~n10159 ;
  assign n12066 = n7598 ^ n7149 ^ x52 ;
  assign n12067 = n12066 ^ n5425 ^ 1'b0 ;
  assign n12068 = ~n3626 & n12067 ;
  assign n12070 = n12069 ^ n12068 ^ 1'b0 ;
  assign n12071 = n5423 & n5481 ;
  assign n12072 = ~n9220 & n9409 ;
  assign n12073 = n3043 & ~n7895 ;
  assign n12074 = n12016 & n12073 ;
  assign n12075 = n2369 | n12074 ;
  assign n12076 = n2327 & n6811 ;
  assign n12077 = n12076 ^ n4711 ^ 1'b0 ;
  assign n12078 = ( n3960 & n7278 ) | ( n3960 & ~n12077 ) | ( n7278 & ~n12077 ) ;
  assign n12079 = x241 | n840 ;
  assign n12080 = n12079 ^ n593 ^ 1'b0 ;
  assign n12081 = n5877 ^ n2431 ^ 1'b0 ;
  assign n12082 = n12080 | n12081 ;
  assign n12083 = n12082 ^ n345 ^ 1'b0 ;
  assign n12084 = n1833 | n10810 ;
  assign n12085 = n12084 ^ n1829 ^ 1'b0 ;
  assign n12086 = n3131 ^ n3120 ^ 1'b0 ;
  assign n12087 = n5805 | n12086 ;
  assign n12088 = n6079 ^ n298 ^ 1'b0 ;
  assign n12089 = n2713 & ~n12088 ;
  assign n12090 = ( n387 & n12087 ) | ( n387 & n12089 ) | ( n12087 & n12089 ) ;
  assign n12093 = n5522 & ~n11805 ;
  assign n12094 = ~n3911 & n12093 ;
  assign n12091 = n9642 ^ n8129 ^ n4099 ;
  assign n12092 = n5783 & n12091 ;
  assign n12095 = n12094 ^ n12092 ^ 1'b0 ;
  assign n12096 = ~n467 & n12095 ;
  assign n12097 = n9246 & n12096 ;
  assign n12098 = ~n3055 & n11937 ;
  assign n12099 = n12098 ^ n2471 ^ 1'b0 ;
  assign n12100 = n2885 & n10204 ;
  assign n12101 = ~n4135 & n12100 ;
  assign n12102 = n4592 | n12101 ;
  assign n12103 = ~n1152 & n12102 ;
  assign n12104 = n5081 | n8750 ;
  assign n12105 = n12104 ^ n8512 ^ 1'b0 ;
  assign n12106 = ( ~n3979 & n10845 ) | ( ~n3979 & n12105 ) | ( n10845 & n12105 ) ;
  assign n12107 = n1666 & ~n2698 ;
  assign n12108 = n12107 ^ n3798 ^ 1'b0 ;
  assign n12109 = n7639 ^ n365 ^ 1'b0 ;
  assign n12110 = n12108 & ~n12109 ;
  assign n12111 = ~n5992 & n12110 ;
  assign n12112 = n12111 ^ n9630 ^ 1'b0 ;
  assign n12113 = n10447 ^ n3365 ^ 1'b0 ;
  assign n12114 = n12113 ^ n10837 ^ n7429 ;
  assign n12115 = ( ~x63 & n4284 ) | ( ~x63 & n8386 ) | ( n4284 & n8386 ) ;
  assign n12116 = n10692 ^ n9490 ^ n6869 ;
  assign n12117 = n12116 ^ n4957 ^ 1'b0 ;
  assign n12118 = n4385 ^ n1508 ^ 1'b0 ;
  assign n12119 = n2807 | n12118 ;
  assign n12120 = n2176 | n6400 ;
  assign n12121 = n12120 ^ n9541 ^ 1'b0 ;
  assign n12122 = n12121 ^ n3447 ^ 1'b0 ;
  assign n12123 = ~n1572 & n12122 ;
  assign n12124 = ~n12119 & n12123 ;
  assign n12125 = n5708 ^ n1780 ^ n1364 ;
  assign n12130 = ~n10313 & n10624 ;
  assign n12126 = ( n1202 & ~n2406 ) | ( n1202 & n2956 ) | ( ~n2406 & n2956 ) ;
  assign n12127 = n1393 & n12126 ;
  assign n12128 = n12127 ^ n4967 ^ 1'b0 ;
  assign n12129 = ~n6423 & n12128 ;
  assign n12131 = n12130 ^ n12129 ^ 1'b0 ;
  assign n12132 = n4724 | n10640 ;
  assign n12135 = n4654 ^ n2057 ^ n1848 ;
  assign n12133 = n2952 & ~n3757 ;
  assign n12134 = ( n3072 & ~n10480 ) | ( n3072 & n12133 ) | ( ~n10480 & n12133 ) ;
  assign n12136 = n12135 ^ n12134 ^ n5720 ;
  assign n12137 = x233 & ~n626 ;
  assign n12138 = n12137 ^ n997 ^ 1'b0 ;
  assign n12139 = n12138 ^ n11019 ^ 1'b0 ;
  assign n12140 = ~n6602 & n12139 ;
  assign n12144 = n6849 ^ n2096 ^ 1'b0 ;
  assign n12141 = n6276 & ~n9230 ;
  assign n12142 = n12141 ^ n3588 ^ 1'b0 ;
  assign n12143 = n3218 & ~n12142 ;
  assign n12145 = n12144 ^ n12143 ^ 1'b0 ;
  assign n12146 = n2449 & n12145 ;
  assign n12147 = ~n3689 & n12146 ;
  assign n12148 = ~n2230 & n7346 ;
  assign n12149 = n12148 ^ n918 ^ 1'b0 ;
  assign n12150 = n12147 | n12149 ;
  assign n12151 = ~n3635 & n4105 ;
  assign n12152 = n5652 ^ n1509 ^ 1'b0 ;
  assign n12153 = ( n269 & ~n9259 ) | ( n269 & n12152 ) | ( ~n9259 & n12152 ) ;
  assign n12154 = n1235 ^ n780 ^ 1'b0 ;
  assign n12155 = ~n12153 & n12154 ;
  assign n12156 = n2218 & ~n10221 ;
  assign n12157 = n12156 ^ n6307 ^ 1'b0 ;
  assign n12158 = n11374 ^ n9437 ^ 1'b0 ;
  assign n12159 = n8572 & n11587 ;
  assign n12160 = n12159 ^ n2922 ^ 1'b0 ;
  assign n12161 = n4615 ^ n759 ^ 1'b0 ;
  assign n12162 = ( n1173 & n1869 ) | ( n1173 & n7462 ) | ( n1869 & n7462 ) ;
  assign n12163 = n12161 & n12162 ;
  assign n12164 = n2497 | n12163 ;
  assign n12165 = n12164 ^ x160 ^ 1'b0 ;
  assign n12166 = x120 & ~n9854 ;
  assign n12167 = n12166 ^ n9467 ^ 1'b0 ;
  assign n12168 = n12167 ^ n8528 ^ n4534 ;
  assign n12169 = n2036 ^ n1791 ^ 1'b0 ;
  assign n12170 = n1869 & ~n12169 ;
  assign n12171 = n12170 ^ n4232 ^ 1'b0 ;
  assign n12172 = n12171 ^ n9912 ^ n4154 ;
  assign n12173 = n1362 & n5422 ;
  assign n12174 = n12173 ^ n3360 ^ 1'b0 ;
  assign n12175 = n5303 | n12174 ;
  assign n12176 = n12175 ^ n6602 ^ n952 ;
  assign n12177 = n9759 ^ n4802 ^ n3277 ;
  assign n12178 = n12177 ^ n9484 ^ n8698 ;
  assign n12179 = n8301 | n10036 ;
  assign n12180 = n12179 ^ n5461 ^ 1'b0 ;
  assign n12181 = x139 & n3229 ;
  assign n12182 = n4647 & n12181 ;
  assign n12183 = ~n5945 & n10777 ;
  assign n12184 = n12183 ^ n4196 ^ 1'b0 ;
  assign n12185 = n12184 ^ n9253 ^ 1'b0 ;
  assign n12186 = ( x111 & n12182 ) | ( x111 & ~n12185 ) | ( n12182 & ~n12185 ) ;
  assign n12187 = ~n3654 & n3720 ;
  assign n12188 = n1418 | n2322 ;
  assign n12189 = n2282 | n12188 ;
  assign n12190 = n600 & n12189 ;
  assign n12191 = ( n3104 & n3142 ) | ( n3104 & ~n5176 ) | ( n3142 & ~n5176 ) ;
  assign n12192 = n7709 ^ n2048 ^ 1'b0 ;
  assign n12193 = ~n12191 & n12192 ;
  assign n12194 = n8901 & ~n12193 ;
  assign n12195 = n5264 & ~n12194 ;
  assign n12196 = n6607 & n9477 ;
  assign n12197 = n12196 ^ n11309 ^ 1'b0 ;
  assign n12198 = n7110 | n12189 ;
  assign n12199 = n3312 ^ n1040 ^ 1'b0 ;
  assign n12200 = n12199 ^ n4760 ^ 1'b0 ;
  assign n12201 = ~n9561 & n12200 ;
  assign n12202 = n12201 ^ n7480 ^ 1'b0 ;
  assign n12203 = n4966 ^ n3138 ^ 1'b0 ;
  assign n12204 = ~n5797 & n12203 ;
  assign n12205 = ~n5359 & n5684 ;
  assign n12206 = n607 & ~n1762 ;
  assign n12207 = n12206 ^ n840 ^ 1'b0 ;
  assign n12208 = n12207 ^ n2623 ^ 1'b0 ;
  assign n12209 = n1758 | n10794 ;
  assign n12210 = ( n353 & n2658 ) | ( n353 & ~n4917 ) | ( n2658 & ~n4917 ) ;
  assign n12211 = n405 & n12210 ;
  assign n12212 = n12211 ^ n6142 ^ 1'b0 ;
  assign n12213 = n12209 & n12212 ;
  assign n12214 = x87 & ~n604 ;
  assign n12215 = n12214 ^ n879 ^ 1'b0 ;
  assign n12216 = n4719 ^ n2102 ^ 1'b0 ;
  assign n12217 = n10907 & ~n12216 ;
  assign n12218 = n12215 & n12217 ;
  assign n12219 = n12218 ^ n11907 ^ 1'b0 ;
  assign n12220 = n2959 & ~n9128 ;
  assign n12221 = n5731 & n12220 ;
  assign n12222 = n11767 ^ n6327 ^ 1'b0 ;
  assign n12223 = ~n12221 & n12222 ;
  assign n12225 = n2212 | n11191 ;
  assign n12226 = n12225 ^ n2882 ^ 1'b0 ;
  assign n12224 = n598 & n3062 ;
  assign n12227 = n12226 ^ n12224 ^ 1'b0 ;
  assign n12228 = n12227 ^ n8545 ^ 1'b0 ;
  assign n12229 = n12228 ^ n1763 ^ 1'b0 ;
  assign n12230 = ~n1712 & n2399 ;
  assign n12231 = n12229 & n12230 ;
  assign n12232 = n1777 | n4148 ;
  assign n12233 = n5295 & ~n12232 ;
  assign n12234 = n753 & ~n7000 ;
  assign n12235 = n12234 ^ n6149 ^ 1'b0 ;
  assign n12236 = n11533 ^ n4310 ^ 1'b0 ;
  assign n12237 = n380 & ~n11603 ;
  assign n12240 = ~n2869 & n5115 ;
  assign n12241 = n1657 & n12240 ;
  assign n12238 = n1058 ^ x36 ^ 1'b0 ;
  assign n12239 = n8865 | n12238 ;
  assign n12242 = n12241 ^ n12239 ^ 1'b0 ;
  assign n12243 = ~n9155 & n9822 ;
  assign n12244 = n2801 & ~n3430 ;
  assign n12245 = n12244 ^ n6885 ^ 1'b0 ;
  assign n12246 = n6096 ^ n1913 ^ 1'b0 ;
  assign n12247 = n6630 | n12246 ;
  assign n12248 = n5170 | n11426 ;
  assign n12252 = x25 & x187 ;
  assign n12253 = n12252 ^ n2875 ^ 1'b0 ;
  assign n12251 = x130 & n509 ;
  assign n12249 = n3803 & ~n4563 ;
  assign n12250 = n12249 ^ n5828 ^ 1'b0 ;
  assign n12254 = n12253 ^ n12251 ^ n12250 ;
  assign n12255 = n12254 ^ n4662 ^ 1'b0 ;
  assign n12256 = ( n6920 & ~n7463 ) | ( n6920 & n12255 ) | ( ~n7463 & n12255 ) ;
  assign n12257 = n12256 ^ n7535 ^ n6731 ;
  assign n12258 = n6021 & n12257 ;
  assign n12259 = ~n371 & n7128 ;
  assign n12260 = n12259 ^ n533 ^ 1'b0 ;
  assign n12261 = n3798 | n12260 ;
  assign n12262 = x195 & n2884 ;
  assign n12263 = n12262 ^ n3208 ^ 1'b0 ;
  assign n12264 = n3947 | n12263 ;
  assign n12265 = n12261 | n12264 ;
  assign n12266 = n2012 & ~n7540 ;
  assign n12267 = n7377 & n12266 ;
  assign n12268 = ~n1525 & n12267 ;
  assign n12269 = ( x120 & n4102 ) | ( x120 & n5623 ) | ( n4102 & n5623 ) ;
  assign n12270 = n12269 ^ n7531 ^ 1'b0 ;
  assign n12271 = n2939 & n12270 ;
  assign n12272 = n12271 ^ n2262 ^ 1'b0 ;
  assign n12273 = n12268 | n12272 ;
  assign n12274 = x5 & n9731 ;
  assign n12275 = n1254 & n12274 ;
  assign n12276 = n1868 & ~n7965 ;
  assign n12277 = n5598 & n12276 ;
  assign n12278 = ( ~n3318 & n3725 ) | ( ~n3318 & n12277 ) | ( n3725 & n12277 ) ;
  assign n12279 = n1793 & n3743 ;
  assign n12280 = n1801 | n5271 ;
  assign n12281 = x221 | n12280 ;
  assign n12285 = n7480 ^ n4086 ^ 1'b0 ;
  assign n12282 = n2437 ^ n700 ^ 1'b0 ;
  assign n12283 = n12282 ^ n740 ^ 1'b0 ;
  assign n12284 = ~n10615 & n12283 ;
  assign n12286 = n12285 ^ n12284 ^ 1'b0 ;
  assign n12295 = ~n2028 & n4442 ;
  assign n12296 = n5621 & n12295 ;
  assign n12289 = n1660 & ~n2054 ;
  assign n12287 = x31 & ~n3296 ;
  assign n12288 = n12287 ^ n4066 ^ 1'b0 ;
  assign n12290 = n12289 ^ n12288 ^ 1'b0 ;
  assign n12291 = n3880 & ~n12290 ;
  assign n12292 = n3556 & n6430 ;
  assign n12293 = ~n12291 & n12292 ;
  assign n12294 = n12021 & ~n12293 ;
  assign n12297 = n12296 ^ n12294 ^ 1'b0 ;
  assign n12298 = x85 & n3989 ;
  assign n12299 = n12298 ^ n3374 ^ 1'b0 ;
  assign n12300 = n12299 ^ n8900 ^ n4349 ;
  assign n12301 = n10548 ^ n5075 ^ 1'b0 ;
  assign n12302 = n4807 & n12301 ;
  assign n12303 = n5264 | n6846 ;
  assign n12304 = n12303 ^ n3332 ^ 1'b0 ;
  assign n12305 = n10313 ^ n8639 ^ 1'b0 ;
  assign n12321 = n3103 ^ n529 ^ 1'b0 ;
  assign n12316 = n1679 & ~n1804 ;
  assign n12317 = n3915 & n12316 ;
  assign n12318 = n12317 ^ x110 ^ 1'b0 ;
  assign n12319 = n10311 | n12318 ;
  assign n12307 = n5384 ^ n4160 ^ 1'b0 ;
  assign n12308 = n8949 & n12307 ;
  assign n12309 = ~n690 & n1683 ;
  assign n12310 = ~n12308 & n12309 ;
  assign n12311 = ~n1162 & n3053 ;
  assign n12312 = n12311 ^ n1336 ^ 1'b0 ;
  assign n12313 = n12312 ^ n10530 ^ n2942 ;
  assign n12314 = ~n5226 & n12313 ;
  assign n12315 = n12310 & n12314 ;
  assign n12320 = n12319 ^ n12315 ^ 1'b0 ;
  assign n12306 = n5666 & n9614 ;
  assign n12322 = n12321 ^ n12320 ^ n12306 ;
  assign n12323 = n2440 & n6966 ;
  assign n12324 = n329 | n12323 ;
  assign n12325 = n1419 | n9827 ;
  assign n12326 = n3517 ^ n3174 ^ 1'b0 ;
  assign n12327 = n6192 & n12326 ;
  assign n12328 = ~n12325 & n12327 ;
  assign n12329 = ~n8236 & n12328 ;
  assign n12330 = n2963 & ~n5671 ;
  assign n12331 = n12330 ^ n3993 ^ 1'b0 ;
  assign n12332 = n7088 & ~n12331 ;
  assign n12333 = n12332 ^ x149 ^ 1'b0 ;
  assign n12334 = n4981 | n12333 ;
  assign n12335 = ~n4525 & n11457 ;
  assign n12336 = n10122 & ~n12335 ;
  assign n12337 = ~n647 & n12336 ;
  assign n12338 = n8770 | n9120 ;
  assign n12339 = n3464 & ~n12338 ;
  assign n12340 = ( n1140 & ~n2564 ) | ( n1140 & n4298 ) | ( ~n2564 & n4298 ) ;
  assign n12341 = ( ~n3871 & n9383 ) | ( ~n3871 & n12340 ) | ( n9383 & n12340 ) ;
  assign n12342 = ( n347 & n4208 ) | ( n347 & ~n9088 ) | ( n4208 & ~n9088 ) ;
  assign n12343 = ~n8592 & n10534 ;
  assign n12344 = n11961 ^ n11517 ^ n5295 ;
  assign n12345 = n363 | n2530 ;
  assign n12346 = n2004 | n12345 ;
  assign n12352 = ~n1093 & n2031 ;
  assign n12353 = ~n3196 & n12352 ;
  assign n12354 = n12353 ^ n2959 ^ 1'b0 ;
  assign n12355 = n4641 & ~n12354 ;
  assign n12347 = ( n2824 & ~n3926 ) | ( n2824 & n5684 ) | ( ~n3926 & n5684 ) ;
  assign n12348 = n930 ^ x180 ^ x103 ;
  assign n12349 = ~n4907 & n12348 ;
  assign n12350 = n5949 & n12349 ;
  assign n12351 = ( n12299 & n12347 ) | ( n12299 & ~n12350 ) | ( n12347 & ~n12350 ) ;
  assign n12356 = n12355 ^ n12351 ^ 1'b0 ;
  assign n12357 = n5107 ^ n3374 ^ n2146 ;
  assign n12358 = n9099 ^ n1253 ^ 1'b0 ;
  assign n12359 = ~n3366 & n12358 ;
  assign n12360 = ~n12357 & n12359 ;
  assign n12361 = ~n6673 & n10114 ;
  assign n12362 = n5680 & n12361 ;
  assign n12363 = ( n6590 & ~n7753 ) | ( n6590 & n9831 ) | ( ~n7753 & n9831 ) ;
  assign n12364 = n11312 ^ n6853 ^ 1'b0 ;
  assign n12365 = ~n2950 & n12364 ;
  assign n12366 = ( n489 & n3583 ) | ( n489 & ~n12365 ) | ( n3583 & ~n12365 ) ;
  assign n12367 = n12366 ^ n11859 ^ 1'b0 ;
  assign n12368 = n12363 & ~n12367 ;
  assign n12369 = n7954 & ~n10469 ;
  assign n12370 = n12369 ^ n6430 ^ 1'b0 ;
  assign n12372 = x43 | n2052 ;
  assign n12373 = n3681 & ~n12372 ;
  assign n12371 = ~n2941 & n7403 ;
  assign n12374 = n12373 ^ n12371 ^ 1'b0 ;
  assign n12375 = n10577 & n12374 ;
  assign n12376 = n9065 ^ n2169 ^ n1679 ;
  assign n12381 = n3185 ^ n2061 ^ 1'b0 ;
  assign n12382 = n2851 & ~n12381 ;
  assign n12383 = x205 & n12382 ;
  assign n12384 = n12383 ^ n7294 ^ 1'b0 ;
  assign n12377 = n2832 ^ n2165 ^ 1'b0 ;
  assign n12378 = n1059 | n12377 ;
  assign n12379 = n12378 ^ n773 ^ 1'b0 ;
  assign n12380 = ~n9054 & n12379 ;
  assign n12385 = n12384 ^ n12380 ^ 1'b0 ;
  assign n12388 = n8773 ^ n7863 ^ n5790 ;
  assign n12386 = n8398 ^ n5800 ^ 1'b0 ;
  assign n12387 = n527 | n12386 ;
  assign n12389 = n12388 ^ n12387 ^ 1'b0 ;
  assign n12390 = n2651 ^ n1959 ^ n950 ;
  assign n12391 = n5456 & n12390 ;
  assign n12392 = n12391 ^ x81 ^ 1'b0 ;
  assign n12393 = n12389 | n12392 ;
  assign n12394 = n5639 & ~n12393 ;
  assign n12395 = n8924 | n9977 ;
  assign n12396 = n1559 | n12395 ;
  assign n12397 = n9950 ^ n6682 ^ 1'b0 ;
  assign n12398 = n4704 & ~n12397 ;
  assign n12399 = n2148 | n12398 ;
  assign n12400 = n7426 ^ n7219 ^ n2796 ;
  assign n12401 = n12400 ^ n8352 ^ 1'b0 ;
  assign n12402 = n10567 & n12401 ;
  assign n12403 = n8388 ^ n7041 ^ 1'b0 ;
  assign n12404 = n5164 | n10429 ;
  assign n12405 = n3556 | n12404 ;
  assign n12406 = ( n1330 & ~n2831 ) | ( n1330 & n3175 ) | ( ~n2831 & n3175 ) ;
  assign n12407 = n12406 ^ n10707 ^ 1'b0 ;
  assign n12408 = n10891 & n12407 ;
  assign n12409 = n462 & ~n5613 ;
  assign n12410 = n5059 & n12409 ;
  assign n12411 = n12365 | n12410 ;
  assign n12412 = n12411 ^ n271 ^ 1'b0 ;
  assign n12413 = n4927 & n12412 ;
  assign n12414 = ( n894 & ~n2419 ) | ( n894 & n3963 ) | ( ~n2419 & n3963 ) ;
  assign n12415 = n12414 ^ n960 ^ 1'b0 ;
  assign n12416 = n12415 ^ n5484 ^ 1'b0 ;
  assign n12417 = n12413 & ~n12416 ;
  assign n12418 = x28 & n1785 ;
  assign n12419 = n12418 ^ n1099 ^ 1'b0 ;
  assign n12420 = n12419 ^ n8056 ^ n4638 ;
  assign n12421 = n11956 | n11974 ;
  assign n12422 = ~n1325 & n4918 ;
  assign n12423 = ~n4918 & n12422 ;
  assign n12424 = n4086 | n7245 ;
  assign n12425 = n12423 & ~n12424 ;
  assign n12426 = n12425 ^ n4644 ^ 1'b0 ;
  assign n12429 = n1156 & ~n1878 ;
  assign n12427 = n6909 ^ n995 ^ 1'b0 ;
  assign n12428 = n6910 & n12427 ;
  assign n12430 = n12429 ^ n12428 ^ 1'b0 ;
  assign n12431 = n4039 | n12430 ;
  assign n12432 = n4828 | n12431 ;
  assign n12433 = ~n4015 & n9150 ;
  assign n12434 = n12433 ^ n3048 ^ 1'b0 ;
  assign n12435 = n12161 & n12434 ;
  assign n12436 = ( n2601 & ~n7381 ) | ( n2601 & n12435 ) | ( ~n7381 & n12435 ) ;
  assign n12437 = n8234 | n10688 ;
  assign n12442 = n7040 ^ n5694 ^ 1'b0 ;
  assign n12443 = n5285 & n12442 ;
  assign n12444 = n7795 & n12443 ;
  assign n12438 = n3877 | n11421 ;
  assign n12439 = ~n9269 & n12438 ;
  assign n12440 = n12439 ^ n9534 ^ 1'b0 ;
  assign n12441 = n11924 & ~n12440 ;
  assign n12445 = n12444 ^ n12441 ^ 1'b0 ;
  assign n12446 = n4707 & ~n8866 ;
  assign n12447 = n12391 & ~n12446 ;
  assign n12448 = n12447 ^ n3832 ^ 1'b0 ;
  assign n12449 = ~n4506 & n4954 ;
  assign n12450 = ~n6215 & n7037 ;
  assign n12451 = n12450 ^ n983 ^ 1'b0 ;
  assign n12452 = n10443 ^ n4286 ^ 1'b0 ;
  assign n12453 = n12451 & ~n12452 ;
  assign n12454 = n968 | n8756 ;
  assign n12455 = n5085 & n6529 ;
  assign n12456 = ( n3396 & n7802 ) | ( n3396 & ~n12455 ) | ( n7802 & ~n12455 ) ;
  assign n12461 = n2564 | n3673 ;
  assign n12462 = n12461 ^ n3063 ^ 1'b0 ;
  assign n12463 = n12462 ^ n1442 ^ 1'b0 ;
  assign n12464 = n8708 | n12463 ;
  assign n12457 = n2534 & n4969 ;
  assign n12458 = n12457 ^ n3256 ^ 1'b0 ;
  assign n12459 = ~n4945 & n12458 ;
  assign n12460 = n4726 & n12459 ;
  assign n12465 = n12464 ^ n12460 ^ 1'b0 ;
  assign n12466 = ~n4990 & n12465 ;
  assign n12467 = n3531 & ~n6279 ;
  assign n12468 = ~n598 & n12467 ;
  assign n12469 = n8128 | n12468 ;
  assign n12470 = ~n2202 & n4597 ;
  assign n12471 = n10620 & ~n11920 ;
  assign n12472 = n495 | n4677 ;
  assign n12473 = n5135 & n12472 ;
  assign n12474 = ( n5257 & n5977 ) | ( n5257 & n12473 ) | ( n5977 & n12473 ) ;
  assign n12479 = n5765 ^ n449 ^ x87 ;
  assign n12475 = n8908 ^ n259 ^ 1'b0 ;
  assign n12476 = n1277 & n3369 ;
  assign n12477 = n12475 & n12476 ;
  assign n12478 = ~n6762 & n12477 ;
  assign n12480 = n12479 ^ n12478 ^ 1'b0 ;
  assign n12481 = n12480 ^ n10001 ^ 1'b0 ;
  assign n12482 = n3068 & n7157 ;
  assign n12483 = n12482 ^ n5432 ^ 1'b0 ;
  assign n12484 = ( ~n6797 & n11769 ) | ( ~n6797 & n12483 ) | ( n11769 & n12483 ) ;
  assign n12485 = ~n1782 & n6755 ;
  assign n12486 = n12485 ^ n6522 ^ 1'b0 ;
  assign n12487 = n3869 & ~n12486 ;
  assign n12488 = n12487 ^ n11160 ^ 1'b0 ;
  assign n12489 = x67 & n10788 ;
  assign n12490 = n12489 ^ n3466 ^ 1'b0 ;
  assign n12491 = ~n2054 & n2253 ;
  assign n12492 = n5735 & ~n12491 ;
  assign n12493 = n12492 ^ x38 ^ 1'b0 ;
  assign n12494 = ( x214 & n5671 ) | ( x214 & ~n8598 ) | ( n5671 & ~n8598 ) ;
  assign n12495 = n12494 ^ n7583 ^ 1'b0 ;
  assign n12496 = n5588 ^ n2869 ^ 1'b0 ;
  assign n12497 = n12495 & n12496 ;
  assign n12498 = n1550 & ~n2741 ;
  assign n12499 = n2440 | n12498 ;
  assign n12500 = n12499 ^ n4531 ^ 1'b0 ;
  assign n12501 = n7398 | n12500 ;
  assign n12502 = n12501 ^ n5830 ^ n1271 ;
  assign n12503 = n2214 & ~n8461 ;
  assign n12504 = n2347 ^ x87 ^ 1'b0 ;
  assign n12505 = n4499 & ~n12504 ;
  assign n12506 = ~n3890 & n12505 ;
  assign n12507 = ~n12505 & n12506 ;
  assign n12508 = n5141 | n12507 ;
  assign n12509 = n12507 & ~n12508 ;
  assign n12510 = n5276 ^ n3666 ^ n1358 ;
  assign n12511 = n12509 | n12510 ;
  assign n12512 = n12511 ^ n3150 ^ 1'b0 ;
  assign n12513 = ~n1980 & n2546 ;
  assign n12514 = n6246 & n12513 ;
  assign n12515 = n6552 & ~n12514 ;
  assign n12516 = n489 & n12515 ;
  assign n12517 = n12516 ^ n8957 ^ 1'b0 ;
  assign n12518 = n3702 & n12517 ;
  assign n12520 = n1769 | n7293 ;
  assign n12521 = n7074 & ~n12520 ;
  assign n12519 = n6450 ^ n2070 ^ 1'b0 ;
  assign n12522 = n12521 ^ n12519 ^ 1'b0 ;
  assign n12523 = n1228 & ~n5114 ;
  assign n12524 = x23 & ~n9826 ;
  assign n12525 = n3133 & n4355 ;
  assign n12526 = n12525 ^ n305 ^ 1'b0 ;
  assign n12527 = ( ~n6466 & n12524 ) | ( ~n6466 & n12526 ) | ( n12524 & n12526 ) ;
  assign n12528 = n10905 ^ n8445 ^ n981 ;
  assign n12529 = n6233 & n12528 ;
  assign n12530 = n826 & n3640 ;
  assign n12531 = ( n5476 & n11866 ) | ( n5476 & ~n12530 ) | ( n11866 & ~n12530 ) ;
  assign n12532 = n12531 ^ n5979 ^ n4606 ;
  assign n12533 = n4736 | n12532 ;
  assign n12534 = n11268 & ~n11292 ;
  assign n12535 = n397 & n3333 ;
  assign n12536 = n12535 ^ n3320 ^ 1'b0 ;
  assign n12537 = n5463 & n12536 ;
  assign n12538 = n1746 & ~n12537 ;
  assign n12539 = ~n5081 & n9997 ;
  assign n12540 = n12539 ^ n2216 ^ 1'b0 ;
  assign n12541 = n2832 & ~n5257 ;
  assign n12542 = n12541 ^ n6159 ^ 1'b0 ;
  assign n12543 = n4024 | n5261 ;
  assign n12544 = n12543 ^ n4852 ^ 1'b0 ;
  assign n12545 = n2276 & n12544 ;
  assign n12546 = ~n12542 & n12545 ;
  assign n12547 = n12546 ^ n6754 ^ 1'b0 ;
  assign n12548 = n301 | n3924 ;
  assign n12549 = n7887 ^ n1725 ^ 1'b0 ;
  assign n12550 = n1665 & ~n12549 ;
  assign n12551 = n12550 ^ n3449 ^ 1'b0 ;
  assign n12552 = n12551 ^ n1228 ^ 1'b0 ;
  assign n12553 = n5246 ^ n1005 ^ 1'b0 ;
  assign n12554 = ~n5271 & n12553 ;
  assign n12555 = n12554 ^ n3326 ^ x103 ;
  assign n12561 = n4281 & n6888 ;
  assign n12562 = n6115 & n12561 ;
  assign n12558 = ~n2743 & n5837 ;
  assign n12556 = x28 & ~n7942 ;
  assign n12557 = n12556 ^ n6781 ^ 1'b0 ;
  assign n12559 = n12558 ^ n12557 ^ n5652 ;
  assign n12560 = n1679 & n12559 ;
  assign n12563 = n12562 ^ n12560 ^ 1'b0 ;
  assign n12565 = n11531 ^ n2284 ^ 1'b0 ;
  assign n12566 = n11930 & ~n12565 ;
  assign n12564 = n3725 ^ n883 ^ 1'b0 ;
  assign n12567 = n12566 ^ n12564 ^ n9483 ;
  assign n12568 = ~x137 & n6739 ;
  assign n12570 = n7804 ^ n6508 ^ 1'b0 ;
  assign n12571 = n7494 & ~n12570 ;
  assign n12572 = ( n3439 & n10624 ) | ( n3439 & ~n12571 ) | ( n10624 & ~n12571 ) ;
  assign n12573 = n4878 | n12572 ;
  assign n12569 = n1273 & ~n5598 ;
  assign n12574 = n12573 ^ n12569 ^ 1'b0 ;
  assign n12575 = n12574 ^ n4567 ^ 1'b0 ;
  assign n12577 = n5269 | n5352 ;
  assign n12578 = n12577 ^ n10425 ^ 1'b0 ;
  assign n12576 = n341 | n2341 ;
  assign n12579 = n12578 ^ n12576 ^ 1'b0 ;
  assign n12580 = n5978 & ~n6227 ;
  assign n12581 = ~n5648 & n7231 ;
  assign n12582 = n12581 ^ n2293 ^ 1'b0 ;
  assign n12586 = ~n5194 & n11531 ;
  assign n12587 = ~n1246 & n12586 ;
  assign n12583 = ~n1453 & n7585 ;
  assign n12584 = n12583 ^ n8474 ^ 1'b0 ;
  assign n12585 = ~n9742 & n12584 ;
  assign n12588 = n12587 ^ n12585 ^ 1'b0 ;
  assign n12589 = n2807 ^ n2302 ^ 1'b0 ;
  assign n12590 = n4378 | n12589 ;
  assign n12591 = n12590 ^ n2907 ^ 1'b0 ;
  assign n12592 = n7515 & ~n8535 ;
  assign n12593 = n12592 ^ n6464 ^ 1'b0 ;
  assign n12594 = ~n12591 & n12593 ;
  assign n12595 = ( n3420 & ~n4932 ) | ( n3420 & n10760 ) | ( ~n4932 & n10760 ) ;
  assign n12596 = n4289 | n9341 ;
  assign n12597 = n12596 ^ x154 ^ 1'b0 ;
  assign n12598 = ( n9139 & n12595 ) | ( n9139 & n12597 ) | ( n12595 & n12597 ) ;
  assign n12599 = n8618 ^ n803 ^ 1'b0 ;
  assign n12600 = ~n1023 & n12599 ;
  assign n12601 = n12600 ^ x115 ^ 1'b0 ;
  assign n12602 = n11920 ^ n8639 ^ 1'b0 ;
  assign n12603 = n12601 | n12602 ;
  assign n12604 = n12603 ^ n2523 ^ 1'b0 ;
  assign n12605 = n9222 ^ n4376 ^ 1'b0 ;
  assign n12606 = n1603 & n12605 ;
  assign n12607 = ~x200 & n3172 ;
  assign n12608 = ( n7514 & ~n12606 ) | ( n7514 & n12607 ) | ( ~n12606 & n12607 ) ;
  assign n12609 = ~n1202 & n9484 ;
  assign n12610 = n5923 ^ n1401 ^ 1'b0 ;
  assign n12611 = n600 | n12610 ;
  assign n12612 = n4142 & n4818 ;
  assign n12613 = x13 & ~n1879 ;
  assign n12614 = ( ~n4550 & n12612 ) | ( ~n4550 & n12613 ) | ( n12612 & n12613 ) ;
  assign n12615 = n1620 & ~n3927 ;
  assign n12616 = n12615 ^ n2097 ^ 1'b0 ;
  assign n12617 = n4651 & n12616 ;
  assign n12618 = ~n4001 & n10761 ;
  assign n12619 = n12618 ^ n1937 ^ 1'b0 ;
  assign n12620 = n12619 ^ n3890 ^ 1'b0 ;
  assign n12621 = n1004 & n8821 ;
  assign n12622 = ~n2743 & n12621 ;
  assign n12626 = n6285 ^ n2839 ^ 1'b0 ;
  assign n12627 = ( n5279 & n6625 ) | ( n5279 & ~n12626 ) | ( n6625 & ~n12626 ) ;
  assign n12623 = x212 & n3551 ;
  assign n12624 = n12623 ^ n3218 ^ 1'b0 ;
  assign n12625 = ( x247 & n2849 ) | ( x247 & n12624 ) | ( n2849 & n12624 ) ;
  assign n12628 = n12627 ^ n12625 ^ 1'b0 ;
  assign n12629 = ~n9674 & n12628 ;
  assign n12630 = n8765 ^ n4761 ^ 1'b0 ;
  assign n12631 = n12630 ^ n1674 ^ 1'b0 ;
  assign n12632 = n657 & n3480 ;
  assign n12633 = ~x30 & n12632 ;
  assign n12634 = n12633 ^ n4912 ^ 1'b0 ;
  assign n12635 = n12631 & n12634 ;
  assign n12636 = n3326 & n12635 ;
  assign n12637 = n12636 ^ n8662 ^ 1'b0 ;
  assign n12638 = ~n5573 & n12637 ;
  assign n12646 = n5732 | n7887 ;
  assign n12647 = n7534 & ~n12646 ;
  assign n12639 = n984 & n3124 ;
  assign n12640 = n9977 ^ n9415 ^ x217 ;
  assign n12641 = n4021 ^ n2275 ^ 1'b0 ;
  assign n12642 = n4931 & n12641 ;
  assign n12643 = n12642 ^ n12624 ^ 1'b0 ;
  assign n12644 = n12640 & ~n12643 ;
  assign n12645 = ~n12639 & n12644 ;
  assign n12648 = n12647 ^ n12645 ^ 1'b0 ;
  assign n12649 = ~n1125 & n10319 ;
  assign n12650 = x252 & ~n585 ;
  assign n12651 = n5400 & n12650 ;
  assign n12652 = n3277 & ~n12651 ;
  assign n12653 = n12649 & n12652 ;
  assign n12654 = n3193 ^ n3071 ^ n2197 ;
  assign n12655 = n12654 ^ n6556 ^ n5264 ;
  assign n12656 = ( n1865 & ~n3145 ) | ( n1865 & n8642 ) | ( ~n3145 & n8642 ) ;
  assign n12657 = n5890 & n6686 ;
  assign n12658 = n10650 | n10897 ;
  assign n12659 = n12658 ^ n1415 ^ 1'b0 ;
  assign n12660 = n1152 & ~n7391 ;
  assign n12661 = n1625 ^ x78 ^ 1'b0 ;
  assign n12662 = n10543 ^ n5244 ^ n3398 ;
  assign n12663 = n4620 & n8024 ;
  assign n12664 = n706 | n12663 ;
  assign n12665 = n5676 | n12664 ;
  assign n12666 = n1707 & ~n2401 ;
  assign n12667 = n12666 ^ n7369 ^ 1'b0 ;
  assign n12668 = n399 & n12667 ;
  assign n12669 = n1233 ^ n432 ^ 1'b0 ;
  assign n12670 = n12669 ^ n3947 ^ 1'b0 ;
  assign n12671 = ~n5019 & n12670 ;
  assign n12672 = ~n5379 & n12671 ;
  assign n12673 = n1177 & n4388 ;
  assign n12674 = n3480 | n12673 ;
  assign n12675 = n2641 | n11889 ;
  assign n12676 = n12674 | n12675 ;
  assign n12677 = ~n1340 & n11158 ;
  assign n12678 = n4806 ^ n4020 ^ 1'b0 ;
  assign n12679 = n5376 ^ n4969 ^ n1064 ;
  assign n12680 = n9786 & n12679 ;
  assign n12681 = ( x233 & n3552 ) | ( x233 & ~n5277 ) | ( n3552 & ~n5277 ) ;
  assign n12682 = n12681 ^ n12571 ^ 1'b0 ;
  assign n12683 = ~n7007 & n12682 ;
  assign n12684 = n3515 | n11102 ;
  assign n12685 = n12684 ^ n1486 ^ 1'b0 ;
  assign n12686 = n5830 | n12685 ;
  assign n12687 = n12686 ^ n3804 ^ 1'b0 ;
  assign n12688 = n6732 | n11053 ;
  assign n12689 = n4300 & ~n11446 ;
  assign n12690 = n1168 | n7199 ;
  assign n12691 = n12169 ^ n11951 ^ 1'b0 ;
  assign n12692 = n1192 & n5977 ;
  assign n12693 = ( n3975 & n7423 ) | ( n3975 & ~n12692 ) | ( n7423 & ~n12692 ) ;
  assign n12694 = n6607 & ~n11504 ;
  assign n12695 = n4848 ^ n3090 ^ 1'b0 ;
  assign n12696 = n10405 | n12695 ;
  assign n12697 = n1404 ^ n1253 ^ 1'b0 ;
  assign n12698 = n10225 & n12697 ;
  assign n12699 = ~n2481 & n4562 ;
  assign n12700 = n12699 ^ n956 ^ n455 ;
  assign n12701 = n4231 ^ n3029 ^ 1'b0 ;
  assign n12702 = n3359 ^ n3142 ^ 1'b0 ;
  assign n12703 = n4312 | n12702 ;
  assign n12706 = n6798 ^ n6023 ^ 1'b0 ;
  assign n12707 = n4764 & n12706 ;
  assign n12708 = n12707 ^ n3283 ^ 1'b0 ;
  assign n12704 = n736 & ~n9862 ;
  assign n12705 = n12704 ^ x163 ^ 1'b0 ;
  assign n12709 = n12708 ^ n12705 ^ 1'b0 ;
  assign n12710 = n5763 ^ n1853 ^ 1'b0 ;
  assign n12711 = n1535 & n7925 ;
  assign n12712 = ~n6919 & n12483 ;
  assign n12713 = n11438 ^ n9795 ^ n7665 ;
  assign n12714 = n7632 ^ n4887 ^ n4070 ;
  assign n12715 = n12714 ^ n12163 ^ 1'b0 ;
  assign n12716 = n2359 ^ n666 ^ 1'b0 ;
  assign n12717 = n2377 & n12716 ;
  assign n12718 = n8953 ^ n6307 ^ n3788 ;
  assign n12719 = n12718 ^ n9292 ^ 1'b0 ;
  assign n12720 = n5397 & n12719 ;
  assign n12721 = ( n4493 & n10454 ) | ( n4493 & n11472 ) | ( n10454 & n11472 ) ;
  assign n12723 = n11859 ^ n5578 ^ 1'b0 ;
  assign n12722 = ( n8343 & ~n10592 ) | ( n8343 & n10607 ) | ( ~n10592 & n10607 ) ;
  assign n12724 = n12723 ^ n12722 ^ n10558 ;
  assign n12725 = n8190 ^ n1535 ^ 1'b0 ;
  assign n12726 = n12009 | n12725 ;
  assign n12727 = n12726 ^ n4931 ^ 1'b0 ;
  assign n12728 = n371 & n1072 ;
  assign n12729 = n12728 ^ n9244 ^ 1'b0 ;
  assign n12730 = ~n5094 & n12729 ;
  assign n12731 = n12727 & n12730 ;
  assign n12732 = n4652 ^ x41 ^ 1'b0 ;
  assign n12733 = n560 & ~n12732 ;
  assign n12736 = ~n1769 & n3781 ;
  assign n12737 = n8866 & n12736 ;
  assign n12738 = n2827 | n12737 ;
  assign n12739 = n12738 ^ n5449 ^ 1'b0 ;
  assign n12740 = n12739 ^ n10796 ^ 1'b0 ;
  assign n12734 = n9950 ^ n383 ^ 1'b0 ;
  assign n12735 = n1233 & n12734 ;
  assign n12741 = n12740 ^ n12735 ^ 1'b0 ;
  assign n12742 = ~n4611 & n4806 ;
  assign n12743 = n12742 ^ n7222 ^ 1'b0 ;
  assign n12744 = n5079 ^ n1102 ^ 1'b0 ;
  assign n12745 = ~n8465 & n12744 ;
  assign n12746 = n1840 | n9747 ;
  assign n12747 = n7802 ^ n4272 ^ n407 ;
  assign n12748 = n896 | n12747 ;
  assign n12749 = n9255 ^ n7923 ^ 1'b0 ;
  assign n12750 = ~n646 & n7013 ;
  assign n12751 = n9612 & n12750 ;
  assign n12752 = n12749 & n12751 ;
  assign n12753 = n2274 | n2519 ;
  assign n12754 = n11547 & ~n12753 ;
  assign n12755 = n2670 ^ n1630 ^ 1'b0 ;
  assign n12756 = n5137 & ~n12755 ;
  assign n12757 = n1658 ^ x28 ^ 1'b0 ;
  assign n12758 = n342 & ~n12757 ;
  assign n12759 = n12758 ^ n1122 ^ 1'b0 ;
  assign n12760 = n1739 & n12759 ;
  assign n12761 = ( n1728 & ~n4488 ) | ( n1728 & n12760 ) | ( ~n4488 & n12760 ) ;
  assign n12762 = n12756 & n12761 ;
  assign n12763 = n12346 & n12762 ;
  assign n12767 = n2064 ^ n1295 ^ 1'b0 ;
  assign n12764 = ~n1666 & n3008 ;
  assign n12765 = ~n11357 & n12764 ;
  assign n12766 = n514 | n12765 ;
  assign n12768 = n12767 ^ n12766 ^ 1'b0 ;
  assign n12769 = n3989 & n12768 ;
  assign n12770 = ~n989 & n2963 ;
  assign n12771 = ~n4651 & n12770 ;
  assign n12772 = ( ~n2509 & n7971 ) | ( ~n2509 & n12771 ) | ( n7971 & n12771 ) ;
  assign n12773 = ~n4852 & n8262 ;
  assign n12774 = n8522 ^ n1897 ^ 1'b0 ;
  assign n12775 = n12774 ^ n11521 ^ 1'b0 ;
  assign n12776 = ( n6964 & n8167 ) | ( n6964 & n11705 ) | ( n8167 & n11705 ) ;
  assign n12777 = n3524 & ~n4272 ;
  assign n12778 = ~n9880 & n12777 ;
  assign n12779 = n425 | n12778 ;
  assign n12780 = n12776 | n12779 ;
  assign n12781 = n4207 ^ n2870 ^ n826 ;
  assign n12782 = n4421 ^ n1136 ^ 1'b0 ;
  assign n12783 = ~n12781 & n12782 ;
  assign n12784 = n12783 ^ n10450 ^ 1'b0 ;
  assign n12785 = ~n2946 & n12784 ;
  assign n12786 = n1838 & ~n12785 ;
  assign n12787 = ~n2783 & n9861 ;
  assign n12788 = n4455 & n12787 ;
  assign n12789 = ~n7437 & n11906 ;
  assign n12790 = n12789 ^ n1719 ^ 1'b0 ;
  assign n12791 = n7033 & n12790 ;
  assign n12792 = ~n12788 & n12791 ;
  assign n12793 = n12792 ^ n8497 ^ 1'b0 ;
  assign n12795 = n8035 ^ n4796 ^ 1'b0 ;
  assign n12796 = n7587 & n12795 ;
  assign n12794 = n5683 ^ n3275 ^ n3066 ;
  assign n12797 = n12796 ^ n12794 ^ 1'b0 ;
  assign n12798 = n12793 | n12797 ;
  assign n12799 = n3360 & ~n10464 ;
  assign n12800 = ( n5098 & ~n6506 ) | ( n5098 & n6724 ) | ( ~n6506 & n6724 ) ;
  assign n12801 = n12800 ^ n3378 ^ 1'b0 ;
  assign n12802 = n4493 & n12801 ;
  assign n12803 = n3617 & n5288 ;
  assign n12804 = n12803 ^ n6403 ^ n3984 ;
  assign n12805 = n4135 ^ n599 ^ 1'b0 ;
  assign n12806 = n9976 & n12805 ;
  assign n12807 = n7667 ^ n3013 ^ 1'b0 ;
  assign n12808 = n11191 | n12807 ;
  assign n12809 = ( n704 & n8122 ) | ( n704 & ~n8465 ) | ( n8122 & ~n8465 ) ;
  assign n12810 = n1033 & ~n3947 ;
  assign n12811 = n8984 & ~n12810 ;
  assign n12812 = ~n8573 & n12811 ;
  assign n12813 = n10673 ^ n6164 ^ 1'b0 ;
  assign n12814 = n7723 & ~n12813 ;
  assign n12815 = n12814 ^ n10298 ^ 1'b0 ;
  assign n12816 = n558 | n11267 ;
  assign n12817 = n3106 & n5207 ;
  assign n12818 = n12817 ^ n2162 ^ 1'b0 ;
  assign n12819 = n12818 ^ n7349 ^ n7316 ;
  assign n12820 = n12819 ^ n9539 ^ 1'b0 ;
  assign n12826 = n5512 ^ n3885 ^ 1'b0 ;
  assign n12827 = n1166 & ~n12826 ;
  assign n12821 = n681 | n9221 ;
  assign n12822 = n9470 ^ n2774 ^ n2608 ;
  assign n12823 = n4448 & n12822 ;
  assign n12824 = ( n4638 & n12821 ) | ( n4638 & n12823 ) | ( n12821 & n12823 ) ;
  assign n12825 = n843 & ~n12824 ;
  assign n12828 = n12827 ^ n12825 ^ 1'b0 ;
  assign n12829 = n4833 ^ n1029 ^ 1'b0 ;
  assign n12830 = ~n2161 & n12829 ;
  assign n12831 = n3240 | n5608 ;
  assign n12832 = n12831 ^ n3413 ^ 1'b0 ;
  assign n12833 = n9925 ^ n8623 ^ 1'b0 ;
  assign n12834 = ~n5081 & n12833 ;
  assign n12835 = n11845 & ~n12834 ;
  assign n12836 = n2834 & n4677 ;
  assign n12837 = n9365 & n11105 ;
  assign n12838 = ~n6400 & n12837 ;
  assign n12839 = ~n11667 & n12838 ;
  assign n12840 = n12836 | n12839 ;
  assign n12841 = n7376 & ~n12840 ;
  assign n12842 = n3556 & n6365 ;
  assign n12843 = n12842 ^ n9367 ^ 1'b0 ;
  assign n12844 = n10629 ^ n4343 ^ 1'b0 ;
  assign n12845 = ~n719 & n12844 ;
  assign n12846 = n12845 ^ n648 ^ 1'b0 ;
  assign n12847 = ~n3431 & n9870 ;
  assign n12848 = n12847 ^ n8264 ^ 1'b0 ;
  assign n12849 = n4344 ^ n4236 ^ 1'b0 ;
  assign n12850 = n12848 & n12849 ;
  assign n12851 = n6663 | n12850 ;
  assign n12852 = n6611 & n8544 ;
  assign n12853 = n12852 ^ n1194 ^ 1'b0 ;
  assign n12854 = x244 & n4549 ;
  assign n12855 = n12853 & n12854 ;
  assign n12856 = n9330 ^ n6063 ^ 1'b0 ;
  assign n12857 = n7543 ^ n2341 ^ 1'b0 ;
  assign n12858 = n12856 & n12857 ;
  assign n12859 = n10897 ^ n1218 ^ 1'b0 ;
  assign n12860 = n12858 & ~n12859 ;
  assign n12861 = ~n2213 & n9535 ;
  assign n12862 = ~n7128 & n12861 ;
  assign n12863 = n1793 & ~n4030 ;
  assign n12864 = n12077 ^ n7260 ^ 1'b0 ;
  assign n12865 = n12864 ^ n6788 ^ 1'b0 ;
  assign n12866 = n4184 | n5840 ;
  assign n12867 = n5953 ^ n3352 ^ 1'b0 ;
  assign n12869 = n6857 ^ n2949 ^ n2509 ;
  assign n12868 = n3213 & n6584 ;
  assign n12870 = n12869 ^ n12868 ^ 1'b0 ;
  assign n12871 = ( n6758 & n12867 ) | ( n6758 & n12870 ) | ( n12867 & n12870 ) ;
  assign n12872 = n1378 | n12871 ;
  assign n12873 = n6921 | n12872 ;
  assign n12874 = n12873 ^ n5812 ^ n3467 ;
  assign n12875 = n4196 ^ n1957 ^ 1'b0 ;
  assign n12876 = n3245 & ~n12875 ;
  assign n12877 = ( n5048 & ~n6364 ) | ( n5048 & n12876 ) | ( ~n6364 & n12876 ) ;
  assign n12878 = ~n5188 & n9058 ;
  assign n12879 = ~n12877 & n12878 ;
  assign n12880 = ~n5782 & n11425 ;
  assign n12881 = ~n4604 & n12880 ;
  assign n12882 = n12881 ^ n11706 ^ n8102 ;
  assign n12883 = n3554 & n12882 ;
  assign n12884 = ~n697 & n12883 ;
  assign n12885 = n3261 | n7534 ;
  assign n12886 = ~n5535 & n12885 ;
  assign n12887 = ~n4086 & n12886 ;
  assign n12888 = n585 | n10284 ;
  assign n12889 = n3422 | n4583 ;
  assign n12890 = n8842 & ~n12889 ;
  assign n12891 = n6161 & ~n12890 ;
  assign n12892 = n12891 ^ n9586 ^ 1'b0 ;
  assign n12893 = ~n5369 & n9935 ;
  assign n12894 = ~n1622 & n12893 ;
  assign n12895 = n2543 | n12894 ;
  assign n12899 = n6027 ^ n2378 ^ 1'b0 ;
  assign n12896 = n4460 ^ n4455 ^ 1'b0 ;
  assign n12897 = ~n2942 & n12896 ;
  assign n12898 = ~n9365 & n12897 ;
  assign n12900 = n12899 ^ n12898 ^ 1'b0 ;
  assign n12901 = n3382 ^ n3287 ^ n3259 ;
  assign n12902 = ( n9490 & n12900 ) | ( n9490 & ~n12901 ) | ( n12900 & ~n12901 ) ;
  assign n12903 = ~n1105 & n5242 ;
  assign n12904 = n4463 | n5319 ;
  assign n12905 = n12903 | n12904 ;
  assign n12908 = n590 & ~n743 ;
  assign n12909 = n12908 ^ n12221 ^ 1'b0 ;
  assign n12906 = ( n1186 & n3599 ) | ( n1186 & n5052 ) | ( n3599 & n5052 ) ;
  assign n12907 = ( x82 & ~n1160 ) | ( x82 & n12906 ) | ( ~n1160 & n12906 ) ;
  assign n12910 = n12909 ^ n12907 ^ 1'b0 ;
  assign n12911 = n3981 & ~n5921 ;
  assign n12912 = ~n6063 & n12911 ;
  assign n12913 = n1525 & n5628 ;
  assign n12914 = n2197 & n12913 ;
  assign n12915 = ( n2404 & ~n12912 ) | ( n2404 & n12914 ) | ( ~n12912 & n12914 ) ;
  assign n12916 = n11175 | n12915 ;
  assign n12917 = n4923 ^ n4509 ^ n1197 ;
  assign n12918 = n10582 & ~n12917 ;
  assign n12920 = n3424 ^ n410 ^ 1'b0 ;
  assign n12921 = ~n8695 & n12920 ;
  assign n12922 = n12921 ^ n10658 ^ n1082 ;
  assign n12919 = n400 | n8029 ;
  assign n12923 = n12922 ^ n12919 ^ 1'b0 ;
  assign n12924 = n967 | n12923 ;
  assign n12925 = n8500 & ~n12924 ;
  assign n12926 = n6661 | n12925 ;
  assign n12927 = n7138 | n12926 ;
  assign n12931 = ~n2218 & n2351 ;
  assign n12932 = n4263 | n12931 ;
  assign n12929 = n8466 | n8519 ;
  assign n12928 = ~n798 & n3270 ;
  assign n12930 = n12929 ^ n12928 ^ 1'b0 ;
  assign n12933 = n12932 ^ n12930 ^ n7221 ;
  assign n12934 = n12805 ^ n11031 ^ n4195 ;
  assign n12935 = ~n1706 & n2066 ;
  assign n12936 = ~n8308 & n12935 ;
  assign n12937 = n2521 ^ n1365 ^ n1291 ;
  assign n12938 = n12937 ^ n4518 ^ 1'b0 ;
  assign n12939 = ~n1232 & n12938 ;
  assign n12940 = n12939 ^ n8057 ^ 1'b0 ;
  assign n12941 = n1491 & ~n2337 ;
  assign n12942 = n12941 ^ n1401 ^ 1'b0 ;
  assign n12943 = n5208 & n5707 ;
  assign n12944 = n12942 & n12943 ;
  assign n12945 = n3328 ^ n2337 ^ 1'b0 ;
  assign n12946 = n12945 ^ n6344 ^ n4827 ;
  assign n12947 = n4953 ^ n3671 ^ n2431 ;
  assign n12948 = ~n10818 & n12947 ;
  assign n12949 = n10926 & ~n12948 ;
  assign n12950 = n11090 & n12949 ;
  assign n12951 = x86 & ~n11212 ;
  assign n12952 = n12951 ^ n1102 ^ 1'b0 ;
  assign n12953 = n2266 & n7277 ;
  assign n12954 = n832 & ~n12953 ;
  assign n12955 = n4907 & n12954 ;
  assign n12956 = n7161 ^ n4223 ^ n4120 ;
  assign n12957 = ( x196 & n4746 ) | ( x196 & n12956 ) | ( n4746 & n12956 ) ;
  assign n12958 = n6085 & n12957 ;
  assign n12959 = n3600 | n7097 ;
  assign n12960 = n12739 ^ n10363 ^ 1'b0 ;
  assign n12961 = n8194 & ~n12960 ;
  assign n12962 = n3992 & ~n7408 ;
  assign n12963 = ~n8351 & n12962 ;
  assign n12964 = n5802 & ~n6049 ;
  assign n12965 = n12964 ^ n7923 ^ 1'b0 ;
  assign n12966 = ~n1058 & n7823 ;
  assign n12967 = n7587 & ~n12966 ;
  assign n12968 = n3975 & n12967 ;
  assign n12969 = n12965 & ~n12968 ;
  assign n12970 = ~n5264 & n12969 ;
  assign n12971 = ( ~n538 & n946 ) | ( ~n538 & n7429 ) | ( n946 & n7429 ) ;
  assign n12972 = n9141 | n12562 ;
  assign n12973 = n4087 | n12972 ;
  assign n12974 = n5846 ^ n4684 ^ 1'b0 ;
  assign n12975 = n12600 & n12974 ;
  assign n12976 = n7127 & n12975 ;
  assign n12977 = n5071 & n5939 ;
  assign n12978 = n4455 ^ n1949 ^ 1'b0 ;
  assign n12979 = ~n12603 & n12978 ;
  assign n12981 = n6761 ^ n3005 ^ n1934 ;
  assign n12980 = n4565 ^ n4407 ^ n3728 ;
  assign n12982 = n12981 ^ n12980 ^ 1'b0 ;
  assign n12983 = n12979 & n12982 ;
  assign n12984 = n1671 | n4686 ;
  assign n12985 = n12984 ^ n4289 ^ 1'b0 ;
  assign n12986 = n9515 & n12985 ;
  assign n12987 = n12986 ^ n11442 ^ n5597 ;
  assign n12988 = n12987 ^ n4126 ^ 1'b0 ;
  assign n12989 = n4279 & ~n12988 ;
  assign n12990 = n12989 ^ n8152 ^ 1'b0 ;
  assign n12991 = ~n984 & n7844 ;
  assign n12992 = n1535 & ~n6327 ;
  assign n12993 = ~n9212 & n12992 ;
  assign n12994 = ~n6795 & n9720 ;
  assign n12996 = n3023 & ~n11975 ;
  assign n12997 = n6298 & n12996 ;
  assign n12995 = n1265 & ~n2853 ;
  assign n12998 = n12997 ^ n12995 ^ 1'b0 ;
  assign n12999 = n2076 | n2084 ;
  assign n13000 = n12999 ^ n4984 ^ 1'b0 ;
  assign n13001 = n3641 ^ n2057 ^ 1'b0 ;
  assign n13002 = n1500 & n13001 ;
  assign n13003 = ~n1246 & n13002 ;
  assign n13004 = n13000 & n13003 ;
  assign n13005 = ~n6409 & n12539 ;
  assign n13006 = n2548 & n13005 ;
  assign n13007 = ( n2746 & n9724 ) | ( n2746 & n13006 ) | ( n9724 & n13006 ) ;
  assign n13010 = n3077 ^ n1657 ^ n1010 ;
  assign n13008 = n4276 ^ n3272 ^ n2791 ;
  assign n13009 = n12347 | n13008 ;
  assign n13011 = n13010 ^ n13009 ^ 1'b0 ;
  assign n13012 = n11219 ^ n880 ^ 1'b0 ;
  assign n13013 = ~n6227 & n12606 ;
  assign n13014 = n8077 ^ n6891 ^ 1'b0 ;
  assign n13015 = ~n13013 & n13014 ;
  assign n13016 = n342 & ~n9716 ;
  assign n13017 = n13016 ^ n451 ^ 1'b0 ;
  assign n13018 = n3441 & ~n13017 ;
  assign n13019 = n13018 ^ n5807 ^ 1'b0 ;
  assign n13020 = ( n458 & n4328 ) | ( n458 & ~n13019 ) | ( n4328 & ~n13019 ) ;
  assign n13021 = ( n1186 & n1889 ) | ( n1186 & ~n2513 ) | ( n1889 & ~n2513 ) ;
  assign n13022 = n13021 ^ n1685 ^ 1'b0 ;
  assign n13023 = n5660 & n13022 ;
  assign n13024 = ~n5357 & n13023 ;
  assign n13025 = n13020 & ~n13024 ;
  assign n13026 = n13025 ^ n3769 ^ 1'b0 ;
  assign n13027 = n4501 & n7369 ;
  assign n13028 = ~n4366 & n13027 ;
  assign n13029 = n1108 & n10548 ;
  assign n13030 = n13029 ^ n1372 ^ 1'b0 ;
  assign n13031 = ( n3236 & ~n5853 ) | ( n3236 & n13030 ) | ( ~n5853 & n13030 ) ;
  assign n13032 = n8663 | n13031 ;
  assign n13033 = n13032 ^ n12456 ^ 1'b0 ;
  assign n13036 = n2455 | n8290 ;
  assign n13034 = n4797 & ~n8306 ;
  assign n13035 = ~n1403 & n13034 ;
  assign n13037 = n13036 ^ n13035 ^ 1'b0 ;
  assign n13038 = n4267 ^ x151 ^ 1'b0 ;
  assign n13039 = n6751 | n13038 ;
  assign n13040 = n13039 ^ n5729 ^ 1'b0 ;
  assign n13041 = n13023 ^ n3975 ^ n1253 ;
  assign n13042 = n908 | n13041 ;
  assign n13043 = n13040 & ~n13042 ;
  assign n13044 = ( n6259 & n12170 ) | ( n6259 & ~n13043 ) | ( n12170 & ~n13043 ) ;
  assign n13045 = n2151 & n3942 ;
  assign n13046 = n13045 ^ n327 ^ 1'b0 ;
  assign n13047 = n601 & ~n2337 ;
  assign n13048 = ~n538 & n13047 ;
  assign n13049 = n13046 | n13048 ;
  assign n13050 = n9793 | n13049 ;
  assign n13051 = ( n4109 & ~n5070 ) | ( n4109 & n9456 ) | ( ~n5070 & n9456 ) ;
  assign n13052 = n13051 ^ n2368 ^ 1'b0 ;
  assign n13053 = ~n10820 & n13052 ;
  assign n13054 = n768 | n5397 ;
  assign n13055 = ~n7278 & n13054 ;
  assign n13056 = ~n4731 & n12894 ;
  assign n13057 = ~n4749 & n10447 ;
  assign n13058 = n7063 ^ n5296 ^ 1'b0 ;
  assign n13059 = n1272 | n13058 ;
  assign n13060 = n5502 & ~n13059 ;
  assign n13061 = ~n3149 & n13060 ;
  assign n13062 = n1306 | n5261 ;
  assign n13063 = n13062 ^ n5708 ^ 1'b0 ;
  assign n13064 = n13063 ^ n9108 ^ n8235 ;
  assign n13071 = n3516 ^ n3435 ^ 1'b0 ;
  assign n13072 = n1604 | n13071 ;
  assign n13073 = n3651 | n13072 ;
  assign n13074 = n13073 ^ n3664 ^ 1'b0 ;
  assign n13070 = n2560 ^ n2418 ^ 1'b0 ;
  assign n13065 = n1604 | n9206 ;
  assign n13066 = n5057 & ~n13065 ;
  assign n13067 = n2091 & n4900 ;
  assign n13068 = n13066 & n13067 ;
  assign n13069 = n5248 & ~n13068 ;
  assign n13075 = n13074 ^ n13070 ^ n13069 ;
  assign n13076 = n5731 ^ n4910 ^ 1'b0 ;
  assign n13077 = ~n7460 & n13076 ;
  assign n13078 = n13077 ^ n8839 ^ 1'b0 ;
  assign n13079 = ~n4001 & n13078 ;
  assign n13080 = n12184 ^ n8287 ^ 1'b0 ;
  assign n13081 = n2141 & ~n6397 ;
  assign n13082 = n5710 ^ n4580 ^ 1'b0 ;
  assign n13083 = n13081 & n13082 ;
  assign n13087 = n1195 & n4996 ;
  assign n13088 = n13087 ^ n4404 ^ 1'b0 ;
  assign n13084 = n10076 ^ n6428 ^ 1'b0 ;
  assign n13085 = n5426 | n13084 ;
  assign n13086 = n13085 ^ n8503 ^ 1'b0 ;
  assign n13089 = n13088 ^ n13086 ^ 1'b0 ;
  assign n13090 = n13083 & ~n13089 ;
  assign n13091 = n5879 ^ n5493 ^ 1'b0 ;
  assign n13092 = n6036 & ~n13091 ;
  assign n13093 = n13092 ^ n535 ^ 1'b0 ;
  assign n13094 = n6330 & n13093 ;
  assign n13095 = ~n418 & n1902 ;
  assign n13096 = n5841 ^ n417 ^ 1'b0 ;
  assign n13100 = n2225 & ~n3523 ;
  assign n13101 = n3523 & n13100 ;
  assign n13102 = x27 & ~n6246 ;
  assign n13103 = n593 & n13102 ;
  assign n13104 = n1286 & ~n13103 ;
  assign n13105 = n13101 & n13104 ;
  assign n13097 = x22 | n2910 ;
  assign n13098 = x22 & ~n13097 ;
  assign n13099 = n7743 & ~n13098 ;
  assign n13106 = n13105 ^ n13099 ^ 1'b0 ;
  assign n13107 = ~n3055 & n4240 ;
  assign n13108 = n3055 & n13107 ;
  assign n13109 = n3523 | n13108 ;
  assign n13110 = n5166 & ~n11400 ;
  assign n13111 = ~n5166 & n13110 ;
  assign n13112 = n13109 | n13111 ;
  assign n13113 = n13106 | n13112 ;
  assign n13114 = n3456 & ~n5477 ;
  assign n13115 = ( n3750 & n7264 ) | ( n3750 & ~n10949 ) | ( n7264 & ~n10949 ) ;
  assign n13116 = ~n2278 & n13115 ;
  assign n13117 = ~n4544 & n11904 ;
  assign n13118 = n908 | n3651 ;
  assign n13119 = n9247 & ~n13118 ;
  assign n13120 = n10863 ^ n5014 ^ 1'b0 ;
  assign n13121 = n13120 ^ n8914 ^ 1'b0 ;
  assign n13122 = n6035 | n7955 ;
  assign n13123 = n5648 | n13122 ;
  assign n13124 = n2577 | n5027 ;
  assign n13125 = n13124 ^ n11771 ^ 1'b0 ;
  assign n13127 = ( x250 & n1455 ) | ( x250 & n12118 ) | ( n1455 & n12118 ) ;
  assign n13126 = ~n5742 & n8109 ;
  assign n13128 = n13127 ^ n13126 ^ n8183 ;
  assign n13130 = n2358 ^ n1025 ^ 1'b0 ;
  assign n13131 = n2979 & ~n13130 ;
  assign n13129 = n3548 & ~n5977 ;
  assign n13132 = n13131 ^ n13129 ^ 1'b0 ;
  assign n13133 = n3456 & n4996 ;
  assign n13134 = n13132 & n13133 ;
  assign n13135 = n3220 ^ n1406 ^ 1'b0 ;
  assign n13136 = n3975 | n9213 ;
  assign n13137 = ( n512 & ~n3405 ) | ( n512 & n11080 ) | ( ~n3405 & n11080 ) ;
  assign n13138 = n8154 & ~n13137 ;
  assign n13139 = ~n13136 & n13138 ;
  assign n13140 = n2093 ^ n1752 ^ 1'b0 ;
  assign n13141 = n13140 ^ n5408 ^ 1'b0 ;
  assign n13142 = n7789 ^ n3234 ^ n2914 ;
  assign n13143 = n12832 & n13142 ;
  assign n13144 = n13141 & n13143 ;
  assign n13145 = n5074 | n7225 ;
  assign n13146 = ( n790 & ~n2376 ) | ( n790 & n13145 ) | ( ~n2376 & n13145 ) ;
  assign n13147 = n3094 ^ n1239 ^ 1'b0 ;
  assign n13148 = n1806 | n13147 ;
  assign n13149 = n1800 | n13148 ;
  assign n13150 = n12668 & ~n13149 ;
  assign n13151 = n1865 & n13150 ;
  assign n13152 = n2054 | n4211 ;
  assign n13153 = n13152 ^ n6389 ^ 1'b0 ;
  assign n13154 = n13153 ^ x243 ^ 1'b0 ;
  assign n13155 = ~n4352 & n13154 ;
  assign n13156 = x183 & ~n4768 ;
  assign n13157 = ~n822 & n9117 ;
  assign n13158 = n13157 ^ n4970 ^ 1'b0 ;
  assign n13159 = n1993 | n13158 ;
  assign n13160 = n13156 | n13159 ;
  assign n13161 = n3550 & ~n9775 ;
  assign n13164 = n4189 ^ n2226 ^ x2 ;
  assign n13162 = n6112 ^ n5934 ^ 1'b0 ;
  assign n13163 = n11466 | n13162 ;
  assign n13165 = n13164 ^ n13163 ^ 1'b0 ;
  assign n13166 = n6131 ^ n4036 ^ 1'b0 ;
  assign n13167 = n12047 | n13166 ;
  assign n13168 = n13165 & ~n13167 ;
  assign n13169 = ~n13161 & n13168 ;
  assign n13170 = n4415 ^ n2399 ^ 1'b0 ;
  assign n13171 = n2085 & ~n13170 ;
  assign n13172 = n13171 ^ n11175 ^ 1'b0 ;
  assign n13173 = n1877 | n2261 ;
  assign n13174 = n3286 & ~n13173 ;
  assign n13175 = n4626 | n12024 ;
  assign n13176 = ( ~n411 & n3598 ) | ( ~n411 & n11930 ) | ( n3598 & n11930 ) ;
  assign n13177 = n9941 ^ n8039 ^ 1'b0 ;
  assign n13178 = n13177 ^ n698 ^ 1'b0 ;
  assign n13179 = n322 | n13178 ;
  assign n13180 = n13179 ^ n4915 ^ 1'b0 ;
  assign n13181 = n2574 & n13180 ;
  assign n13182 = n12800 ^ n12452 ^ n6096 ;
  assign n13183 = ( x222 & n740 ) | ( x222 & n1724 ) | ( n740 & n1724 ) ;
  assign n13184 = n2146 & n13183 ;
  assign n13185 = n13184 ^ n1346 ^ 1'b0 ;
  assign n13186 = n7474 & ~n12639 ;
  assign n13187 = n13186 ^ n5870 ^ 1'b0 ;
  assign n13188 = n8927 & n13187 ;
  assign n13189 = ~n1060 & n8675 ;
  assign n13190 = n13189 ^ n3794 ^ 1'b0 ;
  assign n13191 = n13190 ^ n5850 ^ 1'b0 ;
  assign n13192 = n8026 ^ n2376 ^ n790 ;
  assign n13193 = ~n428 & n5313 ;
  assign n13194 = n1453 & n13193 ;
  assign n13195 = n2527 | n13194 ;
  assign n13196 = ( n7723 & n11457 ) | ( n7723 & ~n13195 ) | ( n11457 & ~n13195 ) ;
  assign n13197 = n11376 | n13196 ;
  assign n13198 = n13197 ^ n11930 ^ n2384 ;
  assign n13199 = n5980 & n10628 ;
  assign n13200 = n659 & ~n11227 ;
  assign n13201 = n972 | n13200 ;
  assign n13202 = n13201 ^ n6947 ^ 1'b0 ;
  assign n13203 = ~n2008 & n6463 ;
  assign n13204 = ~n1685 & n6798 ;
  assign n13205 = n12733 ^ n11152 ^ 1'b0 ;
  assign n13206 = n6921 & ~n13205 ;
  assign n13207 = n1587 & ~n1930 ;
  assign n13208 = n723 | n6152 ;
  assign n13209 = n3059 & ~n13208 ;
  assign n13210 = n7509 ^ n2556 ^ 1'b0 ;
  assign n13211 = n13209 | n13210 ;
  assign n13212 = n11915 ^ n7164 ^ 1'b0 ;
  assign n13213 = n997 & n13212 ;
  assign n13214 = ~n5306 & n13213 ;
  assign n13215 = ~n3363 & n7444 ;
  assign n13216 = n2836 & ~n6204 ;
  assign n13217 = ~n924 & n13216 ;
  assign n13218 = ( n1127 & n3481 ) | ( n1127 & ~n11872 ) | ( n3481 & ~n11872 ) ;
  assign n13219 = n12753 ^ n3481 ^ 1'b0 ;
  assign n13220 = n9205 & ~n13219 ;
  assign n13221 = n13220 ^ n11361 ^ 1'b0 ;
  assign n13222 = n1145 & n8299 ;
  assign n13223 = ~n5795 & n13222 ;
  assign n13224 = n3380 | n8026 ;
  assign n13225 = n13223 & ~n13224 ;
  assign n13226 = n6543 & ~n11742 ;
  assign n13227 = ~n1690 & n13226 ;
  assign n13228 = n1349 & ~n4310 ;
  assign n13229 = n13228 ^ n1285 ^ 1'b0 ;
  assign n13230 = n3030 ^ n2055 ^ 1'b0 ;
  assign n13231 = n13230 ^ n1960 ^ 1'b0 ;
  assign n13232 = ( n1177 & ~n10935 ) | ( n1177 & n13231 ) | ( ~n10935 & n13231 ) ;
  assign n13233 = n13229 & n13232 ;
  assign n13234 = ~n4651 & n13233 ;
  assign n13235 = n1943 & ~n4043 ;
  assign n13236 = n1444 & n5550 ;
  assign n13237 = n6988 ^ n4086 ^ n2711 ;
  assign n13238 = ( ~n2793 & n4828 ) | ( ~n2793 & n10501 ) | ( n4828 & n10501 ) ;
  assign n13239 = n8747 ^ n646 ^ x156 ;
  assign n13240 = n11599 ^ n5423 ^ n984 ;
  assign n13241 = n13240 ^ n3172 ^ 1'b0 ;
  assign n13242 = n2203 & n13241 ;
  assign n13243 = n6622 ^ n4876 ^ 1'b0 ;
  assign n13244 = ( ~n13239 & n13242 ) | ( ~n13239 & n13243 ) | ( n13242 & n13243 ) ;
  assign n13245 = ~n4385 & n6496 ;
  assign n13246 = n3904 | n13245 ;
  assign n13247 = n9862 & ~n13246 ;
  assign n13248 = n1173 & n13247 ;
  assign n13249 = n13248 ^ n8458 ^ x114 ;
  assign n13250 = n1064 | n10023 ;
  assign n13251 = n9566 & ~n13250 ;
  assign n13252 = ( n2686 & n10558 ) | ( n2686 & n13251 ) | ( n10558 & n13251 ) ;
  assign n13253 = ( n423 & n4002 ) | ( n423 & n13252 ) | ( n4002 & n13252 ) ;
  assign n13254 = n1358 & ~n12195 ;
  assign n13255 = n13141 ^ n8336 ^ 1'b0 ;
  assign n13256 = n9200 ^ n4158 ^ n1192 ;
  assign n13257 = n13256 ^ n11901 ^ 1'b0 ;
  assign n13258 = n2676 & ~n9175 ;
  assign n13259 = ~n4300 & n13258 ;
  assign n13260 = n13259 ^ n2395 ^ 1'b0 ;
  assign n13261 = n13260 ^ n1899 ^ 1'b0 ;
  assign n13262 = n9112 & n13261 ;
  assign n13263 = n7386 ^ n1073 ^ 1'b0 ;
  assign n13264 = n13263 ^ n6704 ^ n6544 ;
  assign n13265 = ( n8137 & n8752 ) | ( n8137 & n10089 ) | ( n8752 & n10089 ) ;
  assign n13266 = n1589 | n1744 ;
  assign n13267 = n5511 & ~n13266 ;
  assign n13268 = ~x189 & n13267 ;
  assign n13269 = n3375 ^ n1225 ^ 1'b0 ;
  assign n13270 = n538 & ~n13269 ;
  assign n13271 = n13270 ^ n2509 ^ 1'b0 ;
  assign n13272 = n1130 & ~n1631 ;
  assign n13273 = n13272 ^ n6079 ^ 1'b0 ;
  assign n13274 = n6730 & ~n13273 ;
  assign n13275 = n10203 ^ n9192 ^ 1'b0 ;
  assign n13276 = n9033 & ~n13275 ;
  assign n13277 = n4383 ^ n1698 ^ n1279 ;
  assign n13278 = n7630 & n13277 ;
  assign n13279 = n5033 | n10071 ;
  assign n13280 = n10840 ^ n1234 ^ n1151 ;
  assign n13281 = n13279 & n13280 ;
  assign n13282 = ( n1712 & n3296 ) | ( n1712 & ~n13281 ) | ( n3296 & ~n13281 ) ;
  assign n13283 = n1708 | n3019 ;
  assign n13284 = n11743 | n13283 ;
  assign n13285 = n13284 ^ n7213 ^ 1'b0 ;
  assign n13286 = n5006 & n13285 ;
  assign n13287 = n1808 & n9614 ;
  assign n13288 = ~n11389 & n13287 ;
  assign n13289 = n13288 ^ x183 ^ 1'b0 ;
  assign n13290 = n1680 | n7948 ;
  assign n13291 = n12223 & n13290 ;
  assign n13292 = ( ~n768 & n6403 ) | ( ~n768 & n12061 ) | ( n6403 & n12061 ) ;
  assign n13293 = n5211 ^ n694 ^ 1'b0 ;
  assign n13294 = n4160 & ~n13293 ;
  assign n13295 = n3953 & n13294 ;
  assign n13296 = n13295 ^ n5022 ^ 1'b0 ;
  assign n13297 = n8997 ^ n601 ^ 1'b0 ;
  assign n13298 = ~n3683 & n13297 ;
  assign n13299 = n13298 ^ n3695 ^ 1'b0 ;
  assign n13301 = n1374 & ~n5067 ;
  assign n13302 = n13301 ^ n952 ^ 1'b0 ;
  assign n13300 = ~n5188 & n6443 ;
  assign n13303 = n13302 ^ n13300 ^ 1'b0 ;
  assign n13304 = ~n7746 & n11425 ;
  assign n13305 = n13303 & n13304 ;
  assign n13306 = n1885 | n9279 ;
  assign n13307 = n13305 & ~n13306 ;
  assign n13308 = ( ~x208 & n3112 ) | ( ~x208 & n8313 ) | ( n3112 & n8313 ) ;
  assign n13309 = ( n981 & n5445 ) | ( n981 & ~n13308 ) | ( n5445 & ~n13308 ) ;
  assign n13310 = n13309 ^ n7834 ^ 1'b0 ;
  assign n13311 = n890 & n13310 ;
  assign n13312 = n13311 ^ n6553 ^ 1'b0 ;
  assign n13313 = n9459 & ~n13312 ;
  assign n13314 = n8280 ^ n402 ^ 1'b0 ;
  assign n13315 = n3815 | n3833 ;
  assign n13316 = n5656 & ~n13315 ;
  assign n13317 = n6760 | n7714 ;
  assign n13318 = n13317 ^ n5259 ^ 1'b0 ;
  assign n13319 = n13316 | n13318 ;
  assign n13320 = n9198 ^ n8071 ^ 1'b0 ;
  assign n13321 = ~n7809 & n12681 ;
  assign n13322 = n12130 ^ n6197 ^ 1'b0 ;
  assign n13323 = n9548 ^ n8161 ^ 1'b0 ;
  assign n13324 = ~n13322 & n13323 ;
  assign n13325 = ~n13321 & n13324 ;
  assign n13326 = ~n5809 & n11072 ;
  assign n13327 = n3852 & n13326 ;
  assign n13328 = ( ~n2765 & n4049 ) | ( ~n2765 & n10311 ) | ( n4049 & n10311 ) ;
  assign n13329 = n8398 & n10969 ;
  assign n13330 = ~n451 & n13329 ;
  assign n13331 = n13330 ^ n8173 ^ 1'b0 ;
  assign n13332 = n13328 | n13331 ;
  assign n13333 = n1236 ^ n1164 ^ n258 ;
  assign n13334 = n2711 | n11431 ;
  assign n13335 = n13333 & n13334 ;
  assign n13336 = n13335 ^ n4339 ^ 1'b0 ;
  assign n13337 = n13336 ^ n12653 ^ 1'b0 ;
  assign n13338 = n10744 & n13337 ;
  assign n13339 = n13338 ^ n12429 ^ n9589 ;
  assign n13340 = n6588 & ~n9618 ;
  assign n13341 = n8513 & ~n9261 ;
  assign n13342 = n13341 ^ n7554 ^ 1'b0 ;
  assign n13343 = n5514 ^ n3594 ^ n1803 ;
  assign n13344 = n11668 | n13343 ;
  assign n13346 = n791 & n2503 ;
  assign n13347 = n13346 ^ n513 ^ 1'b0 ;
  assign n13348 = n6669 | n13347 ;
  assign n13349 = n13348 ^ n404 ^ 1'b0 ;
  assign n13350 = ( n3659 & n6069 ) | ( n3659 & ~n13349 ) | ( n6069 & ~n13349 ) ;
  assign n13345 = n1188 | n1419 ;
  assign n13351 = n13350 ^ n13345 ^ 1'b0 ;
  assign n13352 = ~n1073 & n11521 ;
  assign n13353 = n13352 ^ n10279 ^ 1'b0 ;
  assign n13354 = ( n9468 & n10551 ) | ( n9468 & n11764 ) | ( n10551 & n11764 ) ;
  assign n13356 = n10141 ^ n7963 ^ 1'b0 ;
  assign n13357 = n13356 ^ n4688 ^ 1'b0 ;
  assign n13355 = n760 | n7567 ;
  assign n13358 = n13357 ^ n13355 ^ 1'b0 ;
  assign n13359 = ~n5094 & n13358 ;
  assign n13360 = n909 & ~n13088 ;
  assign n13361 = ~n4232 & n4792 ;
  assign n13362 = n13361 ^ n3407 ^ 1'b0 ;
  assign n13363 = n1785 | n13362 ;
  assign n13364 = n3773 & ~n13363 ;
  assign n13365 = ~n10187 & n13364 ;
  assign n13366 = n13365 ^ n7206 ^ 1'b0 ;
  assign n13367 = n13360 | n13366 ;
  assign n13368 = n2819 & ~n6722 ;
  assign n13369 = ~n7535 & n13368 ;
  assign n13370 = n13369 ^ n4597 ^ 1'b0 ;
  assign n13371 = n1427 & n13370 ;
  assign n13372 = ( n4433 & n4870 ) | ( n4433 & ~n6651 ) | ( n4870 & ~n6651 ) ;
  assign n13373 = ( n574 & n2182 ) | ( n574 & n5989 ) | ( n2182 & n5989 ) ;
  assign n13374 = n5398 ^ n3825 ^ 1'b0 ;
  assign n13375 = n13373 | n13374 ;
  assign n13376 = n2325 ^ x209 ^ 1'b0 ;
  assign n13377 = ~n753 & n13376 ;
  assign n13378 = ( n5603 & n6723 ) | ( n5603 & ~n13377 ) | ( n6723 & ~n13377 ) ;
  assign n13379 = n3195 | n5116 ;
  assign n13380 = n10503 | n13379 ;
  assign n13381 = n13380 ^ n11127 ^ 1'b0 ;
  assign n13382 = n5302 | n8747 ;
  assign n13383 = x222 & ~n3625 ;
  assign n13384 = n5019 ^ n2854 ^ 1'b0 ;
  assign n13385 = n13383 & ~n13384 ;
  assign n13386 = ~n13382 & n13385 ;
  assign n13387 = n5672 | n13386 ;
  assign n13388 = n13387 ^ n4668 ^ 1'b0 ;
  assign n13389 = n8555 ^ n2765 ^ 1'b0 ;
  assign n13390 = n13388 | n13389 ;
  assign n13391 = n6272 & n8785 ;
  assign n13392 = n9551 ^ n7000 ^ 1'b0 ;
  assign n13393 = ( n1847 & ~n8737 ) | ( n1847 & n13392 ) | ( ~n8737 & n13392 ) ;
  assign n13394 = ( ~n6383 & n13391 ) | ( ~n6383 & n13393 ) | ( n13391 & n13393 ) ;
  assign n13395 = n11993 ^ n3422 ^ 1'b0 ;
  assign n13396 = n8558 | n13395 ;
  assign n13397 = n8058 & ~n8694 ;
  assign n13399 = ~n1803 & n3608 ;
  assign n13398 = ~n2721 & n3556 ;
  assign n13400 = n13399 ^ n13398 ^ 1'b0 ;
  assign n13401 = n13400 ^ n12620 ^ 1'b0 ;
  assign n13402 = n5094 | n13401 ;
  assign n13403 = n2181 & ~n4042 ;
  assign n13404 = ~n5572 & n13403 ;
  assign n13405 = n617 | n7063 ;
  assign n13406 = n13404 & ~n13405 ;
  assign n13407 = n13406 ^ n9895 ^ n1987 ;
  assign n13408 = n326 & n6003 ;
  assign n13409 = n706 | n7552 ;
  assign n13410 = n12856 ^ n7846 ^ 1'b0 ;
  assign n13411 = n11396 | n13410 ;
  assign n13412 = n8754 ^ n3738 ^ 1'b0 ;
  assign n13413 = n10127 | n13412 ;
  assign n13414 = ~n2212 & n5643 ;
  assign n13415 = n8912 & n13414 ;
  assign n13416 = n8717 ^ n6392 ^ 1'b0 ;
  assign n13417 = n3148 & ~n5620 ;
  assign n13418 = n13416 & n13417 ;
  assign n13419 = ~n683 & n4137 ;
  assign n13420 = n1129 | n3671 ;
  assign n13421 = n13419 | n13420 ;
  assign n13427 = x200 & ~n2340 ;
  assign n13428 = n2340 & n13427 ;
  assign n13429 = n3598 & ~n13428 ;
  assign n13430 = ~n3598 & n13429 ;
  assign n13431 = n13430 ^ n2539 ^ 1'b0 ;
  assign n13432 = n9222 & ~n13431 ;
  assign n13422 = n4891 ^ n3747 ^ 1'b0 ;
  assign n13423 = ~n9375 & n13422 ;
  assign n13424 = n1199 | n13423 ;
  assign n13425 = n11728 & ~n13424 ;
  assign n13426 = n13425 ^ n11167 ^ 1'b0 ;
  assign n13433 = n13432 ^ n13426 ^ 1'b0 ;
  assign n13434 = n6031 ^ n4881 ^ 1'b0 ;
  assign n13435 = n4375 & n13434 ;
  assign n13436 = ( x63 & ~n6907 ) | ( x63 & n9639 ) | ( ~n6907 & n9639 ) ;
  assign n13437 = n13435 & ~n13436 ;
  assign n13438 = n5055 & ~n6831 ;
  assign n13439 = ~n13437 & n13438 ;
  assign n13440 = x15 & ~n12915 ;
  assign n13441 = n4018 & ~n13440 ;
  assign n13442 = n5341 ^ n1910 ^ x232 ;
  assign n13443 = n13442 ^ n2794 ^ 1'b0 ;
  assign n13444 = n13441 & ~n13443 ;
  assign n13445 = n13444 ^ n2105 ^ 1'b0 ;
  assign n13446 = n3720 & ~n5060 ;
  assign n13447 = n13446 ^ n8691 ^ n1411 ;
  assign n13448 = n8837 ^ x252 ^ 1'b0 ;
  assign n13449 = n3245 & n13448 ;
  assign n13450 = n13449 ^ n785 ^ 1'b0 ;
  assign n13451 = n5762 | n8689 ;
  assign n13452 = n13451 ^ n5006 ^ 1'b0 ;
  assign n13453 = n13452 ^ n3363 ^ x145 ;
  assign n13454 = ( ~n6500 & n13450 ) | ( ~n6500 & n13453 ) | ( n13450 & n13453 ) ;
  assign n13459 = ~n5216 & n6317 ;
  assign n13460 = n13459 ^ n4926 ^ 1'b0 ;
  assign n13455 = n10070 ^ n8471 ^ 1'b0 ;
  assign n13456 = ~n5327 & n13455 ;
  assign n13457 = n1486 & n13456 ;
  assign n13458 = n13457 ^ n3523 ^ 1'b0 ;
  assign n13461 = n13460 ^ n13458 ^ 1'b0 ;
  assign n13462 = x225 & n13461 ;
  assign n13463 = n513 & ~n7703 ;
  assign n13464 = ~n9964 & n13463 ;
  assign n13465 = n3317 & ~n13464 ;
  assign n13466 = ~n9466 & n13465 ;
  assign n13467 = n7643 ^ n7431 ^ n7028 ;
  assign n13468 = n4410 ^ n3003 ^ 1'b0 ;
  assign n13469 = n13468 ^ n4496 ^ n1024 ;
  assign n13470 = n13469 ^ n10655 ^ 1'b0 ;
  assign n13471 = n13467 & ~n13470 ;
  assign n13472 = n5621 ^ n3617 ^ 1'b0 ;
  assign n13473 = ~n488 & n13472 ;
  assign n13474 = n13473 ^ n6023 ^ 1'b0 ;
  assign n13475 = n809 | n10582 ;
  assign n13476 = n13475 ^ x19 ^ 1'b0 ;
  assign n13477 = n4470 | n13476 ;
  assign n13478 = n8861 ^ n3007 ^ 1'b0 ;
  assign n13479 = n4506 | n13478 ;
  assign n13480 = n12021 ^ n8917 ^ 1'b0 ;
  assign n13481 = n13480 ^ n5175 ^ 1'b0 ;
  assign n13482 = n8310 & ~n13481 ;
  assign n13483 = n3543 | n10689 ;
  assign n13484 = n13483 ^ n4901 ^ 1'b0 ;
  assign n13485 = n7177 ^ n1377 ^ 1'b0 ;
  assign n13486 = n7137 & n13485 ;
  assign n13487 = ( ~n6000 & n9842 ) | ( ~n6000 & n13486 ) | ( n9842 & n13486 ) ;
  assign n13488 = n13487 ^ n10481 ^ 1'b0 ;
  assign n13489 = n5508 | n11235 ;
  assign n13490 = n12385 & ~n13489 ;
  assign n13491 = n13490 ^ n2694 ^ 1'b0 ;
  assign n13492 = ~n469 & n5388 ;
  assign n13493 = n13492 ^ n1418 ^ 1'b0 ;
  assign n13494 = n9714 & n13493 ;
  assign n13495 = n4410 ^ n1897 ^ 1'b0 ;
  assign n13496 = x100 & n2744 ;
  assign n13497 = n13495 & n13496 ;
  assign n13498 = n3038 | n4945 ;
  assign n13499 = n7556 & ~n13498 ;
  assign n13500 = n13499 ^ n686 ^ 1'b0 ;
  assign n13501 = ~n3501 & n13500 ;
  assign n13502 = n6123 ^ n2378 ^ 1'b0 ;
  assign n13503 = ~n1858 & n13502 ;
  assign n13504 = ~n1871 & n3933 ;
  assign n13505 = n6232 & n13504 ;
  assign n13506 = n13503 | n13505 ;
  assign n13507 = n13506 ^ n11321 ^ 1'b0 ;
  assign n13508 = n13501 | n13507 ;
  assign n13509 = n3856 & ~n5824 ;
  assign n13510 = n3373 & n11309 ;
  assign n13511 = n8427 ^ n8216 ^ 1'b0 ;
  assign n13512 = n8662 | n13511 ;
  assign n13513 = n4615 & ~n13512 ;
  assign n13514 = n13510 & ~n13513 ;
  assign n13515 = n13514 ^ x137 ^ 1'b0 ;
  assign n13516 = ( n2555 & n3737 ) | ( n2555 & n8579 ) | ( n3737 & n8579 ) ;
  assign n13517 = n13516 ^ n9856 ^ 1'b0 ;
  assign n13518 = n13517 ^ n1372 ^ 1'b0 ;
  assign n13519 = n713 | n852 ;
  assign n13520 = n13519 ^ n3903 ^ 1'b0 ;
  assign n13521 = n13520 ^ n2971 ^ 1'b0 ;
  assign n13522 = n7913 ^ n1470 ^ 1'b0 ;
  assign n13523 = n5428 | n13522 ;
  assign n13524 = n13523 ^ n11572 ^ 1'b0 ;
  assign n13525 = n5982 | n13524 ;
  assign n13526 = n13521 | n13525 ;
  assign n13527 = n13526 ^ n9486 ^ 1'b0 ;
  assign n13528 = n13518 & n13527 ;
  assign n13529 = x221 & n4852 ;
  assign n13530 = n13529 ^ n371 ^ 1'b0 ;
  assign n13531 = x227 & n13530 ;
  assign n13532 = n6393 ^ n3530 ^ 1'b0 ;
  assign n13533 = ~n6170 & n13532 ;
  assign n13534 = n10453 ^ n7325 ^ 1'b0 ;
  assign n13535 = n13533 & n13534 ;
  assign n13536 = n11426 ^ n9371 ^ 1'b0 ;
  assign n13537 = x104 & ~n11242 ;
  assign n13538 = ~n5645 & n5923 ;
  assign n13539 = n10516 ^ n1321 ^ 1'b0 ;
  assign n13540 = ~n13538 & n13539 ;
  assign n13541 = n2034 & ~n5720 ;
  assign n13542 = n3691 & n13541 ;
  assign n13543 = n1472 & ~n10155 ;
  assign n13544 = ( n1302 & n5259 ) | ( n1302 & n13543 ) | ( n5259 & n13543 ) ;
  assign n13545 = n5695 | n13544 ;
  assign n13546 = n13545 ^ n10162 ^ 1'b0 ;
  assign n13547 = ~n1199 & n6279 ;
  assign n13548 = ~n3198 & n3716 ;
  assign n13549 = n3507 & n13548 ;
  assign n13550 = n13547 | n13549 ;
  assign n13551 = n1782 & ~n2714 ;
  assign n13552 = n13030 ^ n7703 ^ n7317 ;
  assign n13553 = n12475 ^ n5767 ^ n4662 ;
  assign n13554 = n2493 ^ n650 ^ 1'b0 ;
  assign n13555 = n13553 | n13554 ;
  assign n13556 = ( n7760 & n13552 ) | ( n7760 & ~n13555 ) | ( n13552 & ~n13555 ) ;
  assign n13557 = n11067 & n13556 ;
  assign n13558 = n8046 & n13557 ;
  assign n13559 = ~n2250 & n3598 ;
  assign n13560 = n8833 ^ n8270 ^ n2719 ;
  assign n13562 = n7654 ^ n4323 ^ n3806 ;
  assign n13561 = n4432 | n7732 ;
  assign n13563 = n13562 ^ n13561 ^ 1'b0 ;
  assign n13564 = n8125 ^ n7810 ^ n7632 ;
  assign n13565 = n7339 & n11471 ;
  assign n13566 = n8722 ^ n8525 ^ n6555 ;
  assign n13567 = n13566 ^ n10014 ^ 1'b0 ;
  assign n13568 = n13567 ^ n7520 ^ 1'b0 ;
  assign n13569 = n4862 & n8612 ;
  assign n13570 = ~n5968 & n13569 ;
  assign n13571 = n4967 | n13570 ;
  assign n13572 = n10628 & n10935 ;
  assign n13573 = n7088 ^ n3501 ^ 1'b0 ;
  assign n13574 = n399 & n13573 ;
  assign n13575 = n11111 | n13574 ;
  assign n13576 = ~n1830 & n7627 ;
  assign n13577 = n13576 ^ n8310 ^ 1'b0 ;
  assign n13578 = n13577 ^ n13278 ^ 1'b0 ;
  assign n13579 = n5491 & ~n10020 ;
  assign n13580 = ~n2537 & n8661 ;
  assign n13581 = n13580 ^ n11725 ^ n7531 ;
  assign n13582 = n559 & n8829 ;
  assign n13583 = n13582 ^ n743 ^ 1'b0 ;
  assign n13584 = ( ~n1520 & n12573 ) | ( ~n1520 & n13583 ) | ( n12573 & n13583 ) ;
  assign n13585 = n13584 ^ n4342 ^ 1'b0 ;
  assign n13586 = n3089 | n7263 ;
  assign n13587 = n13585 & ~n13586 ;
  assign n13588 = ~n2795 & n13587 ;
  assign n13595 = n2737 ^ x76 ^ 1'b0 ;
  assign n13596 = n2558 & n13595 ;
  assign n13594 = ~n3202 & n3700 ;
  assign n13597 = n13596 ^ n13594 ^ 1'b0 ;
  assign n13589 = ( n1890 & n4074 ) | ( n1890 & n4868 ) | ( n4074 & n4868 ) ;
  assign n13590 = n8437 | n13589 ;
  assign n13591 = n13590 ^ n3439 ^ 1'b0 ;
  assign n13592 = n7370 | n13591 ;
  assign n13593 = n13592 ^ n7680 ^ 1'b0 ;
  assign n13598 = n13597 ^ n13593 ^ n8202 ;
  assign n13599 = n9115 ^ n3209 ^ 1'b0 ;
  assign n13600 = n9625 & n13599 ;
  assign n13601 = n13600 ^ n13141 ^ n9320 ;
  assign n13602 = n3955 & ~n5531 ;
  assign n13603 = ~n13584 & n13602 ;
  assign n13604 = n13603 ^ n13421 ^ 1'b0 ;
  assign n13605 = ( n3175 & n3274 ) | ( n3175 & n9431 ) | ( n3274 & n9431 ) ;
  assign n13606 = n516 | n5538 ;
  assign n13607 = ( x17 & ~n12044 ) | ( x17 & n13605 ) | ( ~n12044 & n13605 ) ;
  assign n13612 = ( x248 & n387 ) | ( x248 & n5261 ) | ( n387 & n5261 ) ;
  assign n13608 = ( n1129 & n4793 ) | ( n1129 & ~n6228 ) | ( n4793 & ~n6228 ) ;
  assign n13609 = n13608 ^ n7421 ^ n1210 ;
  assign n13610 = n13609 ^ n4864 ^ 1'b0 ;
  assign n13611 = ( ~n1619 & n3415 ) | ( ~n1619 & n13610 ) | ( n3415 & n13610 ) ;
  assign n13613 = n13612 ^ n13611 ^ 1'b0 ;
  assign n13628 = n7853 & n12767 ;
  assign n13629 = n13628 ^ n6422 ^ 1'b0 ;
  assign n13630 = ~n2785 & n13629 ;
  assign n13614 = n13333 ^ n2780 ^ 1'b0 ;
  assign n13615 = x120 & n10867 ;
  assign n13616 = n4009 & n13615 ;
  assign n13620 = x38 & n5474 ;
  assign n13621 = n13620 ^ n3922 ^ 1'b0 ;
  assign n13617 = ~x135 & n446 ;
  assign n13618 = n4969 & n13617 ;
  assign n13619 = n13618 ^ n2305 ^ 1'b0 ;
  assign n13622 = n13621 ^ n13619 ^ 1'b0 ;
  assign n13623 = n13616 | n13622 ;
  assign n13624 = n13614 | n13623 ;
  assign n13625 = n10893 & n13624 ;
  assign n13626 = ~n9680 & n13625 ;
  assign n13627 = n11988 & n13626 ;
  assign n13631 = n13630 ^ n13627 ^ 1'b0 ;
  assign n13632 = ~n4462 & n5590 ;
  assign n13633 = n8310 | n12810 ;
  assign n13634 = n6227 | n13633 ;
  assign n13635 = n2799 ^ n1054 ^ 1'b0 ;
  assign n13636 = n6835 ^ n5347 ^ 1'b0 ;
  assign n13637 = n6709 & n13636 ;
  assign n13638 = n9569 ^ n6342 ^ 1'b0 ;
  assign n13639 = n13637 & n13638 ;
  assign n13647 = n369 & ~n2318 ;
  assign n13640 = n7801 ^ n1930 ^ 1'b0 ;
  assign n13642 = n727 | n3132 ;
  assign n13643 = n2468 & ~n13642 ;
  assign n13641 = n2352 & ~n8710 ;
  assign n13644 = n13643 ^ n13641 ^ 1'b0 ;
  assign n13645 = n6353 & n13644 ;
  assign n13646 = n13640 & n13645 ;
  assign n13648 = n13647 ^ n13646 ^ 1'b0 ;
  assign n13649 = n9656 & n13648 ;
  assign n13650 = n740 & n2916 ;
  assign n13651 = n1547 & ~n4007 ;
  assign n13652 = n7068 | n9537 ;
  assign n13653 = n13651 & ~n13652 ;
  assign n13657 = n933 & ~n5532 ;
  assign n13654 = n4862 ^ n3493 ^ 1'b0 ;
  assign n13655 = n3099 | n13654 ;
  assign n13656 = n5380 | n13655 ;
  assign n13658 = n13657 ^ n13656 ^ 1'b0 ;
  assign n13659 = ~n1453 & n13658 ;
  assign n13660 = ~n2833 & n13659 ;
  assign n13661 = n13653 & n13660 ;
  assign n13662 = n13661 ^ n13203 ^ n7884 ;
  assign n13663 = n5899 & n9083 ;
  assign n13664 = n3640 | n12747 ;
  assign n13666 = n8630 ^ n4100 ^ n2959 ;
  assign n13667 = ~n7706 & n13666 ;
  assign n13668 = n8080 & n13667 ;
  assign n13669 = n9793 | n13668 ;
  assign n13665 = n6409 | n7374 ;
  assign n13670 = n13669 ^ n13665 ^ 1'b0 ;
  assign n13671 = n11614 ^ n5582 ^ n5425 ;
  assign n13672 = n6510 & ~n13203 ;
  assign n13673 = n13672 ^ n8000 ^ 1'b0 ;
  assign n13674 = ~n3145 & n4978 ;
  assign n13675 = n6726 & ~n12020 ;
  assign n13676 = n13675 ^ n565 ^ 1'b0 ;
  assign n13677 = n13437 ^ n1126 ^ 1'b0 ;
  assign n13678 = n4757 & ~n4758 ;
  assign n13679 = n9986 | n13678 ;
  assign n13680 = n10393 ^ n809 ^ 1'b0 ;
  assign n13681 = n9942 & n13680 ;
  assign n13682 = n13679 & n13681 ;
  assign n13683 = n10639 ^ n7894 ^ n7112 ;
  assign n13684 = n617 & n3682 ;
  assign n13685 = n8138 ^ n604 ^ 1'b0 ;
  assign n13688 = n946 ^ n555 ^ 1'b0 ;
  assign n13687 = n4335 ^ n1210 ^ 1'b0 ;
  assign n13689 = n13688 ^ n13687 ^ 1'b0 ;
  assign n13690 = n1610 & ~n4440 ;
  assign n13691 = n13689 & n13690 ;
  assign n13692 = n13691 ^ n11225 ^ 1'b0 ;
  assign n13686 = n1340 & n4579 ;
  assign n13693 = n13692 ^ n13686 ^ 1'b0 ;
  assign n13694 = n878 | n4903 ;
  assign n13695 = ~n418 & n1458 ;
  assign n13696 = ( n6364 & ~n13694 ) | ( n6364 & n13695 ) | ( ~n13694 & n13695 ) ;
  assign n13697 = n13696 ^ n12568 ^ 1'b0 ;
  assign n13698 = n2797 & n13697 ;
  assign n13699 = n9640 ^ n6739 ^ 1'b0 ;
  assign n13700 = n6931 & ~n13699 ;
  assign n13702 = n11792 ^ n9026 ^ 1'b0 ;
  assign n13701 = ~n4203 & n12973 ;
  assign n13703 = n13702 ^ n13701 ^ 1'b0 ;
  assign n13704 = n6700 | n12608 ;
  assign n13705 = n1429 & ~n1477 ;
  assign n13706 = ( n5343 & n9767 ) | ( n5343 & n13705 ) | ( n9767 & n13705 ) ;
  assign n13707 = ~n2084 & n13706 ;
  assign n13708 = n3610 ^ n727 ^ 1'b0 ;
  assign n13709 = n8886 ^ n7325 ^ 1'b0 ;
  assign n13710 = n7008 | n8717 ;
  assign n13711 = n12666 | n13710 ;
  assign n13712 = n8702 ^ n1064 ^ 1'b0 ;
  assign n13713 = n13711 & ~n13712 ;
  assign n13714 = n7598 ^ n692 ^ 1'b0 ;
  assign n13715 = n928 | n13714 ;
  assign n13716 = n4480 | n13715 ;
  assign n13717 = ( n1985 & ~n2523 ) | ( n1985 & n9618 ) | ( ~n2523 & n9618 ) ;
  assign n13718 = ~n13716 & n13717 ;
  assign n13719 = ~n852 & n9670 ;
  assign n13720 = n13719 ^ n1610 ^ 1'b0 ;
  assign n13721 = n12341 ^ n1117 ^ 1'b0 ;
  assign n13722 = n5269 | n13721 ;
  assign n13723 = n10323 | n13140 ;
  assign n13724 = ~n10707 & n12213 ;
  assign n13725 = n9247 & n13724 ;
  assign n13726 = n13725 ^ n12480 ^ n1944 ;
  assign n13727 = n3098 & ~n6442 ;
  assign n13728 = n13727 ^ n13362 ^ 1'b0 ;
  assign n13729 = x15 & ~n13728 ;
  assign n13730 = n1775 & n10999 ;
  assign n13731 = n7002 ^ n4438 ^ 1'b0 ;
  assign n13732 = n6166 & ~n13731 ;
  assign n13733 = n5138 & n13732 ;
  assign n13734 = n13733 ^ n12500 ^ 1'b0 ;
  assign n13735 = x1 & ~n13734 ;
  assign n13736 = n13735 ^ n7282 ^ 1'b0 ;
  assign n13737 = n2160 | n13736 ;
  assign n13738 = ( n3829 & ~n8586 ) | ( n3829 & n8588 ) | ( ~n8586 & n8588 ) ;
  assign n13739 = n13738 ^ n7965 ^ n6868 ;
  assign n13740 = n2100 & n2648 ;
  assign n13741 = n13740 ^ n7926 ^ n7799 ;
  assign n13746 = n3257 & ~n3487 ;
  assign n13742 = n2967 & ~n3089 ;
  assign n13743 = n471 | n5045 ;
  assign n13744 = n13742 & ~n13743 ;
  assign n13745 = n9429 & ~n13744 ;
  assign n13747 = n13746 ^ n13745 ^ 1'b0 ;
  assign n13748 = ( n1518 & n1880 ) | ( n1518 & n3293 ) | ( n1880 & n3293 ) ;
  assign n13749 = n1453 & ~n4840 ;
  assign n13750 = n13748 | n13749 ;
  assign n13751 = ~n6424 & n13750 ;
  assign n13752 = ~n8533 & n13751 ;
  assign n13753 = n723 & n9962 ;
  assign n13754 = n2746 & n13753 ;
  assign n13755 = x94 & ~n4073 ;
  assign n13756 = n13755 ^ n897 ^ 1'b0 ;
  assign n13757 = n13756 ^ n4765 ^ 1'b0 ;
  assign n13758 = ~n10516 & n13757 ;
  assign n13759 = n1266 | n11641 ;
  assign n13760 = ( n2192 & n4902 ) | ( n2192 & ~n5667 ) | ( n4902 & ~n5667 ) ;
  assign n13761 = n13760 ^ x158 ^ 1'b0 ;
  assign n13762 = n13759 & ~n13761 ;
  assign n13763 = n8494 ^ n3658 ^ 1'b0 ;
  assign n13764 = n3551 ^ n1036 ^ 1'b0 ;
  assign n13765 = n13763 & n13764 ;
  assign n13766 = ( n8415 & ~n10690 ) | ( n8415 & n13674 ) | ( ~n10690 & n13674 ) ;
  assign n13767 = n8309 ^ n1072 ^ 1'b0 ;
  assign n13768 = n7852 & n13767 ;
  assign n13769 = n2101 | n10114 ;
  assign n13770 = n6501 ^ n2651 ^ 1'b0 ;
  assign n13771 = ~n13194 & n13770 ;
  assign n13772 = n13771 ^ n8315 ^ 1'b0 ;
  assign n13773 = n2029 & ~n6045 ;
  assign n13774 = n9961 & n13773 ;
  assign n13775 = n13774 ^ n8532 ^ 1'b0 ;
  assign n13776 = n4328 ^ n2433 ^ 1'b0 ;
  assign n13777 = n13775 & ~n13776 ;
  assign n13778 = ( x211 & n4921 ) | ( x211 & ~n13488 ) | ( n4921 & ~n13488 ) ;
  assign n13779 = n5989 | n10479 ;
  assign n13780 = n5051 & ~n13779 ;
  assign n13781 = n5518 ^ n1296 ^ 1'b0 ;
  assign n13782 = n5260 | n10625 ;
  assign n13783 = n13781 & ~n13782 ;
  assign n13784 = n4458 ^ n1212 ^ 1'b0 ;
  assign n13785 = n984 & n10010 ;
  assign n13786 = n5882 & n13785 ;
  assign n13787 = n13786 ^ n4719 ^ 1'b0 ;
  assign n13788 = n11297 & ~n13787 ;
  assign n13789 = ~n13784 & n13788 ;
  assign n13790 = n5834 ^ n4966 ^ 1'b0 ;
  assign n13791 = n6938 | n7424 ;
  assign n13792 = n3376 & ~n11357 ;
  assign n13793 = n3479 & ~n13792 ;
  assign n13794 = ~n9261 & n13793 ;
  assign n13795 = ~n10344 & n13794 ;
  assign n13796 = n2095 & n11670 ;
  assign n13797 = n8510 ^ n8329 ^ 1'b0 ;
  assign n13798 = n831 & ~n4626 ;
  assign n13799 = ~x11 & n13798 ;
  assign n13800 = n4279 & ~n13799 ;
  assign n13801 = ~n3103 & n13800 ;
  assign n13802 = n13801 ^ n4505 ^ 1'b0 ;
  assign n13803 = n3414 & ~n13802 ;
  assign n13804 = n13715 ^ n2471 ^ 1'b0 ;
  assign n13805 = n8100 & n13804 ;
  assign n13806 = n952 | n13805 ;
  assign n13807 = n10922 ^ n747 ^ 1'b0 ;
  assign n13808 = ~n2362 & n11764 ;
  assign n13809 = n13808 ^ n3600 ^ 1'b0 ;
  assign n13810 = n4378 ^ n1985 ^ 1'b0 ;
  assign n13811 = n6406 & n13810 ;
  assign n13812 = n13811 ^ x77 ^ 1'b0 ;
  assign n13813 = n6042 & n11906 ;
  assign n13814 = n2555 | n4677 ;
  assign n13815 = n3775 & n13814 ;
  assign n13816 = ~n13813 & n13815 ;
  assign n13817 = n3048 | n3402 ;
  assign n13818 = ( n5762 & ~n13816 ) | ( n5762 & n13817 ) | ( ~n13816 & n13817 ) ;
  assign n13819 = ( ~n6671 & n11039 ) | ( ~n6671 & n12172 ) | ( n11039 & n12172 ) ;
  assign n13820 = n4123 | n10768 ;
  assign n13821 = n420 & ~n13820 ;
  assign n13822 = n4639 | n5095 ;
  assign n13823 = n13822 ^ n3650 ^ 1'b0 ;
  assign n13824 = n13823 ^ n3808 ^ 1'b0 ;
  assign n13825 = ~n6470 & n8721 ;
  assign n13826 = ~n2567 & n13825 ;
  assign n13827 = n13826 ^ n8957 ^ n5496 ;
  assign n13829 = n4210 & ~n6202 ;
  assign n13828 = n3062 & ~n11471 ;
  assign n13830 = n13829 ^ n13828 ^ 1'b0 ;
  assign n13831 = n6535 ^ n3738 ^ 1'b0 ;
  assign n13832 = n6766 & n13831 ;
  assign n13833 = n2601 & ~n10359 ;
  assign n13834 = ~n13832 & n13833 ;
  assign n13835 = n10713 ^ n2877 ^ 1'b0 ;
  assign n13836 = n5451 ^ n1477 ^ 1'b0 ;
  assign n13837 = n5496 | n13836 ;
  assign n13838 = n3716 & ~n9011 ;
  assign n13839 = n13837 & n13838 ;
  assign n13840 = n12085 | n13040 ;
  assign n13841 = n13839 & ~n13840 ;
  assign n13842 = n5469 ^ n3222 ^ 1'b0 ;
  assign n13843 = n6401 ^ n1088 ^ 1'b0 ;
  assign n13844 = ~n854 & n13843 ;
  assign n13845 = n4990 ^ n3118 ^ 1'b0 ;
  assign n13846 = n5329 & ~n13845 ;
  assign n13847 = n10288 ^ n2619 ^ 1'b0 ;
  assign n13848 = n7976 ^ n4223 ^ x189 ;
  assign n13849 = n2578 & ~n13848 ;
  assign n13850 = n13849 ^ x86 ^ 1'b0 ;
  assign n13851 = n7752 | n12152 ;
  assign n13852 = n13851 ^ n9332 ^ 1'b0 ;
  assign n13853 = n10975 ^ n9501 ^ 1'b0 ;
  assign n13854 = n3413 | n10536 ;
  assign n13857 = n1843 & ~n2800 ;
  assign n13855 = n732 & ~n3051 ;
  assign n13856 = n9295 & n13855 ;
  assign n13858 = n13857 ^ n13856 ^ 1'b0 ;
  assign n13859 = n3691 | n13858 ;
  assign n13860 = n10451 ^ n4212 ^ 1'b0 ;
  assign n13861 = x32 & n13860 ;
  assign n13862 = ~n3205 & n6182 ;
  assign n13863 = n337 & n13862 ;
  assign n13864 = n3216 & n9067 ;
  assign n13865 = n13752 ^ n2055 ^ 1'b0 ;
  assign n13866 = ~n13864 & n13865 ;
  assign n13867 = n13866 ^ n11133 ^ 1'b0 ;
  assign n13876 = n1339 ^ x58 ^ 1'b0 ;
  assign n13877 = n1113 & ~n13876 ;
  assign n13874 = n11884 ^ n506 ^ 1'b0 ;
  assign n13875 = n3315 | n13874 ;
  assign n13868 = ~n2881 & n3023 ;
  assign n13869 = ~x0 & n1097 ;
  assign n13870 = n10749 & n13869 ;
  assign n13871 = n10675 & ~n13870 ;
  assign n13872 = n13868 & n13871 ;
  assign n13873 = n3430 & n13872 ;
  assign n13878 = n13877 ^ n13875 ^ n13873 ;
  assign n13879 = n1007 | n7580 ;
  assign n13880 = n3487 ^ n2374 ^ 1'b0 ;
  assign n13881 = n7943 & n13880 ;
  assign n13882 = n5618 & n13881 ;
  assign n13883 = n13882 ^ n7658 ^ 1'b0 ;
  assign n13884 = n2262 ^ n1963 ^ 1'b0 ;
  assign n13885 = n7175 | n13884 ;
  assign n13886 = n13885 ^ n4019 ^ 1'b0 ;
  assign n13887 = n1869 & n13886 ;
  assign n13888 = n13887 ^ n9195 ^ 1'b0 ;
  assign n13889 = n9718 & ~n13888 ;
  assign n13890 = ( n6893 & n11499 ) | ( n6893 & n13889 ) | ( n11499 & n13889 ) ;
  assign n13891 = n1470 & n13122 ;
  assign n13892 = n13891 ^ n1781 ^ 1'b0 ;
  assign n13893 = ( x114 & n998 ) | ( x114 & ~n13892 ) | ( n998 & ~n13892 ) ;
  assign n13894 = n5315 ^ n2953 ^ 1'b0 ;
  assign n13895 = ( n1993 & n9108 ) | ( n1993 & ~n13894 ) | ( n9108 & ~n13894 ) ;
  assign n13896 = ( ~n3709 & n7190 ) | ( ~n3709 & n13895 ) | ( n7190 & n13895 ) ;
  assign n13897 = n13896 ^ n10610 ^ 1'b0 ;
  assign n13898 = n2406 | n2808 ;
  assign n13899 = n13898 ^ n8889 ^ 1'b0 ;
  assign n13900 = n9974 ^ n9954 ^ n1041 ;
  assign n13901 = n8739 | n13900 ;
  assign n13902 = n13899 & ~n13901 ;
  assign n13903 = n13897 & ~n13902 ;
  assign n13904 = ~n5205 & n11064 ;
  assign n13905 = n2141 & ~n9170 ;
  assign n13906 = n13905 ^ n11149 ^ 1'b0 ;
  assign n13907 = n7622 ^ n614 ^ 1'b0 ;
  assign n13908 = n13907 ^ n1233 ^ 1'b0 ;
  assign n13909 = ~n11945 & n13908 ;
  assign n13910 = n8354 ^ n1886 ^ 1'b0 ;
  assign n13911 = n8130 & ~n13910 ;
  assign n13912 = ~n5806 & n13911 ;
  assign n13913 = ~n11931 & n13912 ;
  assign n13914 = n6203 | n9623 ;
  assign n13915 = n13914 ^ n906 ^ 1'b0 ;
  assign n13916 = ~n13913 & n13915 ;
  assign n13917 = n2518 & n5636 ;
  assign n13918 = n10990 | n13917 ;
  assign n13919 = n13916 | n13918 ;
  assign n13920 = n514 | n4023 ;
  assign n13921 = n13920 ^ n10411 ^ n2518 ;
  assign n13922 = n10445 ^ n2637 ^ 1'b0 ;
  assign n13923 = n4980 & n13922 ;
  assign n13928 = n5610 ^ n2507 ^ 1'b0 ;
  assign n13929 = n2337 & ~n2915 ;
  assign n13930 = n13928 & n13929 ;
  assign n13926 = ~n8266 & n8663 ;
  assign n13924 = n4298 ^ n2682 ^ 1'b0 ;
  assign n13925 = n13924 ^ n2151 ^ n1932 ;
  assign n13927 = n13926 ^ n13925 ^ n5271 ;
  assign n13931 = n13930 ^ n13927 ^ 1'b0 ;
  assign n13932 = ( ~n5833 & n8340 ) | ( ~n5833 & n13144 ) | ( n8340 & n13144 ) ;
  assign n13933 = n7930 & ~n11681 ;
  assign n13934 = n9341 & n13933 ;
  assign n13935 = n6526 ^ x48 ^ 1'b0 ;
  assign n13936 = n4428 & n13935 ;
  assign n13937 = n2787 | n13936 ;
  assign n13938 = n3218 & ~n8189 ;
  assign n13944 = n13774 ^ n1265 ^ 1'b0 ;
  assign n13939 = ( ~n407 & n3363 ) | ( ~n407 & n7095 ) | ( n3363 & n7095 ) ;
  assign n13940 = n565 & ~n6963 ;
  assign n13941 = ~x170 & n13940 ;
  assign n13942 = n13939 & ~n13941 ;
  assign n13943 = x165 & n13942 ;
  assign n13945 = n13944 ^ n13943 ^ 1'b0 ;
  assign n13946 = n13945 ^ n1025 ^ 1'b0 ;
  assign n13947 = n13946 ^ n10209 ^ n288 ;
  assign n13948 = n2497 | n3413 ;
  assign n13949 = n5172 | n7987 ;
  assign n13950 = n6359 ^ n2959 ^ 1'b0 ;
  assign n13951 = n1029 & ~n2783 ;
  assign n13952 = ~n13950 & n13951 ;
  assign n13953 = n1258 | n7765 ;
  assign n13954 = n13952 & ~n13953 ;
  assign n13955 = x169 & n13954 ;
  assign n13956 = n1034 & ~n13543 ;
  assign n13957 = n10122 ^ n2449 ^ 1'b0 ;
  assign n13958 = x34 & n10548 ;
  assign n13959 = ~n10548 & n13958 ;
  assign n13960 = n13959 ^ n8453 ^ 1'b0 ;
  assign n13961 = n4423 & ~n9126 ;
  assign n13962 = ~n4423 & n13961 ;
  assign n13963 = n13962 ^ n13364 ^ 1'b0 ;
  assign n13964 = ( n8065 & n13960 ) | ( n8065 & n13963 ) | ( n13960 & n13963 ) ;
  assign n13965 = n6726 & ~n10720 ;
  assign n13966 = ~n5579 & n13965 ;
  assign n13967 = n8020 ^ n2357 ^ 1'b0 ;
  assign n13968 = ( n6455 & n13966 ) | ( n6455 & n13967 ) | ( n13966 & n13967 ) ;
  assign n13969 = x248 & n6216 ;
  assign n13970 = n13969 ^ n3118 ^ 1'b0 ;
  assign n13971 = n13970 ^ n1518 ^ 1'b0 ;
  assign n13972 = n2668 & n13971 ;
  assign n13973 = n557 & ~n13915 ;
  assign n13974 = n5942 | n6894 ;
  assign n13975 = n13974 ^ n3599 ^ 1'b0 ;
  assign n13976 = n13975 ^ n13183 ^ 1'b0 ;
  assign n13977 = n9076 ^ n7204 ^ 1'b0 ;
  assign n13978 = n6682 | n13977 ;
  assign n13979 = n13978 ^ n13666 ^ 1'b0 ;
  assign n13980 = ~n1103 & n13979 ;
  assign n13981 = n2598 ^ n1869 ^ 1'b0 ;
  assign n13982 = ( n387 & n1729 ) | ( n387 & ~n13981 ) | ( n1729 & ~n13981 ) ;
  assign n13983 = n8007 | n13982 ;
  assign n13985 = n5040 ^ n2061 ^ x135 ;
  assign n13986 = n5825 & ~n13985 ;
  assign n13987 = n5085 | n13986 ;
  assign n13988 = n13987 ^ n8539 ^ 1'b0 ;
  assign n13989 = n13988 ^ n1189 ^ 1'b0 ;
  assign n13984 = x7 | n1312 ;
  assign n13990 = n13989 ^ n13984 ^ 1'b0 ;
  assign n13991 = n13990 ^ n1272 ^ 1'b0 ;
  assign n13992 = n13983 | n13991 ;
  assign n13993 = n7211 ^ n6138 ^ 1'b0 ;
  assign n13994 = ~n11642 & n13993 ;
  assign n13995 = n5379 ^ n5116 ^ 1'b0 ;
  assign n13996 = n438 & n4493 ;
  assign n13997 = n3039 & ~n13996 ;
  assign n13998 = n1486 & n13997 ;
  assign n13999 = n10159 | n13998 ;
  assign n14000 = n13999 ^ n518 ^ 1'b0 ;
  assign n14001 = ~n12329 & n14000 ;
  assign n14002 = ~n13995 & n14001 ;
  assign n14007 = n2786 ^ n395 ^ 1'b0 ;
  assign n14008 = n14007 ^ n10164 ^ n5016 ;
  assign n14005 = n9320 ^ n7645 ^ 1'b0 ;
  assign n14006 = n14005 ^ n11756 ^ 1'b0 ;
  assign n14003 = ( n2428 & ~n2773 ) | ( n2428 & n12011 ) | ( ~n2773 & n12011 ) ;
  assign n14004 = n6054 & ~n14003 ;
  assign n14009 = n14008 ^ n14006 ^ n14004 ;
  assign n14010 = n5996 ^ n5425 ^ 1'b0 ;
  assign n14011 = n14010 ^ n11459 ^ 1'b0 ;
  assign n14012 = n3419 & n14011 ;
  assign n14013 = n14012 ^ n7646 ^ 1'b0 ;
  assign n14014 = n326 & ~n14013 ;
  assign n14015 = n13217 ^ n7645 ^ 1'b0 ;
  assign n14016 = n2135 & n6980 ;
  assign n14017 = n14016 ^ n7556 ^ n4907 ;
  assign n14018 = n2610 ^ n1795 ^ 1'b0 ;
  assign n14019 = n8539 | n14018 ;
  assign n14020 = ( x7 & n2081 ) | ( x7 & n4312 ) | ( n2081 & n4312 ) ;
  assign n14021 = n14019 & ~n14020 ;
  assign n14022 = ~n14017 & n14021 ;
  assign n14023 = ~n1033 & n1155 ;
  assign n14024 = ~n9457 & n14023 ;
  assign n14025 = n14022 & n14024 ;
  assign n14026 = n1865 | n14025 ;
  assign n14027 = n14026 ^ n9757 ^ 1'b0 ;
  assign n14028 = n1437 & ~n8314 ;
  assign n14029 = n1550 & n7863 ;
  assign n14030 = ~n5464 & n14029 ;
  assign n14031 = n14030 ^ n1011 ^ 1'b0 ;
  assign n14032 = n14028 & n14031 ;
  assign n14033 = n10016 ^ n4602 ^ 1'b0 ;
  assign n14034 = n9645 & n14033 ;
  assign n14035 = n5915 & n13239 ;
  assign n14036 = n335 | n14035 ;
  assign n14037 = n3443 & n5414 ;
  assign n14038 = ~n14036 & n14037 ;
  assign n14039 = n14038 ^ n2463 ^ 1'b0 ;
  assign n14040 = ~n904 & n14039 ;
  assign n14041 = ~n10326 & n11749 ;
  assign n14042 = n1520 & ~n3662 ;
  assign n14043 = n8393 ^ n8064 ^ 1'b0 ;
  assign n14044 = n14042 | n14043 ;
  assign n14045 = n9059 | n14044 ;
  assign n14046 = n10268 ^ n3287 ^ 1'b0 ;
  assign n14047 = n14046 ^ n1969 ^ 1'b0 ;
  assign n14048 = n14047 ^ n1255 ^ 1'b0 ;
  assign n14049 = ( ~n1963 & n3058 ) | ( ~n1963 & n7443 ) | ( n3058 & n7443 ) ;
  assign n14050 = n2368 & ~n14049 ;
  assign n14051 = n5503 & n14050 ;
  assign n14052 = n2186 & ~n14051 ;
  assign n14053 = n9068 ^ n2002 ^ 1'b0 ;
  assign n14054 = n2937 & ~n14053 ;
  assign n14055 = n11719 ^ n10815 ^ 1'b0 ;
  assign n14056 = n11383 & n12415 ;
  assign n14057 = n14056 ^ n3328 ^ 1'b0 ;
  assign n14058 = n6292 & n14057 ;
  assign n14059 = n6642 ^ x223 ^ 1'b0 ;
  assign n14060 = n14059 ^ n301 ^ 1'b0 ;
  assign n14061 = n9995 | n14060 ;
  assign n14062 = n3808 ^ n1231 ^ 1'b0 ;
  assign n14063 = n14062 ^ n6792 ^ n645 ;
  assign n14064 = n14063 ^ n3291 ^ 1'b0 ;
  assign n14065 = n12998 & ~n14064 ;
  assign n14067 = n2230 | n10862 ;
  assign n14066 = x197 & ~n2907 ;
  assign n14068 = n14067 ^ n14066 ^ 1'b0 ;
  assign n14069 = n12921 ^ n1281 ^ 1'b0 ;
  assign n14070 = n12785 & ~n14069 ;
  assign n14071 = n961 & ~n11810 ;
  assign n14072 = ~n9542 & n14071 ;
  assign n14073 = ~n1760 & n14072 ;
  assign n14074 = n3171 | n14073 ;
  assign n14075 = n14074 ^ n8515 ^ 1'b0 ;
  assign n14076 = n12148 ^ n5685 ^ n2299 ;
  assign n14080 = n4339 ^ n2212 ^ n840 ;
  assign n14078 = n5537 & n9874 ;
  assign n14079 = n11361 & n14078 ;
  assign n14077 = n2762 ^ n2192 ^ 1'b0 ;
  assign n14081 = n14080 ^ n14079 ^ n14077 ;
  assign n14082 = n7495 ^ n7436 ^ 1'b0 ;
  assign n14083 = n4600 & ~n14082 ;
  assign n14084 = n14083 ^ n5047 ^ n1015 ;
  assign n14085 = n10114 ^ n4511 ^ n1443 ;
  assign n14086 = n14085 ^ n11310 ^ n1281 ;
  assign n14087 = n14086 ^ n10661 ^ 1'b0 ;
  assign n14088 = n14084 & ~n14087 ;
  assign n14089 = n14046 ^ n8908 ^ 1'b0 ;
  assign n14090 = n8651 | n14089 ;
  assign n14091 = n14090 ^ n274 ^ 1'b0 ;
  assign n14092 = ~n10978 & n14091 ;
  assign n14093 = ~n1980 & n3922 ;
  assign n14094 = n2543 ^ n1571 ^ 1'b0 ;
  assign n14095 = n1490 & ~n14094 ;
  assign n14096 = ~n3431 & n14095 ;
  assign n14097 = n14096 ^ n317 ^ 1'b0 ;
  assign n14098 = ( n2561 & n14093 ) | ( n2561 & ~n14097 ) | ( n14093 & ~n14097 ) ;
  assign n14099 = n10690 ^ n8212 ^ 1'b0 ;
  assign n14100 = n5729 & n14099 ;
  assign n14101 = ~n6853 & n14100 ;
  assign n14102 = n14101 ^ n11921 ^ 1'b0 ;
  assign n14103 = n11357 & n11725 ;
  assign n14104 = n14103 ^ n2384 ^ 1'b0 ;
  assign n14106 = n6405 ^ n5953 ^ n1577 ;
  assign n14107 = n8256 & n14106 ;
  assign n14108 = n7515 & n14107 ;
  assign n14105 = n11149 ^ n3882 ^ 1'b0 ;
  assign n14109 = n14108 ^ n14105 ^ 1'b0 ;
  assign n14110 = n13399 & n14109 ;
  assign n14111 = ( ~n6348 & n10493 ) | ( ~n6348 & n14110 ) | ( n10493 & n14110 ) ;
  assign n14112 = ( n2448 & n5680 ) | ( n2448 & ~n6295 ) | ( n5680 & ~n6295 ) ;
  assign n14113 = n2630 | n10043 ;
  assign n14114 = n7362 ^ n5420 ^ 1'b0 ;
  assign n14115 = n3995 & n14114 ;
  assign n14116 = n9490 ^ n5840 ^ 1'b0 ;
  assign n14117 = n14116 ^ n4195 ^ 1'b0 ;
  assign n14118 = n637 | n3369 ;
  assign n14119 = n11425 | n14118 ;
  assign n14120 = n2519 | n9918 ;
  assign n14121 = n2118 & ~n3647 ;
  assign n14122 = n14121 ^ n5223 ^ 1'b0 ;
  assign n14123 = ~n5050 & n14122 ;
  assign n14124 = n14123 ^ n2248 ^ 1'b0 ;
  assign n14125 = n8655 & n14124 ;
  assign n14126 = n828 | n2380 ;
  assign n14127 = n7188 & ~n14126 ;
  assign n14128 = ~n9319 & n14127 ;
  assign n14129 = n631 | n14128 ;
  assign n14130 = n2127 | n2862 ;
  assign n14131 = n14130 ^ n4520 ^ 1'b0 ;
  assign n14132 = n2514 | n14131 ;
  assign n14133 = n14132 ^ n6668 ^ 1'b0 ;
  assign n14134 = ~n2543 & n14133 ;
  assign n14135 = n14134 ^ n2303 ^ 1'b0 ;
  assign n14136 = n8136 | n14135 ;
  assign n14137 = n4560 & n8681 ;
  assign n14138 = ( n286 & n10781 ) | ( n286 & ~n13563 ) | ( n10781 & ~n13563 ) ;
  assign n14139 = n7080 & ~n7118 ;
  assign n14140 = ( ~n6188 & n9788 ) | ( ~n6188 & n14139 ) | ( n9788 & n14139 ) ;
  assign n14141 = ( ~n2221 & n7075 ) | ( ~n2221 & n7303 ) | ( n7075 & n7303 ) ;
  assign n14142 = ~n522 & n926 ;
  assign n14143 = ( ~n1814 & n3423 ) | ( ~n1814 & n14142 ) | ( n3423 & n14142 ) ;
  assign n14144 = n14143 ^ n7593 ^ n4434 ;
  assign n14145 = n14144 ^ n2611 ^ 1'b0 ;
  assign n14146 = ( ~n11058 & n12126 ) | ( ~n11058 & n14145 ) | ( n12126 & n14145 ) ;
  assign n14147 = n4813 | n14146 ;
  assign n14148 = ~n3749 & n7063 ;
  assign n14149 = n14148 ^ n8041 ^ 1'b0 ;
  assign n14152 = n8394 ^ n5153 ^ n3910 ;
  assign n14150 = n1156 | n3183 ;
  assign n14151 = n7112 & n14150 ;
  assign n14153 = n14152 ^ n14151 ^ 1'b0 ;
  assign n14154 = ~n3742 & n14153 ;
  assign n14155 = n14154 ^ n3393 ^ 1'b0 ;
  assign n14156 = n3118 & n4476 ;
  assign n14157 = n674 & n14156 ;
  assign n14158 = n3968 | n4672 ;
  assign n14159 = ~n7041 & n14158 ;
  assign n14160 = ~n3158 & n14159 ;
  assign n14161 = n12055 & n14160 ;
  assign n14162 = n6501 ^ n3330 ^ 1'b0 ;
  assign n14163 = n4380 & n14162 ;
  assign n14164 = n8214 & n9401 ;
  assign n14165 = ~n14163 & n14164 ;
  assign n14166 = n1188 | n10198 ;
  assign n14169 = n1737 & ~n8538 ;
  assign n14167 = ( n2483 & n3072 ) | ( n2483 & ~n5029 ) | ( n3072 & ~n5029 ) ;
  assign n14168 = n14167 ^ n269 ^ 1'b0 ;
  assign n14170 = n14169 ^ n14168 ^ n4100 ;
  assign n14171 = ~n1958 & n3196 ;
  assign n14172 = n9771 ^ n4540 ^ 1'b0 ;
  assign n14173 = n14171 | n14172 ;
  assign n14174 = ~n5400 & n12193 ;
  assign n14175 = n7484 & n14174 ;
  assign n14176 = n14175 ^ n7489 ^ 1'b0 ;
  assign n14177 = n11645 ^ n4973 ^ n2466 ;
  assign n14180 = n539 | n984 ;
  assign n14181 = n14180 ^ n3239 ^ 1'b0 ;
  assign n14182 = n14181 ^ n5634 ^ n4415 ;
  assign n14178 = n2114 ^ n1069 ^ 1'b0 ;
  assign n14179 = n14178 ^ n7646 ^ n6804 ;
  assign n14183 = n14182 ^ n14179 ^ 1'b0 ;
  assign n14184 = n2144 & n10178 ;
  assign n14185 = ~n6207 & n14184 ;
  assign n14186 = n4654 ^ n2766 ^ 1'b0 ;
  assign n14187 = n3430 & ~n14186 ;
  assign n14188 = n14187 ^ n4191 ^ 1'b0 ;
  assign n14189 = n13456 ^ n1124 ^ 1'b0 ;
  assign n14190 = n1451 & ~n14189 ;
  assign n14191 = ~n755 & n8060 ;
  assign n14192 = n14191 ^ n2272 ^ 1'b0 ;
  assign n14193 = n4746 ^ n887 ^ 1'b0 ;
  assign n14194 = n3439 & ~n14193 ;
  assign n14195 = ( n1678 & n5471 ) | ( n1678 & ~n14194 ) | ( n5471 & ~n14194 ) ;
  assign n14196 = ( n4585 & n8306 ) | ( n4585 & ~n14195 ) | ( n8306 & ~n14195 ) ;
  assign n14197 = n13998 ^ n13486 ^ n9709 ;
  assign n14198 = ~n926 & n3267 ;
  assign n14199 = n8029 ^ n1631 ^ 1'b0 ;
  assign n14200 = n8503 | n14199 ;
  assign n14201 = n2846 | n3212 ;
  assign n14202 = ~n5463 & n14201 ;
  assign n14203 = ~x48 & n14202 ;
  assign n14204 = n4342 & n14203 ;
  assign n14205 = n14204 ^ n8912 ^ n8590 ;
  assign n14206 = n9607 | n14205 ;
  assign n14207 = n13631 ^ n8860 ^ 1'b0 ;
  assign n14208 = n5166 ^ n1871 ^ 1'b0 ;
  assign n14209 = n10985 & ~n14208 ;
  assign n14210 = n14209 ^ n6152 ^ 1'b0 ;
  assign n14211 = n9614 ^ n4829 ^ 1'b0 ;
  assign n14212 = ~n12094 & n14211 ;
  assign n14213 = n8977 ^ n3126 ^ 1'b0 ;
  assign n14214 = n14212 & n14213 ;
  assign n14215 = n14214 ^ n11499 ^ 1'b0 ;
  assign n14216 = n9172 | n14215 ;
  assign n14217 = n11398 ^ n4894 ^ n3935 ;
  assign n14218 = x0 & ~n8287 ;
  assign n14219 = ~n12944 & n13649 ;
  assign n14223 = n8054 & n9752 ;
  assign n14220 = x228 | n9201 ;
  assign n14221 = n2058 & n14220 ;
  assign n14222 = n14221 ^ n11861 ^ 1'b0 ;
  assign n14224 = n14223 ^ n14222 ^ n458 ;
  assign n14225 = ~n11056 & n12711 ;
  assign n14226 = n14225 ^ n10326 ^ 1'b0 ;
  assign n14227 = n1546 | n4840 ;
  assign n14228 = n5984 & ~n14227 ;
  assign n14235 = n5099 & n7362 ;
  assign n14236 = ~n6525 & n14235 ;
  assign n14229 = n9196 ^ n6030 ^ 1'b0 ;
  assign n14230 = n14229 ^ n548 ^ 1'b0 ;
  assign n14231 = n4990 | n14230 ;
  assign n14232 = n1648 | n14231 ;
  assign n14233 = n14232 ^ n10761 ^ 1'b0 ;
  assign n14234 = n13229 & n14233 ;
  assign n14237 = n14236 ^ n14234 ^ 1'b0 ;
  assign n14238 = n5629 ^ n1860 ^ 1'b0 ;
  assign n14239 = ~n1851 & n14238 ;
  assign n14240 = n2836 ^ n2618 ^ 1'b0 ;
  assign n14241 = n14240 ^ n502 ^ 1'b0 ;
  assign n14242 = ( n1924 & ~n14239 ) | ( n1924 & n14241 ) | ( ~n14239 & n14241 ) ;
  assign n14243 = x197 ^ x156 ^ 1'b0 ;
  assign n14244 = n14243 ^ n6851 ^ 1'b0 ;
  assign n14245 = n5707 ^ n526 ^ 1'b0 ;
  assign n14246 = n14245 ^ n6719 ^ 1'b0 ;
  assign n14247 = ( n1910 & n7481 ) | ( n1910 & n12070 ) | ( n7481 & n12070 ) ;
  assign n14248 = n2100 & ~n4438 ;
  assign n14249 = n14248 ^ n4582 ^ 1'b0 ;
  assign n14250 = x165 | n14249 ;
  assign n14251 = n5146 ^ n353 ^ 1'b0 ;
  assign n14252 = n274 & ~n11724 ;
  assign n14253 = ~n14251 & n14252 ;
  assign n14254 = n6373 | n13131 ;
  assign n14255 = ( ~n3860 & n4769 ) | ( ~n3860 & n14254 ) | ( n4769 & n14254 ) ;
  assign n14256 = n7016 & ~n9088 ;
  assign n14257 = n10346 & n14256 ;
  assign n14258 = n10932 ^ n692 ^ 1'b0 ;
  assign n14259 = ( n803 & n3413 ) | ( n803 & n14258 ) | ( n3413 & n14258 ) ;
  assign n14266 = n5724 ^ n2882 ^ 1'b0 ;
  assign n14260 = n3695 ^ n480 ^ 1'b0 ;
  assign n14261 = n12723 | n14260 ;
  assign n14262 = ( n7211 & ~n8847 ) | ( n7211 & n13195 ) | ( ~n8847 & n13195 ) ;
  assign n14263 = ~n14261 & n14262 ;
  assign n14264 = ~x193 & n14263 ;
  assign n14265 = n2961 | n14264 ;
  assign n14267 = n14266 ^ n14265 ^ 1'b0 ;
  assign n14268 = n11060 ^ n590 ^ 1'b0 ;
  assign n14269 = n14268 ^ n4173 ^ 1'b0 ;
  assign n14270 = ~n4719 & n5079 ;
  assign n14271 = n5020 & ~n6214 ;
  assign n14272 = ~n2774 & n14271 ;
  assign n14273 = n14272 ^ n5285 ^ 1'b0 ;
  assign n14274 = n7487 ^ n6785 ^ n1997 ;
  assign n14275 = n8821 ^ x204 ^ 1'b0 ;
  assign n14276 = n2585 & n14275 ;
  assign n14277 = n14276 ^ n9281 ^ 1'b0 ;
  assign n14278 = ~n14274 & n14277 ;
  assign n14279 = n11039 ^ n9618 ^ 1'b0 ;
  assign n14280 = ~n6460 & n14279 ;
  assign n14281 = n14280 ^ n752 ^ 1'b0 ;
  assign n14282 = n259 & ~n9451 ;
  assign n14283 = n9451 & n14282 ;
  assign n14284 = n14283 ^ n10548 ^ 1'b0 ;
  assign n14285 = n2542 ^ n1263 ^ n301 ;
  assign n14286 = ( n2138 & n9297 ) | ( n2138 & ~n14285 ) | ( n9297 & ~n14285 ) ;
  assign n14287 = n2320 | n4402 ;
  assign n14288 = n14287 ^ n2071 ^ 1'b0 ;
  assign n14289 = ( x241 & n7177 ) | ( x241 & ~n14288 ) | ( n7177 & ~n14288 ) ;
  assign n14290 = n8965 & n14289 ;
  assign n14291 = n14290 ^ n8472 ^ 1'b0 ;
  assign n14292 = n14291 ^ n14025 ^ 1'b0 ;
  assign n14293 = n14286 | n14292 ;
  assign n14294 = n3981 & ~n7539 ;
  assign n14295 = x189 & n4257 ;
  assign n14296 = n13986 & n14295 ;
  assign n14297 = n4380 & n11420 ;
  assign n14298 = n14297 ^ n4549 ^ 1'b0 ;
  assign n14299 = n14298 ^ n3077 ^ 1'b0 ;
  assign n14300 = n14299 ^ n7439 ^ 1'b0 ;
  assign n14301 = n1678 & n3410 ;
  assign n14302 = n14301 ^ n4446 ^ 1'b0 ;
  assign n14303 = n5952 ^ n2991 ^ 1'b0 ;
  assign n14304 = n14303 ^ n2465 ^ n1501 ;
  assign n14305 = n8352 | n14304 ;
  assign n14306 = n14302 | n14305 ;
  assign n14307 = ~n267 & n14306 ;
  assign n14308 = ~n3737 & n14307 ;
  assign n14309 = n7325 ^ n1233 ^ 1'b0 ;
  assign n14310 = n3671 ^ n704 ^ 1'b0 ;
  assign n14311 = n1073 | n14310 ;
  assign n14312 = n14309 & ~n14311 ;
  assign n14313 = n2781 & n6401 ;
  assign n14314 = n2793 & ~n2806 ;
  assign n14315 = n14314 ^ n7398 ^ 1'b0 ;
  assign n14316 = n851 & n14315 ;
  assign n14317 = n8252 & n14316 ;
  assign n14318 = n14317 ^ n4194 ^ 1'b0 ;
  assign n14319 = n5903 & n9169 ;
  assign n14320 = n4672 & n11201 ;
  assign n14321 = n967 & n2738 ;
  assign n14322 = n2194 | n14321 ;
  assign n14323 = n14322 ^ n3951 ^ 1'b0 ;
  assign n14324 = ~n2463 & n14323 ;
  assign n14325 = n851 & n4776 ;
  assign n14326 = n7016 & n14325 ;
  assign n14327 = n2307 | n9802 ;
  assign n14328 = n14327 ^ n5232 ^ 1'b0 ;
  assign n14331 = n1750 | n4018 ;
  assign n14329 = n3278 & n9363 ;
  assign n14330 = n13424 & n14329 ;
  assign n14332 = n14331 ^ n14330 ^ 1'b0 ;
  assign n14333 = n7029 ^ n1260 ^ 1'b0 ;
  assign n14334 = n4356 & ~n14333 ;
  assign n14335 = ~n13487 & n13867 ;
  assign n14337 = n1571 | n3233 ;
  assign n14336 = ~n3207 & n3738 ;
  assign n14338 = n14337 ^ n14336 ^ 1'b0 ;
  assign n14339 = n2836 & n11573 ;
  assign n14340 = n14339 ^ n13801 ^ n2858 ;
  assign n14341 = ( n647 & n1944 ) | ( n647 & n7519 ) | ( n1944 & n7519 ) ;
  assign n14342 = ~n14340 & n14341 ;
  assign n14343 = n3889 & n5770 ;
  assign n14344 = ( n1312 & ~n2486 ) | ( n1312 & n14343 ) | ( ~n2486 & n14343 ) ;
  assign n14345 = n8942 & ~n14344 ;
  assign n14346 = n14345 ^ n7259 ^ 1'b0 ;
  assign n14347 = n1315 & ~n9804 ;
  assign n14349 = n1037 | n5457 ;
  assign n14348 = n3843 & n8100 ;
  assign n14350 = n14349 ^ n14348 ^ 1'b0 ;
  assign n14351 = n5102 & n5649 ;
  assign n14352 = ~n9209 & n14351 ;
  assign n14353 = ~n5672 & n10824 ;
  assign n14354 = ~n3218 & n14353 ;
  assign n14355 = n6303 & ~n6502 ;
  assign n14356 = ~n5660 & n14355 ;
  assign n14357 = n4817 & n11316 ;
  assign n14358 = n4655 ^ n1726 ^ 1'b0 ;
  assign n14359 = ~n1532 & n14358 ;
  assign n14360 = n6526 & n14359 ;
  assign n14361 = n12080 & n14360 ;
  assign n14362 = n8834 | n14361 ;
  assign n14363 = n2497 & ~n11127 ;
  assign n14364 = n9367 & n14363 ;
  assign n14365 = n11062 ^ n5469 ^ 1'b0 ;
  assign n14366 = ~n4633 & n14365 ;
  assign n14367 = n14366 ^ n10185 ^ n7068 ;
  assign n14368 = ( n3747 & n4580 ) | ( n3747 & ~n6153 ) | ( n4580 & ~n6153 ) ;
  assign n14369 = ~n4194 & n14368 ;
  assign n14370 = n14369 ^ n704 ^ 1'b0 ;
  assign n14371 = n10503 ^ n9848 ^ 1'b0 ;
  assign n14372 = n1636 & ~n14371 ;
  assign n14373 = n7013 ^ n6594 ^ n685 ;
  assign n14374 = ( ~n467 & n5799 ) | ( ~n467 & n5976 ) | ( n5799 & n5976 ) ;
  assign n14375 = n5063 & n14374 ;
  assign n14376 = ~n2860 & n6134 ;
  assign n14377 = n14376 ^ n11326 ^ 1'b0 ;
  assign n14378 = ~n8159 & n14377 ;
  assign n14379 = n1068 | n14378 ;
  assign n14380 = n12456 ^ n7139 ^ 1'b0 ;
  assign n14381 = n13024 ^ n8833 ^ 1'b0 ;
  assign n14382 = n3962 & n14381 ;
  assign n14383 = ( n7409 & n13793 ) | ( n7409 & n14382 ) | ( n13793 & n14382 ) ;
  assign n14384 = n12184 ^ n4664 ^ 1'b0 ;
  assign n14385 = n7418 & ~n14384 ;
  assign n14386 = n1256 & n14385 ;
  assign n14387 = n9034 & n14386 ;
  assign n14388 = n2243 & n5519 ;
  assign n14389 = n8803 ^ n5982 ^ 1'b0 ;
  assign n14390 = ~n14388 & n14389 ;
  assign n14391 = n14390 ^ n4029 ^ 1'b0 ;
  assign n14392 = n14387 | n14391 ;
  assign n14393 = n3239 ^ n2715 ^ 1'b0 ;
  assign n14394 = n8187 & ~n14393 ;
  assign n14395 = n12671 ^ n2807 ^ 1'b0 ;
  assign n14396 = ( n886 & n7068 ) | ( n886 & ~n7690 ) | ( n7068 & ~n7690 ) ;
  assign n14397 = n14396 ^ n12550 ^ n7670 ;
  assign n14398 = n987 & n14397 ;
  assign n14399 = n14395 & n14398 ;
  assign n14400 = n9390 & ~n14399 ;
  assign n14401 = n14400 ^ n12400 ^ 1'b0 ;
  assign n14402 = n773 & ~n9858 ;
  assign n14403 = n14402 ^ n2751 ^ 1'b0 ;
  assign n14404 = n14403 ^ n8886 ^ 1'b0 ;
  assign n14405 = n6337 & n14404 ;
  assign n14406 = ~n9540 & n14405 ;
  assign n14407 = n8544 & ~n11640 ;
  assign n14408 = n14407 ^ n11986 ^ 1'b0 ;
  assign n14409 = n1907 & ~n13230 ;
  assign n14410 = n14409 ^ n5133 ^ 1'b0 ;
  assign n14411 = ( n1225 & n3201 ) | ( n1225 & n14410 ) | ( n3201 & n14410 ) ;
  assign n14412 = n14411 ^ n13941 ^ 1'b0 ;
  assign n14413 = ~n6827 & n7637 ;
  assign n14414 = n3808 & n14413 ;
  assign n14415 = x111 & ~n14414 ;
  assign n14416 = ~n2698 & n14415 ;
  assign n14417 = n14416 ^ n8320 ^ 1'b0 ;
  assign n14418 = ( n1705 & n2824 ) | ( n1705 & n6081 ) | ( n2824 & n6081 ) ;
  assign n14419 = n4064 | n14418 ;
  assign n14420 = n5226 | n9375 ;
  assign n14421 = n14420 ^ n4809 ^ 1'b0 ;
  assign n14422 = ( n1589 & n11897 ) | ( n1589 & ~n14421 ) | ( n11897 & ~n14421 ) ;
  assign n14423 = x115 & ~n4613 ;
  assign n14424 = n14423 ^ n11461 ^ 1'b0 ;
  assign n14425 = ( n5045 & ~n9207 ) | ( n5045 & n11287 ) | ( ~n9207 & n11287 ) ;
  assign n14426 = n4247 & ~n7314 ;
  assign n14427 = ~x241 & n14426 ;
  assign n14428 = n14321 & ~n14427 ;
  assign n14429 = n14428 ^ n3978 ^ 1'b0 ;
  assign n14430 = n7429 ^ n351 ^ 1'b0 ;
  assign n14431 = ~n749 & n6352 ;
  assign n14432 = n2292 & n14431 ;
  assign n14433 = n932 & ~n14432 ;
  assign n14434 = n14433 ^ n790 ^ 1'b0 ;
  assign n14435 = n14434 ^ n4887 ^ 1'b0 ;
  assign n14436 = n5899 | n9236 ;
  assign n14437 = n14436 ^ n5556 ^ 1'b0 ;
  assign n14438 = ~n291 & n14437 ;
  assign n14439 = ~n2687 & n14438 ;
  assign n14440 = n2578 ^ n504 ^ 1'b0 ;
  assign n14441 = n4300 | n14440 ;
  assign n14442 = n14441 ^ n1553 ^ 1'b0 ;
  assign n14443 = n1993 | n14442 ;
  assign n14444 = n4081 & ~n4548 ;
  assign n14445 = n14444 ^ n14258 ^ 1'b0 ;
  assign n14446 = n14445 ^ n5211 ^ n4558 ;
  assign n14447 = n14446 ^ n326 ^ 1'b0 ;
  assign n14448 = n14446 & n14447 ;
  assign n14449 = n14448 ^ n10406 ^ n8921 ;
  assign n14450 = n13981 ^ n8239 ^ n3225 ;
  assign n14451 = n5051 & ~n14450 ;
  assign n14452 = ~n583 & n1197 ;
  assign n14453 = n4852 ^ n2463 ^ 1'b0 ;
  assign n14454 = n14452 | n14453 ;
  assign n14455 = n6409 | n8654 ;
  assign n14456 = n14454 & ~n14455 ;
  assign n14457 = n14451 & ~n14456 ;
  assign n14458 = n10443 & n14457 ;
  assign n14459 = n12251 ^ n5131 ^ 1'b0 ;
  assign n14460 = n14458 | n14459 ;
  assign n14461 = n3256 ^ n1951 ^ 1'b0 ;
  assign n14462 = n5832 & n14461 ;
  assign n14463 = n11438 & n14462 ;
  assign n14464 = ~n1762 & n8655 ;
  assign n14465 = n14463 & n14464 ;
  assign n14466 = n14465 ^ n2155 ^ 1'b0 ;
  assign n14467 = ~n10501 & n14466 ;
  assign n14468 = n13467 ^ n6398 ^ n2055 ;
  assign n14469 = n10109 ^ n9322 ^ 1'b0 ;
  assign n14470 = n6565 & ~n14469 ;
  assign n14471 = n271 & ~n5695 ;
  assign n14472 = n12373 ^ n4920 ^ 1'b0 ;
  assign n14473 = n1433 & ~n14472 ;
  assign n14474 = n2548 & ~n11596 ;
  assign n14475 = n2895 & n14474 ;
  assign n14476 = ~n3056 & n14475 ;
  assign n14477 = n14476 ^ n9995 ^ 1'b0 ;
  assign n14478 = n4729 & n7863 ;
  assign n14479 = ~n13212 & n14478 ;
  assign n14480 = n14479 ^ n6111 ^ 1'b0 ;
  assign n14481 = n11458 & n14480 ;
  assign n14482 = n2525 ^ n1630 ^ n338 ;
  assign n14483 = n14482 ^ n2002 ^ 1'b0 ;
  assign n14485 = x78 | n1253 ;
  assign n14486 = n14485 ^ n4312 ^ 1'b0 ;
  assign n14484 = n451 & ~n6820 ;
  assign n14487 = n14486 ^ n14484 ^ 1'b0 ;
  assign n14488 = n9556 & ~n14487 ;
  assign n14489 = ~n14483 & n14488 ;
  assign n14490 = n14489 ^ n9529 ^ n1887 ;
  assign n14491 = n6458 & ~n9957 ;
  assign n14492 = n5772 | n14491 ;
  assign n14493 = n2221 | n14492 ;
  assign n14494 = ~n6292 & n9118 ;
  assign n14495 = n14494 ^ x138 ^ 1'b0 ;
  assign n14496 = n2823 | n5605 ;
  assign n14497 = n14496 ^ n4349 ^ 1'b0 ;
  assign n14498 = ~n4298 & n14497 ;
  assign n14499 = n14498 ^ n286 ^ 1'b0 ;
  assign n14500 = n10089 | n14499 ;
  assign n14501 = x144 & n7230 ;
  assign n14502 = n14501 ^ n3740 ^ 1'b0 ;
  assign n14503 = n14502 ^ n2227 ^ 1'b0 ;
  assign n14504 = n9011 & n14503 ;
  assign n14505 = n14504 ^ n1712 ^ 1'b0 ;
  assign n14506 = n11772 ^ n8244 ^ n5372 ;
  assign n14507 = n2081 & ~n4860 ;
  assign n14508 = n1728 | n14507 ;
  assign n14509 = ( ~n6982 & n14506 ) | ( ~n6982 & n14508 ) | ( n14506 & n14508 ) ;
  assign n14510 = n1330 & ~n5321 ;
  assign n14511 = n1957 | n7321 ;
  assign n14512 = n1213 & n14511 ;
  assign n14513 = n14512 ^ n372 ^ 1'b0 ;
  assign n14514 = n14510 | n14513 ;
  assign n14515 = n14514 ^ n6069 ^ 1'b0 ;
  assign n14516 = ~n2401 & n4012 ;
  assign n14517 = n14516 ^ n6630 ^ 1'b0 ;
  assign n14518 = ~n7917 & n14517 ;
  assign n14519 = n3322 & n6435 ;
  assign n14520 = n7607 & n14519 ;
  assign n14521 = n14520 ^ n6191 ^ n6019 ;
  assign n14522 = n288 | n5411 ;
  assign n14523 = n4508 & ~n14522 ;
  assign n14524 = n4828 & ~n14523 ;
  assign n14525 = ~n11577 & n14524 ;
  assign n14526 = n7558 & ~n8567 ;
  assign n14527 = ~n4180 & n14526 ;
  assign n14528 = n6370 ^ n3548 ^ 1'b0 ;
  assign n14529 = n7342 ^ n3300 ^ 1'b0 ;
  assign n14530 = n10498 & n14529 ;
  assign n14531 = ~x56 & n14530 ;
  assign n14532 = n14528 & n14531 ;
  assign n14533 = ~n11417 & n14532 ;
  assign n14534 = ~n3927 & n14417 ;
  assign n14537 = n14310 ^ n2737 ^ 1'b0 ;
  assign n14535 = n1961 & ~n9640 ;
  assign n14536 = ~n2243 & n14535 ;
  assign n14538 = n14537 ^ n14536 ^ 1'b0 ;
  assign n14539 = n14538 ^ n589 ^ 1'b0 ;
  assign n14540 = n8690 ^ n2365 ^ 1'b0 ;
  assign n14541 = n4764 & ~n13549 ;
  assign n14542 = ~n9932 & n14541 ;
  assign n14543 = n5720 & n14542 ;
  assign n14544 = n1246 & ~n11786 ;
  assign n14545 = n14544 ^ n3734 ^ 1'b0 ;
  assign n14546 = n14545 ^ n3645 ^ 1'b0 ;
  assign n14547 = ~n14543 & n14546 ;
  assign n14548 = ( n1519 & ~n6766 ) | ( n1519 & n9600 ) | ( ~n6766 & n9600 ) ;
  assign n14549 = ( n328 & n6297 ) | ( n328 & n7322 ) | ( n6297 & n7322 ) ;
  assign n14550 = n4652 | n14549 ;
  assign n14551 = n3291 & n7338 ;
  assign n14552 = n14551 ^ n413 ^ 1'b0 ;
  assign n14553 = n6432 & n14552 ;
  assign n14554 = n420 | n5162 ;
  assign n14555 = n6194 | n14554 ;
  assign n14556 = n13744 | n14555 ;
  assign n14557 = n1782 ^ x52 ^ 1'b0 ;
  assign n14558 = n2173 | n14557 ;
  assign n14559 = ~n2950 & n14558 ;
  assign n14560 = n758 & n14559 ;
  assign n14564 = n2286 | n12766 ;
  assign n14565 = n7049 & ~n14564 ;
  assign n14566 = ~n9880 & n14565 ;
  assign n14561 = ~n5972 & n7170 ;
  assign n14562 = ~n8306 & n14561 ;
  assign n14563 = n14562 ^ n6468 ^ 1'b0 ;
  assign n14567 = n14566 ^ n14563 ^ 1'b0 ;
  assign n14568 = n5685 | n11947 ;
  assign n14569 = n14568 ^ n4764 ^ 1'b0 ;
  assign n14572 = n1996 ^ n258 ^ 1'b0 ;
  assign n14570 = n2133 ^ n322 ^ 1'b0 ;
  assign n14571 = ( ~n5468 & n11976 ) | ( ~n5468 & n14570 ) | ( n11976 & n14570 ) ;
  assign n14573 = n14572 ^ n14571 ^ 1'b0 ;
  assign n14574 = n13013 | n14573 ;
  assign n14575 = n11262 & ~n12386 ;
  assign n14576 = ~n5628 & n14575 ;
  assign n14577 = n10992 | n14576 ;
  assign n14578 = n14574 & ~n14577 ;
  assign n14579 = n6686 & ~n8951 ;
  assign n14580 = n9067 & n14579 ;
  assign n14581 = n14580 ^ x230 ^ 1'b0 ;
  assign n14582 = n1024 & n1072 ;
  assign n14583 = n14582 ^ n5327 ^ 1'b0 ;
  assign n14584 = n3128 & ~n14583 ;
  assign n14585 = ~n6672 & n14584 ;
  assign n14586 = n11989 & n14585 ;
  assign n14591 = n12004 ^ n11160 ^ n10019 ;
  assign n14587 = n2959 & n7458 ;
  assign n14588 = ~n3850 & n9731 ;
  assign n14589 = n14588 ^ n4703 ^ 1'b0 ;
  assign n14590 = ~n14587 & n14589 ;
  assign n14592 = n14591 ^ n14590 ^ 1'b0 ;
  assign n14593 = n7370 & n8737 ;
  assign n14594 = ( ~n3170 & n7945 ) | ( ~n3170 & n12382 ) | ( n7945 & n12382 ) ;
  assign n14595 = n6141 | n8828 ;
  assign n14596 = n12756 | n14595 ;
  assign n14597 = ~n2538 & n9822 ;
  assign n14598 = n14597 ^ n5544 ^ 1'b0 ;
  assign n14602 = n6694 & ~n8956 ;
  assign n14603 = n3369 ^ n385 ^ 1'b0 ;
  assign n14604 = n14602 & ~n14603 ;
  assign n14599 = n463 & ~n12853 ;
  assign n14600 = ~n681 & n14599 ;
  assign n14601 = n14600 ^ n10112 ^ 1'b0 ;
  assign n14605 = n14604 ^ n14601 ^ n11705 ;
  assign n14606 = n743 ^ n581 ^ 1'b0 ;
  assign n14607 = n14606 ^ n14477 ^ 1'b0 ;
  assign n14608 = n8913 & ~n9748 ;
  assign n14609 = n14608 ^ n11103 ^ 1'b0 ;
  assign n14610 = n1168 | n3093 ;
  assign n14611 = n14610 ^ n11610 ^ 1'b0 ;
  assign n14612 = n14609 & n14611 ;
  assign n14613 = n7336 ^ n7271 ^ 1'b0 ;
  assign n14615 = n1401 & ~n1742 ;
  assign n14616 = n14615 ^ n2608 ^ 1'b0 ;
  assign n14617 = n2521 & ~n14616 ;
  assign n14614 = x73 & n2527 ;
  assign n14618 = n14617 ^ n14614 ^ 1'b0 ;
  assign n14619 = n7128 | n14618 ;
  assign n14620 = n1807 ^ n1153 ^ 1'b0 ;
  assign n14621 = n14619 | n14620 ;
  assign n14622 = n6147 ^ n5235 ^ 1'b0 ;
  assign n14623 = n8016 & ~n14622 ;
  assign n14624 = n14623 ^ n2896 ^ 1'b0 ;
  assign n14625 = n4829 & n9715 ;
  assign n14626 = ~n4981 & n6091 ;
  assign n14627 = ~n14625 & n14626 ;
  assign n14628 = n7861 ^ n3467 ^ 1'b0 ;
  assign n14629 = ~n12160 & n14628 ;
  assign n14630 = ~n3362 & n4670 ;
  assign n14631 = n12080 ^ n5830 ^ 1'b0 ;
  assign n14632 = n14631 ^ n10851 ^ 1'b0 ;
  assign n14633 = n3542 | n6214 ;
  assign n14634 = n1590 & ~n14633 ;
  assign n14635 = n14634 ^ n8262 ^ 1'b0 ;
  assign n14636 = n11878 ^ n10989 ^ 1'b0 ;
  assign n14637 = n399 | n1982 ;
  assign n14638 = n14637 ^ n8880 ^ 1'b0 ;
  assign n14639 = n14638 ^ n4423 ^ 1'b0 ;
  assign n14640 = n14636 | n14639 ;
  assign n14641 = n14640 ^ n6029 ^ 1'b0 ;
  assign n14642 = n14641 ^ n5169 ^ 1'b0 ;
  assign n14643 = n2935 | n6480 ;
  assign n14644 = n4996 | n14643 ;
  assign n14645 = n14644 ^ n861 ^ 1'b0 ;
  assign n14646 = n5675 ^ n2298 ^ n856 ;
  assign n14647 = ~n1233 & n14646 ;
  assign n14648 = n5680 & n14647 ;
  assign n14649 = n2829 | n14648 ;
  assign n14650 = n14649 ^ n13740 ^ 1'b0 ;
  assign n14654 = n2556 & ~n2868 ;
  assign n14655 = n1851 & n14654 ;
  assign n14656 = n14655 ^ n2673 ^ 1'b0 ;
  assign n14657 = n14656 ^ x206 ^ 1'b0 ;
  assign n14658 = n14657 ^ n2890 ^ 1'b0 ;
  assign n14659 = n4711 & ~n14658 ;
  assign n14651 = n4065 & ~n12315 ;
  assign n14652 = ~n6954 & n14651 ;
  assign n14653 = n2907 | n14652 ;
  assign n14660 = n14659 ^ n14653 ^ 1'b0 ;
  assign n14661 = n11477 ^ n5182 ^ 1'b0 ;
  assign n14662 = n10129 & n14661 ;
  assign n14663 = ~n6589 & n6775 ;
  assign n14664 = n14663 ^ n6502 ^ 1'b0 ;
  assign n14665 = ~n4976 & n14664 ;
  assign n14666 = ~n3447 & n5393 ;
  assign n14668 = n14410 ^ n3672 ^ 1'b0 ;
  assign n14667 = n1679 ^ n616 ^ 1'b0 ;
  assign n14669 = n14668 ^ n14667 ^ 1'b0 ;
  assign n14670 = n4573 ^ n3043 ^ 1'b0 ;
  assign n14671 = n2058 & n14670 ;
  assign n14672 = n14671 ^ n12678 ^ n11212 ;
  assign n14673 = n6937 ^ n1166 ^ 1'b0 ;
  assign n14674 = n4463 | n11175 ;
  assign n14675 = n13039 & ~n14674 ;
  assign n14676 = n3051 | n14675 ;
  assign n14677 = n1044 | n14676 ;
  assign n14678 = ~n1608 & n10015 ;
  assign n14679 = ~n9380 & n14678 ;
  assign n14680 = n1512 & n10884 ;
  assign n14681 = n14680 ^ n7035 ^ 1'b0 ;
  assign n14682 = n2165 ^ n1455 ^ 1'b0 ;
  assign n14683 = n3032 & n14682 ;
  assign n14684 = n14683 ^ x2 ^ 1'b0 ;
  assign n14685 = ~n3985 & n14684 ;
  assign n14686 = ~n4238 & n6881 ;
  assign n14687 = n14686 ^ n5922 ^ 1'b0 ;
  assign n14688 = n14687 ^ n11413 ^ 1'b0 ;
  assign n14689 = n14685 & n14688 ;
  assign n14693 = ~n1291 & n5970 ;
  assign n14690 = n1130 & n6174 ;
  assign n14691 = n14480 ^ n10880 ^ n4072 ;
  assign n14692 = n14690 & n14691 ;
  assign n14694 = n14693 ^ n14692 ^ 1'b0 ;
  assign n14695 = n8630 | n8969 ;
  assign n14696 = n14695 ^ n685 ^ 1'b0 ;
  assign n14700 = n9496 & n10872 ;
  assign n14701 = n8125 & n14700 ;
  assign n14702 = n13357 | n14701 ;
  assign n14703 = n14702 ^ n8608 ^ 1'b0 ;
  assign n14697 = n2853 ^ n919 ^ 1'b0 ;
  assign n14698 = n14697 ^ n6397 ^ 1'b0 ;
  assign n14699 = ~n13043 & n14698 ;
  assign n14704 = n14703 ^ n14699 ^ 1'b0 ;
  assign n14705 = n14704 ^ n5217 ^ 1'b0 ;
  assign n14706 = ~n14696 & n14705 ;
  assign n14707 = n3982 & ~n7149 ;
  assign n14708 = ~x88 & n14707 ;
  assign n14709 = n14708 ^ n9029 ^ 1'b0 ;
  assign n14710 = n5680 ^ n4626 ^ 1'b0 ;
  assign n14711 = n4448 ^ n1611 ^ n629 ;
  assign n14712 = n13596 & n14711 ;
  assign n14713 = n14712 ^ n10777 ^ 1'b0 ;
  assign n14714 = n7756 ^ n4471 ^ n1236 ;
  assign n14715 = n14714 ^ n9975 ^ n4066 ;
  assign n14716 = ( n7386 & n14713 ) | ( n7386 & ~n14715 ) | ( n14713 & ~n14715 ) ;
  assign n14717 = n1808 | n2209 ;
  assign n14718 = n7316 | n14717 ;
  assign n14719 = n3511 ^ n2684 ^ 1'b0 ;
  assign n14720 = ( n5151 & ~n14718 ) | ( n5151 & n14719 ) | ( ~n14718 & n14719 ) ;
  assign n14721 = n5773 & n8783 ;
  assign n14722 = n6041 & n14721 ;
  assign n14723 = n14722 ^ n5531 ^ 1'b0 ;
  assign n14724 = ~n2033 & n5980 ;
  assign n14725 = n12102 ^ n1866 ^ 1'b0 ;
  assign n14726 = n9084 | n14725 ;
  assign n14727 = n6379 | n10790 ;
  assign n14728 = n1031 & ~n14727 ;
  assign n14729 = n9200 & ~n14728 ;
  assign n14730 = n14729 ^ n9475 ^ 1'b0 ;
  assign n14731 = n14730 ^ n9032 ^ n4036 ;
  assign n14732 = n1525 & ~n7880 ;
  assign n14733 = n14732 ^ n882 ^ 1'b0 ;
  assign n14734 = n5271 & ~n6553 ;
  assign n14735 = n5961 | n14734 ;
  assign n14736 = n9518 ^ n4587 ^ 1'b0 ;
  assign n14737 = n5751 & n14736 ;
  assign n14738 = ~n7861 & n14737 ;
  assign n14739 = ( n427 & ~n6146 ) | ( n427 & n14738 ) | ( ~n6146 & n14738 ) ;
  assign n14740 = n8642 ^ n2518 ^ 1'b0 ;
  assign n14741 = n979 & n14740 ;
  assign n14742 = ~n10593 & n14741 ;
  assign n14743 = n9003 ^ n8011 ^ n5463 ;
  assign n14744 = n2902 & n14743 ;
  assign n14745 = n7570 & ~n9367 ;
  assign n14746 = n14745 ^ n3517 ^ 1'b0 ;
  assign n14747 = n7044 & ~n9666 ;
  assign n14748 = n14062 ^ n1001 ^ 1'b0 ;
  assign n14749 = ( n1067 & n14747 ) | ( n1067 & ~n14748 ) | ( n14747 & ~n14748 ) ;
  assign n14750 = n3976 ^ n1679 ^ 1'b0 ;
  assign n14751 = n14750 ^ n4000 ^ 1'b0 ;
  assign n14752 = n12580 ^ n11308 ^ 1'b0 ;
  assign n14753 = n4128 & ~n4832 ;
  assign n14754 = n7833 ^ x236 ^ 1'b0 ;
  assign n14763 = n3274 & ~n4096 ;
  assign n14764 = n14763 ^ n4261 ^ 1'b0 ;
  assign n14759 = n2326 & n9374 ;
  assign n14760 = ~n6232 & n14759 ;
  assign n14755 = n432 | n1258 ;
  assign n14756 = n14755 ^ n8516 ^ 1'b0 ;
  assign n14757 = x143 & ~n14756 ;
  assign n14758 = n14757 ^ n1072 ^ 1'b0 ;
  assign n14761 = n14760 ^ n14758 ^ 1'b0 ;
  assign n14762 = ~n1411 & n14761 ;
  assign n14765 = n14764 ^ n14762 ^ 1'b0 ;
  assign n14766 = n2153 & n13477 ;
  assign n14767 = ~n1993 & n4604 ;
  assign n14768 = n8606 & n14767 ;
  assign n14769 = n5649 | n6241 ;
  assign n14770 = ( ~n2113 & n2275 ) | ( ~n2113 & n14769 ) | ( n2275 & n14769 ) ;
  assign n14771 = n14770 ^ n9919 ^ n9865 ;
  assign n14772 = n14771 ^ n9986 ^ n3077 ;
  assign n14773 = n1101 | n4371 ;
  assign n14774 = n3924 | n7226 ;
  assign n14775 = n14774 ^ n6448 ^ 1'b0 ;
  assign n14776 = ~n5735 & n10064 ;
  assign n14777 = n3483 & ~n6531 ;
  assign n14778 = n14777 ^ n14205 ^ 1'b0 ;
  assign n14779 = n5324 & ~n10193 ;
  assign n14780 = ~n5065 & n14779 ;
  assign n14781 = n14780 ^ n10248 ^ 1'b0 ;
  assign n14782 = n11149 & n14781 ;
  assign n14786 = n3782 | n11701 ;
  assign n14783 = ( n2224 & n3041 ) | ( n2224 & n8377 ) | ( n3041 & n8377 ) ;
  assign n14784 = n9820 & ~n14783 ;
  assign n14785 = x251 & n14784 ;
  assign n14787 = n14786 ^ n14785 ^ 1'b0 ;
  assign n14788 = n6141 & n14787 ;
  assign n14789 = ~n9800 & n14788 ;
  assign n14790 = ~n690 & n1806 ;
  assign n14791 = n14790 ^ n7859 ^ 1'b0 ;
  assign n14792 = x9 & ~n14791 ;
  assign n14793 = n11454 & ~n14792 ;
  assign n14794 = n14793 ^ n11189 ^ 1'b0 ;
  assign n14795 = n8471 & ~n14794 ;
  assign n14796 = n2650 ^ n2436 ^ 1'b0 ;
  assign n14797 = n13211 ^ n8627 ^ 1'b0 ;
  assign n14798 = ~n354 & n14797 ;
  assign n14799 = n9694 ^ n3709 ^ 1'b0 ;
  assign n14800 = n7015 & ~n12678 ;
  assign n14801 = n14800 ^ n9128 ^ 1'b0 ;
  assign n14802 = ( n4966 & n5143 ) | ( n4966 & ~n9144 ) | ( n5143 & ~n9144 ) ;
  assign n14803 = n6945 & n14802 ;
  assign n14804 = n928 | n5800 ;
  assign n14805 = x228 | n7033 ;
  assign n14806 = n6565 | n6606 ;
  assign n14807 = n4480 & ~n14806 ;
  assign n14808 = n6732 | n14807 ;
  assign n14809 = n14805 & ~n14808 ;
  assign n14810 = n1813 | n14809 ;
  assign n14811 = n7924 & ~n14810 ;
  assign n14812 = n9786 ^ n5836 ^ 1'b0 ;
  assign n14813 = n12256 & n14812 ;
  assign n14814 = n7380 ^ n397 ^ x246 ;
  assign n14815 = n4608 ^ n3806 ^ 1'b0 ;
  assign n14816 = n8078 ^ n4620 ^ n3498 ;
  assign n14818 = n5127 & ~n10221 ;
  assign n14817 = n12974 ^ n5981 ^ 1'b0 ;
  assign n14819 = n14818 ^ n14817 ^ 1'b0 ;
  assign n14820 = x159 & n14819 ;
  assign n14821 = ~n14816 & n14820 ;
  assign n14827 = x16 & x234 ;
  assign n14828 = n3872 & n14827 ;
  assign n14822 = ~n2262 & n5302 ;
  assign n14823 = n2262 & n14822 ;
  assign n14824 = n4100 & ~n14823 ;
  assign n14825 = ~n4100 & n14824 ;
  assign n14826 = n6766 | n14825 ;
  assign n14829 = n14828 ^ n14826 ^ n12053 ;
  assign n14830 = ~n2336 & n8197 ;
  assign n14831 = n14437 ^ n10767 ^ 1'b0 ;
  assign n14832 = n12867 ^ n2787 ^ 1'b0 ;
  assign n14833 = ~n5793 & n14832 ;
  assign n14834 = n9541 & ~n14833 ;
  assign n14835 = ~n1932 & n14834 ;
  assign n14836 = n588 | n4981 ;
  assign n14837 = n2839 & ~n14836 ;
  assign n14838 = ~n5194 & n13006 ;
  assign n14839 = n610 | n7146 ;
  assign n14840 = n12725 ^ n261 ^ 1'b0 ;
  assign n14841 = n5439 & n14840 ;
  assign n14842 = x41 | n1717 ;
  assign n14843 = n12931 ^ n10863 ^ 1'b0 ;
  assign n14844 = n6944 & ~n14843 ;
  assign n14845 = n12614 ^ n7866 ^ n1965 ;
  assign n14846 = n7113 ^ n1486 ^ 1'b0 ;
  assign n14848 = n2664 ^ n1930 ^ 1'b0 ;
  assign n14847 = n1544 & ~n11532 ;
  assign n14849 = n14848 ^ n14847 ^ 1'b0 ;
  assign n14850 = n14849 ^ n11723 ^ 1'b0 ;
  assign n14851 = n14846 & n14850 ;
  assign n14852 = n1944 | n5037 ;
  assign n14853 = n1625 ^ n425 ^ 1'b0 ;
  assign n14854 = n14852 & n14853 ;
  assign n14855 = n1098 & ~n1680 ;
  assign n14856 = n5098 ^ n1223 ^ 1'b0 ;
  assign n14857 = ~n8592 & n14856 ;
  assign n14858 = n14857 ^ x237 ^ 1'b0 ;
  assign n14859 = n14855 & ~n14858 ;
  assign n14860 = n10428 ^ n6829 ^ n3286 ;
  assign n14861 = n1880 & n2372 ;
  assign n14862 = n14861 ^ n7670 ^ 1'b0 ;
  assign n14863 = n14862 ^ n10250 ^ 1'b0 ;
  assign n14864 = n3024 & n7184 ;
  assign n14865 = n3666 & n14864 ;
  assign n14866 = n5558 | n14865 ;
  assign n14867 = n14866 ^ n988 ^ 1'b0 ;
  assign n14869 = ( n854 & n1910 ) | ( n854 & ~n12308 ) | ( n1910 & ~n12308 ) ;
  assign n14868 = n302 | n3777 ;
  assign n14870 = n14869 ^ n14868 ^ n12185 ;
  assign n14871 = n6448 & ~n9930 ;
  assign n14872 = n14871 ^ n14733 ^ 1'b0 ;
  assign n14873 = ( ~n6203 & n6319 ) | ( ~n6203 & n9026 ) | ( n6319 & n9026 ) ;
  assign n14874 = n14873 ^ n8602 ^ 1'b0 ;
  assign n14875 = n7004 & ~n14874 ;
  assign n14876 = n758 & ~n5127 ;
  assign n14877 = ( x139 & ~n6035 ) | ( x139 & n14876 ) | ( ~n6035 & n14876 ) ;
  assign n14878 = n13189 ^ n6075 ^ 1'b0 ;
  assign n14879 = n8328 & ~n14878 ;
  assign n14880 = ~n2649 & n10560 ;
  assign n14881 = n14880 ^ n13708 ^ 1'b0 ;
  assign n14882 = n4056 & ~n12788 ;
  assign n14883 = ~n1932 & n14882 ;
  assign n14884 = n7602 ^ n7374 ^ 1'b0 ;
  assign n14885 = n14884 ^ n8930 ^ 1'b0 ;
  assign n14886 = n3450 & ~n14885 ;
  assign n14892 = n14790 ^ n4135 ^ 1'b0 ;
  assign n14887 = n4561 | n5724 ;
  assign n14888 = n10941 & n14887 ;
  assign n14889 = n14888 ^ n3369 ^ 1'b0 ;
  assign n14890 = n5772 | n14889 ;
  assign n14891 = n14890 ^ n1177 ^ 1'b0 ;
  assign n14893 = n14892 ^ n14891 ^ 1'b0 ;
  assign n14894 = n5861 & ~n14893 ;
  assign n14895 = n14212 & ~n14894 ;
  assign n14896 = n5536 ^ n3759 ^ n2882 ;
  assign n14897 = n14896 ^ n3647 ^ 1'b0 ;
  assign n14898 = n8632 & n14897 ;
  assign n14899 = ~n9566 & n11319 ;
  assign n14900 = n341 & n14899 ;
  assign n14901 = n2078 ^ n623 ^ 1'b0 ;
  assign n14902 = n5805 ^ n2807 ^ 1'b0 ;
  assign n14903 = n12169 & ~n14902 ;
  assign n14904 = n14903 ^ n1473 ^ 1'b0 ;
  assign n14905 = n2575 ^ n2036 ^ 1'b0 ;
  assign n14906 = n9987 ^ n4319 ^ 1'b0 ;
  assign n14907 = n14905 & n14906 ;
  assign n14908 = n1943 & ~n2986 ;
  assign n14914 = n11237 ^ n7554 ^ n2473 ;
  assign n14909 = x10 & ~n1922 ;
  assign n14910 = n1069 | n4029 ;
  assign n14911 = n14910 ^ n8430 ^ 1'b0 ;
  assign n14912 = n502 | n14911 ;
  assign n14913 = n14909 & ~n14912 ;
  assign n14915 = n14914 ^ n14913 ^ 1'b0 ;
  assign n14918 = ~n5644 & n6985 ;
  assign n14919 = n14918 ^ n1590 ^ n1000 ;
  assign n14916 = n7466 ^ n3399 ^ 1'b0 ;
  assign n14917 = n14916 ^ n13787 ^ n11119 ;
  assign n14920 = n14919 ^ n14917 ^ 1'b0 ;
  assign n14921 = n6385 & ~n9522 ;
  assign n14922 = n14921 ^ n7838 ^ 1'b0 ;
  assign n14923 = n1613 | n11305 ;
  assign n14928 = ~n535 & n5324 ;
  assign n14929 = n4518 | n14928 ;
  assign n14924 = n9388 ^ n2434 ^ 1'b0 ;
  assign n14925 = n14924 ^ n7847 ^ n5759 ;
  assign n14926 = n7598 & ~n14925 ;
  assign n14927 = ~n5949 & n14926 ;
  assign n14930 = n14929 ^ n14927 ^ 1'b0 ;
  assign n14931 = n489 & n6501 ;
  assign n14932 = ( n1255 & n1571 ) | ( n1255 & ~n14931 ) | ( n1571 & ~n14931 ) ;
  assign n14933 = n5489 | n14932 ;
  assign n14935 = ~x182 & n1223 ;
  assign n14934 = n1998 & n12031 ;
  assign n14936 = n14935 ^ n14934 ^ 1'b0 ;
  assign n14937 = n7353 ^ n6244 ^ 1'b0 ;
  assign n14938 = n5766 & n14937 ;
  assign n14939 = n7013 & n12505 ;
  assign n14940 = n14939 ^ n2618 ^ 1'b0 ;
  assign n14941 = ( ~n13580 & n14704 ) | ( ~n13580 & n14940 ) | ( n14704 & n14940 ) ;
  assign n14942 = n14938 & n14941 ;
  assign n14943 = n14942 ^ n4282 ^ 1'b0 ;
  assign n14944 = n10596 & ~n14715 ;
  assign n14945 = n14943 & n14944 ;
  assign n14946 = n10063 ^ n2548 ^ 1'b0 ;
  assign n14947 = n4895 & ~n14946 ;
  assign n14948 = n14947 ^ n6798 ^ 1'b0 ;
  assign n14949 = ( n3804 & n6096 ) | ( n3804 & n14730 ) | ( n6096 & n14730 ) ;
  assign n14953 = ~n1495 & n4982 ;
  assign n14954 = ~n1478 & n14953 ;
  assign n14950 = n1084 | n4995 ;
  assign n14951 = n14950 ^ n11041 ^ 1'b0 ;
  assign n14952 = n10189 & n14951 ;
  assign n14955 = n14954 ^ n14952 ^ 1'b0 ;
  assign n14959 = n1813 ^ n780 ^ 1'b0 ;
  assign n14960 = n4722 & ~n14959 ;
  assign n14956 = n8404 ^ n6169 ^ 1'b0 ;
  assign n14957 = n7088 & ~n14956 ;
  assign n14958 = n14569 & n14957 ;
  assign n14961 = n14960 ^ n14958 ^ 1'b0 ;
  assign n14962 = n10908 ^ n1808 ^ 1'b0 ;
  assign n14963 = n14962 ^ n11728 ^ 1'b0 ;
  assign n14964 = ~n3984 & n4570 ;
  assign n14965 = ~n13748 & n14964 ;
  assign n14966 = ( n5426 & n9813 ) | ( n5426 & n14965 ) | ( n9813 & n14965 ) ;
  assign n14967 = n14629 ^ n9467 ^ n3010 ;
  assign n14968 = n3136 | n10618 ;
  assign n14969 = n4867 & ~n14300 ;
  assign n14970 = n14969 ^ n5305 ^ n4363 ;
  assign n14971 = n7785 ^ n6250 ^ n998 ;
  assign n14972 = n8314 | n14971 ;
  assign n14973 = n4038 | n6669 ;
  assign n14974 = n3643 & ~n7443 ;
  assign n14975 = n3120 | n14974 ;
  assign n14976 = n14973 & n14975 ;
  assign n14977 = n9950 | n13952 ;
  assign n14978 = n7817 & ~n14977 ;
  assign n14979 = n9607 & ~n14978 ;
  assign n14980 = ( n5725 & ~n7724 ) | ( n5725 & n10405 ) | ( ~n7724 & n10405 ) ;
  assign n14981 = ~n13694 & n14980 ;
  assign n14982 = n8114 & ~n14981 ;
  assign n14983 = n4041 ^ n1565 ^ 1'b0 ;
  assign n14984 = n5305 ^ n1471 ^ 1'b0 ;
  assign n14985 = n6309 | n14984 ;
  assign n14986 = ~n8125 & n14985 ;
  assign n14987 = n13915 | n14986 ;
  assign n14988 = n14983 | n14987 ;
  assign n14989 = n4873 & ~n10649 ;
  assign n14990 = n13571 ^ n1265 ^ 1'b0 ;
  assign n14991 = n14142 ^ n2853 ^ 1'b0 ;
  assign n14992 = n1147 & ~n7824 ;
  assign n14993 = n5313 & ~n14992 ;
  assign n14994 = n4211 | n10534 ;
  assign n14995 = ( n4483 & n5623 ) | ( n4483 & ~n14994 ) | ( n5623 & ~n14994 ) ;
  assign n14996 = n14995 ^ n10262 ^ 1'b0 ;
  assign n14997 = ( ~n883 & n4389 ) | ( ~n883 & n10867 ) | ( n4389 & n10867 ) ;
  assign n14998 = n14997 ^ n3738 ^ n2235 ;
  assign n14999 = n10028 ^ n1671 ^ 1'b0 ;
  assign n15000 = n6506 | n12273 ;
  assign n15001 = n15000 ^ n7070 ^ 1'b0 ;
  assign n15002 = ( x85 & ~n6668 ) | ( x85 & n7612 ) | ( ~n6668 & n7612 ) ;
  assign n15003 = ~n557 & n15002 ;
  assign n15004 = n15003 ^ n4460 ^ 1'b0 ;
  assign n15005 = ~n5172 & n8772 ;
  assign n15006 = n1397 | n15005 ;
  assign n15008 = n3997 & ~n8968 ;
  assign n15009 = n5635 & n15008 ;
  assign n15010 = n8999 & n15009 ;
  assign n15007 = n896 & n8231 ;
  assign n15011 = n15010 ^ n15007 ^ 1'b0 ;
  assign n15012 = n2081 | n7698 ;
  assign n15013 = n2046 & ~n4693 ;
  assign n15014 = ( n10237 & ~n15012 ) | ( n10237 & n15013 ) | ( ~n15012 & n15013 ) ;
  assign n15015 = ~n7697 & n8809 ;
  assign n15016 = n15015 ^ n3910 ^ 1'b0 ;
  assign n15017 = ~n3554 & n7560 ;
  assign n15018 = n1967 & n15017 ;
  assign n15019 = n5057 & n13264 ;
  assign n15026 = n3514 ^ n1291 ^ 1'b0 ;
  assign n15027 = n6597 | n15026 ;
  assign n15028 = ( x73 & ~n922 ) | ( x73 & n5172 ) | ( ~n922 & n5172 ) ;
  assign n15029 = n3803 & n15028 ;
  assign n15030 = ~n15027 & n15029 ;
  assign n15023 = n4271 & n11709 ;
  assign n15024 = n15023 ^ n412 ^ 1'b0 ;
  assign n15020 = ~n2590 & n3145 ;
  assign n15021 = n4899 & n13239 ;
  assign n15022 = ~n15020 & n15021 ;
  assign n15025 = n15024 ^ n15022 ^ 1'b0 ;
  assign n15031 = n15030 ^ n15025 ^ 1'b0 ;
  assign n15032 = ~n8567 & n12648 ;
  assign n15033 = n3147 | n11259 ;
  assign n15034 = n592 ^ x107 ^ 1'b0 ;
  assign n15035 = n13171 & ~n15034 ;
  assign n15036 = n15035 ^ n6286 ^ 1'b0 ;
  assign n15037 = ( n1489 & ~n3949 ) | ( n1489 & n15036 ) | ( ~n3949 & n15036 ) ;
  assign n15038 = ~n11910 & n15037 ;
  assign n15039 = ~n3790 & n15038 ;
  assign n15040 = n7346 | n15039 ;
  assign n15041 = n4117 ^ n1138 ^ n967 ;
  assign n15042 = ~n1727 & n15041 ;
  assign n15043 = n15042 ^ n11807 ^ 1'b0 ;
  assign n15044 = n9334 ^ n5021 ^ 1'b0 ;
  assign n15045 = n2023 & ~n10305 ;
  assign n15046 = ~n9261 & n15045 ;
  assign n15047 = n15046 ^ x235 ^ 1'b0 ;
  assign n15048 = n3720 & n4731 ;
  assign n15049 = n15048 ^ n2144 ^ 1'b0 ;
  assign n15050 = ~n2718 & n5264 ;
  assign n15051 = ~n15049 & n15050 ;
  assign n15052 = n3869 ^ x241 ^ 1'b0 ;
  assign n15053 = n3288 | n15052 ;
  assign n15054 = n5504 | n15053 ;
  assign n15055 = ~n3251 & n15054 ;
  assign n15056 = ( n5861 & n6546 ) | ( n5861 & ~n11303 ) | ( n6546 & ~n11303 ) ;
  assign n15057 = n3047 ^ n2209 ^ 1'b0 ;
  assign n15058 = n6723 & ~n15057 ;
  assign n15059 = n1639 & ~n7447 ;
  assign n15060 = n15059 ^ n12057 ^ 1'b0 ;
  assign n15061 = n12288 ^ n785 ^ 1'b0 ;
  assign n15062 = n2411 | n15061 ;
  assign n15063 = ( n1475 & n2325 ) | ( n1475 & n2445 ) | ( n2325 & n2445 ) ;
  assign n15064 = n15063 ^ n1501 ^ 1'b0 ;
  assign n15065 = n13260 ^ n4056 ^ 1'b0 ;
  assign n15066 = n13294 & ~n14471 ;
  assign n15067 = n15066 ^ n1951 ^ 1'b0 ;
  assign n15068 = n7413 | n12414 ;
  assign n15069 = n3255 & ~n10363 ;
  assign n15070 = n15069 ^ n7342 ^ 1'b0 ;
  assign n15071 = n15070 ^ n4724 ^ 1'b0 ;
  assign n15072 = n3102 & n15071 ;
  assign n15073 = n1959 & ~n14860 ;
  assign n15074 = n9021 ^ n8829 ^ n3875 ;
  assign n15075 = n5056 & ~n8585 ;
  assign n15076 = n10293 & n15075 ;
  assign n15077 = n15074 & n15076 ;
  assign n15078 = n5321 ^ n395 ^ 1'b0 ;
  assign n15079 = n15078 ^ n4267 ^ x52 ;
  assign n15080 = n5544 ^ n3330 ^ 1'b0 ;
  assign n15081 = ~n12083 & n15080 ;
  assign n15082 = n12103 & ~n15081 ;
  assign n15083 = n15082 ^ n2610 ^ 1'b0 ;
  assign n15084 = ~n4820 & n9632 ;
  assign n15085 = ( n3957 & n9279 ) | ( n3957 & ~n10890 ) | ( n9279 & ~n10890 ) ;
  assign n15086 = n6584 | n15085 ;
  assign n15087 = n12253 ^ n7866 ^ 1'b0 ;
  assign n15088 = n2824 & n5621 ;
  assign n15089 = ( ~n2345 & n7497 ) | ( ~n2345 & n15088 ) | ( n7497 & n15088 ) ;
  assign n15090 = n1972 | n7403 ;
  assign n15091 = n5768 & ~n15090 ;
  assign n15092 = n6818 | n9849 ;
  assign n15093 = n13184 & ~n15092 ;
  assign n15094 = ~n3773 & n5179 ;
  assign n15095 = n15094 ^ x125 ^ 1'b0 ;
  assign n15096 = ~n3891 & n15095 ;
  assign n15097 = ~n7303 & n15096 ;
  assign n15098 = n15097 ^ n3027 ^ 1'b0 ;
  assign n15099 = n15098 ^ n6272 ^ 1'b0 ;
  assign n15100 = ~x121 & n4010 ;
  assign n15101 = n7381 & ~n8413 ;
  assign n15102 = ~x136 & n15101 ;
  assign n15103 = n15100 | n15102 ;
  assign n15104 = n15103 ^ n7953 ^ 1'b0 ;
  assign n15105 = n8688 ^ n5877 ^ 1'b0 ;
  assign n15106 = n10070 & ~n15105 ;
  assign n15107 = n15106 ^ n11621 ^ 1'b0 ;
  assign n15108 = n15107 ^ n11163 ^ 1'b0 ;
  assign n15109 = n15104 & n15108 ;
  assign n15110 = n2224 & n15109 ;
  assign n15111 = n15110 ^ n395 ^ 1'b0 ;
  assign n15112 = n15111 ^ n4194 ^ 1'b0 ;
  assign n15113 = ~n15099 & n15112 ;
  assign n15114 = n7363 | n13640 ;
  assign n15115 = ( ~n1904 & n2272 ) | ( ~n1904 & n4229 ) | ( n2272 & n4229 ) ;
  assign n15116 = n15115 ^ n6379 ^ 1'b0 ;
  assign n15117 = ~n11608 & n15116 ;
  assign n15118 = n2950 | n3251 ;
  assign n15119 = n1115 & ~n15118 ;
  assign n15120 = n725 & n3332 ;
  assign n15121 = n15120 ^ n11493 ^ 1'b0 ;
  assign n15122 = ~n9351 & n15121 ;
  assign n15123 = n5685 | n8129 ;
  assign n15124 = ( n8067 & n15122 ) | ( n8067 & ~n15123 ) | ( n15122 & ~n15123 ) ;
  assign n15127 = n1166 | n4661 ;
  assign n15128 = n15127 ^ n8747 ^ 1'b0 ;
  assign n15125 = n5289 ^ n5170 ^ 1'b0 ;
  assign n15126 = ~n7688 & n15125 ;
  assign n15129 = n15128 ^ n15126 ^ 1'b0 ;
  assign n15130 = n463 | n15129 ;
  assign n15131 = n5984 | n10130 ;
  assign n15132 = n7431 & ~n9982 ;
  assign n15133 = n1827 & ~n3263 ;
  assign n15134 = n5529 ^ n258 ^ 1'b0 ;
  assign n15135 = ~n1111 & n3905 ;
  assign n15136 = n2653 & n15135 ;
  assign n15137 = ~n9175 & n15136 ;
  assign n15138 = n8751 ^ n6764 ^ 1'b0 ;
  assign n15139 = n14486 ^ n2597 ^ 1'b0 ;
  assign n15140 = n1095 & ~n15139 ;
  assign n15141 = n1029 & ~n14309 ;
  assign n15142 = n15141 ^ n7389 ^ 1'b0 ;
  assign n15143 = n15142 ^ n4666 ^ 1'b0 ;
  assign n15144 = n11850 | n15143 ;
  assign n15145 = n5025 ^ n3306 ^ 1'b0 ;
  assign n15146 = ~n2640 & n15145 ;
  assign n15147 = n15146 ^ n11144 ^ 1'b0 ;
  assign n15148 = n3889 & n7707 ;
  assign n15149 = n15148 ^ n5624 ^ 1'b0 ;
  assign n15150 = n13066 ^ n9987 ^ n9919 ;
  assign n15151 = n15150 ^ n1304 ^ 1'b0 ;
  assign n15152 = n15151 ^ n3462 ^ 1'b0 ;
  assign n15157 = n6700 ^ n4835 ^ 1'b0 ;
  assign n15158 = ~n1066 & n15157 ;
  assign n15153 = n1613 & ~n12788 ;
  assign n15154 = n3895 & ~n13386 ;
  assign n15155 = n15153 & n15154 ;
  assign n15156 = n5770 | n15155 ;
  assign n15159 = n15158 ^ n15156 ^ 1'b0 ;
  assign n15160 = n11041 ^ n8101 ^ 1'b0 ;
  assign n15161 = n15159 & n15160 ;
  assign n15162 = ~n3947 & n15161 ;
  assign n15165 = n10209 ^ n7023 ^ 1'b0 ;
  assign n15163 = n3332 & ~n14771 ;
  assign n15164 = n12191 & n15163 ;
  assign n15166 = n15165 ^ n15164 ^ n5098 ;
  assign n15167 = n1666 & n1983 ;
  assign n15168 = n15167 ^ n14599 ^ 1'b0 ;
  assign n15169 = ( ~n12070 & n12588 ) | ( ~n12070 & n15168 ) | ( n12588 & n15168 ) ;
  assign n15170 = n6923 ^ n3911 ^ 1'b0 ;
  assign n15171 = n5304 & ~n12740 ;
  assign n15172 = ~n15170 & n15171 ;
  assign n15173 = n1054 | n15172 ;
  assign n15174 = n12816 | n15173 ;
  assign n15175 = n3826 | n13194 ;
  assign n15176 = n8222 ^ n2393 ^ 1'b0 ;
  assign n15177 = n4415 | n7086 ;
  assign n15178 = n15177 ^ n8152 ^ 1'b0 ;
  assign n15181 = ~n756 & n7329 ;
  assign n15179 = n1275 ^ n1172 ^ 1'b0 ;
  assign n15180 = n3821 | n15179 ;
  assign n15182 = n15181 ^ n15180 ^ 1'b0 ;
  assign n15183 = n15182 ^ n2442 ^ 1'b0 ;
  assign n15184 = ~n11786 & n15183 ;
  assign n15185 = ~n2791 & n7060 ;
  assign n15186 = ~n3423 & n15185 ;
  assign n15187 = n7403 | n15186 ;
  assign n15188 = n6686 & ~n15187 ;
  assign n15189 = n15188 ^ n12704 ^ 1'b0 ;
  assign n15190 = ( n2819 & ~n3910 ) | ( n2819 & n15189 ) | ( ~n3910 & n15189 ) ;
  assign n15191 = n6047 ^ x65 ^ 1'b0 ;
  assign n15192 = n4496 & n12554 ;
  assign n15193 = n15192 ^ n2231 ^ 1'b0 ;
  assign n15194 = n10601 ^ n2002 ^ 1'b0 ;
  assign n15195 = n8318 | n12041 ;
  assign n15196 = n15194 | n15195 ;
  assign n15197 = n15196 ^ n2907 ^ 1'b0 ;
  assign n15198 = ( n14208 & n15193 ) | ( n14208 & n15197 ) | ( n15193 & n15197 ) ;
  assign n15199 = n12128 ^ n5043 ^ n3940 ;
  assign n15200 = n11874 | n14491 ;
  assign n15201 = n9112 & n15200 ;
  assign n15202 = n15201 ^ n1136 ^ 1'b0 ;
  assign n15206 = n451 & ~n753 ;
  assign n15207 = ~n451 & n15206 ;
  assign n15208 = n904 | n2420 ;
  assign n15209 = n904 & ~n15208 ;
  assign n15210 = n2235 | n12372 ;
  assign n15211 = n15209 | n15210 ;
  assign n15212 = n15207 & ~n15211 ;
  assign n15203 = n7552 ^ n4194 ^ 1'b0 ;
  assign n15204 = n14496 | n15203 ;
  assign n15205 = n4911 & n15204 ;
  assign n15213 = n15212 ^ n15205 ^ 1'b0 ;
  assign n15214 = n1344 & ~n1530 ;
  assign n15215 = n1530 & n15214 ;
  assign n15216 = n983 | n15215 ;
  assign n15217 = n15213 | n15216 ;
  assign n15218 = n15018 ^ n5780 ^ 1'b0 ;
  assign n15220 = n516 ^ x105 ^ 1'b0 ;
  assign n15219 = n2186 ^ x154 ^ 1'b0 ;
  assign n15221 = n15220 ^ n15219 ^ 1'b0 ;
  assign n15222 = ~n7926 & n12613 ;
  assign n15223 = ~n3504 & n10164 ;
  assign n15224 = ~n2187 & n10070 ;
  assign n15225 = n15224 ^ n1328 ^ 1'b0 ;
  assign n15226 = n12595 ^ n10166 ^ 1'b0 ;
  assign n15227 = n2826 | n4460 ;
  assign n15228 = n11137 & n11482 ;
  assign n15229 = ~n15227 & n15228 ;
  assign n15234 = n1317 | n4228 ;
  assign n15230 = n6830 ^ n2669 ^ 1'b0 ;
  assign n15231 = ( n2084 & n3271 ) | ( n2084 & ~n15230 ) | ( n3271 & ~n15230 ) ;
  assign n15232 = n10421 & ~n15231 ;
  assign n15233 = n15232 ^ n704 ^ 1'b0 ;
  assign n15235 = n15234 ^ n15233 ^ 1'b0 ;
  assign n15236 = n6114 & n15235 ;
  assign n15237 = n15122 ^ n11486 ^ 1'b0 ;
  assign n15238 = ~n6807 & n10796 ;
  assign n15239 = n755 | n3295 ;
  assign n15240 = n8944 ^ n8602 ^ n4797 ;
  assign n15241 = n4423 ^ n2041 ^ x179 ;
  assign n15242 = ( n11631 & ~n15240 ) | ( n11631 & n15241 ) | ( ~n15240 & n15241 ) ;
  assign n15243 = x100 & n15242 ;
  assign n15244 = ~n15239 & n15243 ;
  assign n15245 = n8662 | n8760 ;
  assign n15246 = n3126 | n15245 ;
  assign n15247 = n10274 | n15246 ;
  assign n15248 = n12483 ^ n9336 ^ n2797 ;
  assign n15249 = n8256 ^ n5155 ^ 1'b0 ;
  assign n15250 = ~n3027 & n3506 ;
  assign n15252 = ( n6038 & n6286 ) | ( n6038 & ~n9515 ) | ( n6286 & ~n9515 ) ;
  assign n15251 = n7521 ^ n488 ^ 1'b0 ;
  assign n15253 = n15252 ^ n15251 ^ n8778 ;
  assign n15254 = n8366 ^ n1228 ^ 1'b0 ;
  assign n15255 = ~n12310 & n15254 ;
  assign n15256 = n15255 ^ n10935 ^ n6484 ;
  assign n15257 = n5736 ^ n4859 ^ 1'b0 ;
  assign n15258 = ~n6889 & n15257 ;
  assign n15259 = n8435 & n15258 ;
  assign n15260 = n11290 ^ n713 ^ 1'b0 ;
  assign n15267 = n7269 ^ n3447 ^ 1'b0 ;
  assign n15268 = n7839 & ~n15267 ;
  assign n15269 = n824 | n1980 ;
  assign n15270 = n15268 | n15269 ;
  assign n15271 = n15270 ^ n5720 ^ 1'b0 ;
  assign n15261 = n4245 & n6892 ;
  assign n15262 = ~n8295 & n15261 ;
  assign n15263 = ~n581 & n2164 ;
  assign n15264 = ~n10824 & n15263 ;
  assign n15265 = ( ~n569 & n15262 ) | ( ~n569 & n15264 ) | ( n15262 & n15264 ) ;
  assign n15266 = n1304 | n15265 ;
  assign n15272 = n15271 ^ n15266 ^ 1'b0 ;
  assign n15275 = n1031 & ~n9838 ;
  assign n15274 = n4503 & n11321 ;
  assign n15276 = n15275 ^ n15274 ^ 1'b0 ;
  assign n15273 = ~n331 & n7128 ;
  assign n15277 = n15276 ^ n15273 ^ 1'b0 ;
  assign n15278 = n2573 & n10845 ;
  assign n15279 = n15277 & n15278 ;
  assign n15280 = n6877 ^ n3895 ^ 1'b0 ;
  assign n15281 = n5195 & n6352 ;
  assign n15282 = n15281 ^ n329 ^ 1'b0 ;
  assign n15283 = n6155 & n15282 ;
  assign n15284 = n15283 ^ n5339 ^ 1'b0 ;
  assign n15285 = n5882 & ~n15284 ;
  assign n15286 = n15285 ^ n6630 ^ 1'b0 ;
  assign n15287 = ~n2951 & n5094 ;
  assign n15288 = n7714 ^ n2916 ^ 1'b0 ;
  assign n15289 = n1643 & ~n6844 ;
  assign n15290 = ( ~n13220 & n15288 ) | ( ~n13220 & n15289 ) | ( n15288 & n15289 ) ;
  assign n15291 = n2433 | n5283 ;
  assign n15292 = n3554 | n15291 ;
  assign n15293 = n13448 ^ n4927 ^ 1'b0 ;
  assign n15294 = n1177 & n15293 ;
  assign n15295 = ( n5988 & n7453 ) | ( n5988 & ~n15294 ) | ( n7453 & ~n15294 ) ;
  assign n15296 = n15295 ^ n4808 ^ 1'b0 ;
  assign n15297 = n2778 & ~n9802 ;
  assign n15298 = n15297 ^ x64 ^ 1'b0 ;
  assign n15299 = n4460 | n11382 ;
  assign n15300 = ( n9365 & ~n9694 ) | ( n9365 & n15299 ) | ( ~n9694 & n15299 ) ;
  assign n15301 = n11039 & ~n15300 ;
  assign n15302 = n1882 ^ n1145 ^ 1'b0 ;
  assign n15303 = n15302 ^ n2380 ^ 1'b0 ;
  assign n15304 = n9953 & n15303 ;
  assign n15305 = n15304 ^ n6810 ^ 1'b0 ;
  assign n15306 = n10891 & n15305 ;
  assign n15307 = ( n8795 & n11772 ) | ( n8795 & n12266 ) | ( n11772 & n12266 ) ;
  assign n15308 = n3586 & ~n12446 ;
  assign n15309 = ~n1237 & n15308 ;
  assign n15310 = n9070 ^ n4433 ^ 1'b0 ;
  assign n15311 = n1598 | n5694 ;
  assign n15312 = ( n2647 & ~n8911 ) | ( n2647 & n9997 ) | ( ~n8911 & n9997 ) ;
  assign n15313 = n4148 | n15312 ;
  assign n15314 = n15311 & ~n15313 ;
  assign n15315 = ~n2547 & n3477 ;
  assign n15316 = n592 & n15315 ;
  assign n15317 = n1813 | n15316 ;
  assign n15318 = n15317 ^ n6775 ^ 1'b0 ;
  assign n15319 = n7008 | n15318 ;
  assign n15320 = ( ~n1477 & n8115 ) | ( ~n1477 & n8491 ) | ( n8115 & n8491 ) ;
  assign n15321 = ~n1995 & n15320 ;
  assign n15322 = n6105 ^ n5892 ^ n5671 ;
  assign n15323 = n15322 ^ n4216 ^ 1'b0 ;
  assign n15324 = n13123 | n15323 ;
  assign n15325 = ~n7969 & n8218 ;
  assign n15326 = n6822 & n15325 ;
  assign n15327 = n7731 & ~n15326 ;
  assign n15328 = n15327 ^ n3029 ^ 1'b0 ;
  assign n15329 = n4990 | n13006 ;
  assign n15330 = n14141 & ~n15329 ;
  assign n15331 = n15330 ^ n4547 ^ 1'b0 ;
  assign n15332 = n15328 & n15331 ;
  assign n15333 = n6250 ^ n5582 ^ n4626 ;
  assign n15334 = n9011 ^ n2761 ^ 1'b0 ;
  assign n15335 = n3546 & n15334 ;
  assign n15336 = n15335 ^ n950 ^ 1'b0 ;
  assign n15337 = n9925 | n15336 ;
  assign n15338 = n15337 ^ n8845 ^ 1'b0 ;
  assign n15339 = ~n4506 & n13712 ;
  assign n15340 = n10130 ^ x65 ^ 1'b0 ;
  assign n15341 = ~n3834 & n15340 ;
  assign n15342 = ~n9539 & n15341 ;
  assign n15343 = ~n2350 & n15342 ;
  assign n15344 = n11404 ^ n645 ^ 1'b0 ;
  assign n15345 = ~n6327 & n15344 ;
  assign n15346 = n3438 & n5877 ;
  assign n15347 = n15346 ^ n9656 ^ 1'b0 ;
  assign n15348 = n15347 ^ n10070 ^ n981 ;
  assign n15350 = n9693 ^ n8522 ^ 1'b0 ;
  assign n15349 = n6440 | n9203 ;
  assign n15351 = n15350 ^ n15349 ^ 1'b0 ;
  assign n15352 = n15351 ^ n2612 ^ 1'b0 ;
  assign n15353 = n13343 | n15352 ;
  assign n15359 = ~n5991 & n9275 ;
  assign n15360 = n15359 ^ n10600 ^ 1'b0 ;
  assign n15361 = n4882 | n8795 ;
  assign n15362 = n15360 | n15361 ;
  assign n15354 = n2284 | n7200 ;
  assign n15355 = n7381 & ~n15354 ;
  assign n15356 = n6334 | n15355 ;
  assign n15357 = n15356 ^ n4757 ^ 1'b0 ;
  assign n15358 = n6904 & n15357 ;
  assign n15363 = n15362 ^ n15358 ^ 1'b0 ;
  assign n15364 = ~n648 & n8026 ;
  assign n15365 = n15364 ^ n13948 ^ 1'b0 ;
  assign n15366 = n2538 ^ n1667 ^ 1'b0 ;
  assign n15367 = n6915 & n15366 ;
  assign n15368 = n15367 ^ n13897 ^ 1'b0 ;
  assign n15369 = n3723 & ~n10361 ;
  assign n15373 = n1865 | n2951 ;
  assign n15374 = n15373 ^ n6352 ^ 1'b0 ;
  assign n15370 = n2241 & ~n3389 ;
  assign n15371 = n15370 ^ n7102 ^ 1'b0 ;
  assign n15372 = n5828 & n15371 ;
  assign n15375 = n15374 ^ n15372 ^ 1'b0 ;
  assign n15376 = n15369 | n15375 ;
  assign n15377 = ~n1404 & n3410 ;
  assign n15378 = n15377 ^ n2654 ^ 1'b0 ;
  assign n15379 = ~n12974 & n15378 ;
  assign n15380 = n13566 ^ n8664 ^ 1'b0 ;
  assign n15381 = ~n2160 & n15380 ;
  assign n15382 = ~n3696 & n6825 ;
  assign n15383 = ~n2522 & n15382 ;
  assign n15384 = n10125 | n15383 ;
  assign n15385 = x193 | n15384 ;
  assign n15386 = n9858 ^ n1317 ^ 1'b0 ;
  assign n15387 = n2862 & ~n15386 ;
  assign n15388 = n15387 ^ n7233 ^ 1'b0 ;
  assign n15389 = n9261 ^ n5033 ^ 1'b0 ;
  assign n15390 = n10763 | n10920 ;
  assign n15391 = n8719 ^ n1210 ^ 1'b0 ;
  assign n15392 = n15391 ^ x167 ^ 1'b0 ;
  assign n15393 = n6967 | n15392 ;
  assign n15394 = n15393 ^ n2292 ^ 1'b0 ;
  assign n15395 = n14743 ^ n3322 ^ 1'b0 ;
  assign n15396 = ( ~n3096 & n11383 ) | ( ~n3096 & n14214 ) | ( n11383 & n14214 ) ;
  assign n15397 = n15396 ^ n5179 ^ 1'b0 ;
  assign n15398 = n2394 & n15397 ;
  assign n15399 = n15398 ^ n6443 ^ 1'b0 ;
  assign n15400 = n15395 & n15399 ;
  assign n15401 = n1455 & n4191 ;
  assign n15402 = n3464 | n8793 ;
  assign n15403 = n8058 | n15402 ;
  assign n15404 = n8035 & n15403 ;
  assign n15405 = n1473 & ~n6288 ;
  assign n15406 = n15405 ^ n3363 ^ 1'b0 ;
  assign n15407 = n15406 ^ n7552 ^ 1'b0 ;
  assign n15408 = n401 | n15407 ;
  assign n15409 = n1049 & n3599 ;
  assign n15410 = n4099 ^ n3508 ^ 1'b0 ;
  assign n15411 = n15410 ^ n8087 ^ 1'b0 ;
  assign n15412 = n7603 ^ n4724 ^ 1'b0 ;
  assign n15413 = n10648 ^ n4460 ^ n3723 ;
  assign n15414 = n12377 ^ n10137 ^ 1'b0 ;
  assign n15415 = n15413 | n15414 ;
  assign n15416 = n15415 ^ n12765 ^ 1'b0 ;
  assign n15417 = n4004 ^ x239 ^ 1'b0 ;
  assign n15418 = n4731 ^ x53 ^ 1'b0 ;
  assign n15419 = n14306 & n15418 ;
  assign n15420 = n15417 & n15419 ;
  assign n15421 = n681 ^ x194 ^ 1'b0 ;
  assign n15422 = ~n2965 & n6539 ;
  assign n15423 = n4001 & n5036 ;
  assign n15424 = n5172 ^ n436 ^ 1'b0 ;
  assign n15425 = n271 & n15424 ;
  assign n15426 = n7655 & n15425 ;
  assign n15427 = ( n11242 & ~n15423 ) | ( n11242 & n15426 ) | ( ~n15423 & n15426 ) ;
  assign n15428 = n9975 ^ n7940 ^ 1'b0 ;
  assign n15429 = n11872 ^ n8929 ^ 1'b0 ;
  assign n15430 = ~n15428 & n15429 ;
  assign n15431 = ~n5482 & n8614 ;
  assign n15432 = n15431 ^ n10155 ^ n9369 ;
  assign n15433 = n6360 | n14261 ;
  assign n15434 = n5918 ^ n5192 ^ 1'b0 ;
  assign n15435 = n15434 ^ n4929 ^ 1'b0 ;
  assign n15436 = n2509 & n15435 ;
  assign n15437 = n3714 ^ n2531 ^ 1'b0 ;
  assign n15438 = n9319 & n12288 ;
  assign n15439 = n304 | n840 ;
  assign n15440 = n15439 ^ n1019 ^ 1'b0 ;
  assign n15441 = n15440 ^ n13998 ^ 1'b0 ;
  assign n15442 = n594 | n11895 ;
  assign n15443 = ~n6194 & n6651 ;
  assign n15444 = ( n4064 & n8086 ) | ( n4064 & ~n15443 ) | ( n8086 & ~n15443 ) ;
  assign n15445 = n12902 & ~n15240 ;
  assign n15446 = n6470 & n15445 ;
  assign n15447 = n15444 & n15446 ;
  assign n15448 = ~n2860 & n6365 ;
  assign n15449 = ~n7701 & n15448 ;
  assign n15450 = n11552 ^ n3701 ^ 1'b0 ;
  assign n15451 = n15450 ^ n8974 ^ n1213 ;
  assign n15452 = n706 | n6292 ;
  assign n15453 = n7866 ^ n7099 ^ 1'b0 ;
  assign n15454 = n985 & n14662 ;
  assign n15455 = n5431 & ~n8490 ;
  assign n15456 = n15455 ^ n9682 ^ 1'b0 ;
  assign n15457 = n7732 ^ n1991 ^ 1'b0 ;
  assign n15458 = ~n755 & n15457 ;
  assign n15459 = n10062 ^ n3844 ^ n852 ;
  assign n15460 = x21 & n6465 ;
  assign n15462 = n6179 ^ n5795 ^ 1'b0 ;
  assign n15463 = n15462 ^ n9651 ^ 1'b0 ;
  assign n15461 = x30 & x120 ;
  assign n15464 = n15463 ^ n15461 ^ 1'b0 ;
  assign n15467 = n1919 & ~n14506 ;
  assign n15465 = n4231 & ~n6366 ;
  assign n15466 = n8477 & ~n15465 ;
  assign n15468 = n15467 ^ n15466 ^ 1'b0 ;
  assign n15469 = n10882 ^ n9119 ^ 1'b0 ;
  assign n15470 = n6863 ^ n1515 ^ 1'b0 ;
  assign n15471 = n12921 & ~n15470 ;
  assign n15472 = n15471 ^ n6768 ^ 1'b0 ;
  assign n15473 = ~n4749 & n15472 ;
  assign n15474 = ( ~n2345 & n6808 ) | ( ~n2345 & n15473 ) | ( n6808 & n15473 ) ;
  assign n15481 = n4169 ^ n2081 ^ n1033 ;
  assign n15482 = ~n5205 & n15481 ;
  assign n15475 = n5491 ^ n2708 ^ 1'b0 ;
  assign n15476 = n8455 ^ n7984 ^ 1'b0 ;
  assign n15477 = n15475 | n15476 ;
  assign n15478 = n5373 & ~n15477 ;
  assign n15479 = ~n3912 & n15478 ;
  assign n15480 = n5958 & ~n15479 ;
  assign n15483 = n15482 ^ n15480 ^ 1'b0 ;
  assign n15484 = n13527 & n15483 ;
  assign n15485 = ( n4802 & n4976 ) | ( n4802 & n15484 ) | ( n4976 & n15484 ) ;
  assign n15490 = n5006 & n8022 ;
  assign n15487 = n11563 ^ n8342 ^ 1'b0 ;
  assign n15488 = n5232 & ~n15487 ;
  assign n15489 = n6413 & n15488 ;
  assign n15486 = n3133 ^ n2844 ^ 1'b0 ;
  assign n15491 = n15490 ^ n15489 ^ n15486 ;
  assign n15492 = n13981 ^ n12341 ^ 1'b0 ;
  assign n15493 = ~n3744 & n15492 ;
  assign n15494 = ~n2601 & n14410 ;
  assign n15495 = ( n588 & n989 ) | ( n588 & ~n2100 ) | ( n989 & ~n2100 ) ;
  assign n15496 = n5641 | n13906 ;
  assign n15497 = n3879 ^ n1225 ^ 1'b0 ;
  assign n15498 = n8894 & ~n9067 ;
  assign n15505 = ~n5535 & n12947 ;
  assign n15506 = ~n4458 & n15505 ;
  assign n15499 = n478 ^ x68 ^ 1'b0 ;
  assign n15500 = n2756 & ~n15499 ;
  assign n15501 = n5336 & n6091 ;
  assign n15502 = n15501 ^ n7371 ^ 1'b0 ;
  assign n15503 = n15502 ^ n2405 ^ 1'b0 ;
  assign n15504 = n15500 & n15503 ;
  assign n15507 = n15506 ^ n15504 ^ 1'b0 ;
  assign n15508 = n8409 ^ n1323 ^ n821 ;
  assign n15509 = n15508 ^ n1981 ^ 1'b0 ;
  assign n15510 = n2437 & ~n14538 ;
  assign n15511 = n15510 ^ n14881 ^ 1'b0 ;
  assign n15512 = n6766 ^ n5776 ^ 1'b0 ;
  assign n15513 = x4 & ~n15512 ;
  assign n15521 = n3234 & n5092 ;
  assign n15522 = n15521 ^ n5742 ^ 1'b0 ;
  assign n15523 = n15522 ^ n6820 ^ 1'b0 ;
  assign n15524 = n4887 & ~n15523 ;
  assign n15525 = ~n1046 & n15524 ;
  assign n15518 = n3013 | n6351 ;
  assign n15519 = n13547 & ~n15518 ;
  assign n15514 = n6541 | n7413 ;
  assign n15515 = n5623 | n15514 ;
  assign n15516 = ~n2147 & n15515 ;
  assign n15517 = n1809 & n15516 ;
  assign n15520 = n15519 ^ n15517 ^ n14278 ;
  assign n15526 = n15525 ^ n15520 ^ 1'b0 ;
  assign n15527 = n15513 & n15526 ;
  assign n15528 = n4380 & ~n7569 ;
  assign n15529 = n1378 & n15528 ;
  assign n15530 = n1066 | n11305 ;
  assign n15531 = n7080 ^ n3126 ^ 1'b0 ;
  assign n15532 = n10198 & ~n15531 ;
  assign n15533 = n8381 ^ n5400 ^ n2816 ;
  assign n15534 = ~n2626 & n15533 ;
  assign n15535 = n7745 ^ n1255 ^ 1'b0 ;
  assign n15536 = n15535 ^ n6432 ^ n1176 ;
  assign n15537 = n1567 & ~n15536 ;
  assign n15538 = n15537 ^ n2614 ^ 1'b0 ;
  assign n15539 = n5404 ^ n3729 ^ n3228 ;
  assign n15540 = n15539 ^ n11372 ^ n5905 ;
  assign n15541 = ~n9875 & n15540 ;
  assign n15542 = n3427 ^ x75 ^ 1'b0 ;
  assign n15543 = n10236 & ~n14469 ;
  assign n15544 = ~n6284 & n15543 ;
  assign n15545 = n6259 ^ n1679 ^ 1'b0 ;
  assign n15546 = n9583 & ~n15545 ;
  assign n15547 = n5711 ^ n1651 ^ 1'b0 ;
  assign n15548 = n3611 & ~n15547 ;
  assign n15549 = ~n1156 & n15548 ;
  assign n15550 = n8352 & n15549 ;
  assign n15551 = n7407 ^ n6098 ^ 1'b0 ;
  assign n15552 = ( n15546 & n15550 ) | ( n15546 & n15551 ) | ( n15550 & n15551 ) ;
  assign n15553 = ~n3043 & n3242 ;
  assign n15554 = n15553 ^ n14733 ^ 1'b0 ;
  assign n15555 = x186 & ~n3291 ;
  assign n15556 = n529 | n11457 ;
  assign n15557 = n15556 ^ n9118 ^ 1'b0 ;
  assign n15558 = ( ~n1732 & n6442 ) | ( ~n1732 & n6671 ) | ( n6442 & n6671 ) ;
  assign n15559 = n15557 & n15558 ;
  assign n15560 = n14909 & n15559 ;
  assign n15561 = ( n2096 & n6146 ) | ( n2096 & ~n7014 ) | ( n6146 & ~n7014 ) ;
  assign n15562 = n15561 ^ n6797 ^ 1'b0 ;
  assign n15563 = n3600 ^ n847 ^ 1'b0 ;
  assign n15564 = ( n481 & n1753 ) | ( n481 & ~n15563 ) | ( n1753 & ~n15563 ) ;
  assign n15565 = n5221 ^ n1667 ^ x248 ;
  assign n15566 = ( n2782 & n6049 ) | ( n2782 & ~n15565 ) | ( n6049 & ~n15565 ) ;
  assign n15567 = n8625 ^ n7433 ^ 1'b0 ;
  assign n15568 = n2937 & n10346 ;
  assign n15569 = n15568 ^ n4615 ^ 1'b0 ;
  assign n15570 = ~n7109 & n10070 ;
  assign n15571 = ~n8531 & n15570 ;
  assign n15572 = ( n3960 & n4083 ) | ( n3960 & ~n15571 ) | ( n4083 & ~n15571 ) ;
  assign n15573 = n11963 | n15572 ;
  assign n15574 = n15569 | n15573 ;
  assign n15575 = n3008 ^ n2544 ^ x228 ;
  assign n15576 = n15575 ^ n9942 ^ x111 ;
  assign n15577 = n6381 | n15576 ;
  assign n15578 = n12020 ^ n8101 ^ 1'b0 ;
  assign n15580 = n5187 ^ n1168 ^ 1'b0 ;
  assign n15581 = n15580 ^ n5832 ^ 1'b0 ;
  assign n15582 = ~n3860 & n15581 ;
  assign n15583 = n800 & n15582 ;
  assign n15579 = n2187 | n9857 ;
  assign n15584 = n15583 ^ n15579 ^ 1'b0 ;
  assign n15585 = n5379 & n7674 ;
  assign n15586 = ( ~n2748 & n7267 ) | ( ~n2748 & n15585 ) | ( n7267 & n15585 ) ;
  assign n15587 = n10888 ^ n6299 ^ 1'b0 ;
  assign n15588 = x239 & ~n15587 ;
  assign n15589 = n7519 ^ n3586 ^ n1625 ;
  assign n15592 = n4705 & n10185 ;
  assign n15593 = ~n11368 & n15592 ;
  assign n15590 = n11187 ^ n5417 ^ 1'b0 ;
  assign n15591 = n14226 & ~n15590 ;
  assign n15594 = n15593 ^ n15591 ^ 1'b0 ;
  assign n15595 = n10300 ^ n1082 ^ n307 ;
  assign n15596 = n1880 | n4132 ;
  assign n15597 = n15595 | n15596 ;
  assign n15598 = n9045 & n15597 ;
  assign n15599 = n10782 & n15598 ;
  assign n15600 = ~n4799 & n5303 ;
  assign n15601 = n15600 ^ n2258 ^ 1'b0 ;
  assign n15602 = n15601 ^ n2715 ^ 1'b0 ;
  assign n15603 = n15602 ^ n13146 ^ 1'b0 ;
  assign n15604 = n5556 & ~n15603 ;
  assign n15605 = n15599 & n15604 ;
  assign n15606 = ~n2952 & n9286 ;
  assign n15607 = n7724 & n15606 ;
  assign n15608 = ~n11141 & n15607 ;
  assign n15609 = ~n3915 & n13857 ;
  assign n15610 = n2733 & ~n13243 ;
  assign n15611 = n4573 | n15610 ;
  assign n15612 = n4455 & ~n15611 ;
  assign n15613 = n10935 & ~n15612 ;
  assign n15614 = n6198 & n15613 ;
  assign n15615 = n10006 ^ n895 ^ 1'b0 ;
  assign n15616 = ~n681 & n15615 ;
  assign n15617 = n7814 | n13127 ;
  assign n15618 = n15617 ^ n3678 ^ 1'b0 ;
  assign n15619 = n15618 ^ n10434 ^ 1'b0 ;
  assign n15620 = n15616 & ~n15619 ;
  assign n15621 = n9480 ^ n6375 ^ 1'b0 ;
  assign n15622 = ( n7402 & n10555 ) | ( n7402 & n15621 ) | ( n10555 & n15621 ) ;
  assign n15623 = n15622 ^ n12261 ^ 1'b0 ;
  assign n15624 = n14868 ^ n13941 ^ n12633 ;
  assign n15625 = n15150 ^ n1025 ^ 1'b0 ;
  assign n15626 = n6893 & ~n13086 ;
  assign n15627 = n3822 & n15626 ;
  assign n15628 = ( n6294 & ~n6683 ) | ( n6294 & n9211 ) | ( ~n6683 & n9211 ) ;
  assign n15629 = n15628 ^ n15158 ^ 1'b0 ;
  assign n15630 = n5415 & ~n15219 ;
  assign n15631 = ~n15629 & n15630 ;
  assign n15632 = n6319 & n15140 ;
  assign n15633 = n8109 | n12903 ;
  assign n15634 = n15633 ^ n831 ^ 1'b0 ;
  assign n15635 = ( n5540 & n10175 ) | ( n5540 & ~n10405 ) | ( n10175 & ~n10405 ) ;
  assign n15636 = n15635 ^ x137 ^ 1'b0 ;
  assign n15637 = n2404 ^ n2033 ^ n1234 ;
  assign n15638 = n8930 | n12216 ;
  assign n15639 = n15638 ^ n7158 ^ 1'b0 ;
  assign n15640 = ( n7915 & n15637 ) | ( n7915 & ~n15639 ) | ( n15637 & ~n15639 ) ;
  assign n15641 = n935 & n5839 ;
  assign n15642 = n5295 & n15641 ;
  assign n15643 = n9319 ^ n2892 ^ 1'b0 ;
  assign n15644 = ~n15642 & n15643 ;
  assign n15645 = n2361 & n15644 ;
  assign n15649 = n5025 ^ n340 ^ 1'b0 ;
  assign n15646 = n1145 & ~n11920 ;
  assign n15647 = ~n3534 & n8303 ;
  assign n15648 = n15646 & n15647 ;
  assign n15650 = n15649 ^ n15648 ^ 1'b0 ;
  assign n15652 = n5116 ^ n2019 ^ 1'b0 ;
  assign n15653 = ~n8731 & n15652 ;
  assign n15651 = n13980 ^ x201 ^ 1'b0 ;
  assign n15654 = n15653 ^ n15651 ^ 1'b0 ;
  assign n15655 = x70 & ~n15654 ;
  assign n15656 = n15317 ^ n4152 ^ 1'b0 ;
  assign n15657 = n15656 ^ n4679 ^ 1'b0 ;
  assign n15658 = ~n1176 & n3435 ;
  assign n15659 = n15658 ^ n13453 ^ 1'b0 ;
  assign n15660 = ~n8756 & n14698 ;
  assign n15661 = n802 & n15660 ;
  assign n15662 = n8882 & n11929 ;
  assign n15663 = n15662 ^ n12124 ^ 1'b0 ;
  assign n15664 = ~n5303 & n9157 ;
  assign n15665 = n15664 ^ n9562 ^ 1'b0 ;
  assign n15666 = ~n7748 & n15665 ;
  assign n15667 = n8194 & n15666 ;
  assign n15668 = n10443 & n15667 ;
  assign n15669 = n15668 ^ n3590 ^ 1'b0 ;
  assign n15670 = n2703 | n3261 ;
  assign n15671 = n15670 ^ n12131 ^ n9729 ;
  assign n15672 = ( n366 & n6093 ) | ( n366 & ~n12167 ) | ( n6093 & ~n12167 ) ;
  assign n15673 = n3779 ^ n3311 ^ 1'b0 ;
  assign n15674 = n12744 | n15673 ;
  assign n15675 = n5675 | n15674 ;
  assign n15676 = ~n11633 & n15675 ;
  assign n15677 = n14773 ^ n7170 ^ 1'b0 ;
  assign n15678 = x156 & ~n562 ;
  assign n15679 = ~n1543 & n15678 ;
  assign n15680 = ( n4536 & n14603 ) | ( n4536 & n15679 ) | ( n14603 & n15679 ) ;
  assign n15681 = n8130 ^ n4089 ^ 1'b0 ;
  assign n15682 = n15680 & ~n15681 ;
  assign n15683 = n6686 & ~n9174 ;
  assign n15684 = n4493 & ~n5732 ;
  assign n15685 = n5732 & n15684 ;
  assign n15686 = n15685 ^ n14248 ^ 1'b0 ;
  assign n15687 = n13239 & n15686 ;
  assign n15688 = n15687 ^ x248 ^ 1'b0 ;
  assign n15689 = n6926 & ~n15443 ;
  assign n15690 = n6355 & ~n13153 ;
  assign n15691 = n15690 ^ n12607 ^ 1'b0 ;
  assign n15692 = n3957 | n15691 ;
  assign n15693 = n7124 ^ n909 ^ 1'b0 ;
  assign n15694 = n6496 & ~n15693 ;
  assign n15695 = n9988 & n15694 ;
  assign n15696 = n13584 ^ n2278 ^ 1'b0 ;
  assign n15697 = n15696 ^ n14016 ^ n10121 ;
  assign n15698 = ~n1462 & n15697 ;
  assign n15699 = n15698 ^ n4656 ^ 1'b0 ;
  assign n15702 = x162 & ~n9237 ;
  assign n15703 = n2797 & n15702 ;
  assign n15701 = n11225 ^ n3095 ^ 1'b0 ;
  assign n15700 = ~n537 & n4731 ;
  assign n15704 = n15703 ^ n15701 ^ n15700 ;
  assign n15705 = n9942 ^ n753 ^ 1'b0 ;
  assign n15706 = n10771 & ~n15705 ;
  assign n15707 = n6734 & ~n15179 ;
  assign n15708 = n6754 & n14584 ;
  assign n15709 = n2761 | n4405 ;
  assign n15710 = n5137 ^ n718 ^ 1'b0 ;
  assign n15711 = n15710 ^ n7721 ^ 1'b0 ;
  assign n15712 = n5250 | n15711 ;
  assign n15713 = n11112 | n15712 ;
  assign n15718 = n6225 ^ n3671 ^ 1'b0 ;
  assign n15719 = n2509 | n15718 ;
  assign n15716 = n1231 & ~n2275 ;
  assign n15717 = ~n4065 & n15716 ;
  assign n15720 = n15719 ^ n15717 ^ 1'b0 ;
  assign n15721 = n6888 & n15720 ;
  assign n15715 = n7413 | n10275 ;
  assign n15714 = n9394 & n14236 ;
  assign n15722 = n15721 ^ n15715 ^ n15714 ;
  assign n15723 = n15722 ^ n2332 ^ 1'b0 ;
  assign n15724 = ( n15709 & n15713 ) | ( n15709 & n15723 ) | ( n15713 & n15723 ) ;
  assign n15725 = n15724 ^ n3940 ^ 1'b0 ;
  assign n15726 = n4696 | n15725 ;
  assign n15727 = n601 | n4852 ;
  assign n15728 = ( n7766 & n14896 ) | ( n7766 & ~n15727 ) | ( n14896 & ~n15727 ) ;
  assign n15729 = n15575 ^ n5912 ^ 1'b0 ;
  assign n15730 = n13807 & ~n14744 ;
  assign n15731 = ~n6330 & n10360 ;
  assign n15732 = n3915 & n15731 ;
  assign n15733 = n15732 ^ n3251 ^ 1'b0 ;
  assign n15734 = n11840 ^ n11572 ^ 1'b0 ;
  assign n15735 = n3551 & ~n4440 ;
  assign n15736 = ~n15734 & n15735 ;
  assign n15737 = n8281 ^ n3119 ^ 1'b0 ;
  assign n15738 = n7673 & n15737 ;
  assign n15739 = n6092 & n15738 ;
  assign n15740 = n15739 ^ n6161 ^ 1'b0 ;
  assign n15741 = n10092 & ~n15740 ;
  assign n15742 = n6681 ^ n3551 ^ 1'b0 ;
  assign n15743 = n8899 & ~n15742 ;
  assign n15744 = x36 & n3209 ;
  assign n15745 = ( n5049 & ~n6677 ) | ( n5049 & n9415 ) | ( ~n6677 & n9415 ) ;
  assign n15746 = ( ~x199 & n13114 ) | ( ~x199 & n15745 ) | ( n13114 & n15745 ) ;
  assign n15747 = n5103 & n8223 ;
  assign n15748 = n3806 | n14262 ;
  assign n15749 = n15747 | n15748 ;
  assign n15750 = ~n9345 & n15749 ;
  assign n15751 = n10982 & n12519 ;
  assign n15752 = n1279 & ~n3198 ;
  assign n15753 = ~n5432 & n15752 ;
  assign n15754 = n4742 & n15753 ;
  assign n15755 = n10760 ^ n1499 ^ 1'b0 ;
  assign n15756 = n3213 | n14743 ;
  assign n15757 = n15756 ^ n10969 ^ n10579 ;
  assign n15758 = ~n1768 & n5049 ;
  assign n15759 = n15758 ^ n7488 ^ n6719 ;
  assign n15760 = n1097 & ~n15759 ;
  assign n15761 = n7051 & ~n14854 ;
  assign n15762 = n12598 ^ n4686 ^ 1'b0 ;
  assign n15763 = ~n2275 & n5783 ;
  assign n15764 = n3058 & n15763 ;
  assign n15765 = n15764 ^ n9375 ^ 1'b0 ;
  assign n15766 = n13744 ^ n12637 ^ 1'b0 ;
  assign n15767 = x241 & ~n15766 ;
  assign n15768 = n1506 ^ x181 ^ 1'b0 ;
  assign n15769 = n4703 | n7080 ;
  assign n15770 = n15769 ^ n2266 ^ 1'b0 ;
  assign n15771 = n3269 | n15770 ;
  assign n15772 = n15771 ^ n3292 ^ 1'b0 ;
  assign n15773 = n6411 & n12002 ;
  assign n15774 = ( n3877 & n4852 ) | ( n3877 & ~n15773 ) | ( n4852 & ~n15773 ) ;
  assign n15775 = n4213 & n9394 ;
  assign n15776 = n15775 ^ n5242 ^ 1'b0 ;
  assign n15777 = n15776 ^ n1555 ^ 1'b0 ;
  assign n15778 = n1144 | n15777 ;
  assign n15779 = n2862 ^ x223 ^ 1'b0 ;
  assign n15780 = ~n3236 & n15779 ;
  assign n15781 = n7700 & n15780 ;
  assign n15782 = n6249 ^ n1746 ^ 1'b0 ;
  assign n15783 = n6865 & n10444 ;
  assign n15784 = ~n5179 & n15783 ;
  assign n15785 = n11181 & ~n15784 ;
  assign n15786 = n15785 ^ n6336 ^ n1107 ;
  assign n15787 = n15782 & ~n15786 ;
  assign n15788 = ~n3126 & n4471 ;
  assign n15789 = n563 ^ x32 ^ 1'b0 ;
  assign n15790 = n5226 | n15789 ;
  assign n15791 = ( n10404 & n15788 ) | ( n10404 & ~n15790 ) | ( n15788 & ~n15790 ) ;
  assign n15792 = n11885 ^ n6674 ^ 1'b0 ;
  assign n15793 = n13767 ^ n4370 ^ 1'b0 ;
  assign n15794 = n11879 | n14145 ;
  assign n15795 = n15793 | n15794 ;
  assign n15796 = n5279 & ~n10312 ;
  assign n15797 = ~n3980 & n15796 ;
  assign n15798 = n6734 | n15797 ;
  assign n15799 = n15798 ^ n6517 ^ 1'b0 ;
  assign n15800 = n14281 ^ n4034 ^ 1'b0 ;
  assign n15801 = n14908 ^ n8117 ^ 1'b0 ;
  assign n15802 = ~n1423 & n15801 ;
  assign n15803 = ~n4505 & n4929 ;
  assign n15804 = n905 & n11601 ;
  assign n15805 = n15804 ^ n4639 ^ 1'b0 ;
  assign n15806 = n2162 ^ n351 ^ 1'b0 ;
  assign n15807 = n15806 ^ n8455 ^ x189 ;
  assign n15808 = n15807 ^ n3866 ^ n2418 ;
  assign n15809 = n4664 & n7721 ;
  assign n15810 = n15809 ^ n4638 ^ 1'b0 ;
  assign n15811 = ~n15808 & n15810 ;
  assign n15814 = n7448 ^ n1913 ^ 1'b0 ;
  assign n15812 = ( n2131 & ~n7873 ) | ( n2131 & n8770 ) | ( ~n7873 & n8770 ) ;
  assign n15813 = n15812 ^ n6904 ^ 1'b0 ;
  assign n15815 = n15814 ^ n15813 ^ n14538 ;
  assign n15816 = ~n11887 & n12144 ;
  assign n15818 = n2668 & ~n4024 ;
  assign n15817 = ~n3557 & n7097 ;
  assign n15819 = n15818 ^ n15817 ^ 1'b0 ;
  assign n15820 = n10867 | n15806 ;
  assign n15821 = n459 & n6600 ;
  assign n15822 = n15820 & n15821 ;
  assign n15823 = n15819 | n15822 ;
  assign n15824 = n1520 & ~n15823 ;
  assign n15825 = n15824 ^ n6645 ^ 1'b0 ;
  assign n15826 = n8167 & ~n12190 ;
  assign n15827 = n15826 ^ n14816 ^ 1'b0 ;
  assign n15828 = n15825 & ~n15827 ;
  assign n15829 = n10368 ^ n8026 ^ 1'b0 ;
  assign n15830 = n1856 | n14865 ;
  assign n15831 = n15830 ^ n14861 ^ 1'b0 ;
  assign n15832 = n2561 ^ n2024 ^ 1'b0 ;
  assign n15833 = n15832 ^ n1932 ^ 1'b0 ;
  assign n15836 = n1620 & n4083 ;
  assign n15834 = n3924 ^ n1330 ^ 1'b0 ;
  assign n15835 = n15834 ^ n4723 ^ n1686 ;
  assign n15837 = n15836 ^ n15835 ^ 1'b0 ;
  assign n15838 = ( ~n10250 & n10450 ) | ( ~n10250 & n15837 ) | ( n10450 & n15837 ) ;
  assign n15839 = n14204 ^ n7928 ^ 1'b0 ;
  assign n15840 = n15107 & n15839 ;
  assign n15841 = n13832 ^ n13156 ^ n2547 ;
  assign n15842 = n8041 ^ n1976 ^ 1'b0 ;
  assign n15843 = n1957 | n2995 ;
  assign n15844 = n8931 ^ n3796 ^ 1'b0 ;
  assign n15845 = n15843 | n15844 ;
  assign n15846 = n1000 & ~n3136 ;
  assign n15847 = n8674 ^ n2754 ^ 1'b0 ;
  assign n15848 = n15847 ^ n5383 ^ 1'b0 ;
  assign n15849 = n15846 & ~n15848 ;
  assign n15850 = n6961 & ~n8661 ;
  assign n15851 = n15850 ^ n7145 ^ 1'b0 ;
  assign n15852 = n15851 ^ n8762 ^ 1'b0 ;
  assign n15855 = n3770 ^ n506 ^ 1'b0 ;
  assign n15856 = n14599 & n15855 ;
  assign n15857 = n15856 ^ n12479 ^ 1'b0 ;
  assign n15853 = n10568 ^ n3220 ^ 1'b0 ;
  assign n15854 = n1340 & n15853 ;
  assign n15858 = n15857 ^ n15854 ^ 1'b0 ;
  assign n15859 = ~n9785 & n15858 ;
  assign n15860 = n14905 ^ n6975 ^ 1'b0 ;
  assign n15861 = ~n5298 & n15860 ;
  assign n15862 = ~n3123 & n8944 ;
  assign n15863 = n3396 & ~n8570 ;
  assign n15864 = n15863 ^ n4195 ^ 1'b0 ;
  assign n15865 = ( n643 & ~n6485 ) | ( n643 & n15864 ) | ( ~n6485 & n15864 ) ;
  assign n15866 = ~n3927 & n8197 ;
  assign n15867 = ~n668 & n15866 ;
  assign n15868 = ( n2996 & ~n4180 ) | ( n2996 & n5260 ) | ( ~n4180 & n5260 ) ;
  assign n15869 = n15868 ^ n385 ^ 1'b0 ;
  assign n15870 = ( n1275 & n15867 ) | ( n1275 & n15869 ) | ( n15867 & n15869 ) ;
  assign n15871 = n7047 | n9733 ;
  assign n15873 = n2868 & n15194 ;
  assign n15872 = n1631 & n11979 ;
  assign n15874 = n15873 ^ n15872 ^ 1'b0 ;
  assign n15875 = ~n3248 & n5359 ;
  assign n15876 = ~n8328 & n15875 ;
  assign n15877 = n5420 ^ n2712 ^ 1'b0 ;
  assign n15878 = ~n15876 & n15877 ;
  assign n15879 = n7960 | n8005 ;
  assign n15880 = n15879 ^ n9346 ^ 1'b0 ;
  assign n15881 = n1313 ^ n1208 ^ 1'b0 ;
  assign n15882 = ( n1023 & n5566 ) | ( n1023 & ~n15881 ) | ( n5566 & ~n15881 ) ;
  assign n15883 = n2956 & ~n10159 ;
  assign n15884 = n15883 ^ x213 ^ 1'b0 ;
  assign n15885 = n14742 | n15884 ;
  assign n15886 = n562 & ~n15885 ;
  assign n15887 = ( n8856 & ~n15882 ) | ( n8856 & n15886 ) | ( ~n15882 & n15886 ) ;
  assign n15888 = n3091 & ~n6080 ;
  assign n15889 = ~n3091 & n15888 ;
  assign n15890 = n954 | n15889 ;
  assign n15891 = n954 & ~n15890 ;
  assign n15892 = n4369 | n4379 ;
  assign n15893 = n15892 ^ n800 ^ 1'b0 ;
  assign n15894 = n2325 & ~n15893 ;
  assign n15895 = n15893 & n15894 ;
  assign n15896 = n15895 ^ n5592 ^ 1'b0 ;
  assign n15897 = n15891 | n15896 ;
  assign n15898 = ( n3613 & n5934 ) | ( n3613 & n15897 ) | ( n5934 & n15897 ) ;
  assign n15899 = ~n5839 & n10935 ;
  assign n15900 = ~n11657 & n15899 ;
  assign n15901 = n8062 & n15900 ;
  assign n15902 = n5663 ^ n2910 ^ n1024 ;
  assign n15903 = ( n5267 & ~n6807 ) | ( n5267 & n15902 ) | ( ~n6807 & n15902 ) ;
  assign n15904 = n15903 ^ n9215 ^ 1'b0 ;
  assign n15905 = n8378 | n10028 ;
  assign n15908 = n5205 | n7867 ;
  assign n15906 = n478 | n6757 ;
  assign n15907 = n4950 & ~n15906 ;
  assign n15909 = n15908 ^ n15907 ^ 1'b0 ;
  assign n15910 = n11100 & n15909 ;
  assign n15911 = n14231 ^ n6651 ^ 1'b0 ;
  assign n15912 = ( ~n2710 & n5923 ) | ( ~n2710 & n15911 ) | ( n5923 & n15911 ) ;
  assign n15913 = n12501 ^ n3271 ^ 1'b0 ;
  assign n15914 = n1000 & ~n3374 ;
  assign n15915 = n3705 ^ n2057 ^ 1'b0 ;
  assign n15916 = n15915 ^ n4325 ^ 1'b0 ;
  assign n15917 = n15914 & n15916 ;
  assign n15918 = n3431 | n12344 ;
  assign n15919 = n1134 & ~n15918 ;
  assign n15926 = n3907 & ~n3968 ;
  assign n15920 = n2000 & n7474 ;
  assign n15921 = n7783 ^ n4779 ^ 1'b0 ;
  assign n15922 = n15920 & n15921 ;
  assign n15923 = n15922 ^ n14764 ^ 1'b0 ;
  assign n15924 = x204 & ~n15923 ;
  assign n15925 = n12733 & n15924 ;
  assign n15927 = n15926 ^ n15925 ^ 1'b0 ;
  assign n15928 = n8167 ^ n7277 ^ 1'b0 ;
  assign n15929 = n7402 & ~n9591 ;
  assign n15930 = ~n1584 & n15929 ;
  assign n15931 = n7986 & ~n15930 ;
  assign n15932 = n15931 ^ n12771 ^ n9636 ;
  assign n15933 = ( n3359 & ~n6698 ) | ( n3359 & n12231 ) | ( ~n6698 & n12231 ) ;
  assign n15934 = n4521 & ~n15933 ;
  assign n15935 = n15934 ^ n838 ^ 1'b0 ;
  assign n15936 = n10791 ^ n10640 ^ 1'b0 ;
  assign n15938 = ( n1840 & n3157 ) | ( n1840 & n14655 ) | ( n3157 & n14655 ) ;
  assign n15937 = n6286 ^ n3476 ^ 1'b0 ;
  assign n15939 = n15938 ^ n15937 ^ n4844 ;
  assign n15940 = ~n3107 & n15939 ;
  assign n15941 = ~n15936 & n15940 ;
  assign n15942 = ~n13870 & n15941 ;
  assign n15943 = n635 & n10223 ;
  assign n15944 = ~n15942 & n15943 ;
  assign n15945 = n12749 ^ n7531 ^ n5861 ;
  assign n15946 = ~n3272 & n4398 ;
  assign n15947 = n4538 ^ n1558 ^ 1'b0 ;
  assign n15948 = n4174 & n5739 ;
  assign n15949 = n836 & ~n7071 ;
  assign n15950 = n15949 ^ n357 ^ 1'b0 ;
  assign n15951 = n15948 & ~n15950 ;
  assign n15952 = n15590 & ~n15951 ;
  assign n15953 = n764 | n11772 ;
  assign n15954 = ~n404 & n4154 ;
  assign n15955 = ~n5773 & n15954 ;
  assign n15956 = n2815 | n3265 ;
  assign n15957 = ( n13624 & n15955 ) | ( n13624 & ~n15956 ) | ( n15955 & ~n15956 ) ;
  assign n15958 = n1396 | n9355 ;
  assign n15959 = n15958 ^ n6873 ^ 1'b0 ;
  assign n15960 = n15959 ^ n8463 ^ 1'b0 ;
  assign n15961 = n14212 & n15960 ;
  assign n15962 = n15961 ^ n9879 ^ 1'b0 ;
  assign n15970 = n1843 ^ n1736 ^ 1'b0 ;
  assign n15971 = n15970 ^ n6010 ^ 1'b0 ;
  assign n15965 = n9639 ^ n6553 ^ 1'b0 ;
  assign n15966 = n8065 & ~n15965 ;
  assign n15967 = ~n13196 & n15966 ;
  assign n15963 = x22 & ~n4146 ;
  assign n15964 = n15963 ^ n3043 ^ 1'b0 ;
  assign n15968 = n15967 ^ n15964 ^ 1'b0 ;
  assign n15969 = n3096 & n15968 ;
  assign n15972 = n15971 ^ n15969 ^ 1'b0 ;
  assign n15973 = n13748 & n15972 ;
  assign n15974 = n14634 ^ n5140 ^ 1'b0 ;
  assign n15975 = n6645 & ~n15974 ;
  assign n15976 = n15975 ^ n4083 ^ 1'b0 ;
  assign n15977 = n7260 & ~n9938 ;
  assign n15978 = n15977 ^ n980 ^ 1'b0 ;
  assign n15979 = ( n1381 & ~n13920 ) | ( n1381 & n15978 ) | ( ~n13920 & n15978 ) ;
  assign n15980 = n12767 ^ n881 ^ 1'b0 ;
  assign n15982 = x94 & ~n8484 ;
  assign n15983 = n15982 ^ n1110 ^ 1'b0 ;
  assign n15981 = n9475 ^ n7668 ^ x176 ;
  assign n15984 = n15983 ^ n15981 ^ n3473 ;
  assign n15985 = ~n9242 & n11638 ;
  assign n15986 = ( n486 & n7532 ) | ( n486 & n12044 ) | ( n7532 & n12044 ) ;
  assign n15987 = n4998 ^ n4815 ^ n1411 ;
  assign n15988 = n15987 ^ n6287 ^ 1'b0 ;
  assign n15989 = n11157 & ~n15988 ;
  assign n15990 = n15989 ^ n4015 ^ 1'b0 ;
  assign n15991 = ~n15986 & n15990 ;
  assign n15992 = n4183 & n4308 ;
  assign n15993 = n15992 ^ n5901 ^ 1'b0 ;
  assign n16000 = n11508 | n11615 ;
  assign n15994 = n3716 & ~n5213 ;
  assign n15995 = n15994 ^ n3667 ^ 1'b0 ;
  assign n15996 = n1091 & ~n15995 ;
  assign n15997 = n9950 ^ n4774 ^ 1'b0 ;
  assign n15998 = n15996 & ~n15997 ;
  assign n15999 = x158 & n15998 ;
  assign n16001 = n16000 ^ n15999 ^ 1'b0 ;
  assign n16002 = ~n2176 & n2462 ;
  assign n16003 = n2935 | n16002 ;
  assign n16004 = n9695 ^ n4215 ^ 1'b0 ;
  assign n16005 = n2374 & n16004 ;
  assign n16006 = n16003 | n16005 ;
  assign n16007 = n2751 | n2921 ;
  assign n16008 = n3000 | n16007 ;
  assign n16009 = ~x94 & n587 ;
  assign n16010 = ( n9267 & n10746 ) | ( n9267 & n15130 ) | ( n10746 & n15130 ) ;
  assign n16011 = n3587 & n6318 ;
  assign n16012 = ~n1689 & n16011 ;
  assign n16013 = n16012 ^ n14012 ^ 1'b0 ;
  assign n16014 = n10385 & ~n16013 ;
  assign n16015 = n16014 ^ n4873 ^ 1'b0 ;
  assign n16016 = n8121 ^ n1130 ^ 1'b0 ;
  assign n16017 = n9612 ^ n4521 ^ 1'b0 ;
  assign n16018 = n2272 & n16017 ;
  assign n16019 = n8659 & n16018 ;
  assign n16020 = n513 & ~n11213 ;
  assign n16021 = ~n16019 & n16020 ;
  assign n16022 = n5907 ^ n2134 ^ 1'b0 ;
  assign n16023 = ( n2640 & n2877 ) | ( n2640 & n3506 ) | ( n2877 & n3506 ) ;
  assign n16024 = n5884 ^ n963 ^ 1'b0 ;
  assign n16025 = n326 & ~n16024 ;
  assign n16026 = ~n13600 & n16025 ;
  assign n16027 = n2704 | n7381 ;
  assign n16028 = n2704 & ~n16027 ;
  assign n16029 = ( n1406 & n1453 ) | ( n1406 & n2553 ) | ( n1453 & n2553 ) ;
  assign n16030 = ~n16028 & n16029 ;
  assign n16031 = n16028 & n16030 ;
  assign n16032 = n3326 | n16031 ;
  assign n16033 = n3326 & ~n16032 ;
  assign n16034 = x130 & ~n16033 ;
  assign n16035 = n16033 & n16034 ;
  assign n16036 = n16035 ^ n13377 ^ 1'b0 ;
  assign n16037 = n14468 & ~n16036 ;
  assign n16038 = n12544 ^ n9595 ^ 1'b0 ;
  assign n16039 = ~n7799 & n16038 ;
  assign n16040 = n6962 ^ n5988 ^ n1786 ;
  assign n16041 = n6607 ^ n1571 ^ 1'b0 ;
  assign n16042 = ~x135 & n8526 ;
  assign n16043 = n15141 ^ n1851 ^ 1'b0 ;
  assign n16044 = n7587 & ~n7726 ;
  assign n16045 = n8990 & n16044 ;
  assign n16046 = n15422 & n16045 ;
  assign n16047 = n1900 | n2355 ;
  assign n16048 = n495 | n16047 ;
  assign n16049 = n8259 | n16048 ;
  assign n16050 = n14620 ^ n10662 ^ 1'b0 ;
  assign n16051 = n5159 & ~n16050 ;
  assign n16052 = n8613 & ~n10984 ;
  assign n16053 = n9112 ^ n1988 ^ 1'b0 ;
  assign n16054 = n4284 & n16053 ;
  assign n16055 = ( n7788 & n16052 ) | ( n7788 & n16054 ) | ( n16052 & n16054 ) ;
  assign n16057 = n395 & ~n604 ;
  assign n16058 = n12514 & n16057 ;
  assign n16059 = n16058 ^ n365 ^ 1'b0 ;
  assign n16060 = ~n9399 & n16059 ;
  assign n16061 = n15150 & n16060 ;
  assign n16056 = n1712 | n5445 ;
  assign n16062 = n16061 ^ n16056 ^ 1'b0 ;
  assign n16063 = ( x184 & n926 ) | ( x184 & ~n5175 ) | ( n926 & ~n5175 ) ;
  assign n16064 = n9873 & n16063 ;
  assign n16065 = n5413 & ~n13375 ;
  assign n16066 = n16065 ^ n15465 ^ 1'b0 ;
  assign n16067 = n13893 ^ n4481 ^ 1'b0 ;
  assign n16068 = n13630 & n16067 ;
  assign n16069 = n6337 ^ n4241 ^ 1'b0 ;
  assign n16070 = x211 & ~n16069 ;
  assign n16071 = n8235 | n16070 ;
  assign n16072 = n13742 ^ n7705 ^ 1'b0 ;
  assign n16073 = n16071 & ~n16072 ;
  assign n16074 = ~n3894 & n13023 ;
  assign n16075 = n16074 ^ x168 ^ 1'b0 ;
  assign n16076 = n16075 ^ n555 ^ 1'b0 ;
  assign n16077 = n16073 & ~n16076 ;
  assign n16078 = n16077 ^ n606 ^ 1'b0 ;
  assign n16079 = n16078 ^ n2922 ^ 1'b0 ;
  assign n16080 = n16079 ^ n6058 ^ n5477 ;
  assign n16081 = n5912 & ~n8972 ;
  assign n16082 = n16081 ^ n7649 ^ 1'b0 ;
  assign n16083 = n7046 & ~n16082 ;
  assign n16084 = n6543 ^ n5600 ^ 1'b0 ;
  assign n16085 = n6523 | n16084 ;
  assign n16086 = n8729 | n16085 ;
  assign n16087 = n14856 | n16086 ;
  assign n16088 = n11543 ^ n5663 ^ 1'b0 ;
  assign n16089 = n5922 & n6926 ;
  assign n16090 = n16089 ^ n5029 ^ 1'b0 ;
  assign n16091 = n16090 ^ n874 ^ 1'b0 ;
  assign n16092 = n16091 ^ n1791 ^ 1'b0 ;
  assign n16093 = n16088 | n16092 ;
  assign n16094 = ( n14142 & ~n16087 ) | ( n14142 & n16093 ) | ( ~n16087 & n16093 ) ;
  assign n16095 = ~n4455 & n16094 ;
  assign n16096 = n9154 ^ n3152 ^ 1'b0 ;
  assign n16097 = ( n2286 & ~n9295 ) | ( n2286 & n16096 ) | ( ~n9295 & n16096 ) ;
  assign n16098 = n15846 ^ n1879 ^ 1'b0 ;
  assign n16099 = n16098 ^ n13137 ^ 1'b0 ;
  assign n16100 = n7794 ^ n5725 ^ 1'b0 ;
  assign n16101 = n10162 ^ x118 ^ 1'b0 ;
  assign n16102 = n1022 & n16101 ;
  assign n16103 = n16100 & n16102 ;
  assign n16104 = n5967 & ~n16103 ;
  assign n16105 = ( n1281 & n7532 ) | ( n1281 & ~n12178 ) | ( n7532 & ~n12178 ) ;
  assign n16106 = n1153 ^ n300 ^ 1'b0 ;
  assign n16107 = ~n12436 & n16106 ;
  assign n16110 = n12372 ^ x40 ^ 1'b0 ;
  assign n16108 = n2698 ^ n1203 ^ 1'b0 ;
  assign n16109 = n5319 | n16108 ;
  assign n16111 = n16110 ^ n16109 ^ n8712 ;
  assign n16112 = n5653 | n7791 ;
  assign n16113 = n14613 ^ n12029 ^ n9157 ;
  assign n16114 = ~n5155 & n5262 ;
  assign n16115 = n13223 & n16114 ;
  assign n16116 = n8432 & ~n14085 ;
  assign n16129 = n4516 & ~n14388 ;
  assign n16127 = n4684 ^ n749 ^ 1'b0 ;
  assign n16128 = n16127 ^ n11105 ^ n5140 ;
  assign n16130 = n16129 ^ n16128 ^ 1'b0 ;
  assign n16117 = n9508 ^ n4985 ^ 1'b0 ;
  assign n16118 = n16002 & ~n16117 ;
  assign n16121 = n2441 ^ n2153 ^ 1'b0 ;
  assign n16122 = n4039 | n16121 ;
  assign n16119 = n1724 & n6081 ;
  assign n16120 = n3435 & n16119 ;
  assign n16123 = n16122 ^ n16120 ^ 1'b0 ;
  assign n16124 = n16123 ^ n1004 ^ 1'b0 ;
  assign n16125 = n16124 ^ n9501 ^ 1'b0 ;
  assign n16126 = n16118 & n16125 ;
  assign n16131 = n16130 ^ n16126 ^ n7344 ;
  assign n16132 = ~n267 & n6865 ;
  assign n16133 = n15970 & n16132 ;
  assign n16134 = n6623 & ~n16133 ;
  assign n16135 = n12970 ^ n7928 ^ 1'b0 ;
  assign n16136 = n627 & n16135 ;
  assign n16137 = ~n6453 & n12559 ;
  assign n16141 = n3210 & n9403 ;
  assign n16142 = ~x42 & n16141 ;
  assign n16138 = n2791 ^ n2708 ^ 1'b0 ;
  assign n16139 = n6011 & n16138 ;
  assign n16140 = n12072 & ~n16139 ;
  assign n16143 = n16142 ^ n16140 ^ n2212 ;
  assign n16144 = n16143 ^ n2855 ^ 1'b0 ;
  assign n16145 = n15067 ^ n4775 ^ 1'b0 ;
  assign n16146 = n5311 | n16145 ;
  assign n16147 = n8692 ^ n3430 ^ 1'b0 ;
  assign n16148 = n3606 | n4597 ;
  assign n16149 = n13920 ^ n12116 ^ 1'b0 ;
  assign n16150 = n16148 & n16149 ;
  assign n16151 = n16147 & n16150 ;
  assign n16152 = n14632 ^ n14479 ^ 1'b0 ;
  assign n16153 = ~n11045 & n16152 ;
  assign n16154 = n2738 & n11108 ;
  assign n16155 = ~n1798 & n16154 ;
  assign n16156 = n16155 ^ n14138 ^ n1026 ;
  assign n16157 = n11870 ^ n9430 ^ 1'b0 ;
  assign n16158 = n947 & ~n15401 ;
  assign n16159 = n16158 ^ n5217 ^ 1'b0 ;
  assign n16160 = n5927 & ~n16159 ;
  assign n16161 = n16160 ^ n5324 ^ 1'b0 ;
  assign n16162 = ~n2806 & n12289 ;
  assign n16163 = n16162 ^ n3295 ^ 1'b0 ;
  assign n16164 = n13347 ^ n10320 ^ n3720 ;
  assign n16165 = n16164 ^ n7877 ^ 1'b0 ;
  assign n16166 = n10605 ^ x88 ^ 1'b0 ;
  assign n16167 = x118 & ~n5431 ;
  assign n16168 = n16167 ^ n2988 ^ 1'b0 ;
  assign n16169 = n16166 | n16168 ;
  assign n16170 = n3910 ^ n3438 ^ n1880 ;
  assign n16171 = n16170 ^ n12765 ^ n1527 ;
  assign n16172 = n9362 & n16171 ;
  assign n16173 = ~n7423 & n11596 ;
  assign n16174 = n11073 & n11290 ;
  assign n16175 = n5283 & n5590 ;
  assign n16176 = n7267 & n16175 ;
  assign n16177 = x101 & ~n16176 ;
  assign n16179 = n2592 ^ n1144 ^ 1'b0 ;
  assign n16180 = n16179 ^ n10555 ^ 1'b0 ;
  assign n16178 = n4338 & n8356 ;
  assign n16181 = n16180 ^ n16178 ^ 1'b0 ;
  assign n16182 = x216 & ~n8972 ;
  assign n16183 = ~n2552 & n16182 ;
  assign n16184 = n8134 ^ n1006 ^ 1'b0 ;
  assign n16185 = ( x253 & n6007 ) | ( x253 & ~n6278 ) | ( n6007 & ~n6278 ) ;
  assign n16186 = ( n15299 & n16184 ) | ( n15299 & ~n16185 ) | ( n16184 & ~n16185 ) ;
  assign n16187 = n16186 ^ n15793 ^ n5283 ;
  assign n16188 = n10771 ^ n4002 ^ 1'b0 ;
  assign n16189 = n14656 ^ n7087 ^ n2877 ;
  assign n16190 = n16189 ^ n15219 ^ 1'b0 ;
  assign n16191 = n5719 ^ n668 ^ 1'b0 ;
  assign n16192 = n1021 & n16191 ;
  assign n16193 = n15747 & n16192 ;
  assign n16194 = n12044 & n16193 ;
  assign n16195 = n12415 ^ n5028 ^ 1'b0 ;
  assign n16196 = ~n6671 & n16195 ;
  assign n16197 = n16196 ^ n2720 ^ 1'b0 ;
  assign n16198 = n9920 | n16197 ;
  assign n16199 = n16198 ^ n11026 ^ 1'b0 ;
  assign n16200 = ~n5731 & n16199 ;
  assign n16201 = n16194 & n16200 ;
  assign n16202 = n4300 & n4970 ;
  assign n16203 = ~n2363 & n16202 ;
  assign n16204 = n16203 ^ n673 ^ 1'b0 ;
  assign n16205 = n1868 & ~n16204 ;
  assign n16206 = n5365 | n11773 ;
  assign n16207 = n16206 ^ n2609 ^ 1'b0 ;
  assign n16208 = n3085 | n11421 ;
  assign n16209 = n16208 ^ n1473 ^ 1'b0 ;
  assign n16210 = ~n9468 & n16209 ;
  assign n16211 = n16210 ^ n11262 ^ 1'b0 ;
  assign n16212 = n429 & ~n16211 ;
  assign n16213 = n16212 ^ n14146 ^ 1'b0 ;
  assign n16214 = n16207 & n16213 ;
  assign n16215 = ~n16205 & n16214 ;
  assign n16216 = n9232 ^ x216 ^ 1'b0 ;
  assign n16217 = ~n11400 & n16216 ;
  assign n16218 = ( n3891 & ~n10127 ) | ( n3891 & n16217 ) | ( ~n10127 & n16217 ) ;
  assign n16219 = ~n5531 & n13689 ;
  assign n16220 = n16219 ^ n3943 ^ 1'b0 ;
  assign n16221 = n7584 ^ n6141 ^ n5724 ;
  assign n16222 = ~n4286 & n16221 ;
  assign n16223 = n9724 & n12469 ;
  assign n16224 = n6119 ^ n1698 ^ 1'b0 ;
  assign n16225 = ( n880 & ~n4990 ) | ( n880 & n16224 ) | ( ~n4990 & n16224 ) ;
  assign n16226 = n3321 & ~n3435 ;
  assign n16227 = n11895 | n16221 ;
  assign n16228 = ~n6729 & n14097 ;
  assign n16229 = ( n1209 & ~n6604 ) | ( n1209 & n8911 ) | ( ~n6604 & n8911 ) ;
  assign n16230 = n7958 & n14359 ;
  assign n16231 = ( n1996 & n13527 ) | ( n1996 & n13656 ) | ( n13527 & n13656 ) ;
  assign n16232 = n10274 | n13513 ;
  assign n16233 = n16232 ^ x123 ^ 1'b0 ;
  assign n16234 = ( ~n2315 & n7396 ) | ( ~n2315 & n16233 ) | ( n7396 & n16233 ) ;
  assign n16236 = x161 | n2787 ;
  assign n16237 = n16236 ^ n917 ^ 1'b0 ;
  assign n16235 = n4081 ^ n1132 ^ 1'b0 ;
  assign n16238 = n16237 ^ n16235 ^ n7253 ;
  assign n16239 = n5233 & n16238 ;
  assign n16240 = n16239 ^ n10825 ^ 1'b0 ;
  assign n16241 = n14708 ^ n6443 ^ 1'b0 ;
  assign n16242 = n3096 & n16241 ;
  assign n16243 = n15756 ^ n15246 ^ 1'b0 ;
  assign n16244 = n13190 & ~n16243 ;
  assign n16245 = n5146 ^ n4278 ^ 1'b0 ;
  assign n16246 = n10511 ^ n5824 ^ 1'b0 ;
  assign n16247 = ~n3431 & n16246 ;
  assign n16248 = n14625 ^ n6361 ^ 1'b0 ;
  assign n16249 = n16247 & n16248 ;
  assign n16250 = ~n9072 & n16249 ;
  assign n16251 = ( n15390 & ~n16245 ) | ( n15390 & n16250 ) | ( ~n16245 & n16250 ) ;
  assign n16252 = n2108 & n12850 ;
  assign n16253 = ( n3345 & n4976 ) | ( n3345 & n12876 ) | ( n4976 & n12876 ) ;
  assign n16254 = ~x65 & n16253 ;
  assign n16255 = n13570 & n16254 ;
  assign n16258 = x37 & n5958 ;
  assign n16259 = n16258 ^ n11906 ^ 1'b0 ;
  assign n16260 = n6668 ^ x4 ^ 1'b0 ;
  assign n16261 = n16259 | n16260 ;
  assign n16256 = n9661 & ~n12749 ;
  assign n16257 = ~n2754 & n16256 ;
  assign n16262 = n16261 ^ n16257 ^ 1'b0 ;
  assign n16263 = n8562 | n16262 ;
  assign n16264 = n16263 ^ n16129 ^ 1'b0 ;
  assign n16265 = n16264 ^ n12639 ^ n6988 ;
  assign n16266 = n702 & ~n8423 ;
  assign n16267 = n674 | n14042 ;
  assign n16268 = n1798 & n5343 ;
  assign n16269 = ~n5618 & n16268 ;
  assign n16270 = n12557 | n16269 ;
  assign n16271 = n16267 & ~n16270 ;
  assign n16272 = n1188 | n8548 ;
  assign n16273 = n6743 | n16272 ;
  assign n16274 = n16273 ^ n15701 ^ 1'b0 ;
  assign n16275 = n7560 ^ n6295 ^ 1'b0 ;
  assign n16276 = ~n16274 & n16275 ;
  assign n16277 = n6051 ^ n1762 ^ 1'b0 ;
  assign n16278 = x85 & ~n16277 ;
  assign n16279 = x242 | n702 ;
  assign n16280 = ~n4962 & n16279 ;
  assign n16283 = ~n1098 & n3660 ;
  assign n16284 = ~n5720 & n16283 ;
  assign n16281 = n897 & n2945 ;
  assign n16282 = n5523 & n16281 ;
  assign n16285 = n16284 ^ n16282 ^ 1'b0 ;
  assign n16286 = n1478 & ~n14331 ;
  assign n16287 = n16286 ^ n911 ^ 1'b0 ;
  assign n16288 = n12153 & n16287 ;
  assign n16289 = n3685 & n10008 ;
  assign n16290 = ( n16285 & ~n16288 ) | ( n16285 & n16289 ) | ( ~n16288 & n16289 ) ;
  assign n16291 = n1197 & ~n11382 ;
  assign n16292 = n16291 ^ n11966 ^ 1'b0 ;
  assign n16293 = n9361 | n16292 ;
  assign n16294 = n11258 & ~n16293 ;
  assign n16295 = n1900 | n5063 ;
  assign n16296 = n16295 ^ n13500 ^ 1'b0 ;
  assign n16297 = n10215 & ~n16296 ;
  assign n16298 = n8295 ^ n7557 ^ 1'b0 ;
  assign n16299 = n9581 ^ n6241 ^ 1'b0 ;
  assign n16300 = n15395 ^ n5304 ^ 1'b0 ;
  assign n16301 = ~n16299 & n16300 ;
  assign n16302 = ~n6584 & n9165 ;
  assign n16303 = ~n12727 & n14563 ;
  assign n16304 = n1234 & n2489 ;
  assign n16305 = n16304 ^ n1153 ^ 1'b0 ;
  assign n16306 = n4152 ^ n1350 ^ 1'b0 ;
  assign n16307 = n16305 & n16306 ;
  assign n16308 = n16307 ^ n2230 ^ 1'b0 ;
  assign n16309 = n12074 & n16308 ;
  assign n16310 = n13692 ^ n12279 ^ 1'b0 ;
  assign n16311 = ~n10001 & n16310 ;
  assign n16312 = n453 | n12812 ;
  assign n16313 = n13752 & ~n16312 ;
  assign n16314 = n8763 | n13440 ;
  assign n16315 = n3430 | n7171 ;
  assign n16316 = ~x132 & n2081 ;
  assign n16317 = n9157 & ~n16316 ;
  assign n16318 = n16317 ^ n12247 ^ 1'b0 ;
  assign n16319 = n2561 ^ n1315 ^ 1'b0 ;
  assign n16320 = n4994 | n16319 ;
  assign n16321 = n3744 | n13656 ;
  assign n16322 = n16321 ^ n4132 ^ 1'b0 ;
  assign n16323 = n6391 | n14652 ;
  assign n16324 = n16323 ^ n2074 ^ 1'b0 ;
  assign n16325 = ( n755 & ~n2034 ) | ( n755 & n3689 ) | ( ~n2034 & n3689 ) ;
  assign n16326 = ( n1411 & n1667 ) | ( n1411 & n16325 ) | ( n1667 & n16325 ) ;
  assign n16327 = n16326 ^ n11617 ^ 1'b0 ;
  assign n16328 = ~n3201 & n16327 ;
  assign n16329 = n3198 | n16024 ;
  assign n16330 = n16329 ^ n14711 ^ 1'b0 ;
  assign n16331 = n16328 & ~n16330 ;
  assign n16332 = n9648 ^ n9475 ^ 1'b0 ;
  assign n16333 = n3389 & ~n16332 ;
  assign n16334 = n9203 ^ x30 ^ 1'b0 ;
  assign n16335 = n16333 & ~n16334 ;
  assign n16336 = n5508 | n7632 ;
  assign n16337 = n16335 | n16336 ;
  assign n16338 = n1525 ^ x17 ^ 1'b0 ;
  assign n16339 = n12647 & n16338 ;
  assign n16340 = n14332 ^ n1861 ^ 1'b0 ;
  assign n16341 = n12007 | n16340 ;
  assign n16342 = n10965 & ~n12263 ;
  assign n16343 = n10382 & n16342 ;
  assign n16344 = n14985 | n16343 ;
  assign n16345 = n1998 & ~n13662 ;
  assign n16346 = n16345 ^ n4932 ^ 1'b0 ;
  assign n16347 = n11357 ^ n8763 ^ 1'b0 ;
  assign n16348 = n5304 & n16347 ;
  assign n16349 = n8134 | n16348 ;
  assign n16350 = n16237 ^ n7608 ^ 1'b0 ;
  assign n16351 = n3148 & n16350 ;
  assign n16352 = n2259 & n16351 ;
  assign n16353 = n8029 ^ n7820 ^ 1'b0 ;
  assign n16354 = ~n5804 & n16353 ;
  assign n16355 = n16352 & n16354 ;
  assign n16356 = n16355 ^ n1782 ^ 1'b0 ;
  assign n16357 = n13311 | n14648 ;
  assign n16358 = x67 & ~n292 ;
  assign n16359 = n16358 ^ n836 ^ 1'b0 ;
  assign n16360 = n732 ^ x178 ^ 1'b0 ;
  assign n16361 = n16359 | n16360 ;
  assign n16362 = n8107 ^ n5050 ^ 1'b0 ;
  assign n16363 = n16362 ^ n12261 ^ n10760 ;
  assign n16364 = n3338 & n6987 ;
  assign n16365 = n16364 ^ n2465 ^ 1'b0 ;
  assign n16366 = ~n1064 & n11355 ;
  assign n16367 = n16229 ^ n14617 ^ n9102 ;
  assign n16368 = n5209 & n10595 ;
  assign n16369 = n3777 & n16368 ;
  assign n16370 = ~n10847 & n16369 ;
  assign n16371 = n9447 & ~n14359 ;
  assign n16372 = n16371 ^ x135 ^ 1'b0 ;
  assign n16373 = ( n2148 & n12741 ) | ( n2148 & ~n16372 ) | ( n12741 & ~n16372 ) ;
  assign n16374 = n16373 ^ n6917 ^ 1'b0 ;
  assign n16375 = n7312 & n16374 ;
  assign n16376 = n3441 & n7206 ;
  assign n16377 = ~n716 & n16376 ;
  assign n16378 = n16377 ^ n12212 ^ 1'b0 ;
  assign n16379 = n7811 & ~n9136 ;
  assign n16380 = n4732 & ~n16379 ;
  assign n16381 = n6558 & n16380 ;
  assign n16382 = ( ~n6627 & n12963 ) | ( ~n6627 & n16381 ) | ( n12963 & n16381 ) ;
  assign n16383 = n4274 ^ n3160 ^ x247 ;
  assign n16384 = n16383 ^ n3136 ^ 1'b0 ;
  assign n16385 = n4628 ^ n2470 ^ 1'b0 ;
  assign n16386 = n8327 & n16385 ;
  assign n16387 = n16384 & n16386 ;
  assign n16388 = n13877 ^ n2389 ^ 1'b0 ;
  assign n16389 = n10973 & ~n16388 ;
  assign n16391 = n6904 ^ n298 ^ 1'b0 ;
  assign n16390 = n2756 & ~n13083 ;
  assign n16392 = n16391 ^ n16390 ^ n2712 ;
  assign n16393 = n12914 ^ n9226 ^ 1'b0 ;
  assign n16394 = n14886 & n16393 ;
  assign n16395 = n8440 ^ n3081 ^ 1'b0 ;
  assign n16399 = n9759 ^ n7384 ^ 1'b0 ;
  assign n16400 = ~n9678 & n16399 ;
  assign n16401 = n16400 ^ n11309 ^ 1'b0 ;
  assign n16402 = n5598 | n16401 ;
  assign n16403 = n7987 | n8919 ;
  assign n16404 = n6242 ^ n3279 ^ 1'b0 ;
  assign n16405 = n16403 & n16404 ;
  assign n16406 = ~n16402 & n16405 ;
  assign n16407 = n8363 & n16406 ;
  assign n16396 = x222 ^ x124 ^ 1'b0 ;
  assign n16397 = n16396 ^ n8073 ^ 1'b0 ;
  assign n16398 = ~n13091 & n16397 ;
  assign n16408 = n16407 ^ n16398 ^ 1'b0 ;
  assign n16410 = ( n2187 & n3109 ) | ( n2187 & ~n9451 ) | ( n3109 & ~n9451 ) ;
  assign n16409 = ~n7107 & n15651 ;
  assign n16411 = n16410 ^ n16409 ^ n4251 ;
  assign n16414 = n3725 | n10810 ;
  assign n16415 = n3504 | n16414 ;
  assign n16412 = n6711 & n7992 ;
  assign n16413 = ~n2465 & n16412 ;
  assign n16416 = n16415 ^ n16413 ^ n714 ;
  assign n16417 = ~n7764 & n15653 ;
  assign n16418 = n16417 ^ n8690 ^ 1'b0 ;
  assign n16419 = n16416 | n16418 ;
  assign n16420 = ~n11375 & n16419 ;
  assign n16421 = n7765 ^ n1776 ^ 1'b0 ;
  assign n16422 = ~n2961 & n16421 ;
  assign n16423 = n11213 | n14523 ;
  assign n16424 = n16423 ^ n3947 ^ 1'b0 ;
  assign n16425 = n308 | n3202 ;
  assign n16426 = n16425 ^ n1217 ^ 1'b0 ;
  assign n16427 = n16426 ^ n8678 ^ n917 ;
  assign n16429 = n7824 ^ n6607 ^ n3872 ;
  assign n16430 = n13966 & n16429 ;
  assign n16428 = n8126 & n14504 ;
  assign n16431 = n16430 ^ n16428 ^ 1'b0 ;
  assign n16432 = n1995 | n14930 ;
  assign n16433 = n8697 ^ n1328 ^ 1'b0 ;
  assign n16434 = n15473 ^ n773 ^ 1'b0 ;
  assign n16435 = ~n6402 & n16434 ;
  assign n16436 = ~n11391 & n12800 ;
  assign n16437 = n4409 & n16436 ;
  assign n16438 = n12176 ^ n1455 ^ 1'b0 ;
  assign n16439 = n11906 ^ n1253 ^ 1'b0 ;
  assign n16440 = n16439 ^ n13686 ^ n3010 ;
  assign n16441 = n11351 ^ n7305 ^ 1'b0 ;
  assign n16442 = n3450 & ~n16441 ;
  assign n16443 = n16442 ^ n14982 ^ 1'b0 ;
  assign n16444 = n3904 & ~n8707 ;
  assign n16445 = ~n7251 & n8020 ;
  assign n16446 = n16444 & n16445 ;
  assign n16447 = n8404 & n12435 ;
  assign n16448 = n7788 & n16447 ;
  assign n16449 = n2660 | n13801 ;
  assign n16450 = n16426 ^ n10445 ^ n1249 ;
  assign n16451 = ( n2638 & ~n9937 ) | ( n2638 & n16450 ) | ( ~n9937 & n16450 ) ;
  assign n16452 = n9755 ^ n7336 ^ 1'b0 ;
  assign n16453 = n4117 & n16452 ;
  assign n16454 = ~x169 & n16453 ;
  assign n16455 = n16454 ^ n11103 ^ n6015 ;
  assign n16456 = ~n3804 & n8495 ;
  assign n16457 = n8029 & n16456 ;
  assign n16458 = n7369 & ~n16457 ;
  assign n16459 = n11045 & n16458 ;
  assign n16460 = n6295 | n14243 ;
  assign n16461 = n2751 | n7048 ;
  assign n16462 = n15546 | n16461 ;
  assign n16463 = n3794 ^ n2606 ^ 1'b0 ;
  assign n16464 = ~n2873 & n16463 ;
  assign n16465 = n5455 & n16464 ;
  assign n16466 = n7570 & n16465 ;
  assign n16467 = n8515 & n16466 ;
  assign n16468 = n4735 | n13880 ;
  assign n16469 = ( n2996 & n3881 ) | ( n2996 & n9534 ) | ( n3881 & n9534 ) ;
  assign n16470 = ( n1793 & n16468 ) | ( n1793 & ~n16469 ) | ( n16468 & ~n16469 ) ;
  assign n16471 = n4309 & ~n7817 ;
  assign n16472 = n16471 ^ x234 ^ 1'b0 ;
  assign n16473 = n16472 ^ n11956 ^ 1'b0 ;
  assign n16474 = ~n6592 & n16473 ;
  assign n16475 = n10560 & n16474 ;
  assign n16476 = n16475 ^ n1199 ^ 1'b0 ;
  assign n16477 = ~n604 & n2650 ;
  assign n16478 = n12070 & n16477 ;
  assign n16479 = n16478 ^ n1228 ^ 1'b0 ;
  assign n16480 = ~n4344 & n5626 ;
  assign n16481 = n11511 & ~n16480 ;
  assign n16482 = ~n967 & n4207 ;
  assign n16483 = n16482 ^ n7673 ^ n5778 ;
  assign n16484 = n16483 ^ n15350 ^ 1'b0 ;
  assign n16485 = ( x122 & n8516 ) | ( x122 & ~n8923 ) | ( n8516 & ~n8923 ) ;
  assign n16486 = n16485 ^ n15608 ^ 1'b0 ;
  assign n16487 = n9500 ^ n3274 ^ 1'b0 ;
  assign n16488 = n14855 & n16487 ;
  assign n16489 = n3743 ^ x174 ^ 1'b0 ;
  assign n16490 = ( n12133 & n12923 ) | ( n12133 & n16489 ) | ( n12923 & n16489 ) ;
  assign n16491 = ( n674 & n4445 ) | ( n674 & n6088 ) | ( n4445 & n6088 ) ;
  assign n16492 = n5479 & n16491 ;
  assign n16493 = n16492 ^ n8118 ^ 1'b0 ;
  assign n16494 = n1190 | n8174 ;
  assign n16495 = n2582 | n16494 ;
  assign n16496 = n16495 ^ n11201 ^ 1'b0 ;
  assign n16497 = ~n3919 & n12576 ;
  assign n16498 = n16496 & n16497 ;
  assign n16499 = n8671 & ~n13024 ;
  assign n16500 = n11596 & ~n16359 ;
  assign n16501 = n16500 ^ n8409 ^ 1'b0 ;
  assign n16502 = n2749 & n15440 ;
  assign n16503 = ( n6849 & n12130 ) | ( n6849 & n16129 ) | ( n12130 & n16129 ) ;
  assign n16504 = n5375 | n16503 ;
  assign n16505 = n16504 ^ n4174 ^ 1'b0 ;
  assign n16506 = n1142 | n16505 ;
  assign n16507 = n8295 ^ n1442 ^ 1'b0 ;
  assign n16508 = n7028 | n15737 ;
  assign n16509 = n9048 & ~n16508 ;
  assign n16510 = n8708 | n11039 ;
  assign n16511 = ( n6273 & ~n11773 ) | ( n6273 & n14337 ) | ( ~n11773 & n14337 ) ;
  assign n16512 = n9550 ^ n8076 ^ 1'b0 ;
  assign n16513 = n7871 ^ n1967 ^ 1'b0 ;
  assign n16514 = n3239 & n16513 ;
  assign n16515 = ~n16512 & n16514 ;
  assign n16516 = n16001 | n16515 ;
  assign n16517 = n13732 ^ n4405 ^ 1'b0 ;
  assign n16518 = n15565 ^ n9795 ^ 1'b0 ;
  assign n16519 = n16517 & n16518 ;
  assign n16520 = ~n4749 & n6910 ;
  assign n16521 = n16520 ^ n6748 ^ 1'b0 ;
  assign n16522 = n11898 & n16521 ;
  assign n16523 = n16522 ^ n1265 ^ 1'b0 ;
  assign n16524 = ( ~n8405 & n11621 ) | ( ~n8405 & n16523 ) | ( n11621 & n16523 ) ;
  assign n16525 = n16519 & n16524 ;
  assign n16526 = n12319 ^ n3489 ^ 1'b0 ;
  assign n16527 = n16392 & n16526 ;
  assign n16528 = n1750 | n6371 ;
  assign n16529 = n14677 ^ n6488 ^ 1'b0 ;
  assign n16530 = n9995 | n16529 ;
  assign n16531 = n8016 & n12108 ;
  assign n16532 = n16531 ^ n6593 ^ 1'b0 ;
  assign n16533 = ~n2555 & n8549 ;
  assign n16534 = n16533 ^ n2728 ^ 1'b0 ;
  assign n16535 = ~n5738 & n16534 ;
  assign n16536 = n16535 ^ n13715 ^ 1'b0 ;
  assign n16537 = ~n4094 & n16536 ;
  assign n16538 = n16537 ^ x247 ^ 1'b0 ;
  assign n16539 = ( n672 & n11737 ) | ( n672 & n16538 ) | ( n11737 & n16538 ) ;
  assign n16540 = ( n3404 & n14005 ) | ( n3404 & n16539 ) | ( n14005 & n16539 ) ;
  assign n16541 = n16532 & ~n16540 ;
  assign n16542 = ~n14338 & n16541 ;
  assign n16543 = n3419 & ~n6371 ;
  assign n16544 = n698 & n16543 ;
  assign n16545 = n9833 & n16544 ;
  assign n16546 = n4300 & n6745 ;
  assign n16547 = n11821 & n16546 ;
  assign n16548 = ~n5638 & n8340 ;
  assign n16549 = n16548 ^ n1829 ^ 1'b0 ;
  assign n16550 = n7014 & ~n9957 ;
  assign n16551 = n16550 ^ n5519 ^ 1'b0 ;
  assign n16552 = n3133 | n16551 ;
  assign n16553 = n4289 | n10260 ;
  assign n16558 = n6166 & ~n16269 ;
  assign n16554 = n1590 & n3174 ;
  assign n16555 = ~n6098 & n16554 ;
  assign n16556 = n7558 ^ n2829 ^ 1'b0 ;
  assign n16557 = n16555 | n16556 ;
  assign n16559 = n16558 ^ n16557 ^ 1'b0 ;
  assign n16560 = n9407 | n16559 ;
  assign n16561 = ~n9938 & n13347 ;
  assign n16562 = ( n3374 & n5825 ) | ( n3374 & n10565 ) | ( n5825 & n10565 ) ;
  assign n16563 = n10336 | n16562 ;
  assign n16564 = n7405 | n16563 ;
  assign n16565 = n16552 ^ n1148 ^ 1'b0 ;
  assign n16566 = n16564 | n16565 ;
  assign n16571 = n851 | n9927 ;
  assign n16569 = ( n1272 & n2569 ) | ( n1272 & ~n5513 ) | ( n2569 & ~n5513 ) ;
  assign n16568 = n2132 | n9581 ;
  assign n16570 = n16569 ^ n16568 ^ 1'b0 ;
  assign n16567 = n365 | n8410 ;
  assign n16572 = n16571 ^ n16570 ^ n16567 ;
  assign n16573 = n7324 ^ n1086 ^ 1'b0 ;
  assign n16574 = ~n14073 & n16573 ;
  assign n16575 = n16574 ^ n11108 ^ 1'b0 ;
  assign n16576 = ~n5512 & n11124 ;
  assign n16577 = n6586 & ~n9077 ;
  assign n16578 = n3685 ^ n455 ^ 1'b0 ;
  assign n16579 = ( n9961 & n15351 ) | ( n9961 & ~n16578 ) | ( n15351 & ~n16578 ) ;
  assign n16580 = n718 & ~n14655 ;
  assign n16581 = n1677 & ~n8086 ;
  assign n16582 = n12762 ^ n10379 ^ 1'b0 ;
  assign n16583 = n3686 & ~n16582 ;
  assign n16584 = n16583 ^ n1136 ^ 1'b0 ;
  assign n16585 = n5976 | n6732 ;
  assign n16586 = n9358 | n12221 ;
  assign n16587 = n9479 ^ n9148 ^ 1'b0 ;
  assign n16588 = n14596 & ~n16587 ;
  assign n16589 = n16586 & n16588 ;
  assign n16590 = n1250 | n4995 ;
  assign n16591 = n2601 & ~n16590 ;
  assign n16593 = n7578 | n12899 ;
  assign n16594 = n16593 ^ n2850 ^ 1'b0 ;
  assign n16592 = n5637 | n13864 ;
  assign n16595 = n16594 ^ n16592 ^ 1'b0 ;
  assign n16596 = ( ~n505 & n9374 ) | ( ~n505 & n10480 ) | ( n9374 & n10480 ) ;
  assign n16597 = ( n13881 & n14563 ) | ( n13881 & n16596 ) | ( n14563 & n16596 ) ;
  assign n16598 = ( ~n5592 & n16595 ) | ( ~n5592 & n16597 ) | ( n16595 & n16597 ) ;
  assign n16604 = n12011 ^ n8058 ^ n3470 ;
  assign n16602 = n1991 & ~n8828 ;
  assign n16603 = ~n8512 & n16602 ;
  assign n16605 = n16604 ^ n16603 ^ 1'b0 ;
  assign n16599 = n3721 & ~n10785 ;
  assign n16600 = n16599 ^ n3029 ^ 1'b0 ;
  assign n16601 = n6202 | n16600 ;
  assign n16606 = n16605 ^ n16601 ^ n3299 ;
  assign n16607 = ( n1500 & n3504 ) | ( n1500 & ~n7783 ) | ( n3504 & ~n7783 ) ;
  assign n16608 = n9672 & ~n13197 ;
  assign n16609 = n11842 ^ n4054 ^ 1'b0 ;
  assign n16610 = ~n8077 & n16609 ;
  assign n16611 = n16610 ^ n16234 ^ 1'b0 ;
  assign n16612 = ~n16608 & n16611 ;
  assign n16613 = n3976 & ~n6286 ;
  assign n16614 = n3147 & n16613 ;
  assign n16615 = n8900 ^ n2309 ^ 1'b0 ;
  assign n16616 = x43 & ~n16615 ;
  assign n16617 = n2181 | n3678 ;
  assign n16618 = ~n7339 & n16617 ;
  assign n16619 = n4207 ^ n3911 ^ n3241 ;
  assign n16620 = n4891 & n16619 ;
  assign n16621 = n16620 ^ n12121 ^ 1'b0 ;
  assign n16622 = ( n1260 & n16618 ) | ( n1260 & ~n16621 ) | ( n16618 & ~n16621 ) ;
  assign n16623 = n6559 ^ x209 ^ 1'b0 ;
  assign n16624 = n2922 & n7536 ;
  assign n16625 = n12867 ^ n6676 ^ 1'b0 ;
  assign n16626 = ( n3077 & n7093 ) | ( n3077 & ~n9759 ) | ( n7093 & ~n9759 ) ;
  assign n16627 = n11248 ^ n9802 ^ 1'b0 ;
  assign n16628 = n16626 & n16627 ;
  assign n16629 = ( ~n16624 & n16625 ) | ( ~n16624 & n16628 ) | ( n16625 & n16628 ) ;
  assign n16630 = ~n16623 & n16629 ;
  assign n16631 = ( ~n1139 & n5859 ) | ( ~n1139 & n9501 ) | ( n5859 & n9501 ) ;
  assign n16632 = n9097 ^ n4808 ^ n441 ;
  assign n16633 = n16632 ^ n10077 ^ 1'b0 ;
  assign n16635 = n1847 & n6611 ;
  assign n16636 = ~n5317 & n16635 ;
  assign n16634 = n7944 ^ n2708 ^ 1'b0 ;
  assign n16637 = n16636 ^ n16634 ^ 1'b0 ;
  assign n16638 = ~n16633 & n16637 ;
  assign n16639 = n9093 ^ n8264 ^ n601 ;
  assign n16640 = n8971 ^ n7508 ^ 1'b0 ;
  assign n16641 = n16639 & ~n16640 ;
  assign n16642 = n2719 & n12710 ;
  assign n16643 = n13818 ^ n2896 ^ 1'b0 ;
  assign n16644 = n16176 | n16643 ;
  assign n16645 = n13462 ^ n4879 ^ 1'b0 ;
  assign n16646 = n7351 | n16645 ;
  assign n16647 = ~n8720 & n11649 ;
  assign n16648 = n16647 ^ n16070 ^ n8423 ;
  assign n16651 = ( n1804 & n3254 ) | ( n1804 & n6174 ) | ( n3254 & n6174 ) ;
  assign n16649 = ~n2232 & n16477 ;
  assign n16650 = n16649 ^ n10117 ^ 1'b0 ;
  assign n16652 = n16651 ^ n16650 ^ n3302 ;
  assign n16653 = n16652 ^ n9559 ^ 1'b0 ;
  assign n16654 = ( n3937 & n9476 ) | ( n3937 & ~n16653 ) | ( n9476 & ~n16653 ) ;
  assign n16655 = n15827 ^ n6514 ^ 1'b0 ;
  assign n16656 = n3289 & n16655 ;
  assign n16657 = n16656 ^ n12740 ^ 1'b0 ;
  assign n16658 = n11228 ^ n8378 ^ 1'b0 ;
  assign n16659 = n5130 & n16658 ;
  assign n16660 = n11105 ^ n7085 ^ 1'b0 ;
  assign n16661 = ~n3915 & n16660 ;
  assign n16662 = ~n16659 & n16661 ;
  assign n16667 = n533 & ~n5656 ;
  assign n16666 = n5010 & n7584 ;
  assign n16668 = n16667 ^ n16666 ^ 1'b0 ;
  assign n16663 = n6176 & n6805 ;
  assign n16664 = n16663 ^ n581 ^ 1'b0 ;
  assign n16665 = ( ~n1772 & n2374 ) | ( ~n1772 & n16664 ) | ( n2374 & n16664 ) ;
  assign n16669 = n16668 ^ n16665 ^ 1'b0 ;
  assign n16670 = ~n7782 & n9729 ;
  assign n16671 = n16670 ^ n10130 ^ 1'b0 ;
  assign n16672 = n4806 ^ x254 ^ 1'b0 ;
  assign n16673 = ( ~n1139 & n1356 ) | ( ~n1139 & n2246 ) | ( n1356 & n2246 ) ;
  assign n16674 = n13164 & ~n16673 ;
  assign n16675 = ~n16672 & n16674 ;
  assign n16676 = ~n16631 & n16675 ;
  assign n16677 = n16671 & ~n16676 ;
  assign n16678 = ~n3920 & n16677 ;
  assign n16679 = n12417 & ~n16678 ;
  assign n16680 = n463 & n16679 ;
  assign n16681 = n3438 ^ n1861 ^ 1'b0 ;
  assign n16682 = ( n935 & ~n5372 ) | ( n935 & n8531 ) | ( ~n5372 & n8531 ) ;
  assign n16683 = ~n1099 & n7897 ;
  assign n16684 = n16683 ^ n6607 ^ 1'b0 ;
  assign n16685 = n7149 & n16684 ;
  assign n16686 = n12251 & n16685 ;
  assign n16687 = n9111 ^ n8901 ^ 1'b0 ;
  assign n16688 = n2811 | n2846 ;
  assign n16689 = n4026 | n16688 ;
  assign n16690 = n16107 | n16689 ;
  assign n16691 = n5616 & ~n6119 ;
  assign n16692 = n7306 ^ n6111 ^ 1'b0 ;
  assign n16693 = n16691 & ~n16692 ;
  assign n16694 = n9351 ^ n7293 ^ 1'b0 ;
  assign n16695 = n16659 ^ n13386 ^ n11077 ;
  assign n16696 = n2029 & n12816 ;
  assign n16697 = ~n12131 & n16696 ;
  assign n16698 = ~n9752 & n11720 ;
  assign n16699 = n5550 & n6569 ;
  assign n16700 = n16699 ^ x92 ^ 1'b0 ;
  assign n16701 = ~n12039 & n12766 ;
  assign n16702 = ~n1690 & n15230 ;
  assign n16703 = n16702 ^ n9385 ^ 1'b0 ;
  assign n16704 = ( n8865 & n10296 ) | ( n8865 & n13989 ) | ( n10296 & n13989 ) ;
  assign n16705 = n16704 ^ n9885 ^ n6673 ;
  assign n16706 = n16705 ^ n10595 ^ n5060 ;
  assign n16707 = n16706 ^ n2057 ^ 1'b0 ;
  assign n16708 = n13538 | n16707 ;
  assign n16709 = n2991 & n4550 ;
  assign n16710 = ( n445 & n9968 ) | ( n445 & ~n15948 ) | ( n9968 & ~n15948 ) ;
  assign n16711 = n12373 ^ n3328 ^ 1'b0 ;
  assign n16712 = n16711 ^ n4471 ^ 1'b0 ;
  assign n16713 = ( ~n1967 & n8020 ) | ( ~n1967 & n16712 ) | ( n8020 & n16712 ) ;
  assign n16714 = n11829 ^ n5970 ^ 1'b0 ;
  assign n16715 = ~n2614 & n9190 ;
  assign n16716 = n4308 & n4312 ;
  assign n16717 = n843 & n1590 ;
  assign n16718 = n16717 ^ n12460 ^ 1'b0 ;
  assign n16719 = ( ~n7839 & n14769 ) | ( ~n7839 & n15303 ) | ( n14769 & n15303 ) ;
  assign n16720 = n16718 & n16719 ;
  assign n16721 = ~n16716 & n16720 ;
  assign n16722 = n16721 ^ n3572 ^ 1'b0 ;
  assign n16723 = ( n407 & n4604 ) | ( n407 & ~n10336 ) | ( n4604 & ~n10336 ) ;
  assign n16724 = n3251 | n7783 ;
  assign n16725 = n16723 | n16724 ;
  assign n16726 = n9023 & n16725 ;
  assign n16727 = n16726 ^ n296 ^ 1'b0 ;
  assign n16728 = n791 & n3728 ;
  assign n16729 = n16728 ^ n4394 ^ 1'b0 ;
  assign n16730 = n11512 | n16729 ;
  assign n16731 = ~n7611 & n10617 ;
  assign n16732 = n6077 | n8435 ;
  assign n16733 = ~n5175 & n16567 ;
  assign n16734 = x10 & ~n16733 ;
  assign n16735 = n11823 & n12321 ;
  assign n16736 = n13799 & n16735 ;
  assign n16737 = ( n360 & n989 ) | ( n360 & ~n13055 ) | ( n989 & ~n13055 ) ;
  assign n16738 = n8300 ^ n7633 ^ n527 ;
  assign n16739 = n16738 ^ n14326 ^ 1'b0 ;
  assign n16740 = n8197 ^ n6047 ^ 1'b0 ;
  assign n16741 = ~n3383 & n16740 ;
  assign n16742 = ~n1763 & n13630 ;
  assign n16743 = n16742 ^ n10464 ^ 1'b0 ;
  assign n16744 = n4097 & n15463 ;
  assign n16745 = n16744 ^ n8017 ^ 1'b0 ;
  assign n16746 = ~n5772 & n15653 ;
  assign n16747 = n16746 ^ n13873 ^ 1'b0 ;
  assign n16748 = n972 | n1697 ;
  assign n16749 = n1924 & ~n16748 ;
  assign n16750 = n16749 ^ n2937 ^ 1'b0 ;
  assign n16751 = n16750 ^ n11959 ^ n9428 ;
  assign n16752 = n5630 & n5653 ;
  assign n16756 = n10153 & ~n10661 ;
  assign n16753 = n3386 ^ x121 ^ 1'b0 ;
  assign n16754 = n16753 ^ n12987 ^ n2932 ;
  assign n16755 = ~n2127 & n16754 ;
  assign n16757 = n16756 ^ n16755 ^ 1'b0 ;
  assign n16758 = n16757 ^ n12722 ^ 1'b0 ;
  assign n16759 = n14839 | n16758 ;
  assign n16760 = n16759 ^ n13056 ^ 1'b0 ;
  assign n16761 = n6128 ^ n2203 ^ 1'b0 ;
  assign n16762 = n16761 ^ n4769 ^ 1'b0 ;
  assign n16763 = n4193 | n16762 ;
  assign n16764 = n875 | n8677 ;
  assign n16765 = n14907 ^ n13704 ^ n9642 ;
  assign n16766 = n15620 ^ n14316 ^ n9392 ;
  assign n16767 = n8721 ^ n3135 ^ 1'b0 ;
  assign n16768 = n16767 ^ n10846 ^ 1'b0 ;
  assign n16769 = n8281 | n16768 ;
  assign n16770 = n4934 & ~n16769 ;
  assign n16771 = n1827 & n2291 ;
  assign n16772 = ~n353 & n16771 ;
  assign n16773 = n3071 | n16772 ;
  assign n16774 = n2649 | n7225 ;
  assign n16775 = n16774 ^ n13590 ^ 1'b0 ;
  assign n16776 = n8725 ^ n6898 ^ 1'b0 ;
  assign n16777 = ( ~n2144 & n3388 ) | ( ~n2144 & n16776 ) | ( n3388 & n16776 ) ;
  assign n16778 = ~n2098 & n5414 ;
  assign n16779 = n16778 ^ n3459 ^ 1'b0 ;
  assign n16780 = n12023 | n16779 ;
  assign n16781 = n16780 ^ n2547 ^ 1'b0 ;
  assign n16782 = n950 & n10122 ;
  assign n16783 = ~n16781 & n16782 ;
  assign n16784 = ( ~n3749 & n14570 ) | ( ~n3749 & n16783 ) | ( n14570 & n16783 ) ;
  assign n16785 = n1910 & n16280 ;
  assign n16791 = n5117 & n9230 ;
  assign n16792 = n6313 & n16791 ;
  assign n16793 = n16792 ^ n4966 ^ 1'b0 ;
  assign n16786 = x20 & n1095 ;
  assign n16787 = n16786 ^ n471 ^ 1'b0 ;
  assign n16788 = n10682 | n16787 ;
  assign n16789 = ~n15369 & n16788 ;
  assign n16790 = ~n3175 & n16789 ;
  assign n16794 = n16793 ^ n16790 ^ 1'b0 ;
  assign n16795 = n6155 & n13436 ;
  assign n16796 = n3604 & n16795 ;
  assign n16797 = ~n1521 & n9181 ;
  assign n16798 = ~n1961 & n16797 ;
  assign n16799 = n16798 ^ n3450 ^ 1'b0 ;
  assign n16800 = n16796 | n16799 ;
  assign n16801 = n16569 ^ n4501 ^ 1'b0 ;
  assign n16802 = n16800 | n16801 ;
  assign n16803 = ~n2187 & n16802 ;
  assign n16804 = n16803 ^ n12547 ^ 1'b0 ;
  assign n16805 = n4953 | n16804 ;
  assign n16806 = x165 & n8878 ;
  assign n16807 = n9096 & n16806 ;
  assign n16808 = n1473 | n16807 ;
  assign n16809 = n6929 & n16808 ;
  assign n16810 = n11567 & ~n13780 ;
  assign n16811 = ~n3852 & n16810 ;
  assign n16812 = n9154 ^ n8985 ^ 1'b0 ;
  assign n16813 = n16812 ^ n9065 ^ 1'b0 ;
  assign n16814 = n16811 & ~n16813 ;
  assign n16815 = n5666 ^ n3588 ^ 1'b0 ;
  assign n16816 = n2913 & n16815 ;
  assign n16817 = n3228 & n13985 ;
  assign n16818 = ~n16816 & n16817 ;
  assign n16819 = x154 & ~n11621 ;
  assign n16820 = n16819 ^ n4768 ^ 1'b0 ;
  assign n16821 = ~n1766 & n2202 ;
  assign n16822 = ~n4021 & n16821 ;
  assign n16823 = ~n5052 & n16822 ;
  assign n16824 = n16820 & ~n16823 ;
  assign n16825 = n1902 | n7963 ;
  assign n16826 = n14154 & n16825 ;
  assign n16827 = n4800 & n6509 ;
  assign n16828 = n12677 & n16827 ;
  assign n16829 = n11893 & n16828 ;
  assign n16831 = n5164 ^ n2846 ^ 1'b0 ;
  assign n16832 = ( ~n6537 & n9175 ) | ( ~n6537 & n16831 ) | ( n9175 & n16831 ) ;
  assign n16830 = n6470 & ~n7976 ;
  assign n16833 = n16832 ^ n16830 ^ n14035 ;
  assign n16834 = ~n2728 & n3729 ;
  assign n16835 = n15119 ^ n11385 ^ 1'b0 ;
  assign n16836 = n16834 & ~n16835 ;
  assign n16837 = ~n10650 & n16836 ;
  assign n16838 = n16472 & n16837 ;
  assign n16839 = ( n3782 & n10223 ) | ( n3782 & ~n10236 ) | ( n10223 & ~n10236 ) ;
  assign n16842 = ~n11265 & n14769 ;
  assign n16843 = n16842 ^ n10070 ^ 1'b0 ;
  assign n16844 = n9266 | n16843 ;
  assign n16845 = n1404 | n16844 ;
  assign n16840 = n6001 | n7932 ;
  assign n16841 = n3163 & ~n16840 ;
  assign n16846 = n16845 ^ n16841 ^ 1'b0 ;
  assign n16847 = n3833 & ~n15018 ;
  assign n16849 = n2497 ^ x183 ^ 1'b0 ;
  assign n16850 = n3907 & n16849 ;
  assign n16848 = n3899 ^ n2105 ^ 1'b0 ;
  assign n16851 = n16850 ^ n16848 ^ 1'b0 ;
  assign n16853 = n7191 ^ n1004 ^ 1'b0 ;
  assign n16854 = n5381 | n16853 ;
  assign n16852 = ~n2106 & n12642 ;
  assign n16855 = n16854 ^ n16852 ^ 1'b0 ;
  assign n16856 = n10589 ^ n7658 ^ 1'b0 ;
  assign n16857 = n16856 ^ n11719 ^ n4278 ;
  assign n16858 = n5083 | n8569 ;
  assign n16860 = n8105 ^ n7554 ^ n6636 ;
  assign n16861 = n16860 ^ n12391 ^ n10054 ;
  assign n16859 = n4807 ^ n4467 ^ n647 ;
  assign n16862 = n16861 ^ n16859 ^ n9658 ;
  assign n16863 = n6912 | n16862 ;
  assign n16864 = n520 | n16863 ;
  assign n16865 = ~n2376 & n3176 ;
  assign n16866 = ~n7758 & n8820 ;
  assign n16867 = ~n16865 & n16866 ;
  assign n16868 = ( ~n1498 & n4144 ) | ( ~n1498 & n5412 ) | ( n4144 & n5412 ) ;
  assign n16869 = n3982 & n16868 ;
  assign n16870 = ~n12717 & n16869 ;
  assign n16871 = n6927 & ~n14293 ;
  assign n16872 = n13772 ^ n1298 ^ n429 ;
  assign n16876 = ~n4547 & n5487 ;
  assign n16877 = n16876 ^ n4758 ^ 1'b0 ;
  assign n16873 = n1569 & n2358 ;
  assign n16874 = n16873 ^ n7349 ^ 1'b0 ;
  assign n16875 = n8350 & ~n16874 ;
  assign n16878 = n16877 ^ n16875 ^ 1'b0 ;
  assign n16879 = n2743 | n12020 ;
  assign n16880 = n16879 ^ n4064 ^ 1'b0 ;
  assign n16885 = ( n1663 & n3300 ) | ( n1663 & ~n4807 ) | ( n3300 & ~n4807 ) ;
  assign n16883 = n1824 | n13349 ;
  assign n16882 = n2046 & ~n5739 ;
  assign n16884 = n16883 ^ n16882 ^ 1'b0 ;
  assign n16886 = n16885 ^ n16884 ^ n11790 ;
  assign n16881 = ~n752 & n7250 ;
  assign n16887 = n16886 ^ n16881 ^ 1'b0 ;
  assign n16888 = n3779 ^ n1929 ^ 1'b0 ;
  assign n16889 = ~n8503 & n16888 ;
  assign n16890 = n372 & n16889 ;
  assign n16891 = n16890 ^ n6816 ^ 1'b0 ;
  assign n16892 = x212 & ~n1085 ;
  assign n16893 = ~n13621 & n16892 ;
  assign n16894 = n4010 & ~n8402 ;
  assign n16895 = ~n271 & n16894 ;
  assign n16896 = ( ~n1500 & n16893 ) | ( ~n1500 & n16895 ) | ( n16893 & n16895 ) ;
  assign n16897 = x222 & n2647 ;
  assign n16898 = n13081 & ~n16897 ;
  assign n16899 = n16898 ^ n1978 ^ 1'b0 ;
  assign n16900 = n8614 | n12174 ;
  assign n16901 = n16900 ^ n11808 ^ n2047 ;
  assign n16902 = ~n2696 & n8255 ;
  assign n16903 = n14828 ^ n9693 ^ 1'b0 ;
  assign n16904 = n16902 & ~n16903 ;
  assign n16905 = n7253 ^ n7016 ^ 1'b0 ;
  assign n16906 = ~n14728 & n16905 ;
  assign n16907 = n16906 ^ n9482 ^ 1'b0 ;
  assign n16908 = ~n6496 & n10837 ;
  assign n16909 = x179 & n16908 ;
  assign n16910 = n16909 ^ n843 ^ 1'b0 ;
  assign n16911 = n16910 ^ n3776 ^ n2910 ;
  assign n16912 = n12157 | n16911 ;
  assign n16913 = n3885 | n13555 ;
  assign n16914 = n8655 & n10497 ;
  assign n16915 = n16914 ^ n4931 ^ 1'b0 ;
  assign n16916 = n8752 & n16915 ;
  assign n16917 = n2114 & n11628 ;
  assign n16918 = n9548 ^ n6573 ^ 1'b0 ;
  assign n16919 = n15390 & ~n16918 ;
  assign n16920 = n13316 ^ n8836 ^ 1'b0 ;
  assign n16921 = ~n4167 & n9676 ;
  assign n16922 = n16921 ^ n286 ^ 1'b0 ;
  assign n16923 = n16922 ^ n14298 ^ n3191 ;
  assign n16924 = ( n4238 & n7323 ) | ( n4238 & n16650 ) | ( n7323 & n16650 ) ;
  assign n16925 = n14324 | n16133 ;
  assign n16927 = n8578 | n13738 ;
  assign n16926 = n5217 & ~n9925 ;
  assign n16928 = n16927 ^ n16926 ^ 1'b0 ;
  assign n16929 = n12304 ^ n4628 ^ n3232 ;
  assign n16930 = ~n1800 & n2048 ;
  assign n16931 = ~n1119 & n16930 ;
  assign n16932 = n16931 ^ n7007 ^ 1'b0 ;
  assign n16933 = n11692 ^ n10363 ^ n1709 ;
  assign n16934 = n14998 & n16933 ;
  assign n16935 = n10879 ^ n4524 ^ 1'b0 ;
  assign n16936 = n15025 ^ n14158 ^ n11134 ;
  assign n16937 = n2898 & n8084 ;
  assign n16941 = n8167 ^ n3345 ^ 1'b0 ;
  assign n16942 = n9178 & n16941 ;
  assign n16938 = n3392 & n5020 ;
  assign n16939 = ~n5988 & n16938 ;
  assign n16940 = n7957 & ~n16939 ;
  assign n16943 = n16942 ^ n16940 ^ 1'b0 ;
  assign n16944 = n7435 | n9457 ;
  assign n16945 = n9752 ^ n2860 ^ 1'b0 ;
  assign n16946 = ~n2105 & n16945 ;
  assign n16947 = n1233 & n3501 ;
  assign n16948 = ( n1851 & ~n1868 ) | ( n1851 & n3166 ) | ( ~n1868 & n3166 ) ;
  assign n16949 = n11408 ^ n1813 ^ 1'b0 ;
  assign n16950 = n16948 & n16949 ;
  assign n16951 = n449 & n16729 ;
  assign n16952 = n16951 ^ n7627 ^ 1'b0 ;
  assign n16953 = n8621 & ~n16952 ;
  assign n16954 = n8250 ^ n4658 ^ 1'b0 ;
  assign n16955 = ( n9047 & ~n15555 ) | ( n9047 & n16954 ) | ( ~n15555 & n16954 ) ;
  assign n16956 = n10709 ^ n2778 ^ 1'b0 ;
  assign n16957 = n8632 & ~n16956 ;
  assign n16958 = n8778 ^ n4050 ^ 1'b0 ;
  assign n16959 = ( n9244 & ~n15260 ) | ( n9244 & n16958 ) | ( ~n15260 & n16958 ) ;
  assign n16960 = n4857 ^ n617 ^ 1'b0 ;
  assign n16961 = x120 & ~n16960 ;
  assign n16962 = n16961 ^ n7547 ^ 1'b0 ;
  assign n16963 = n7105 & ~n16962 ;
  assign n16964 = n11258 & n16963 ;
  assign n16965 = n2457 & ~n10601 ;
  assign n16966 = n1160 & n1624 ;
  assign n16967 = ( x68 & n12723 ) | ( x68 & n16626 ) | ( n12723 & n16626 ) ;
  assign n16968 = n936 | n12890 ;
  assign n16969 = n2713 ^ n1440 ^ 1'b0 ;
  assign n16970 = n8782 & ~n16969 ;
  assign n16971 = ( x224 & ~n1581 ) | ( x224 & n16970 ) | ( ~n1581 & n16970 ) ;
  assign n16972 = ~n16968 & n16971 ;
  assign n16973 = n16967 & ~n16972 ;
  assign n16974 = n16973 ^ n2225 ^ 1'b0 ;
  assign n16975 = n11885 ^ n5507 ^ 1'b0 ;
  assign n16976 = n6642 | n10535 ;
  assign n16977 = n933 & ~n16976 ;
  assign n16978 = ( n7649 & n13785 ) | ( n7649 & n16977 ) | ( n13785 & n16977 ) ;
  assign n16979 = n14354 ^ n2728 ^ 1'b0 ;
  assign n16980 = ~n16978 & n16979 ;
  assign n16984 = n1974 | n6851 ;
  assign n16985 = n16984 ^ n1066 ^ 1'b0 ;
  assign n16981 = n5594 ^ x15 ^ 1'b0 ;
  assign n16982 = n6341 | n16981 ;
  assign n16983 = n16982 ^ n10716 ^ 1'b0 ;
  assign n16986 = n16985 ^ n16983 ^ n11726 ;
  assign n16987 = n16986 ^ n8811 ^ n1961 ;
  assign n16988 = n12357 & n15334 ;
  assign n16989 = ~n7658 & n16988 ;
  assign n16990 = ( ~n911 & n4628 ) | ( ~n911 & n6391 ) | ( n4628 & n6391 ) ;
  assign n16991 = n6563 | n8453 ;
  assign n16992 = n16991 ^ n1034 ^ 1'b0 ;
  assign n16993 = ~n7348 & n16992 ;
  assign n16994 = n6451 & n16993 ;
  assign n16995 = n12002 & ~n16994 ;
  assign n16996 = n16990 & n16995 ;
  assign n16997 = n16996 ^ n12961 ^ 1'b0 ;
  assign n16998 = n8129 | n16997 ;
  assign n16999 = n14310 | n15343 ;
  assign n17000 = n5947 | n11183 ;
  assign n17001 = n11328 ^ n11055 ^ 1'b0 ;
  assign n17004 = ( ~n1042 & n8372 ) | ( ~n1042 & n8949 ) | ( n8372 & n8949 ) ;
  assign n17002 = n13469 ^ n4615 ^ 1'b0 ;
  assign n17003 = ~n7334 & n17002 ;
  assign n17005 = n17004 ^ n17003 ^ n7317 ;
  assign n17006 = ~n2497 & n5372 ;
  assign n17007 = ( n2775 & n5680 ) | ( n2775 & ~n10969 ) | ( n5680 & ~n10969 ) ;
  assign n17008 = n3378 & ~n17007 ;
  assign n17009 = x178 | n9740 ;
  assign n17010 = n11244 ^ n258 ^ 1'b0 ;
  assign n17011 = n17009 & ~n17010 ;
  assign n17012 = ~n10582 & n17011 ;
  assign n17013 = n4229 & n17012 ;
  assign n17014 = n6938 ^ n3286 ^ 1'b0 ;
  assign n17015 = n3434 | n17014 ;
  assign n17016 = n7073 ^ n3460 ^ 1'b0 ;
  assign n17017 = n8474 ^ n4520 ^ x170 ;
  assign n17018 = x74 | n12410 ;
  assign n17019 = n5617 & n17018 ;
  assign n17020 = ~n17017 & n17019 ;
  assign n17021 = n2785 & ~n6569 ;
  assign n17022 = n7351 ^ x170 ^ 1'b0 ;
  assign n17023 = n8446 & ~n10055 ;
  assign n17024 = n579 | n11597 ;
  assign n17025 = n17024 ^ n16215 ^ n3156 ;
  assign n17026 = n4646 ^ n2893 ^ 1'b0 ;
  assign n17027 = n2532 & ~n5650 ;
  assign n17028 = n17027 ^ n7539 ^ 1'b0 ;
  assign n17029 = n3767 & n17028 ;
  assign n17030 = n6214 & n17029 ;
  assign n17031 = n17026 & n17030 ;
  assign n17032 = n1555 & n10275 ;
  assign n17033 = x103 & n2377 ;
  assign n17034 = ~n4112 & n17033 ;
  assign n17035 = x232 & n10590 ;
  assign n17036 = n17034 & n17035 ;
  assign n17037 = n9437 | n17036 ;
  assign n17038 = n17032 | n17037 ;
  assign n17039 = n8277 & ~n17038 ;
  assign n17040 = ~n6424 & n9356 ;
  assign n17041 = x185 & n4271 ;
  assign n17042 = n17041 ^ n3081 ^ 1'b0 ;
  assign n17043 = ( n4426 & ~n12400 ) | ( n4426 & n17042 ) | ( ~n12400 & n17042 ) ;
  assign n17044 = ( ~n9279 & n15717 ) | ( ~n9279 & n17043 ) | ( n15717 & n17043 ) ;
  assign n17045 = n16980 ^ n8677 ^ n5139 ;
  assign n17060 = ( n2499 & n3697 ) | ( n2499 & ~n5474 ) | ( n3697 & ~n5474 ) ;
  assign n17061 = n2585 & ~n7501 ;
  assign n17062 = ~n9857 & n17061 ;
  assign n17063 = ~n17060 & n17062 ;
  assign n17046 = n13495 ^ n3279 ^ 1'b0 ;
  assign n17047 = n8800 & ~n17046 ;
  assign n17048 = n17047 ^ n9808 ^ 1'b0 ;
  assign n17049 = n17048 ^ n4767 ^ 1'b0 ;
  assign n17050 = ~n4613 & n10579 ;
  assign n17051 = n1312 & n17050 ;
  assign n17052 = n1236 & ~n7161 ;
  assign n17053 = n14587 ^ n1353 ^ 1'b0 ;
  assign n17054 = n12479 & ~n17053 ;
  assign n17055 = ~n17052 & n17054 ;
  assign n17056 = n15034 | n17055 ;
  assign n17057 = n17051 & ~n17056 ;
  assign n17058 = n17049 | n17057 ;
  assign n17059 = n15516 & ~n17058 ;
  assign n17064 = n17063 ^ n17059 ^ 1'b0 ;
  assign n17065 = n845 & ~n17064 ;
  assign n17066 = ( n1819 & ~n11219 ) | ( n1819 & n11459 ) | ( ~n11219 & n11459 ) ;
  assign n17067 = n12208 & n17066 ;
  assign n17068 = ~n4870 & n17067 ;
  assign n17069 = n4743 ^ n3551 ^ 1'b0 ;
  assign n17070 = x233 & ~n5074 ;
  assign n17071 = n17069 & n17070 ;
  assign n17072 = ( n14550 & ~n15333 ) | ( n14550 & n17071 ) | ( ~n15333 & n17071 ) ;
  assign n17073 = n1223 | n16667 ;
  assign n17074 = n4016 ^ n3830 ^ 1'b0 ;
  assign n17075 = n12319 ^ n8739 ^ 1'b0 ;
  assign n17076 = ( n7997 & n16831 ) | ( n7997 & n17075 ) | ( n16831 & n17075 ) ;
  assign n17077 = n17074 | n17076 ;
  assign n17078 = n17077 ^ n7822 ^ 1'b0 ;
  assign n17079 = n5304 & ~n17078 ;
  assign n17080 = n17079 ^ n15020 ^ 1'b0 ;
  assign n17081 = n6282 & ~n6605 ;
  assign n17082 = x195 & n698 ;
  assign n17083 = n17082 ^ n3862 ^ 1'b0 ;
  assign n17085 = ( n3450 & ~n5065 ) | ( n3450 & n7974 ) | ( ~n5065 & n7974 ) ;
  assign n17084 = ( n3697 & n7301 ) | ( n3697 & ~n7317 ) | ( n7301 & ~n7317 ) ;
  assign n17086 = n17085 ^ n17084 ^ 1'b0 ;
  assign n17087 = n8930 | n17086 ;
  assign n17088 = n17087 ^ n3632 ^ 1'b0 ;
  assign n17089 = n1838 & n17088 ;
  assign n17090 = ~n1024 & n9413 ;
  assign n17091 = ~n3817 & n17090 ;
  assign n17093 = n13142 ^ n6853 ^ 1'b0 ;
  assign n17094 = x233 & ~n17093 ;
  assign n17095 = n2916 & ~n11633 ;
  assign n17100 = ~n1323 & n14852 ;
  assign n17101 = n17100 ^ n2968 ^ 1'b0 ;
  assign n17102 = n6683 & ~n17101 ;
  assign n17096 = n1010 & ~n4894 ;
  assign n17097 = n17096 ^ n8841 ^ 1'b0 ;
  assign n17098 = n1126 | n17097 ;
  assign n17099 = n17098 ^ n11304 ^ 1'b0 ;
  assign n17103 = n17102 ^ n17099 ^ 1'b0 ;
  assign n17104 = n17095 & n17103 ;
  assign n17105 = n17104 ^ n3899 ^ 1'b0 ;
  assign n17106 = n17094 & n17105 ;
  assign n17092 = n1784 | n16861 ;
  assign n17107 = n17106 ^ n17092 ^ 1'b0 ;
  assign n17108 = n5791 & n10441 ;
  assign n17109 = ~n6811 & n17108 ;
  assign n17110 = ( n512 & ~n1291 ) | ( n512 & n17109 ) | ( ~n1291 & n17109 ) ;
  assign n17111 = n2547 | n6488 ;
  assign n17112 = n4721 | n17111 ;
  assign n17113 = n8602 & ~n10879 ;
  assign n17114 = ( n4137 & n10720 ) | ( n4137 & n17113 ) | ( n10720 & n17113 ) ;
  assign n17115 = n12514 & n17114 ;
  assign n17116 = n6314 | n6370 ;
  assign n17117 = n1281 & ~n17116 ;
  assign n17118 = ( n1840 & n3439 ) | ( n1840 & n9561 ) | ( n3439 & n9561 ) ;
  assign n17128 = x85 & ~n4052 ;
  assign n17127 = n16861 ^ n4354 ^ 1'b0 ;
  assign n17129 = n17128 ^ n17127 ^ 1'b0 ;
  assign n17130 = n17129 ^ n10095 ^ 1'b0 ;
  assign n17131 = n7225 & ~n17130 ;
  assign n17119 = n4015 ^ n3904 ^ 1'b0 ;
  assign n17120 = x209 & n17119 ;
  assign n17121 = n17120 ^ n15041 ^ 1'b0 ;
  assign n17122 = ~n4405 & n17121 ;
  assign n17123 = n15378 ^ n7338 ^ 1'b0 ;
  assign n17124 = ( n2866 & ~n6384 ) | ( n2866 & n17123 ) | ( ~n6384 & n17123 ) ;
  assign n17125 = n17124 ^ n12019 ^ n9610 ;
  assign n17126 = n17122 & n17125 ;
  assign n17132 = n17131 ^ n17126 ^ 1'b0 ;
  assign n17133 = n8864 ^ n4573 ^ n1228 ;
  assign n17134 = n7160 & ~n9847 ;
  assign n17135 = n3093 & n17134 ;
  assign n17136 = n11939 ^ n2253 ^ 1'b0 ;
  assign n17137 = x71 & n5523 ;
  assign n17138 = n6704 ^ n5116 ^ 1'b0 ;
  assign n17139 = n3464 & ~n17138 ;
  assign n17142 = n4724 | n13127 ;
  assign n17143 = ~n9618 & n17142 ;
  assign n17140 = n7752 ^ n1885 ^ x201 ;
  assign n17141 = n16318 & ~n17140 ;
  assign n17144 = n17143 ^ n17141 ^ 1'b0 ;
  assign n17150 = n2518 & n5354 ;
  assign n17151 = ~n16235 & n17150 ;
  assign n17145 = x94 & n1315 ;
  assign n17146 = n17145 ^ n4300 ^ 1'b0 ;
  assign n17147 = n3126 & ~n17146 ;
  assign n17148 = n2652 & n17147 ;
  assign n17149 = n9181 & ~n17148 ;
  assign n17152 = n17151 ^ n17149 ^ 1'b0 ;
  assign n17153 = ~n538 & n5690 ;
  assign n17154 = n1297 | n3646 ;
  assign n17155 = n17154 ^ n12863 ^ 1'b0 ;
  assign n17156 = n9835 ^ n2789 ^ 1'b0 ;
  assign n17158 = n1821 | n2190 ;
  assign n17159 = ~n9268 & n9518 ;
  assign n17160 = ~n4117 & n17159 ;
  assign n17161 = n17158 | n17160 ;
  assign n17157 = n16885 ^ n12083 ^ 1'b0 ;
  assign n17162 = n17161 ^ n17157 ^ 1'b0 ;
  assign n17163 = n1395 & n5477 ;
  assign n17164 = n413 & ~n6353 ;
  assign n17165 = n17164 ^ n14217 ^ 1'b0 ;
  assign n17166 = n17163 & n17165 ;
  assign n17167 = n15712 ^ n2692 ^ 1'b0 ;
  assign n17168 = n4840 ^ n3714 ^ 1'b0 ;
  assign n17169 = n12353 ^ n5355 ^ 1'b0 ;
  assign n17170 = n6653 ^ n3926 ^ n3305 ;
  assign n17171 = n286 & n1577 ;
  assign n17172 = n10012 & ~n17171 ;
  assign n17173 = n17170 & ~n17172 ;
  assign n17174 = n17173 ^ n3369 ^ 1'b0 ;
  assign n17175 = n17174 ^ n13764 ^ 1'b0 ;
  assign n17176 = n2322 & n5462 ;
  assign n17177 = ~n6271 & n16571 ;
  assign n17178 = n17177 ^ n13342 ^ 1'b0 ;
  assign n17179 = n8632 & n15996 ;
  assign n17180 = n17104 ^ n15571 ^ n5531 ;
  assign n17181 = n11918 | n17180 ;
  assign n17182 = ( x72 & n1731 ) | ( x72 & ~n8241 ) | ( n1731 & ~n8241 ) ;
  assign n17183 = n17182 ^ n3056 ^ 1'b0 ;
  assign n17184 = n11369 & n17183 ;
  assign n17185 = n17184 ^ n15837 ^ n11599 ;
  assign n17186 = ( ~n3443 & n15074 ) | ( ~n3443 & n15818 ) | ( n15074 & n15818 ) ;
  assign n17187 = n6205 & n8457 ;
  assign n17188 = n17187 ^ n4585 ^ 1'b0 ;
  assign n17189 = n15633 ^ n9209 ^ 1'b0 ;
  assign n17190 = ~n16294 & n17189 ;
  assign n17191 = n4235 | n8402 ;
  assign n17192 = n6807 & ~n14861 ;
  assign n17193 = ~n7508 & n14212 ;
  assign n17194 = ~n17192 & n17193 ;
  assign n17195 = n3660 & ~n17194 ;
  assign n17196 = n17195 ^ n16599 ^ 1'b0 ;
  assign n17197 = n14833 ^ n13366 ^ 1'b0 ;
  assign n17198 = n991 | n17197 ;
  assign n17199 = n17198 ^ n11030 ^ 1'b0 ;
  assign n17200 = ~n8993 & n17199 ;
  assign n17201 = ~n13011 & n17200 ;
  assign n17202 = ~n7790 & n17201 ;
  assign n17203 = ~n12737 & n17202 ;
  assign n17204 = n728 | n4808 ;
  assign n17205 = n14907 & ~n17204 ;
  assign n17206 = n17205 ^ n9688 ^ 1'b0 ;
  assign n17207 = n7674 ^ n5090 ^ 1'b0 ;
  assign n17208 = n14680 ^ n6585 ^ 1'b0 ;
  assign n17209 = n6574 | n17208 ;
  assign n17210 = n14329 & ~n17209 ;
  assign n17211 = n15937 ^ n5321 ^ 1'b0 ;
  assign n17212 = n13920 & ~n15260 ;
  assign n17213 = n4560 & n17212 ;
  assign n17214 = n543 & ~n6818 ;
  assign n17215 = ~n1694 & n2327 ;
  assign n17216 = n17215 ^ n9618 ^ 1'b0 ;
  assign n17217 = n17216 ^ n7203 ^ 1'b0 ;
  assign n17218 = ~n7806 & n17217 ;
  assign n17219 = n6123 ^ n3899 ^ n2002 ;
  assign n17220 = n12126 & ~n17219 ;
  assign n17221 = n14719 & n17220 ;
  assign n17222 = n10325 ^ n6193 ^ 1'b0 ;
  assign n17223 = n2374 | n17222 ;
  assign n17224 = n17223 ^ n11291 ^ 1'b0 ;
  assign n17225 = ( n3714 & n11823 ) | ( n3714 & n12189 ) | ( n11823 & n12189 ) ;
  assign n17226 = n1683 & ~n17225 ;
  assign n17227 = x120 & n14665 ;
  assign n17228 = n1382 & n17227 ;
  assign n17229 = ~n5975 & n6645 ;
  assign n17230 = n1767 | n17229 ;
  assign n17231 = n5356 & ~n17230 ;
  assign n17232 = n6736 | n17231 ;
  assign n17233 = ( n5877 & ~n6676 ) | ( n5877 & n6700 ) | ( ~n6676 & n6700 ) ;
  assign n17234 = ~n2511 & n17233 ;
  assign n17235 = ~n3487 & n17234 ;
  assign n17236 = n6995 & ~n17235 ;
  assign n17237 = n17236 ^ n16483 ^ 1'b0 ;
  assign n17238 = n6382 ^ n2307 ^ 1'b0 ;
  assign n17239 = n13198 | n17238 ;
  assign n17240 = n14342 & ~n17239 ;
  assign n17241 = n9074 ^ n8300 ^ 1'b0 ;
  assign n17242 = n17241 ^ n13198 ^ 1'b0 ;
  assign n17243 = n14570 ^ n3757 ^ 1'b0 ;
  assign n17244 = n16602 ^ n12101 ^ 1'b0 ;
  assign n17245 = n17243 & ~n17244 ;
  assign n17246 = n3477 & ~n11532 ;
  assign n17247 = ~n12226 & n17246 ;
  assign n17248 = n1813 & n2053 ;
  assign n17249 = n17248 ^ n2493 ^ 1'b0 ;
  assign n17250 = n5052 & n17249 ;
  assign n17251 = n17250 ^ n7930 ^ 1'b0 ;
  assign n17252 = n17247 & n17251 ;
  assign n17253 = n16629 ^ n8880 ^ 1'b0 ;
  assign n17254 = ~n9796 & n17253 ;
  assign n17255 = n15193 ^ n6536 ^ 1'b0 ;
  assign n17256 = n7994 | n17255 ;
  assign n17257 = n17256 ^ n2641 ^ 1'b0 ;
  assign n17258 = n17257 ^ n3993 ^ 1'b0 ;
  assign n17259 = n5093 ^ n2598 ^ 1'b0 ;
  assign n17260 = ( x114 & ~n13069 ) | ( x114 & n17259 ) | ( ~n13069 & n17259 ) ;
  assign n17261 = ~n1201 & n15147 ;
  assign n17263 = n5177 | n14276 ;
  assign n17262 = n7021 | n9751 ;
  assign n17264 = n17263 ^ n17262 ^ 1'b0 ;
  assign n17265 = n12087 ^ n4396 ^ 1'b0 ;
  assign n17266 = n11819 & ~n17265 ;
  assign n17267 = ( n292 & n513 ) | ( n292 & ~n17266 ) | ( n513 & ~n17266 ) ;
  assign n17268 = ( n7764 & ~n17264 ) | ( n7764 & n17267 ) | ( ~n17264 & n17267 ) ;
  assign n17269 = n17268 ^ n8539 ^ 1'b0 ;
  assign n17270 = n4064 | n17269 ;
  assign n17271 = n1374 & ~n2017 ;
  assign n17272 = n17271 ^ n1346 ^ 1'b0 ;
  assign n17273 = n3889 & ~n16002 ;
  assign n17274 = n5509 | n6805 ;
  assign n17275 = n1200 | n17274 ;
  assign n17276 = n10709 ^ n9115 ^ n7580 ;
  assign n17277 = n627 & ~n17276 ;
  assign n17278 = n787 | n1943 ;
  assign n17279 = n17278 ^ n12899 ^ 1'b0 ;
  assign n17280 = n15629 ^ n14120 ^ 1'b0 ;
  assign n17284 = n1633 & n1694 ;
  assign n17283 = n1222 & ~n7431 ;
  assign n17281 = n14911 ^ n4065 ^ 1'b0 ;
  assign n17282 = n17281 ^ n3940 ^ 1'b0 ;
  assign n17285 = n17284 ^ n17283 ^ n17282 ;
  assign n17286 = n11163 | n17285 ;
  assign n17287 = n8352 & n17286 ;
  assign n17288 = n2793 ^ n2479 ^ n1421 ;
  assign n17289 = n790 & ~n17288 ;
  assign n17290 = n17289 ^ n5599 ^ 1'b0 ;
  assign n17291 = n9398 ^ n9359 ^ n5694 ;
  assign n17292 = ~n17290 & n17291 ;
  assign n17293 = ~n9531 & n17292 ;
  assign n17296 = n11416 ^ n10272 ^ n3465 ;
  assign n17294 = n7029 ^ n991 ^ 1'b0 ;
  assign n17295 = n3074 & n17294 ;
  assign n17297 = n17296 ^ n17295 ^ n8161 ;
  assign n17298 = ~n17293 & n17297 ;
  assign n17299 = n12894 ^ n2621 ^ 1'b0 ;
  assign n17300 = n13435 & ~n17299 ;
  assign n17304 = n4012 ^ n2971 ^ 1'b0 ;
  assign n17305 = n3606 & n17304 ;
  assign n17306 = ~x125 & n17305 ;
  assign n17301 = n1374 & n5420 ;
  assign n17302 = n17301 ^ n5395 ^ 1'b0 ;
  assign n17303 = n17302 ^ n3695 ^ 1'b0 ;
  assign n17307 = n17306 ^ n17303 ^ n2180 ;
  assign n17308 = n1926 ^ n1258 ^ n836 ;
  assign n17309 = n4907 & ~n17308 ;
  assign n17310 = n17309 ^ n4611 ^ 1'b0 ;
  assign n17311 = n4007 & ~n17310 ;
  assign n17312 = n8643 | n11178 ;
  assign n17313 = n5063 & ~n17312 ;
  assign n17314 = n11351 & n17313 ;
  assign n17315 = n8408 | n11050 ;
  assign n17316 = ( ~n5888 & n16289 ) | ( ~n5888 & n17315 ) | ( n16289 & n17315 ) ;
  assign n17317 = n3292 & n9638 ;
  assign n17318 = ~n3103 & n17317 ;
  assign n17319 = n5711 ^ n3583 ^ 1'b0 ;
  assign n17320 = ~n17318 & n17319 ;
  assign n17321 = n2066 & n17320 ;
  assign n17322 = n2192 & n17321 ;
  assign n17323 = ~n15390 & n15990 ;
  assign n17324 = n17323 ^ n2199 ^ 1'b0 ;
  assign n17325 = n4584 ^ n2463 ^ 1'b0 ;
  assign n17326 = ~n1049 & n17325 ;
  assign n17327 = n13510 ^ n4056 ^ 1'b0 ;
  assign n17328 = n17326 & ~n17327 ;
  assign n17329 = n1266 & n13907 ;
  assign n17330 = n13381 ^ n2942 ^ 1'b0 ;
  assign n17331 = n17329 | n17330 ;
  assign n17332 = n17331 ^ n3497 ^ 1'b0 ;
  assign n17333 = n8826 & n17332 ;
  assign n17335 = n10160 ^ n1742 ^ 1'b0 ;
  assign n17336 = n5315 & n17335 ;
  assign n17334 = n2927 & ~n12410 ;
  assign n17337 = n17336 ^ n17334 ^ 1'b0 ;
  assign n17338 = n1563 | n3947 ;
  assign n17339 = n17338 ^ n7977 ^ 1'b0 ;
  assign n17340 = ~n7458 & n17339 ;
  assign n17341 = n8062 ^ n2431 ^ 1'b0 ;
  assign n17342 = ~n2860 & n17341 ;
  assign n17343 = n6382 ^ n3712 ^ 1'b0 ;
  assign n17344 = n17343 ^ n1715 ^ n1026 ;
  assign n17345 = ~n10280 & n17344 ;
  assign n17346 = ~n16839 & n17345 ;
  assign n17347 = n6567 & n10432 ;
  assign n17348 = n17347 ^ n12077 ^ 1'b0 ;
  assign n17349 = n2814 | n6095 ;
  assign n17350 = ( ~n8851 & n16363 ) | ( ~n8851 & n17349 ) | ( n16363 & n17349 ) ;
  assign n17351 = ( n5668 & n7466 ) | ( n5668 & ~n10432 ) | ( n7466 & ~n10432 ) ;
  assign n17352 = n1782 & n10127 ;
  assign n17353 = ( n11226 & n17351 ) | ( n11226 & ~n17352 ) | ( n17351 & ~n17352 ) ;
  assign n17354 = n8369 | n12564 ;
  assign n17355 = ( n8002 & n10042 ) | ( n8002 & ~n12478 ) | ( n10042 & ~n12478 ) ;
  assign n17356 = n3126 & n4308 ;
  assign n17357 = n17356 ^ n3772 ^ x15 ;
  assign n17358 = ~n2516 & n15868 ;
  assign n17359 = n17358 ^ n4328 ^ 1'b0 ;
  assign n17360 = n4833 & n7073 ;
  assign n17361 = ~n15041 & n17360 ;
  assign n17362 = n17361 ^ n9422 ^ n7170 ;
  assign n17363 = n3777 ^ n1194 ^ 1'b0 ;
  assign n17364 = n7338 & ~n17363 ;
  assign n17365 = n4488 | n17198 ;
  assign n17366 = n17364 | n17365 ;
  assign n17367 = n13920 ^ n11853 ^ 1'b0 ;
  assign n17368 = n17366 & n17367 ;
  assign n17369 = n4109 ^ n3289 ^ 1'b0 ;
  assign n17370 = n17369 ^ n1010 ^ 1'b0 ;
  assign n17371 = n17368 & n17370 ;
  assign n17372 = n3511 | n6459 ;
  assign n17373 = n17372 ^ n12108 ^ 1'b0 ;
  assign n17374 = n12080 ^ n4562 ^ n1836 ;
  assign n17375 = n17374 ^ n7788 ^ n6835 ;
  assign n17376 = n17375 ^ n10575 ^ 1'b0 ;
  assign n17377 = n7127 | n17376 ;
  assign n17378 = n14240 ^ n4054 ^ 1'b0 ;
  assign n17379 = n1866 & ~n17378 ;
  assign n17380 = ~n8555 & n17379 ;
  assign n17381 = n12568 & ~n17380 ;
  assign n17382 = n15795 ^ n8577 ^ 1'b0 ;
  assign n17383 = n6866 & n17382 ;
  assign n17384 = n5070 ^ n3055 ^ n562 ;
  assign n17385 = ( ~x55 & n10949 ) | ( ~x55 & n17384 ) | ( n10949 & n17384 ) ;
  assign n17390 = n1444 | n12822 ;
  assign n17391 = n3746 | n17390 ;
  assign n17386 = ~n1346 & n3344 ;
  assign n17387 = n9307 & n17386 ;
  assign n17388 = n17387 ^ n9379 ^ 1'b0 ;
  assign n17389 = n4565 & ~n17388 ;
  assign n17392 = n17391 ^ n17389 ^ 1'b0 ;
  assign n17393 = n15075 & ~n17392 ;
  assign n17397 = n2652 & n3443 ;
  assign n17398 = n17397 ^ n15926 ^ 1'b0 ;
  assign n17394 = n1707 ^ n591 ^ 1'b0 ;
  assign n17395 = n3517 & ~n17394 ;
  assign n17396 = ~n12744 & n17395 ;
  assign n17399 = n17398 ^ n17396 ^ 1'b0 ;
  assign n17400 = n455 ^ n340 ^ 1'b0 ;
  assign n17401 = n9076 | n17400 ;
  assign n17402 = n17401 ^ n3938 ^ 1'b0 ;
  assign n17403 = n17399 | n17402 ;
  assign n17404 = n16184 ^ n9586 ^ 1'b0 ;
  assign n17405 = ~n954 & n17404 ;
  assign n17406 = ( ~n3556 & n7916 ) | ( ~n3556 & n17405 ) | ( n7916 & n17405 ) ;
  assign n17407 = ~n2846 & n3793 ;
  assign n17408 = n7015 ^ n593 ^ 1'b0 ;
  assign n17409 = n17407 & ~n17408 ;
  assign n17410 = n948 | n2423 ;
  assign n17411 = n17410 ^ n1081 ^ 1'b0 ;
  assign n17412 = n17411 ^ n5381 ^ 1'b0 ;
  assign n17413 = n16719 & ~n17412 ;
  assign n17414 = n17357 ^ n6906 ^ 1'b0 ;
  assign n17415 = n8219 & n9404 ;
  assign n17416 = n4160 & n17415 ;
  assign n17417 = n6448 | n17416 ;
  assign n17418 = n1006 & n10935 ;
  assign n17419 = n6907 & n9304 ;
  assign n17420 = n8181 & n17419 ;
  assign n17421 = n2015 | n17420 ;
  assign n17422 = n7849 | n17421 ;
  assign n17423 = n17422 ^ n4284 ^ 1'b0 ;
  assign n17424 = ~n7229 & n17423 ;
  assign n17425 = n13416 ^ n11215 ^ 1'b0 ;
  assign n17426 = n16477 & n17425 ;
  assign n17427 = n17426 ^ n563 ^ 1'b0 ;
  assign n17428 = n5474 & ~n17427 ;
  assign n17429 = n17424 & n17428 ;
  assign n17430 = n17429 ^ n5572 ^ 1'b0 ;
  assign n17431 = n16227 | n17430 ;
  assign n17432 = n16719 | n17431 ;
  assign n17433 = n11167 ^ n8395 ^ 1'b0 ;
  assign n17434 = n6875 & ~n9529 ;
  assign n17435 = n17434 ^ n10391 ^ 1'b0 ;
  assign n17436 = n2127 | n13528 ;
  assign n17437 = n17436 ^ n9976 ^ 1'b0 ;
  assign n17438 = n17437 ^ n11620 ^ 1'b0 ;
  assign n17439 = n17435 & n17438 ;
  assign n17440 = n1703 | n6442 ;
  assign n17441 = n5089 ^ n2120 ^ 1'b0 ;
  assign n17442 = n7536 & ~n17441 ;
  assign n17443 = n9753 | n17442 ;
  assign n17444 = n13458 ^ n1879 ^ 1'b0 ;
  assign n17445 = n5837 | n17274 ;
  assign n17447 = n9317 ^ n1717 ^ 1'b0 ;
  assign n17446 = ( n3332 & n4310 ) | ( n3332 & ~n6899 ) | ( n4310 & ~n6899 ) ;
  assign n17448 = n17447 ^ n17446 ^ n12468 ;
  assign n17449 = n8459 ^ n645 ^ 1'b0 ;
  assign n17450 = ~n8522 & n17449 ;
  assign n17451 = n6142 ^ n1249 ^ 1'b0 ;
  assign n17452 = n17451 ^ n7109 ^ 1'b0 ;
  assign n17453 = ( n2360 & n17450 ) | ( n2360 & n17452 ) | ( n17450 & n17452 ) ;
  assign n17454 = n10258 ^ n10020 ^ 1'b0 ;
  assign n17455 = n5045 ^ n4941 ^ 1'b0 ;
  assign n17456 = ~n8898 & n17455 ;
  assign n17457 = n6361 & n7072 ;
  assign n17458 = n1225 & n17457 ;
  assign n17459 = n17458 ^ n9995 ^ 1'b0 ;
  assign n17461 = n8051 ^ n2626 ^ 1'b0 ;
  assign n17460 = n3310 & n10951 ;
  assign n17462 = n17461 ^ n17460 ^ 1'b0 ;
  assign n17463 = ~n17115 & n17462 ;
  assign n17464 = n8080 & n17463 ;
  assign n17465 = n1334 & n6766 ;
  assign n17466 = n8859 | n11461 ;
  assign n17467 = n17466 ^ n4240 ^ 1'b0 ;
  assign n17468 = n17467 ^ n8941 ^ 1'b0 ;
  assign n17469 = n17468 ^ n2303 ^ 1'b0 ;
  assign n17470 = n7935 | n12353 ;
  assign n17471 = n7552 & ~n17470 ;
  assign n17472 = ~n6408 & n9738 ;
  assign n17473 = n6802 & n17472 ;
  assign n17474 = n3340 & ~n15392 ;
  assign n17475 = n16667 ^ n6122 ^ 1'b0 ;
  assign n17476 = n7336 & ~n9494 ;
  assign n17477 = n2597 | n17476 ;
  assign n17478 = ~n17475 & n17477 ;
  assign n17479 = n17478 ^ n14016 ^ 1'b0 ;
  assign n17480 = n12163 ^ n11143 ^ 1'b0 ;
  assign n17481 = n17480 ^ n14490 ^ 1'b0 ;
  assign n17488 = n3127 ^ x202 ^ 1'b0 ;
  assign n17482 = n6995 ^ n1199 ^ 1'b0 ;
  assign n17483 = ( n2014 & n2916 ) | ( n2014 & n10225 ) | ( n2916 & n10225 ) ;
  assign n17484 = ~n2455 & n17483 ;
  assign n17485 = n17482 & n17484 ;
  assign n17486 = ( n7727 & ~n7988 ) | ( n7727 & n11078 ) | ( ~n7988 & n11078 ) ;
  assign n17487 = ~n17485 & n17486 ;
  assign n17489 = n17488 ^ n17487 ^ 1'b0 ;
  assign n17490 = ~n6830 & n9201 ;
  assign n17491 = n17490 ^ n766 ^ 1'b0 ;
  assign n17492 = n17491 ^ n14612 ^ n2284 ;
  assign n17493 = n547 & ~n9475 ;
  assign n17494 = ~n17343 & n17483 ;
  assign n17495 = n17494 ^ n506 ^ 1'b0 ;
  assign n17496 = n4646 & ~n17495 ;
  assign n17497 = n17496 ^ n563 ^ 1'b0 ;
  assign n17498 = n7435 | n11872 ;
  assign n17499 = n4656 | n17498 ;
  assign n17500 = ( n1478 & n2350 ) | ( n1478 & ~n17499 ) | ( n2350 & ~n17499 ) ;
  assign n17501 = ( ~n2518 & n3220 ) | ( ~n2518 & n17500 ) | ( n3220 & n17500 ) ;
  assign n17502 = ( n7982 & ~n17497 ) | ( n7982 & n17501 ) | ( ~n17497 & n17501 ) ;
  assign n17503 = n17374 ^ n2853 ^ 1'b0 ;
  assign n17504 = ~n5725 & n17503 ;
  assign n17505 = n9502 & n17504 ;
  assign n17506 = n4507 & n17505 ;
  assign n17507 = ( n972 & n4284 ) | ( n972 & n17506 ) | ( n4284 & n17506 ) ;
  assign n17508 = n1129 & ~n11643 ;
  assign n17509 = n14178 & ~n17508 ;
  assign n17510 = ~n921 & n17509 ;
  assign n17511 = ~n2829 & n4844 ;
  assign n17512 = n3450 & n17511 ;
  assign n17514 = n12199 ^ n9672 ^ n2081 ;
  assign n17513 = n14892 ^ n11428 ^ 1'b0 ;
  assign n17515 = n17514 ^ n17513 ^ 1'b0 ;
  assign n17517 = n7950 ^ n7597 ^ n2247 ;
  assign n17518 = n17517 ^ n10822 ^ 1'b0 ;
  assign n17519 = n17518 ^ n3628 ^ n2708 ;
  assign n17516 = n5400 | n10563 ;
  assign n17520 = n17519 ^ n17516 ^ n12503 ;
  assign n17521 = n6218 | n14335 ;
  assign n17522 = n11577 & ~n17521 ;
  assign n17523 = n3318 ^ n1120 ^ 1'b0 ;
  assign n17524 = n4889 & ~n17523 ;
  assign n17525 = n17524 ^ n14067 ^ n5592 ;
  assign n17526 = ( x147 & n3894 ) | ( x147 & ~n6929 ) | ( n3894 & ~n6929 ) ;
  assign n17527 = n1358 | n17526 ;
  assign n17528 = ( n2849 & n11248 ) | ( n2849 & n17527 ) | ( n11248 & n17527 ) ;
  assign n17529 = n3234 | n4676 ;
  assign n17530 = x38 | n17529 ;
  assign n17531 = n3048 ^ x195 ^ 1'b0 ;
  assign n17532 = n5972 & ~n17531 ;
  assign n17533 = n11792 ^ n5017 ^ 1'b0 ;
  assign n17534 = n17532 & ~n17533 ;
  assign n17535 = ~n13802 & n17534 ;
  assign n17536 = n17535 ^ n853 ^ 1'b0 ;
  assign n17537 = n15443 ^ n2519 ^ n1237 ;
  assign n17538 = ~n6035 & n17537 ;
  assign n17539 = n17536 & n17538 ;
  assign n17540 = ( ~n5033 & n9557 ) | ( ~n5033 & n13664 ) | ( n9557 & n13664 ) ;
  assign n17541 = n6493 ^ n4196 ^ 1'b0 ;
  assign n17542 = n2342 | n17541 ;
  assign n17543 = ( n9058 & ~n9783 ) | ( n9058 & n17542 ) | ( ~n9783 & n17542 ) ;
  assign n17544 = ~n1233 & n1989 ;
  assign n17545 = ~n6842 & n17544 ;
  assign n17546 = n17545 ^ n9067 ^ 1'b0 ;
  assign n17547 = n1033 & n1150 ;
  assign n17548 = n17547 ^ n432 ^ 1'b0 ;
  assign n17549 = ( n5799 & n7226 ) | ( n5799 & n17548 ) | ( n7226 & n17548 ) ;
  assign n17550 = n17549 ^ n8148 ^ x200 ;
  assign n17554 = n4701 ^ n2272 ^ 1'b0 ;
  assign n17551 = n10077 ^ n7948 ^ 1'b0 ;
  assign n17552 = n9652 & n17551 ;
  assign n17553 = n7629 & n17552 ;
  assign n17555 = n17554 ^ n17553 ^ 1'b0 ;
  assign n17556 = n2929 & ~n5420 ;
  assign n17557 = n14130 & n17556 ;
  assign n17558 = ( n3723 & n5542 ) | ( n3723 & ~n17557 ) | ( n5542 & ~n17557 ) ;
  assign n17559 = n17558 ^ n8323 ^ 1'b0 ;
  assign n17560 = n3534 | n17559 ;
  assign n17561 = n11357 ^ n4772 ^ 1'b0 ;
  assign n17562 = ~n4622 & n10495 ;
  assign n17563 = n1350 & n17562 ;
  assign n17564 = n2732 ^ n727 ^ 1'b0 ;
  assign n17565 = ~n17563 & n17564 ;
  assign n17566 = n11938 ^ n5081 ^ 1'b0 ;
  assign n17567 = n17565 & n17566 ;
  assign n17568 = ( ~n3708 & n3765 ) | ( ~n3708 & n7622 ) | ( n3765 & n7622 ) ;
  assign n17569 = n1919 & ~n4984 ;
  assign n17570 = n17569 ^ x77 ^ 1'b0 ;
  assign n17571 = n17570 ^ n1581 ^ 1'b0 ;
  assign n17573 = n13799 ^ n7260 ^ 1'b0 ;
  assign n17574 = n4516 & ~n17573 ;
  assign n17572 = n1160 ^ n759 ^ 1'b0 ;
  assign n17575 = n17574 ^ n17572 ^ 1'b0 ;
  assign n17576 = n16905 & n17575 ;
  assign n17577 = n5338 & n7105 ;
  assign n17578 = n12822 & n17577 ;
  assign n17579 = n1687 & n13349 ;
  assign n17580 = n7899 & n17579 ;
  assign n17581 = n4194 & n12339 ;
  assign n17582 = n17581 ^ n11608 ^ 1'b0 ;
  assign n17583 = n17263 ^ n14449 ^ 1'b0 ;
  assign n17584 = n17582 | n17583 ;
  assign n17585 = n5655 ^ n1657 ^ 1'b0 ;
  assign n17586 = x198 & ~n17585 ;
  assign n17587 = n7484 ^ n5832 ^ 1'b0 ;
  assign n17588 = n2521 & ~n17587 ;
  assign n17589 = ~n12152 & n17588 ;
  assign n17590 = n17589 ^ n7647 ^ 1'b0 ;
  assign n17591 = n1958 & ~n12524 ;
  assign n17592 = n13553 | n17591 ;
  assign n17593 = n1768 & ~n13419 ;
  assign n17594 = n7428 & n16373 ;
  assign n17595 = n17594 ^ n3395 ^ 1'b0 ;
  assign n17596 = n5262 & ~n6774 ;
  assign n17597 = n10517 ^ n1081 ^ 1'b0 ;
  assign n17598 = n2012 & ~n11153 ;
  assign n17599 = n7756 ^ n7559 ^ 1'b0 ;
  assign n17600 = n17598 & n17599 ;
  assign n17601 = n3534 & n17600 ;
  assign n17602 = x26 & ~n14417 ;
  assign n17603 = ( n4775 & ~n8752 ) | ( n4775 & n10617 ) | ( ~n8752 & n10617 ) ;
  assign n17604 = n15532 & ~n17603 ;
  assign n17605 = n17604 ^ n5207 ^ 1'b0 ;
  assign n17606 = n3672 ^ n1233 ^ 1'b0 ;
  assign n17607 = ~n11138 & n17606 ;
  assign n17608 = n11014 ^ n2281 ^ 1'b0 ;
  assign n17609 = n17607 & n17608 ;
  assign n17610 = n5022 | n6577 ;
  assign n17611 = n17610 ^ n956 ^ 1'b0 ;
  assign n17612 = n6798 ^ n1930 ^ 1'b0 ;
  assign n17613 = n17611 & ~n17612 ;
  assign n17614 = n17613 ^ n8606 ^ n8410 ;
  assign n17615 = n9772 | n17614 ;
  assign n17616 = n9552 & ~n17615 ;
  assign n17617 = n1306 | n13189 ;
  assign n17618 = n12537 ^ n3769 ^ 1'b0 ;
  assign n17619 = n17618 ^ n10026 ^ n751 ;
  assign n17620 = ( ~x254 & n1152 ) | ( ~x254 & n7367 ) | ( n1152 & n7367 ) ;
  assign n17621 = n17620 ^ n593 ^ 1'b0 ;
  assign n17622 = ~n12191 & n17621 ;
  assign n17623 = n6276 ^ n3371 ^ 1'b0 ;
  assign n17624 = n14450 | n17623 ;
  assign n17625 = n5147 ^ n1097 ^ 1'b0 ;
  assign n17626 = n15034 | n17625 ;
  assign n17627 = n4670 & ~n17626 ;
  assign n17628 = ~n12069 & n17627 ;
  assign n17629 = n10085 | n17628 ;
  assign n17630 = n3013 | n7505 ;
  assign n17631 = n17630 ^ n7488 ^ 1'b0 ;
  assign n17632 = n17631 ^ n3248 ^ 1'b0 ;
  assign n17633 = n1130 & ~n17632 ;
  assign n17634 = ~n7636 & n17633 ;
  assign n17635 = ( ~n2054 & n6665 ) | ( ~n2054 & n17634 ) | ( n6665 & n17634 ) ;
  assign n17636 = n3558 & ~n5554 ;
  assign n17637 = n4703 | n5038 ;
  assign n17638 = n17637 ^ n4821 ^ 1'b0 ;
  assign n17639 = ~n4137 & n8205 ;
  assign n17640 = ~n7937 & n17639 ;
  assign n17641 = n5600 | n13021 ;
  assign n17642 = n12853 & ~n17641 ;
  assign n17643 = n17640 | n17642 ;
  assign n17644 = n17638 & ~n17643 ;
  assign n17645 = ( ~n8488 & n17636 ) | ( ~n8488 & n17644 ) | ( n17636 & n17644 ) ;
  assign n17646 = n17125 ^ n13271 ^ 1'b0 ;
  assign n17647 = ~n758 & n17283 ;
  assign n17648 = n13859 & n17647 ;
  assign n17649 = n1830 | n13452 ;
  assign n17650 = n2829 | n17649 ;
  assign n17651 = n12550 & n17650 ;
  assign n17652 = ~n16933 & n17651 ;
  assign n17653 = n866 | n17652 ;
  assign n17654 = n2302 | n8640 ;
  assign n17655 = n8900 ^ n3632 ^ 1'b0 ;
  assign n17656 = ~n17654 & n17655 ;
  assign n17657 = ~n2925 & n17656 ;
  assign n17658 = n17657 ^ n8428 ^ 1'b0 ;
  assign n17659 = n4858 ^ n2020 ^ 1'b0 ;
  assign n17660 = ~n9491 & n17659 ;
  assign n17661 = n17660 ^ n17235 ^ 1'b0 ;
  assign n17662 = n2359 & ~n17661 ;
  assign n17663 = ( n2204 & n3772 ) | ( n2204 & n4602 ) | ( n3772 & n4602 ) ;
  assign n17664 = n17663 ^ n1124 ^ 1'b0 ;
  assign n17665 = ~n4909 & n17664 ;
  assign n17666 = ( ~n9263 & n17113 ) | ( ~n9263 & n17665 ) | ( n17113 & n17665 ) ;
  assign n17667 = ( n17658 & ~n17662 ) | ( n17658 & n17666 ) | ( ~n17662 & n17666 ) ;
  assign n17668 = n1040 ^ x191 ^ 1'b0 ;
  assign n17669 = n16781 & ~n17668 ;
  assign n17670 = n15721 ^ n4283 ^ 1'b0 ;
  assign n17671 = n17670 ^ n4309 ^ 1'b0 ;
  assign n17672 = ~n17669 & n17671 ;
  assign n17673 = n13383 ^ n3048 ^ 1'b0 ;
  assign n17674 = n3746 & ~n17673 ;
  assign n17675 = n349 | n5141 ;
  assign n17676 = n349 & ~n17675 ;
  assign n17677 = n10675 ^ n10444 ^ n1233 ;
  assign n17678 = n332 | n6584 ;
  assign n17679 = n15666 & n17678 ;
  assign n17680 = n13555 & n17679 ;
  assign n17681 = n1752 | n8078 ;
  assign n17682 = n17681 ^ n14370 ^ 1'b0 ;
  assign n17683 = ~n7374 & n17682 ;
  assign n17684 = n8051 ^ n3156 ^ 1'b0 ;
  assign n17685 = n17684 ^ n4306 ^ 1'b0 ;
  assign n17688 = ~n4726 & n14163 ;
  assign n17689 = n17688 ^ n10288 ^ 1'b0 ;
  assign n17686 = n11807 | n12881 ;
  assign n17687 = n7950 & ~n17686 ;
  assign n17690 = n17689 ^ n17687 ^ n7115 ;
  assign n17691 = n5730 ^ n1666 ^ 1'b0 ;
  assign n17693 = n7215 ^ n2543 ^ 1'b0 ;
  assign n17694 = ~n1210 & n17693 ;
  assign n17692 = n2452 ^ n411 ^ x2 ;
  assign n17695 = n17694 ^ n17692 ^ 1'b0 ;
  assign n17696 = n5428 | n8537 ;
  assign n17697 = n17696 ^ n2757 ^ 1'b0 ;
  assign n17698 = n1961 & n3690 ;
  assign n17699 = n17698 ^ n1804 ^ 1'b0 ;
  assign n17700 = ~n954 & n17699 ;
  assign n17701 = n8647 ^ n1639 ^ 1'b0 ;
  assign n17702 = n2339 | n7664 ;
  assign n17703 = n12539 ^ n3542 ^ 1'b0 ;
  assign n17704 = n5306 & ~n17703 ;
  assign n17705 = n17704 ^ n5601 ^ 1'b0 ;
  assign n17706 = ~n11030 & n17705 ;
  assign n17707 = n17706 ^ n13617 ^ 1'b0 ;
  assign n17708 = ( n3230 & n10975 ) | ( n3230 & ~n17707 ) | ( n10975 & ~n17707 ) ;
  assign n17709 = n4626 | n12194 ;
  assign n17710 = n1321 & ~n17709 ;
  assign n17711 = n3831 & ~n17710 ;
  assign n17712 = n17711 ^ n13094 ^ 1'b0 ;
  assign n17713 = n2530 ^ x242 ^ 1'b0 ;
  assign n17714 = ( n845 & n13293 ) | ( n845 & ~n14557 ) | ( n13293 & ~n14557 ) ;
  assign n17715 = n1991 & ~n7942 ;
  assign n17716 = n2395 & n11369 ;
  assign n17717 = n17716 ^ n7569 ^ n3874 ;
  assign n17718 = n9693 & n17717 ;
  assign n17719 = ~n5550 & n17718 ;
  assign n17721 = n9097 ^ n2708 ^ 1'b0 ;
  assign n17722 = n5608 | n17721 ;
  assign n17720 = n13171 ^ n4977 ^ 1'b0 ;
  assign n17723 = n17722 ^ n17720 ^ n9411 ;
  assign n17724 = ( n4236 & n8261 ) | ( n4236 & ~n10617 ) | ( n8261 & ~n10617 ) ;
  assign n17725 = n17724 ^ n12718 ^ n3141 ;
  assign n17726 = n8352 ^ n593 ^ 1'b0 ;
  assign n17727 = ~n3608 & n17726 ;
  assign n17728 = n8662 ^ n1829 ^ 1'b0 ;
  assign n17729 = n14724 & n17728 ;
  assign n17730 = n14016 ^ n11249 ^ n3202 ;
  assign n17734 = n1890 | n13523 ;
  assign n17735 = n17734 ^ x36 ^ 1'b0 ;
  assign n17731 = ( n5053 & ~n5993 ) | ( n5053 & n10141 ) | ( ~n5993 & n10141 ) ;
  assign n17732 = n8425 & ~n9525 ;
  assign n17733 = ~n17731 & n17732 ;
  assign n17736 = n17735 ^ n17733 ^ 1'b0 ;
  assign n17737 = n6599 | n17736 ;
  assign n17738 = ( n6198 & ~n7145 ) | ( n6198 & n13030 ) | ( ~n7145 & n13030 ) ;
  assign n17739 = n492 & n2282 ;
  assign n17740 = ( n3249 & n5988 ) | ( n3249 & n13695 ) | ( n5988 & n13695 ) ;
  assign n17741 = n17740 ^ n2070 ^ 1'b0 ;
  assign n17742 = ~n17739 & n17741 ;
  assign n17743 = ~n3985 & n16729 ;
  assign n17744 = ~n10982 & n17743 ;
  assign n17745 = n2989 | n7918 ;
  assign n17746 = n5907 ^ x11 ^ 1'b0 ;
  assign n17747 = n7536 & ~n17746 ;
  assign n17748 = ( n5634 & n17745 ) | ( n5634 & ~n17747 ) | ( n17745 & ~n17747 ) ;
  assign n17749 = n17748 ^ n13140 ^ 1'b0 ;
  assign n17751 = n2204 | n9295 ;
  assign n17752 = n6249 & ~n17751 ;
  assign n17750 = n1400 | n7341 ;
  assign n17753 = n17752 ^ n17750 ^ 1'b0 ;
  assign n17754 = n7336 ^ n2332 ^ 1'b0 ;
  assign n17755 = ( ~n11201 & n15423 ) | ( ~n11201 & n17754 ) | ( n15423 & n17754 ) ;
  assign n17756 = n12931 ^ n5942 ^ 1'b0 ;
  assign n17757 = n12333 & ~n17756 ;
  assign n17758 = ~n2420 & n2699 ;
  assign n17759 = n17758 ^ n9513 ^ 1'b0 ;
  assign n17760 = n14266 | n17759 ;
  assign n17761 = n2093 & n8471 ;
  assign n17762 = n17761 ^ n14807 ^ 1'b0 ;
  assign n17763 = ~n12890 & n17762 ;
  assign n17767 = n9178 ^ n2047 ^ 1'b0 ;
  assign n17764 = ~n1553 & n11521 ;
  assign n17765 = n17764 ^ n7805 ^ 1'b0 ;
  assign n17766 = n1293 | n17765 ;
  assign n17768 = n17767 ^ n17766 ^ 1'b0 ;
  assign n17769 = n6605 ^ n2829 ^ 1'b0 ;
  assign n17770 = n933 | n1227 ;
  assign n17771 = n17769 | n17770 ;
  assign n17772 = n17771 ^ n13945 ^ n1144 ;
  assign n17773 = ~n2592 & n17772 ;
  assign n17774 = ~n6601 & n17773 ;
  assign n17775 = n4405 | n5920 ;
  assign n17776 = n4845 & n17775 ;
  assign n17777 = n10997 & ~n17776 ;
  assign n17778 = n17777 ^ n14371 ^ 1'b0 ;
  assign n17782 = ~n5817 & n15508 ;
  assign n17779 = n3907 ^ n1937 ^ 1'b0 ;
  assign n17780 = n2943 & ~n17779 ;
  assign n17781 = n8455 & n17780 ;
  assign n17783 = n17782 ^ n17781 ^ 1'b0 ;
  assign n17784 = ~n7583 & n8945 ;
  assign n17785 = n5584 ^ n3951 ^ 1'b0 ;
  assign n17786 = n17784 | n17785 ;
  assign n17787 = ~n8298 & n13079 ;
  assign n17788 = n11087 & n17787 ;
  assign n17789 = n11048 ^ n9211 ^ n7777 ;
  assign n17790 = ~n14793 & n17789 ;
  assign n17791 = n17788 & n17790 ;
  assign n17792 = ~n385 & n10828 ;
  assign n17793 = n17792 ^ n15829 ^ 1'b0 ;
  assign n17794 = n9309 & ~n17793 ;
  assign n17798 = n626 | n4853 ;
  assign n17799 = n17798 ^ n5613 ^ n5529 ;
  assign n17795 = n11907 ^ n10932 ^ 1'b0 ;
  assign n17796 = ~x177 & n5495 ;
  assign n17797 = n17795 | n17796 ;
  assign n17800 = n17799 ^ n17797 ^ 1'b0 ;
  assign n17801 = n17800 ^ n12489 ^ 1'b0 ;
  assign n17802 = ~n4480 & n17801 ;
  assign n17803 = n2761 & ~n5395 ;
  assign n17804 = n16183 ^ n12454 ^ n11844 ;
  assign n17809 = n3398 & n8320 ;
  assign n17805 = x134 & ~n10749 ;
  assign n17806 = n17805 ^ n494 ^ 1'b0 ;
  assign n17807 = n17806 ^ n7481 ^ 1'b0 ;
  assign n17808 = n17807 ^ x26 ^ 1'b0 ;
  assign n17810 = n17809 ^ n17808 ^ 1'b0 ;
  assign n17811 = n3806 & ~n13707 ;
  assign n17812 = n17811 ^ n12330 ^ 1'b0 ;
  assign n17814 = n8156 ^ n1998 ^ 1'b0 ;
  assign n17815 = n4194 & ~n17814 ;
  assign n17813 = n2690 ^ n1142 ^ 1'b0 ;
  assign n17816 = n17815 ^ n17813 ^ 1'b0 ;
  assign n17817 = n17816 ^ n4726 ^ n1409 ;
  assign n17818 = n17817 ^ n17605 ^ 1'b0 ;
  assign n17819 = ~n2076 & n9651 ;
  assign n17820 = n5070 & n17819 ;
  assign n17821 = n17820 ^ n495 ^ 1'b0 ;
  assign n17822 = n17681 & n17821 ;
  assign n17823 = n13338 ^ n11024 ^ 1'b0 ;
  assign n17824 = n17822 & ~n17823 ;
  assign n17825 = ~n17822 & n17824 ;
  assign n17826 = ~n10179 & n17808 ;
  assign n17827 = ~n5850 & n17826 ;
  assign n17828 = ~n13246 & n17827 ;
  assign n17829 = n9964 ^ n4066 ^ n829 ;
  assign n17830 = n2284 | n16211 ;
  assign n17831 = n17830 ^ n15389 ^ 1'b0 ;
  assign n17832 = n7298 | n17831 ;
  assign n17833 = n17829 & ~n17832 ;
  assign n17834 = n8688 & n17833 ;
  assign n17835 = n7475 & n10217 ;
  assign n17836 = n9077 | n11107 ;
  assign n17837 = n8930 | n17836 ;
  assign n17838 = n17837 ^ n697 ^ 1'b0 ;
  assign n17839 = ~n10728 & n16467 ;
  assign n17840 = ~n4354 & n8087 ;
  assign n17841 = ~n14219 & n17840 ;
  assign n17842 = n17076 ^ n10794 ^ 1'b0 ;
  assign n17843 = n5855 | n17842 ;
  assign n17844 = n11321 ^ n2647 ^ 1'b0 ;
  assign n17845 = n9005 | n17844 ;
  assign n17846 = n17845 ^ n1803 ^ 1'b0 ;
  assign n17847 = n13985 ^ n2230 ^ n1802 ;
  assign n17848 = n17847 ^ n7237 ^ 1'b0 ;
  assign n17849 = n17846 | n17848 ;
  assign n17850 = n17849 ^ n6693 ^ 1'b0 ;
  assign n17851 = n15468 | n17850 ;
  assign n17852 = n2315 & n13894 ;
  assign n17853 = ( n16156 & n16987 ) | ( n16156 & n17852 ) | ( n16987 & n17852 ) ;
  assign n17854 = n11705 ^ n6979 ^ n4853 ;
  assign n17855 = n16278 ^ n4083 ^ 1'b0 ;
  assign n17856 = ( n2041 & n5327 ) | ( n2041 & n14222 ) | ( n5327 & n14222 ) ;
  assign n17857 = n8794 & n17856 ;
  assign n17858 = n1671 | n4436 ;
  assign n17859 = n6348 | n17858 ;
  assign n17860 = n2601 & n17859 ;
  assign n17861 = n17860 ^ n9375 ^ 1'b0 ;
  assign n17862 = n7806 & ~n17861 ;
  assign n17863 = n6421 & ~n7887 ;
  assign n17864 = ~n17862 & n17863 ;
  assign n17865 = n14479 ^ n719 ^ 1'b0 ;
  assign n17866 = ( n2441 & n4105 ) | ( n2441 & ~n13036 ) | ( n4105 & ~n13036 ) ;
  assign n17867 = x234 | n16952 ;
  assign n17870 = ~n1358 & n16464 ;
  assign n17871 = n17870 ^ n6112 ^ 1'b0 ;
  assign n17868 = n8737 & ~n15819 ;
  assign n17869 = n4379 & n17868 ;
  assign n17872 = n17871 ^ n17869 ^ 1'b0 ;
  assign n17873 = ( n17866 & ~n17867 ) | ( n17866 & n17872 ) | ( ~n17867 & n17872 ) ;
  assign n17874 = n17873 ^ n14696 ^ x227 ;
  assign n17875 = n9916 | n11304 ;
  assign n17876 = n17875 ^ n17461 ^ n12959 ;
  assign n17877 = n8836 & n10162 ;
  assign n17878 = n17877 ^ n13349 ^ 1'b0 ;
  assign n17879 = ~n2630 & n9708 ;
  assign n17880 = n17879 ^ n2450 ^ 1'b0 ;
  assign n17881 = ( ~n4343 & n5549 ) | ( ~n4343 & n6241 ) | ( n5549 & n6241 ) ;
  assign n17882 = n17881 ^ n12910 ^ n10585 ;
  assign n17883 = n2255 & ~n4089 ;
  assign n17884 = n17883 ^ n10309 ^ 1'b0 ;
  assign n17885 = n1059 & n5336 ;
  assign n17886 = n11136 & ~n17885 ;
  assign n17887 = ~n17884 & n17886 ;
  assign n17888 = n10129 ^ n4656 ^ 1'b0 ;
  assign n17889 = n4601 & n6227 ;
  assign n17890 = n9101 | n11719 ;
  assign n17891 = n17889 | n17890 ;
  assign n17892 = n7739 ^ n342 ^ 1'b0 ;
  assign n17893 = ~n9831 & n17892 ;
  assign n17894 = ~x210 & n17893 ;
  assign n17895 = n5982 & ~n17894 ;
  assign n17896 = ~n7411 & n9559 ;
  assign n17897 = x57 | n1430 ;
  assign n17898 = n4448 & n17729 ;
  assign n17899 = n13692 & n17898 ;
  assign n17900 = n2913 & n16808 ;
  assign n17901 = n15569 & n17900 ;
  assign n17902 = n5230 & n17901 ;
  assign n17903 = ( n2059 & n3564 ) | ( n2059 & n8351 ) | ( n3564 & n8351 ) ;
  assign n17904 = n5567 & n17903 ;
  assign n17905 = n4325 & n17904 ;
  assign n17906 = ~n6985 & n7673 ;
  assign n17907 = n11688 & n17906 ;
  assign n17908 = n17905 | n17907 ;
  assign n17909 = n17908 ^ n8409 ^ 1'b0 ;
  assign n17910 = ~n4597 & n7031 ;
  assign n17911 = n3686 & ~n6830 ;
  assign n17912 = n17911 ^ n10348 ^ n5681 ;
  assign n17913 = n5025 ^ n1989 ^ 1'b0 ;
  assign n17914 = ( ~n4216 & n7820 ) | ( ~n4216 & n14003 ) | ( n7820 & n14003 ) ;
  assign n17915 = n8760 ^ n7995 ^ 1'b0 ;
  assign n17916 = ~n13347 & n17915 ;
  assign n17917 = n8898 | n10640 ;
  assign n17918 = ~n12304 & n17917 ;
  assign n17919 = n11489 ^ n4585 ^ 1'b0 ;
  assign n17920 = n17919 ^ n15778 ^ 1'b0 ;
  assign n17921 = n11521 & n17920 ;
  assign n17922 = ~n840 & n2502 ;
  assign n17923 = n17922 ^ n14049 ^ 1'b0 ;
  assign n17924 = n2044 & ~n15162 ;
  assign n17925 = ~n12152 & n17924 ;
  assign n17926 = n4957 | n12312 ;
  assign n17927 = n17926 ^ n10766 ^ 1'b0 ;
  assign n17928 = n17927 ^ n15564 ^ 1'b0 ;
  assign n17929 = ( n4264 & ~n6647 ) | ( n4264 & n7206 ) | ( ~n6647 & n7206 ) ;
  assign n17930 = n12089 & n12630 ;
  assign n17931 = n17930 ^ n13589 ^ 1'b0 ;
  assign n17935 = n7492 ^ n7213 ^ 1'b0 ;
  assign n17932 = n7408 ^ n5641 ^ 1'b0 ;
  assign n17933 = n16267 ^ n12405 ^ 1'b0 ;
  assign n17934 = n17932 & ~n17933 ;
  assign n17936 = n17935 ^ n17934 ^ n16879 ;
  assign n17937 = x219 & n3980 ;
  assign n17938 = ~n17467 & n17937 ;
  assign n17939 = n17938 ^ x42 ^ 1'b0 ;
  assign n17940 = n16307 ^ n13799 ^ 1'b0 ;
  assign n17941 = n16344 & n17940 ;
  assign n17942 = n5285 & n7241 ;
  assign n17943 = n5804 & ~n17942 ;
  assign n17944 = n9843 & ~n13695 ;
  assign n17945 = ~n666 & n17944 ;
  assign n17946 = n16625 ^ n6808 ^ 1'b0 ;
  assign n17947 = n12783 & ~n16884 ;
  assign n17948 = n17947 ^ n8997 ^ 1'b0 ;
  assign n17949 = n3336 & n6660 ;
  assign n17950 = n17949 ^ n8908 ^ 1'b0 ;
  assign n17951 = n17948 | n17950 ;
  assign n17954 = ~n6023 & n10227 ;
  assign n17952 = n6414 ^ n1160 ^ 1'b0 ;
  assign n17953 = n9652 & n17952 ;
  assign n17955 = n17954 ^ n17953 ^ 1'b0 ;
  assign n17956 = ~n778 & n17955 ;
  assign n17957 = x31 & n2601 ;
  assign n17958 = n17957 ^ n11599 ^ 1'b0 ;
  assign n17959 = n2081 & ~n9163 ;
  assign n17960 = n17958 & n17959 ;
  assign n17961 = n489 & ~n1521 ;
  assign n17962 = n3348 ^ n289 ^ 1'b0 ;
  assign n17963 = n10715 | n17962 ;
  assign n17964 = n17961 & ~n17963 ;
  assign n17965 = n326 | n5257 ;
  assign n17966 = n9435 | n10633 ;
  assign n17967 = n14399 & ~n17966 ;
  assign n17968 = n10689 ^ n7510 ^ 1'b0 ;
  assign n17969 = n17968 ^ n9081 ^ 1'b0 ;
  assign n17970 = ~n1517 & n1581 ;
  assign n17971 = n17970 ^ n5562 ^ 1'b0 ;
  assign n17972 = n10400 ^ n344 ^ 1'b0 ;
  assign n17973 = ~n17971 & n17972 ;
  assign n17974 = ( n3055 & n8017 ) | ( n3055 & n17958 ) | ( n8017 & n17958 ) ;
  assign n17975 = n17974 ^ n2525 ^ 1'b0 ;
  assign n17976 = ~n2371 & n17975 ;
  assign n17978 = ~n4287 & n16070 ;
  assign n17979 = n480 & n17978 ;
  assign n17980 = ( n14777 & n17628 ) | ( n14777 & ~n17979 ) | ( n17628 & ~n17979 ) ;
  assign n17981 = n9978 & ~n17980 ;
  assign n17982 = ~n9764 & n17981 ;
  assign n17977 = n7349 & n17006 ;
  assign n17983 = n17982 ^ n17977 ^ 1'b0 ;
  assign n17984 = ~n4959 & n16626 ;
  assign n17985 = n17984 ^ n7796 ^ 1'b0 ;
  assign n17986 = n17985 ^ n6541 ^ n3690 ;
  assign n17988 = n3825 & n6360 ;
  assign n17987 = n4170 | n13521 ;
  assign n17989 = n17988 ^ n17987 ^ 1'b0 ;
  assign n17990 = n5850 ^ n1192 ^ 1'b0 ;
  assign n17991 = n17989 & n17990 ;
  assign n17992 = n5914 | n6964 ;
  assign n17993 = n2685 & n11007 ;
  assign n17994 = n8864 & ~n17993 ;
  assign n17995 = n5105 & ~n17994 ;
  assign n17996 = n17992 & n17995 ;
  assign n17997 = n6481 | n13458 ;
  assign n17998 = n17997 ^ n5328 ^ 1'b0 ;
  assign n17999 = ~n6654 & n14926 ;
  assign n18000 = n17999 ^ n11854 ^ 1'b0 ;
  assign n18002 = ~n1233 & n1665 ;
  assign n18003 = n1124 & n18002 ;
  assign n18004 = ~n3926 & n18003 ;
  assign n18001 = n4833 & n8529 ;
  assign n18005 = n18004 ^ n18001 ^ 1'b0 ;
  assign n18006 = ( n4626 & n7890 ) | ( n4626 & n18005 ) | ( n7890 & n18005 ) ;
  assign n18007 = n18006 ^ n2264 ^ 1'b0 ;
  assign n18008 = n1324 ^ n610 ^ 1'b0 ;
  assign n18009 = ( ~n3176 & n7597 ) | ( ~n3176 & n12148 ) | ( n7597 & n12148 ) ;
  assign n18010 = n12555 & ~n18009 ;
  assign n18011 = n13291 & n18010 ;
  assign n18012 = n14625 ^ n1963 ^ 1'b0 ;
  assign n18013 = ~n1873 & n18012 ;
  assign n18014 = ~n10212 & n18013 ;
  assign n18015 = ( n3935 & n4815 ) | ( n3935 & n10097 ) | ( n4815 & n10097 ) ;
  assign n18016 = n10323 ^ n5852 ^ n1186 ;
  assign n18017 = n6422 ^ n3441 ^ 1'b0 ;
  assign n18018 = n18016 & ~n18017 ;
  assign n18019 = n18018 ^ n752 ^ 1'b0 ;
  assign n18020 = n18015 | n18019 ;
  assign n18021 = n18014 & ~n18020 ;
  assign n18022 = n18021 ^ n16420 ^ 1'b0 ;
  assign n18025 = n4346 ^ n2812 ^ 1'b0 ;
  assign n18024 = ( n5489 & n7778 ) | ( n5489 & n13142 ) | ( n7778 & n13142 ) ;
  assign n18026 = n18025 ^ n18024 ^ n4584 ;
  assign n18023 = n6516 & ~n9746 ;
  assign n18027 = n18026 ^ n18023 ^ 1'b0 ;
  assign n18028 = x118 & n11457 ;
  assign n18029 = ( n8194 & n8921 ) | ( n8194 & ~n18028 ) | ( n8921 & ~n18028 ) ;
  assign n18030 = ( n4275 & n5114 ) | ( n4275 & ~n13245 ) | ( n5114 & ~n13245 ) ;
  assign n18031 = n12277 & ~n18030 ;
  assign n18032 = ~n3786 & n5763 ;
  assign n18033 = ~n5581 & n18032 ;
  assign n18034 = n11376 ^ n4383 ^ 1'b0 ;
  assign n18035 = n18033 & ~n18034 ;
  assign n18036 = n2808 | n7945 ;
  assign n18037 = x185 | n18036 ;
  assign n18038 = n18037 ^ n14733 ^ 1'b0 ;
  assign n18039 = n11202 & ~n18038 ;
  assign n18041 = ~n2224 & n12435 ;
  assign n18042 = n6870 & n18041 ;
  assign n18040 = n10368 ^ n8555 ^ n2317 ;
  assign n18043 = n18042 ^ n18040 ^ n14803 ;
  assign n18044 = n17290 ^ n4865 ^ 1'b0 ;
  assign n18045 = n2441 | n18044 ;
  assign n18046 = n18043 & ~n18045 ;
  assign n18047 = n9314 ^ n6618 ^ 1'b0 ;
  assign n18048 = n1107 & ~n18047 ;
  assign n18049 = n18048 ^ n1906 ^ 1'b0 ;
  assign n18050 = n8491 ^ n3650 ^ 1'b0 ;
  assign n18051 = n1863 | n18050 ;
  assign n18052 = n3361 & ~n5586 ;
  assign n18053 = n15915 ^ n567 ^ 1'b0 ;
  assign n18054 = n11942 | n18053 ;
  assign n18058 = n9545 ^ n2149 ^ x58 ;
  assign n18059 = n10888 ^ n6268 ^ 1'b0 ;
  assign n18060 = n18058 & ~n18059 ;
  assign n18061 = ( ~n6131 & n8635 ) | ( ~n6131 & n18060 ) | ( n8635 & n18060 ) ;
  assign n18055 = n4672 ^ n2613 ^ n1724 ;
  assign n18056 = n18055 ^ n12548 ^ 1'b0 ;
  assign n18057 = n4567 & n18056 ;
  assign n18062 = n18061 ^ n18057 ^ 1'b0 ;
  assign n18063 = ~n1934 & n7678 ;
  assign n18064 = n10045 & n18063 ;
  assign n18065 = n11413 | n18064 ;
  assign n18066 = n5264 & ~n18065 ;
  assign n18067 = n3391 | n18066 ;
  assign n18068 = n18067 ^ n14472 ^ 1'b0 ;
  assign n18072 = n791 & n14016 ;
  assign n18073 = n7445 & n18072 ;
  assign n18070 = n6005 & ~n7721 ;
  assign n18071 = n2909 & ~n18070 ;
  assign n18074 = n18073 ^ n18071 ^ 1'b0 ;
  assign n18069 = n12633 ^ n2694 ^ n267 ;
  assign n18075 = n18074 ^ n18069 ^ 1'b0 ;
  assign n18076 = n1506 & ~n7647 ;
  assign n18077 = ~n12160 & n18076 ;
  assign n18078 = ~n4281 & n18077 ;
  assign n18082 = ( n2815 & n4775 ) | ( n2815 & n6938 ) | ( n4775 & n6938 ) ;
  assign n18079 = n428 | n12468 ;
  assign n18080 = n2915 & ~n18079 ;
  assign n18081 = n18080 ^ n317 ^ 1'b0 ;
  assign n18083 = n18082 ^ n18081 ^ 1'b0 ;
  assign n18084 = n1674 | n2528 ;
  assign n18085 = n18084 ^ n5262 ^ 1'b0 ;
  assign n18086 = n18085 ^ n833 ^ 1'b0 ;
  assign n18087 = n2722 | n18086 ;
  assign n18088 = n18087 ^ n9392 ^ 1'b0 ;
  assign n18089 = ~n723 & n18088 ;
  assign n18090 = n18089 ^ n9462 ^ 1'b0 ;
  assign n18091 = ( ~n465 & n5056 ) | ( ~n465 & n9076 ) | ( n5056 & n9076 ) ;
  assign n18092 = n13550 & n18091 ;
  assign n18093 = n3399 | n11773 ;
  assign n18094 = n16665 | n18093 ;
  assign n18095 = ( n1715 & ~n11990 ) | ( n1715 & n18094 ) | ( ~n11990 & n18094 ) ;
  assign n18096 = n6488 ^ n4317 ^ 1'b0 ;
  assign n18097 = ~n3960 & n6295 ;
  assign n18098 = ~n18096 & n18097 ;
  assign n18099 = n681 & ~n6807 ;
  assign n18100 = ~n546 & n16307 ;
  assign n18101 = n3904 | n5491 ;
  assign n18102 = n6047 & n18101 ;
  assign n18103 = n18102 ^ n13617 ^ 1'b0 ;
  assign n18104 = n1897 | n13880 ;
  assign n18105 = n3361 | n18104 ;
  assign n18106 = ~n3003 & n15628 ;
  assign n18107 = n14613 & n18106 ;
  assign n18108 = n12744 ^ n4799 ^ 1'b0 ;
  assign n18109 = n15827 & n17730 ;
  assign n18110 = n15418 ^ n4769 ^ 1'b0 ;
  assign n18111 = n6592 | n6847 ;
  assign n18112 = n3743 & ~n18111 ;
  assign n18113 = ( n7339 & n15774 ) | ( n7339 & n18112 ) | ( n15774 & n18112 ) ;
  assign n18114 = n6719 ^ n5614 ^ 1'b0 ;
  assign n18115 = ( ~n634 & n12597 ) | ( ~n634 & n18114 ) | ( n12597 & n18114 ) ;
  assign n18116 = ( n4705 & ~n6129 ) | ( n4705 & n7969 ) | ( ~n6129 & n7969 ) ;
  assign n18117 = n15930 & ~n18116 ;
  assign n18118 = n18117 ^ n5220 ^ 1'b0 ;
  assign n18119 = n3365 ^ n2518 ^ 1'b0 ;
  assign n18120 = n10396 & ~n18119 ;
  assign n18121 = ~n7844 & n15635 ;
  assign n18122 = n16427 & ~n18121 ;
  assign n18123 = n1692 & ~n12074 ;
  assign n18124 = n18123 ^ n6337 ^ n3282 ;
  assign n18125 = n15026 ^ n7700 ^ 1'b0 ;
  assign n18126 = ~n3059 & n13006 ;
  assign n18127 = n14085 ^ n7148 ^ 1'b0 ;
  assign n18128 = n4855 & n5740 ;
  assign n18129 = ~n2063 & n18128 ;
  assign n18130 = n9187 ^ x57 ^ 1'b0 ;
  assign n18131 = ( n326 & n9594 ) | ( n326 & n11304 ) | ( n9594 & n11304 ) ;
  assign n18132 = n9118 & n14009 ;
  assign n18133 = n8303 & n18132 ;
  assign n18134 = ~n5966 & n18133 ;
  assign n18135 = n18134 ^ n13839 ^ 1'b0 ;
  assign n18136 = ~n18131 & n18135 ;
  assign n18137 = n13608 ^ x99 ^ 1'b0 ;
  assign n18138 = n18137 ^ n1813 ^ 1'b0 ;
  assign n18139 = n17871 & n18138 ;
  assign n18140 = ~n5190 & n7507 ;
  assign n18142 = n1102 | n9866 ;
  assign n18143 = n18142 ^ n4359 ^ 1'b0 ;
  assign n18144 = ( n3436 & n10501 ) | ( n3436 & n18143 ) | ( n10501 & n18143 ) ;
  assign n18145 = n10832 & n18144 ;
  assign n18146 = ~x57 & n18145 ;
  assign n18141 = n12530 ^ n1313 ^ 1'b0 ;
  assign n18147 = n18146 ^ n18141 ^ 1'b0 ;
  assign n18148 = ~n15100 & n15851 ;
  assign n18149 = n2955 & n18148 ;
  assign n18154 = n18003 ^ n17264 ^ 1'b0 ;
  assign n18150 = n5049 ^ n1464 ^ 1'b0 ;
  assign n18151 = ( n11935 & n14905 ) | ( n11935 & ~n18150 ) | ( n14905 & ~n18150 ) ;
  assign n18152 = n267 | n18151 ;
  assign n18153 = n15724 | n18152 ;
  assign n18155 = n18154 ^ n18153 ^ 1'b0 ;
  assign n18156 = n11803 ^ n7335 ^ 1'b0 ;
  assign n18157 = n2936 ^ n2455 ^ n423 ;
  assign n18158 = n3497 & ~n4630 ;
  assign n18159 = n18158 ^ n6833 ^ 1'b0 ;
  assign n18160 = n18157 | n18159 ;
  assign n18163 = n13799 ^ n10246 ^ n9365 ;
  assign n18161 = n7480 ^ n4710 ^ 1'b0 ;
  assign n18162 = n11869 & n18161 ;
  assign n18164 = n18163 ^ n18162 ^ 1'b0 ;
  assign n18165 = n11565 & n18164 ;
  assign n18166 = n18160 & n18165 ;
  assign n18167 = ( ~n1274 & n1797 ) | ( ~n1274 & n10902 ) | ( n1797 & n10902 ) ;
  assign n18168 = n18167 ^ n8702 ^ n1097 ;
  assign n18169 = n6616 ^ n5441 ^ 1'b0 ;
  assign n18170 = n18169 ^ n6932 ^ 1'b0 ;
  assign n18171 = x96 & ~n18170 ;
  assign n18172 = ( ~n7165 & n13230 ) | ( ~n7165 & n18171 ) | ( n13230 & n18171 ) ;
  assign n18173 = n17482 ^ n8013 ^ 1'b0 ;
  assign n18174 = n18173 ^ x182 ^ 1'b0 ;
  assign n18175 = n18172 & ~n18174 ;
  assign n18176 = ~n1236 & n1835 ;
  assign n18177 = n18176 ^ n18156 ^ 1'b0 ;
  assign n18178 = ~n16578 & n18177 ;
  assign n18179 = n18178 ^ n12115 ^ 1'b0 ;
  assign n18180 = n11091 & ~n17638 ;
  assign n18181 = n18180 ^ n1763 ^ 1'b0 ;
  assign n18182 = n14617 ^ n7053 ^ n4030 ;
  assign n18183 = n14551 & ~n18182 ;
  assign n18184 = ( n1655 & ~n4688 ) | ( n1655 & n13091 ) | ( ~n4688 & n13091 ) ;
  assign n18185 = n4937 ^ n1961 ^ 1'b0 ;
  assign n18186 = n1246 & n5354 ;
  assign n18187 = n18186 ^ n935 ^ 1'b0 ;
  assign n18188 = n4196 ^ n2871 ^ n1842 ;
  assign n18189 = ( x229 & n533 ) | ( x229 & ~n18188 ) | ( n533 & ~n18188 ) ;
  assign n18190 = n18187 & n18189 ;
  assign n18191 = n4255 | n10214 ;
  assign n18192 = n13217 & n18191 ;
  assign n18193 = n18190 & n18192 ;
  assign n18194 = n18193 ^ x107 ^ 1'b0 ;
  assign n18195 = ~n7074 & n10572 ;
  assign n18196 = n18195 ^ n10576 ^ 1'b0 ;
  assign n18197 = n18196 ^ x65 ^ 1'b0 ;
  assign n18199 = n17806 ^ n2588 ^ 1'b0 ;
  assign n18200 = n13753 & ~n18199 ;
  assign n18198 = ~n2106 & n11136 ;
  assign n18201 = n18200 ^ n18198 ^ 1'b0 ;
  assign n18205 = n1236 | n2180 ;
  assign n18206 = n18205 ^ n3942 ^ 1'b0 ;
  assign n18207 = x244 & ~n18206 ;
  assign n18202 = n11772 ^ n6569 ^ n3210 ;
  assign n18203 = n18202 ^ n10083 ^ 1'b0 ;
  assign n18204 = n2966 & n18203 ;
  assign n18208 = n18207 ^ n18204 ^ 1'b0 ;
  assign n18209 = n1304 | n16439 ;
  assign n18210 = n14054 ^ n530 ^ 1'b0 ;
  assign n18211 = n18209 & n18210 ;
  assign n18212 = n8318 | n13404 ;
  assign n18213 = n18212 ^ n9365 ^ 1'b0 ;
  assign n18214 = ( n9326 & n15842 ) | ( n9326 & n18213 ) | ( n15842 & n18213 ) ;
  assign n18215 = n7499 | n10565 ;
  assign n18216 = n18215 ^ n4467 ^ 1'b0 ;
  assign n18217 = ~n4950 & n7636 ;
  assign n18218 = n18217 ^ n3523 ^ 1'b0 ;
  assign n18219 = n14926 & n18218 ;
  assign n18220 = n18216 & n18219 ;
  assign n18221 = n271 & ~n504 ;
  assign n18222 = n1069 & n18221 ;
  assign n18223 = n1145 & n3116 ;
  assign n18224 = n18222 & n18223 ;
  assign n18225 = ~n4528 & n6303 ;
  assign n18226 = n18225 ^ n2532 ^ 1'b0 ;
  assign n18227 = ~n10532 & n18226 ;
  assign n18228 = ~n15251 & n18150 ;
  assign n18229 = n5513 & ~n18228 ;
  assign n18230 = ~x168 & n8158 ;
  assign n18231 = ( n5681 & n13708 ) | ( n5681 & ~n18230 ) | ( n13708 & ~n18230 ) ;
  assign n18232 = n2860 | n14331 ;
  assign n18233 = n18232 ^ n12871 ^ 1'b0 ;
  assign n18234 = n6188 | n16517 ;
  assign n18235 = n395 & ~n14557 ;
  assign n18236 = n18235 ^ n2769 ^ 1'b0 ;
  assign n18237 = n18236 ^ n4918 ^ 1'b0 ;
  assign n18238 = ~n8803 & n18237 ;
  assign n18239 = n4593 & n18238 ;
  assign n18240 = n18239 ^ n14760 ^ 1'b0 ;
  assign n18241 = n11753 ^ x22 ^ 1'b0 ;
  assign n18242 = n12776 & ~n18241 ;
  assign n18243 = x175 & n18242 ;
  assign n18244 = n10314 & n18243 ;
  assign n18245 = n18244 ^ n2338 ^ 1'b0 ;
  assign n18246 = ( n2338 & n9394 ) | ( n2338 & n10861 ) | ( n9394 & n10861 ) ;
  assign n18247 = n9190 & n18246 ;
  assign n18248 = n13757 & n18247 ;
  assign n18249 = n5017 & ~n18248 ;
  assign n18250 = n18249 ^ n10116 ^ 1'b0 ;
  assign n18251 = n15364 ^ n13230 ^ 1'b0 ;
  assign n18252 = n12386 | n18251 ;
  assign n18253 = n4833 & ~n5108 ;
  assign n18254 = n5942 & ~n8539 ;
  assign n18255 = n10628 | n18254 ;
  assign n18256 = n18253 & ~n18255 ;
  assign n18259 = n6970 & n9331 ;
  assign n18260 = ~n17462 & n18259 ;
  assign n18257 = ~n9589 & n15653 ;
  assign n18258 = n17766 | n18257 ;
  assign n18261 = n18260 ^ n18258 ^ n6830 ;
  assign n18262 = n17453 ^ n2721 ^ 1'b0 ;
  assign n18263 = n5978 & n9020 ;
  assign n18264 = n18263 ^ n1403 ^ 1'b0 ;
  assign n18265 = n2285 | n4931 ;
  assign n18267 = ~n2787 & n2829 ;
  assign n18266 = ~n3761 & n8310 ;
  assign n18268 = n18267 ^ n18266 ^ 1'b0 ;
  assign n18269 = x121 & ~n2884 ;
  assign n18270 = n3176 & ~n18269 ;
  assign n18271 = n1136 | n9554 ;
  assign n18272 = n8067 & ~n18271 ;
  assign n18273 = n2420 | n18272 ;
  assign n18274 = n18270 & ~n18273 ;
  assign n18275 = n18274 ^ n4331 ^ 1'b0 ;
  assign n18276 = n9892 ^ n7385 ^ n5916 ;
  assign n18287 = n8170 ^ n4872 ^ 1'b0 ;
  assign n18288 = n5519 | n18287 ;
  assign n18281 = n7323 ^ n974 ^ 1'b0 ;
  assign n18282 = n4982 & ~n18281 ;
  assign n18283 = n13732 & ~n18282 ;
  assign n18284 = ~n7994 & n10001 ;
  assign n18285 = n18283 & ~n18284 ;
  assign n18286 = ~n2976 & n18285 ;
  assign n18277 = n13848 ^ n3084 ^ 1'b0 ;
  assign n18278 = n15390 & n18277 ;
  assign n18279 = n18278 ^ n5464 ^ 1'b0 ;
  assign n18280 = n12612 | n18279 ;
  assign n18289 = n18288 ^ n18286 ^ n18280 ;
  assign n18290 = n3161 & ~n14736 ;
  assign n18291 = n18144 ^ n3240 ^ 1'b0 ;
  assign n18292 = n7590 & ~n18291 ;
  assign n18293 = n4292 ^ n2883 ^ 1'b0 ;
  assign n18294 = n17391 ^ n11316 ^ 1'b0 ;
  assign n18295 = n18294 ^ n9585 ^ 1'b0 ;
  assign n18296 = n18293 & ~n18295 ;
  assign n18297 = n11141 | n16932 ;
  assign n18298 = ( n3434 & n4833 ) | ( n3434 & n5481 ) | ( n4833 & n5481 ) ;
  assign n18299 = n16045 | n18298 ;
  assign n18300 = ~n10311 & n18299 ;
  assign n18301 = n1413 | n15301 ;
  assign n18302 = n17270 & ~n18301 ;
  assign n18303 = n516 & ~n9792 ;
  assign n18304 = n14412 ^ n7200 ^ 1'b0 ;
  assign n18305 = n13952 ^ x97 ^ 1'b0 ;
  assign n18306 = n13826 ^ n8491 ^ 1'b0 ;
  assign n18307 = n18306 ^ n16244 ^ 1'b0 ;
  assign n18308 = ~n6400 & n12778 ;
  assign n18309 = n3658 & n6982 ;
  assign n18310 = n18309 ^ n14150 ^ 1'b0 ;
  assign n18311 = n18310 ^ n1255 ^ 1'b0 ;
  assign n18312 = ~n3583 & n18311 ;
  assign n18313 = x92 | n1188 ;
  assign n18314 = n3218 & n7006 ;
  assign n18315 = n18314 ^ n5295 ^ 1'b0 ;
  assign n18316 = n18313 | n18315 ;
  assign n18317 = x178 | n10856 ;
  assign n18318 = x175 & ~n8301 ;
  assign n18319 = n12269 & ~n14612 ;
  assign n18320 = n7547 ^ n1667 ^ 1'b0 ;
  assign n18321 = n8241 & n18320 ;
  assign n18322 = ~n9425 & n18321 ;
  assign n18324 = ( n1079 & n2285 ) | ( n1079 & ~n3937 ) | ( n2285 & ~n3937 ) ;
  assign n18323 = n1105 | n14379 ;
  assign n18325 = n18324 ^ n18323 ^ 1'b0 ;
  assign n18326 = n5355 | n18325 ;
  assign n18327 = n3384 & ~n7753 ;
  assign n18328 = ~n7306 & n7367 ;
  assign n18329 = n18328 ^ n1667 ^ 1'b0 ;
  assign n18330 = n2197 & ~n18329 ;
  assign n18331 = n12574 & n18330 ;
  assign n18332 = ~n18327 & n18331 ;
  assign n18333 = n2380 ^ n2076 ^ 1'b0 ;
  assign n18334 = n7462 | n18333 ;
  assign n18335 = n6408 | n18334 ;
  assign n18336 = n1804 & ~n4563 ;
  assign n18337 = n5993 | n18336 ;
  assign n18338 = n18337 ^ n1342 ^ 1'b0 ;
  assign n18339 = ( n674 & ~n3286 ) | ( n674 & n18338 ) | ( ~n3286 & n18338 ) ;
  assign n18340 = n2120 | n18339 ;
  assign n18341 = ~n1594 & n18340 ;
  assign n18342 = n18341 ^ n5328 ^ 1'b0 ;
  assign n18343 = n8235 ^ n7066 ^ 1'b0 ;
  assign n18344 = n5542 & ~n18343 ;
  assign n18345 = n4889 & n18344 ;
  assign n18346 = n18345 ^ n9330 ^ 1'b0 ;
  assign n18347 = n18346 ^ n3521 ^ 1'b0 ;
  assign n18348 = n4570 & ~n18347 ;
  assign n18349 = n1289 | n10488 ;
  assign n18350 = ~n6241 & n8433 ;
  assign n18351 = ( ~n626 & n1275 ) | ( ~n626 & n4936 ) | ( n1275 & n4936 ) ;
  assign n18352 = n9486 ^ n4845 ^ 1'b0 ;
  assign n18353 = n18351 & n18352 ;
  assign n18354 = ~n5061 & n7909 ;
  assign n18355 = n18354 ^ n15153 ^ 1'b0 ;
  assign n18356 = n13031 ^ n4081 ^ 1'b0 ;
  assign n18357 = n12846 & ~n18356 ;
  assign n18358 = n18355 & ~n18357 ;
  assign n18359 = n11127 | n13349 ;
  assign n18360 = n16952 & ~n18359 ;
  assign n18361 = n3112 | n9475 ;
  assign n18362 = n12808 | n16705 ;
  assign n18363 = n2311 & ~n4081 ;
  assign n18364 = n18363 ^ n13695 ^ 1'b0 ;
  assign n18366 = n1063 | n2064 ;
  assign n18367 = n18366 ^ n13162 ^ 1'b0 ;
  assign n18365 = n1807 & n9700 ;
  assign n18368 = n18367 ^ n18365 ^ 1'b0 ;
  assign n18369 = n15441 & n18368 ;
  assign n18370 = n11587 & n12175 ;
  assign n18371 = n2080 & ~n10911 ;
  assign n18372 = n1298 & n2804 ;
  assign n18373 = ~n18371 & n18372 ;
  assign n18375 = n14119 ^ n13945 ^ 1'b0 ;
  assign n18374 = n1233 | n14667 ;
  assign n18376 = n18375 ^ n18374 ^ 1'b0 ;
  assign n18377 = n18376 ^ n13585 ^ 1'b0 ;
  assign n18378 = n2241 & ~n18377 ;
  assign n18379 = ~n18373 & n18378 ;
  assign n18380 = ~n3371 & n11050 ;
  assign n18381 = n4339 ^ n2390 ^ n363 ;
  assign n18382 = ~n18380 & n18381 ;
  assign n18383 = n1518 & ~n5489 ;
  assign n18384 = n18383 ^ x37 ^ 1'b0 ;
  assign n18385 = ( n3806 & n4413 ) | ( n3806 & n10222 ) | ( n4413 & n10222 ) ;
  assign n18386 = n18385 ^ n14476 ^ n10404 ;
  assign n18387 = ( ~x187 & n3808 ) | ( ~x187 & n13201 ) | ( n3808 & n13201 ) ;
  assign n18388 = n18387 ^ n6572 ^ 1'b0 ;
  assign n18389 = n11427 | n18388 ;
  assign n18390 = n18389 ^ n3797 ^ 1'b0 ;
  assign n18391 = n3555 & n18390 ;
  assign n18392 = n5283 & n18391 ;
  assign n18393 = n18392 ^ n16962 ^ 1'b0 ;
  assign n18394 = n14229 & n18393 ;
  assign n18395 = n12203 ^ n6621 ^ 1'b0 ;
  assign n18396 = x227 & n18395 ;
  assign n18397 = n18396 ^ n13153 ^ 1'b0 ;
  assign n18398 = n4253 & n18397 ;
  assign n18399 = n9437 | n18398 ;
  assign n18400 = ( n5248 & n6127 ) | ( n5248 & ~n18399 ) | ( n6127 & ~n18399 ) ;
  assign n18401 = ~n2389 & n14387 ;
  assign n18402 = x51 | n8350 ;
  assign n18403 = n411 & n18402 ;
  assign n18404 = ~n8220 & n10183 ;
  assign n18405 = n18404 ^ n16996 ^ n15951 ;
  assign n18406 = ~x170 & n1102 ;
  assign n18407 = n7013 & n10717 ;
  assign n18408 = n18407 ^ n3009 ^ 1'b0 ;
  assign n18409 = n18406 | n18408 ;
  assign n18410 = n9271 ^ n7834 ^ n7466 ;
  assign n18411 = n4462 | n11621 ;
  assign n18412 = ~n5813 & n18411 ;
  assign n18413 = n18410 & n18412 ;
  assign n18414 = n7362 | n7406 ;
  assign n18415 = n4784 | n7584 ;
  assign n18416 = ~n15768 & n18415 ;
  assign n18417 = n18392 ^ n16508 ^ n14247 ;
  assign n18418 = n6355 & n8419 ;
  assign n18419 = n1409 | n4824 ;
  assign n18420 = n685 & ~n18419 ;
  assign n18421 = n18420 ^ n17185 ^ 1'b0 ;
  assign n18422 = n18418 & n18421 ;
  assign n18423 = ~n2941 & n18422 ;
  assign n18424 = n17120 ^ n7881 ^ n6023 ;
  assign n18425 = n18424 ^ n14251 ^ n5022 ;
  assign n18426 = n5637 | n18425 ;
  assign n18427 = n1926 ^ n1655 ^ 1'b0 ;
  assign n18428 = n18427 ^ n16090 ^ 1'b0 ;
  assign n18429 = ~n6722 & n18428 ;
  assign n18430 = ( n6529 & n8998 ) | ( n6529 & n18429 ) | ( n8998 & n18429 ) ;
  assign n18433 = n431 | n4148 ;
  assign n18434 = n8438 & ~n18433 ;
  assign n18431 = ~n6548 & n13404 ;
  assign n18432 = n18431 ^ n7399 ^ 1'b0 ;
  assign n18435 = n18434 ^ n18432 ^ n15659 ;
  assign n18436 = n15183 ^ n14817 ^ n7354 ;
  assign n18437 = n18043 ^ n9017 ^ 1'b0 ;
  assign n18438 = n2289 | n7074 ;
  assign n18439 = n11663 ^ n379 ^ 1'b0 ;
  assign n18440 = ( n2108 & n10846 ) | ( n2108 & n15014 ) | ( n10846 & n15014 ) ;
  assign n18441 = ( ~n6111 & n11171 ) | ( ~n6111 & n18440 ) | ( n11171 & n18440 ) ;
  assign n18442 = ( n4517 & n5478 ) | ( n4517 & n5884 ) | ( n5478 & n5884 ) ;
  assign n18443 = n17822 & ~n18442 ;
  assign n18444 = n18443 ^ n13194 ^ 1'b0 ;
  assign n18445 = n8803 ^ n6813 ^ 1'b0 ;
  assign n18446 = n16073 & n16290 ;
  assign n18447 = n18446 ^ n14652 ^ 1'b0 ;
  assign n18448 = n3476 ^ n1210 ^ 1'b0 ;
  assign n18449 = n301 | n18448 ;
  assign n18450 = n892 | n18449 ;
  assign n18451 = n18450 ^ n2015 ^ 1'b0 ;
  assign n18452 = n18451 ^ n2057 ^ 1'b0 ;
  assign n18453 = n18452 ^ n4102 ^ 1'b0 ;
  assign n18454 = ~n3901 & n18453 ;
  assign n18455 = n18454 ^ n7440 ^ 1'b0 ;
  assign n18456 = ~n14264 & n18455 ;
  assign n18457 = n18456 ^ n7975 ^ 1'b0 ;
  assign n18458 = n8763 ^ n7156 ^ 1'b0 ;
  assign n18459 = n6232 | n18458 ;
  assign n18460 = n18459 ^ n4734 ^ 1'b0 ;
  assign n18461 = n960 | n3534 ;
  assign n18462 = n18461 ^ n12087 ^ n4960 ;
  assign n18463 = n18462 ^ n15768 ^ 1'b0 ;
  assign n18464 = n14551 ^ n6445 ^ n2176 ;
  assign n18465 = n10923 ^ n8176 ^ n5614 ;
  assign n18466 = n18465 ^ n4479 ^ 1'b0 ;
  assign n18467 = n16299 | n18466 ;
  assign n18468 = n9581 ^ n9375 ^ 1'b0 ;
  assign n18469 = n18468 ^ n3023 ^ 1'b0 ;
  assign n18470 = ~n15726 & n18469 ;
  assign n18472 = n6522 & ~n7194 ;
  assign n18473 = n4624 & n18472 ;
  assign n18474 = ~n7674 & n10253 ;
  assign n18475 = n18473 & n18474 ;
  assign n18471 = ~n4157 & n16595 ;
  assign n18476 = n18475 ^ n18471 ^ 1'b0 ;
  assign n18485 = n8167 ^ n1147 ^ 1'b0 ;
  assign n18477 = n1071 & n2402 ;
  assign n18478 = n652 & n2836 ;
  assign n18479 = n714 & n18478 ;
  assign n18480 = n4436 & ~n18479 ;
  assign n18481 = ~n647 & n18480 ;
  assign n18482 = ~n5235 & n18481 ;
  assign n18483 = ~n18477 & n18482 ;
  assign n18484 = n13614 & ~n18483 ;
  assign n18486 = n18485 ^ n18484 ^ 1'b0 ;
  assign n18487 = ( n4182 & n7220 ) | ( n4182 & ~n11425 ) | ( n7220 & ~n11425 ) ;
  assign n18488 = n7978 & n16431 ;
  assign n18489 = n8080 & ~n18488 ;
  assign n18490 = ( n14483 & ~n16335 ) | ( n14483 & n17140 ) | ( ~n16335 & n17140 ) ;
  assign n18491 = n9680 & ~n15941 ;
  assign n18492 = n18491 ^ n11063 ^ 1'b0 ;
  assign n18493 = n2598 & n2601 ;
  assign n18494 = ~n18492 & n18493 ;
  assign n18495 = n11663 ^ n8314 ^ n5420 ;
  assign n18496 = ~n8841 & n18495 ;
  assign n18497 = n1060 & ~n10749 ;
  assign n18498 = n18497 ^ n10911 ^ 1'b0 ;
  assign n18499 = n18498 ^ n16739 ^ n12994 ;
  assign n18500 = n7570 ^ n2002 ^ 1'b0 ;
  assign n18501 = n15363 | n18500 ;
  assign n18502 = n1916 | n15797 ;
  assign n18503 = n14848 | n18502 ;
  assign n18504 = n18503 ^ n17001 ^ x60 ;
  assign n18505 = n12566 ^ n10879 ^ 1'b0 ;
  assign n18506 = ( ~n8944 & n10414 ) | ( ~n8944 & n10662 ) | ( n10414 & n10662 ) ;
  assign n18507 = ( x218 & n2965 ) | ( x218 & n5209 ) | ( n2965 & n5209 ) ;
  assign n18508 = ~n4976 & n18507 ;
  assign n18509 = ( ~n4924 & n8215 ) | ( ~n4924 & n10109 ) | ( n8215 & n10109 ) ;
  assign n18510 = n7831 | n18509 ;
  assign n18511 = n18508 | n18510 ;
  assign n18512 = ( n3088 & ~n5195 ) | ( n3088 & n8058 ) | ( ~n5195 & n8058 ) ;
  assign n18513 = n2806 ^ x215 ^ 1'b0 ;
  assign n18514 = n3376 | n18513 ;
  assign n18515 = n18514 ^ n6400 ^ 1'b0 ;
  assign n18516 = ~n8438 & n8511 ;
  assign n18517 = ~n14538 & n18516 ;
  assign n18519 = n9653 ^ n2588 ^ 1'b0 ;
  assign n18520 = ~n6821 & n18519 ;
  assign n18521 = ( n4140 & ~n5519 ) | ( n4140 & n6373 ) | ( ~n5519 & n6373 ) ;
  assign n18522 = n18521 ^ n404 ^ 1'b0 ;
  assign n18523 = n18520 & n18522 ;
  assign n18524 = n18087 | n18523 ;
  assign n18518 = n3023 ^ n847 ^ 1'b0 ;
  assign n18525 = n18524 ^ n18518 ^ n2654 ;
  assign n18526 = n3287 & ~n11564 ;
  assign n18527 = n3526 ^ n1592 ^ 1'b0 ;
  assign n18528 = n3955 & n18527 ;
  assign n18529 = n3995 & ~n6053 ;
  assign n18530 = n13772 & n18529 ;
  assign n18531 = n18530 ^ n7777 ^ 1'b0 ;
  assign n18532 = n13635 ^ n5129 ^ 1'b0 ;
  assign n18533 = n18531 | n18532 ;
  assign n18534 = ~n4553 & n13280 ;
  assign n18535 = n11267 ^ n11007 ^ 1'b0 ;
  assign n18536 = n9902 & ~n18535 ;
  assign n18537 = n9726 ^ n9139 ^ 1'b0 ;
  assign n18538 = n5916 | n18537 ;
  assign n18539 = n10736 ^ n8029 ^ 1'b0 ;
  assign n18540 = n1979 | n9253 ;
  assign n18541 = n6514 | n18540 ;
  assign n18542 = n7126 & ~n18541 ;
  assign n18543 = ~n2168 & n17320 ;
  assign n18544 = n18543 ^ n5776 ^ 1'b0 ;
  assign n18545 = n5446 ^ n5060 ^ n2399 ;
  assign n18546 = n18544 & n18545 ;
  assign n18547 = ~n10990 & n18546 ;
  assign n18548 = n2023 & ~n12176 ;
  assign n18549 = n18548 ^ n9296 ^ 1'b0 ;
  assign n18550 = n18549 ^ n2380 ^ 1'b0 ;
  assign n18551 = ~n18547 & n18550 ;
  assign n18552 = n1550 & n18551 ;
  assign n18553 = n18552 ^ n12672 ^ 1'b0 ;
  assign n18554 = n18553 ^ n3053 ^ 1'b0 ;
  assign n18555 = n1440 & n18554 ;
  assign n18556 = ~n511 & n6103 ;
  assign n18557 = ( n5869 & n12600 ) | ( n5869 & n18556 ) | ( n12600 & n18556 ) ;
  assign n18562 = n6129 | n6241 ;
  assign n18558 = n2893 & n12827 ;
  assign n18559 = n5404 & n18558 ;
  assign n18560 = n13772 & ~n18559 ;
  assign n18561 = n18560 ^ n5716 ^ n1489 ;
  assign n18563 = n18562 ^ n18561 ^ n9221 ;
  assign n18564 = n390 | n1199 ;
  assign n18565 = n18564 ^ n1804 ^ 1'b0 ;
  assign n18566 = x17 | n3844 ;
  assign n18567 = n1795 | n18566 ;
  assign n18568 = ( n17398 & n18565 ) | ( n17398 & ~n18567 ) | ( n18565 & ~n18567 ) ;
  assign n18569 = n18213 ^ n12215 ^ n9648 ;
  assign n18570 = ~n6801 & n10164 ;
  assign n18571 = n17951 ^ n1068 ^ 1'b0 ;
  assign n18572 = n599 & n18571 ;
  assign n18573 = n15193 ^ n14784 ^ 1'b0 ;
  assign n18575 = ( n1072 & n3708 ) | ( n1072 & n8603 ) | ( n3708 & n8603 ) ;
  assign n18574 = n5820 & n14212 ;
  assign n18576 = n18575 ^ n18574 ^ 1'b0 ;
  assign n18577 = n18573 & n18576 ;
  assign n18578 = n1334 & ~n6667 ;
  assign n18579 = n18578 ^ n15970 ^ 1'b0 ;
  assign n18580 = n4937 ^ n3868 ^ 1'b0 ;
  assign n18581 = n18579 & ~n18580 ;
  assign n18585 = n1500 | n3259 ;
  assign n18582 = n2684 & ~n8729 ;
  assign n18583 = n1423 & n18582 ;
  assign n18584 = n1887 & ~n18583 ;
  assign n18586 = n18585 ^ n18584 ^ 1'b0 ;
  assign n18589 = n780 & ~n8964 ;
  assign n18587 = n11149 ^ n8200 ^ n1991 ;
  assign n18588 = ~n11274 & n18587 ;
  assign n18590 = n18589 ^ n18588 ^ n12985 ;
  assign n18591 = ( ~n861 & n2512 ) | ( ~n861 & n6887 ) | ( n2512 & n6887 ) ;
  assign n18592 = n18182 ^ n11227 ^ 1'b0 ;
  assign n18593 = n3723 & ~n18592 ;
  assign n18594 = n7223 | n8632 ;
  assign n18597 = n4160 | n6016 ;
  assign n18595 = x135 & n18387 ;
  assign n18596 = ~n9244 & n18595 ;
  assign n18598 = n18597 ^ n18596 ^ 1'b0 ;
  assign n18599 = n18598 ^ n6352 ^ x102 ;
  assign n18600 = n12624 ^ n4263 ^ n889 ;
  assign n18601 = n18600 ^ n13148 ^ 1'b0 ;
  assign n18602 = n3014 & ~n18601 ;
  assign n18603 = ~n16723 & n18602 ;
  assign n18604 = ( n6540 & ~n13746 ) | ( n6540 & n18603 ) | ( ~n13746 & n18603 ) ;
  assign n18605 = n18604 ^ n7913 ^ 1'b0 ;
  assign n18606 = n16335 ^ x11 ^ 1'b0 ;
  assign n18607 = ~n401 & n18606 ;
  assign n18608 = n9969 & n18607 ;
  assign n18610 = ( ~n7452 & n9367 ) | ( ~n7452 & n13527 ) | ( n9367 & n13527 ) ;
  assign n18611 = n18610 ^ n3164 ^ 1'b0 ;
  assign n18609 = n9465 ^ n5634 ^ 1'b0 ;
  assign n18612 = n18611 ^ n18609 ^ n8075 ;
  assign n18613 = n2024 ^ n612 ^ 1'b0 ;
  assign n18614 = n3382 | n4860 ;
  assign n18615 = x136 | n18614 ;
  assign n18616 = n7155 ^ n1425 ^ 1'b0 ;
  assign n18617 = n11246 | n18616 ;
  assign n18618 = n18615 | n18617 ;
  assign n18619 = n18618 ^ n9029 ^ 1'b0 ;
  assign n18620 = n9890 ^ n5188 ^ 1'b0 ;
  assign n18621 = n18620 ^ n6179 ^ 1'b0 ;
  assign n18623 = n18346 ^ n5599 ^ n1744 ;
  assign n18622 = n6153 ^ n4010 ^ 1'b0 ;
  assign n18624 = n18623 ^ n18622 ^ 1'b0 ;
  assign n18625 = n14268 ^ n1798 ^ 1'b0 ;
  assign n18626 = n18624 & ~n18625 ;
  assign n18627 = n7021 ^ n3116 ^ 1'b0 ;
  assign n18628 = n18545 ^ n11770 ^ n7706 ;
  assign n18629 = n13495 ^ n6973 ^ 1'b0 ;
  assign n18630 = n3800 ^ n456 ^ 1'b0 ;
  assign n18631 = ~n18629 & n18630 ;
  assign n18632 = n2972 | n13400 ;
  assign n18636 = n12280 ^ n4679 ^ x13 ;
  assign n18633 = n7101 & ~n12697 ;
  assign n18634 = n18633 ^ n9866 ^ 1'b0 ;
  assign n18635 = ~n10383 & n18634 ;
  assign n18637 = n18636 ^ n18635 ^ 1'b0 ;
  assign n18638 = n18637 ^ n13394 ^ 1'b0 ;
  assign n18639 = ( n13204 & n14587 ) | ( n13204 & n18638 ) | ( n14587 & n18638 ) ;
  assign n18641 = n2437 & n15646 ;
  assign n18642 = n1073 & n18641 ;
  assign n18640 = n6005 & n8287 ;
  assign n18643 = n18642 ^ n18640 ^ 1'b0 ;
  assign n18644 = n6766 & ~n10306 ;
  assign n18645 = n14388 ^ n13544 ^ n8466 ;
  assign n18646 = ~n2649 & n17500 ;
  assign n18647 = ~n18645 & n18646 ;
  assign n18648 = ( n4510 & n8844 ) | ( n4510 & ~n18647 ) | ( n8844 & ~n18647 ) ;
  assign n18649 = n18451 ^ n12808 ^ n11312 ;
  assign n18650 = ~n4953 & n12140 ;
  assign n18651 = n538 & n6294 ;
  assign n18652 = n8319 & n18651 ;
  assign n18653 = n9087 ^ n6726 ^ 1'b0 ;
  assign n18654 = n11975 ^ n5229 ^ 1'b0 ;
  assign n18655 = n18653 | n18654 ;
  assign n18656 = n6361 ^ n2008 ^ n1071 ;
  assign n18657 = n9146 ^ n2203 ^ 1'b0 ;
  assign n18658 = ( n13418 & n15832 ) | ( n13418 & ~n18657 ) | ( n15832 & ~n18657 ) ;
  assign n18659 = ~n4019 & n7521 ;
  assign n18660 = n1304 & n18659 ;
  assign n18662 = n16465 ^ n7130 ^ 1'b0 ;
  assign n18663 = ~n3504 & n18662 ;
  assign n18664 = n18663 ^ n10397 ^ 1'b0 ;
  assign n18665 = n8616 | n18664 ;
  assign n18661 = n5663 ^ n319 ^ 1'b0 ;
  assign n18666 = n18665 ^ n18661 ^ 1'b0 ;
  assign n18667 = n14105 ^ n7185 ^ 1'b0 ;
  assign n18668 = n18667 ^ n14280 ^ 1'b0 ;
  assign n18669 = ~n1781 & n6091 ;
  assign n18670 = ~n7213 & n18669 ;
  assign n18671 = n18668 | n18670 ;
  assign n18672 = n1813 & n8785 ;
  assign n18673 = n4529 & n18672 ;
  assign n18674 = ( n723 & ~n4016 ) | ( n723 & n18673 ) | ( ~n4016 & n18673 ) ;
  assign n18675 = n11882 ^ n6365 ^ n6001 ;
  assign n18676 = n18675 ^ n4540 ^ 1'b0 ;
  assign n18677 = n12696 | n18676 ;
  assign n18678 = n18677 ^ x41 ^ 1'b0 ;
  assign n18679 = n9544 & ~n16407 ;
  assign n18680 = n997 & ~n16998 ;
  assign n18681 = n8619 ^ n4041 ^ 1'b0 ;
  assign n18682 = n4036 & ~n18681 ;
  assign n18689 = n15186 ^ n10063 ^ 1'b0 ;
  assign n18690 = n9020 & n18689 ;
  assign n18685 = n8914 | n18381 ;
  assign n18686 = n2486 | n18685 ;
  assign n18684 = n13749 | n15988 ;
  assign n18687 = n18686 ^ n18684 ^ 1'b0 ;
  assign n18683 = n10209 ^ x15 ^ 1'b0 ;
  assign n18688 = n18687 ^ n18683 ^ n6986 ;
  assign n18691 = n18690 ^ n18688 ^ n17866 ;
  assign n18692 = n2390 | n11137 ;
  assign n18693 = n17968 & ~n18692 ;
  assign n18694 = ( ~n2541 & n14117 ) | ( ~n2541 & n17247 ) | ( n14117 & n17247 ) ;
  assign n18695 = ~n6585 & n11080 ;
  assign n18696 = n15489 ^ n13355 ^ 1'b0 ;
  assign n18697 = n13571 ^ n9463 ^ 1'b0 ;
  assign n18698 = n2915 | n18697 ;
  assign n18699 = n15697 | n18698 ;
  assign n18700 = n3554 & n9945 ;
  assign n18701 = n18700 ^ n5805 ^ 1'b0 ;
  assign n18702 = ~n1360 & n18701 ;
  assign n18703 = n18702 ^ n9995 ^ 1'b0 ;
  assign n18704 = n1055 | n1595 ;
  assign n18705 = n18703 | n18704 ;
  assign n18706 = ( n8845 & n11583 ) | ( n8845 & ~n13070 ) | ( n11583 & ~n13070 ) ;
  assign n18707 = n14795 ^ n2422 ^ 1'b0 ;
  assign n18708 = ~n4055 & n16190 ;
  assign n18709 = n7787 & n8293 ;
  assign n18710 = n18709 ^ n10718 ^ 1'b0 ;
  assign n18711 = ( n2762 & ~n10525 ) | ( n2762 & n11595 ) | ( ~n10525 & n11595 ) ;
  assign n18712 = ~n17104 & n18711 ;
  assign n18713 = ~n6607 & n15788 ;
  assign n18714 = n18713 ^ n11753 ^ n1113 ;
  assign n18715 = n5713 ^ n4821 ^ 1'b0 ;
  assign n18716 = n18715 ^ n7058 ^ 1'b0 ;
  assign n18720 = n5720 ^ n5359 ^ 1'b0 ;
  assign n18717 = ~n1937 & n15080 ;
  assign n18718 = n3363 & n18717 ;
  assign n18719 = n7130 & ~n18718 ;
  assign n18721 = n18720 ^ n18719 ^ 1'b0 ;
  assign n18722 = ( n9322 & n10035 ) | ( n9322 & n13513 ) | ( n10035 & n13513 ) ;
  assign n18723 = n11857 | n16810 ;
  assign n18725 = n8777 ^ n4252 ^ 1'b0 ;
  assign n18724 = n995 ^ x227 ^ 1'b0 ;
  assign n18726 = n18725 ^ n18724 ^ 1'b0 ;
  assign n18727 = n4417 ^ n2357 ^ 1'b0 ;
  assign n18728 = n8219 & ~n18727 ;
  assign n18729 = n7942 ^ n3749 ^ n2231 ;
  assign n18730 = ~n10155 & n18729 ;
  assign n18731 = ~n1256 & n18730 ;
  assign n18732 = ( n11252 & ~n18728 ) | ( n11252 & n18731 ) | ( ~n18728 & n18731 ) ;
  assign n18733 = ~n9413 & n18732 ;
  assign n18734 = ( ~n365 & n6279 ) | ( ~n365 & n17948 ) | ( n6279 & n17948 ) ;
  assign n18735 = n6406 ^ n4986 ^ 1'b0 ;
  assign n18736 = n11850 ^ n5122 ^ 1'b0 ;
  assign n18737 = n16495 & ~n18736 ;
  assign n18738 = n18737 ^ n2216 ^ 1'b0 ;
  assign n18739 = n14280 & ~n18738 ;
  assign n18740 = n3431 ^ n2728 ^ 1'b0 ;
  assign n18741 = ~n16570 & n18740 ;
  assign n18742 = n8787 ^ n5133 ^ 1'b0 ;
  assign n18743 = n6841 ^ n585 ^ 1'b0 ;
  assign n18744 = n18742 & ~n18743 ;
  assign n18745 = n18744 ^ n17586 ^ 1'b0 ;
  assign n18746 = ~n4860 & n18745 ;
  assign n18747 = n13083 ^ n5021 ^ 1'b0 ;
  assign n18748 = n3267 & n18747 ;
  assign n18749 = n18748 ^ n5124 ^ n3646 ;
  assign n18750 = n18749 ^ n15712 ^ 1'b0 ;
  assign n18751 = ~n7036 & n9208 ;
  assign n18752 = n18751 ^ n5892 ^ 1'b0 ;
  assign n18753 = n8925 & n14322 ;
  assign n18754 = n7360 ^ n1853 ^ 1'b0 ;
  assign n18755 = n12057 | n18507 ;
  assign n18757 = ( ~n817 & n1256 ) | ( ~n817 & n10816 ) | ( n1256 & n10816 ) ;
  assign n18756 = n557 | n10961 ;
  assign n18758 = n18757 ^ n18756 ^ 1'b0 ;
  assign n18759 = n18758 ^ n14117 ^ 1'b0 ;
  assign n18760 = n12805 ^ n6590 ^ 1'b0 ;
  assign n18761 = ~n1475 & n18760 ;
  assign n18762 = n18761 ^ n5701 ^ 1'b0 ;
  assign n18763 = n18762 ^ n3150 ^ 1'b0 ;
  assign n18764 = ~n11689 & n18763 ;
  assign n18765 = n11004 ^ n3030 ^ n1605 ;
  assign n18766 = n1270 & n18765 ;
  assign n18767 = n18766 ^ n13380 ^ 1'b0 ;
  assign n18768 = n18767 ^ n17000 ^ 1'b0 ;
  assign n18769 = n5329 ^ n1894 ^ 1'b0 ;
  assign n18770 = n7087 & ~n8503 ;
  assign n18771 = n2188 & ~n8587 ;
  assign n18772 = n18771 ^ n14028 ^ 1'b0 ;
  assign n18773 = n2815 ^ x144 ^ 1'b0 ;
  assign n18774 = n18773 ^ n1947 ^ 1'b0 ;
  assign n18775 = n3524 & n7172 ;
  assign n18776 = n4161 & ~n18775 ;
  assign n18777 = n7458 & n18776 ;
  assign n18778 = n15670 ^ n1033 ^ n718 ;
  assign n18779 = ( n11136 & n11906 ) | ( n11136 & ~n13950 ) | ( n11906 & ~n13950 ) ;
  assign n18780 = ( ~n449 & n7444 ) | ( ~n449 & n15294 ) | ( n7444 & n15294 ) ;
  assign n18781 = n1097 & n4722 ;
  assign n18782 = n8017 & ~n8919 ;
  assign n18783 = n18782 ^ n10039 ^ 1'b0 ;
  assign n18784 = n18390 ^ n15899 ^ n5850 ;
  assign n18785 = n18783 & ~n18784 ;
  assign n18786 = n18785 ^ n4809 ^ 1'b0 ;
  assign n18787 = n18781 & n18786 ;
  assign n18788 = ~n13550 & n18787 ;
  assign n18789 = ( n1177 & n18780 ) | ( n1177 & ~n18788 ) | ( n18780 & ~n18788 ) ;
  assign n18790 = n18789 ^ n13188 ^ n10552 ;
  assign n18791 = n574 & n1512 ;
  assign n18792 = n13774 | n18791 ;
  assign n18793 = n18792 ^ n13659 ^ 1'b0 ;
  assign n18794 = n16821 ^ n1287 ^ n944 ;
  assign n18795 = n18793 & ~n18794 ;
  assign n18796 = n3362 & n9545 ;
  assign n18797 = ( n4305 & ~n12004 ) | ( n4305 & n18796 ) | ( ~n12004 & n18796 ) ;
  assign n18798 = n842 & n9952 ;
  assign n18799 = n7362 & n18798 ;
  assign n18800 = ~n18797 & n18799 ;
  assign n18801 = n7637 & ~n15508 ;
  assign n18802 = ( n1055 & n1285 ) | ( n1055 & ~n1735 ) | ( n1285 & ~n1735 ) ;
  assign n18803 = n18802 ^ n6451 ^ 1'b0 ;
  assign n18804 = n18803 ^ n5071 ^ 1'b0 ;
  assign n18805 = n18804 ^ n2523 ^ 1'b0 ;
  assign n18806 = n12414 ^ n3274 ^ 1'b0 ;
  assign n18807 = n12321 & ~n18806 ;
  assign n18808 = n18805 & n18807 ;
  assign n18809 = n9447 ^ n4881 ^ 1'b0 ;
  assign n18810 = n10829 & n18809 ;
  assign n18817 = x131 & n1297 ;
  assign n18815 = n12886 ^ n3060 ^ 1'b0 ;
  assign n18816 = n9559 & ~n18815 ;
  assign n18812 = n14914 ^ n5597 ^ 1'b0 ;
  assign n18813 = n12546 & n18812 ;
  assign n18811 = n1491 & n11242 ;
  assign n18814 = n18813 ^ n18811 ^ 1'b0 ;
  assign n18818 = n18817 ^ n18816 ^ n18814 ;
  assign n18819 = n8245 & n11540 ;
  assign n18820 = ( ~n2384 & n10962 ) | ( ~n2384 & n18819 ) | ( n10962 & n18819 ) ;
  assign n18822 = n6693 & ~n7934 ;
  assign n18823 = ~n12669 & n18822 ;
  assign n18821 = n5185 | n6822 ;
  assign n18824 = n18823 ^ n18821 ^ 1'b0 ;
  assign n18825 = n14106 ^ n9416 ^ 1'b0 ;
  assign n18826 = n4127 & n4496 ;
  assign n18827 = n1132 & n18826 ;
  assign n18828 = n6611 & n18827 ;
  assign n18831 = ( ~n1213 & n1551 ) | ( ~n1213 & n11376 ) | ( n1551 & n11376 ) ;
  assign n18829 = ~n559 & n7804 ;
  assign n18830 = n6466 & ~n18829 ;
  assign n18832 = n18831 ^ n18830 ^ 1'b0 ;
  assign n18833 = n6145 | n18832 ;
  assign n18834 = n5127 & ~n9204 ;
  assign n18839 = n4872 & ~n6708 ;
  assign n18840 = n18839 ^ n7952 ^ 1'b0 ;
  assign n18841 = n6535 & ~n18840 ;
  assign n18835 = n12295 ^ n4283 ^ 1'b0 ;
  assign n18836 = ~n6205 & n16914 ;
  assign n18837 = ~n5947 & n18836 ;
  assign n18838 = n18835 | n18837 ;
  assign n18842 = n18841 ^ n18838 ^ 1'b0 ;
  assign n18843 = n2178 & ~n7888 ;
  assign n18844 = n18843 ^ n8019 ^ 1'b0 ;
  assign n18845 = n7225 ^ n2441 ^ 1'b0 ;
  assign n18846 = ~n18844 & n18845 ;
  assign n18847 = ( ~n6539 & n6553 ) | ( ~n6539 & n7074 ) | ( n6553 & n7074 ) ;
  assign n18848 = n18846 & n18847 ;
  assign n18849 = n490 & ~n12282 ;
  assign n18850 = n18849 ^ n15865 ^ 1'b0 ;
  assign n18851 = n9632 ^ n5914 ^ 1'b0 ;
  assign n18852 = n14382 & n18851 ;
  assign n18853 = n1321 & n18852 ;
  assign n18854 = ( x100 & ~n2815 ) | ( x100 & n3979 ) | ( ~n2815 & n3979 ) ;
  assign n18855 = n11155 ^ n7382 ^ 1'b0 ;
  assign n18856 = n18854 & n18855 ;
  assign n18857 = ~n13234 & n18856 ;
  assign n18858 = n14465 ^ n5244 ^ 1'b0 ;
  assign n18859 = n14617 ^ n1228 ^ 1'b0 ;
  assign n18860 = n5591 & n18859 ;
  assign n18861 = n17792 ^ n5054 ^ 1'b0 ;
  assign n18862 = n14551 & n16470 ;
  assign n18863 = n12342 & ~n14818 ;
  assign n18864 = n7567 ^ n2243 ^ 1'b0 ;
  assign n18865 = ~n3530 & n7621 ;
  assign n18866 = n15240 ^ n11467 ^ 1'b0 ;
  assign n18867 = n2441 ^ n1308 ^ 1'b0 ;
  assign n18868 = n16342 & n18867 ;
  assign n18869 = n9534 & ~n18868 ;
  assign n18870 = n11722 ^ n1421 ^ 1'b0 ;
  assign n18871 = n18870 ^ n3551 ^ 1'b0 ;
  assign n18872 = x251 & n7019 ;
  assign n18873 = n10475 ^ n5478 ^ 1'b0 ;
  assign n18874 = n18872 & n18873 ;
  assign n18875 = n16122 | n18874 ;
  assign n18876 = n18875 ^ n11483 ^ 1'b0 ;
  assign n18877 = n10788 ^ n814 ^ 1'b0 ;
  assign n18878 = n5474 & ~n18877 ;
  assign n18879 = n723 & n1042 ;
  assign n18880 = ~n2991 & n11248 ;
  assign n18881 = ~n5810 & n18880 ;
  assign n18882 = ( n4858 & n18879 ) | ( n4858 & ~n18881 ) | ( n18879 & ~n18881 ) ;
  assign n18883 = n18716 ^ n9374 ^ n2063 ;
  assign n18884 = ( n3531 & n6589 ) | ( n3531 & ~n16992 ) | ( n6589 & ~n16992 ) ;
  assign n18885 = n5056 & n18884 ;
  assign n18886 = n18885 ^ n536 ^ 1'b0 ;
  assign n18887 = n5538 ^ n2484 ^ 1'b0 ;
  assign n18888 = n14783 & ~n18887 ;
  assign n18889 = n8318 ^ n3292 ^ 1'b0 ;
  assign n18890 = n6196 & n18889 ;
  assign n18891 = n18890 ^ n875 ^ 1'b0 ;
  assign n18892 = n7112 ^ n2365 ^ 1'b0 ;
  assign n18893 = n781 | n18892 ;
  assign n18894 = n18893 ^ n10423 ^ n4096 ;
  assign n18895 = n18894 ^ n18418 ^ n16482 ;
  assign n18896 = n18891 & ~n18895 ;
  assign n18898 = n10992 ^ n10097 ^ 1'b0 ;
  assign n18897 = ~n6632 & n16966 ;
  assign n18899 = n18898 ^ n18897 ^ 1'b0 ;
  assign n18900 = n3081 & ~n6967 ;
  assign n18901 = n18900 ^ n1504 ^ 1'b0 ;
  assign n18902 = n18901 ^ n12413 ^ n7892 ;
  assign n18903 = n2925 & ~n3647 ;
  assign n18904 = n16470 ^ n1283 ^ 1'b0 ;
  assign n18905 = n18903 & n18904 ;
  assign n18906 = n4890 | n15300 ;
  assign n18907 = ~n2146 & n7653 ;
  assign n18908 = n18907 ^ n3445 ^ 1'b0 ;
  assign n18910 = ( n4590 & n7145 ) | ( n4590 & ~n7632 ) | ( n7145 & ~n7632 ) ;
  assign n18911 = n1601 & n18910 ;
  assign n18909 = n668 & ~n10560 ;
  assign n18912 = n18911 ^ n18909 ^ n10298 ;
  assign n18913 = ~n1437 & n18912 ;
  assign n18914 = n16428 & n18913 ;
  assign n18920 = n4212 & n8474 ;
  assign n18915 = ( n3019 & n6005 ) | ( n3019 & n6837 ) | ( n6005 & n6837 ) ;
  assign n18916 = n657 & n7004 ;
  assign n18917 = n18915 & n18916 ;
  assign n18918 = n12117 | n18917 ;
  assign n18919 = n5865 & n18918 ;
  assign n18921 = n18920 ^ n18919 ^ 1'b0 ;
  assign n18922 = n6461 ^ n4815 ^ 1'b0 ;
  assign n18923 = n1286 & n18922 ;
  assign n18924 = n8316 & ~n8656 ;
  assign n18925 = n16798 ^ n14110 ^ 1'b0 ;
  assign n18926 = n6529 ^ n1468 ^ n471 ;
  assign n18927 = n7464 | n18926 ;
  assign n18928 = n1134 | n12624 ;
  assign n18929 = x170 | n18928 ;
  assign n18930 = n18929 ^ n11138 ^ n2746 ;
  assign n18931 = n18930 ^ n13069 ^ 1'b0 ;
  assign n18932 = ~n5006 & n18931 ;
  assign n18933 = n6646 & ~n8647 ;
  assign n18934 = n18933 ^ n10939 ^ 1'b0 ;
  assign n18935 = n1319 & n8154 ;
  assign n18936 = n2935 | n4455 ;
  assign n18937 = n18935 | n18936 ;
  assign n18938 = n12485 | n18937 ;
  assign n18939 = n3388 & n3664 ;
  assign n18940 = ~n3185 & n10225 ;
  assign n18941 = n7934 | n18940 ;
  assign n18942 = n18941 ^ n4711 ^ 1'b0 ;
  assign n18943 = n18942 ^ n2983 ^ 1'b0 ;
  assign n18944 = n18939 & n18943 ;
  assign n18945 = ~n18938 & n18944 ;
  assign n18946 = ( ~n4229 & n5331 ) | ( ~n4229 & n9606 ) | ( n5331 & n9606 ) ;
  assign n18947 = n5119 & n7313 ;
  assign n18948 = ~n18946 & n18947 ;
  assign n18949 = n2230 & n12258 ;
  assign n18950 = n1772 & n18949 ;
  assign n18951 = n18950 ^ n17316 ^ 1'b0 ;
  assign n18952 = n12773 ^ n1768 ^ 1'b0 ;
  assign n18953 = n1930 & n18952 ;
  assign n18954 = n4187 ^ n3701 ^ 1'b0 ;
  assign n18955 = ~n6250 & n18954 ;
  assign n18956 = n7257 & n17336 ;
  assign n18957 = ~n15914 & n18956 ;
  assign n18958 = ~n482 & n3423 ;
  assign n18959 = n13581 ^ n12033 ^ 1'b0 ;
  assign n18960 = n12869 | n17561 ;
  assign n18961 = n18960 ^ n16735 ^ 1'b0 ;
  assign n18962 = n8356 ^ n7226 ^ 1'b0 ;
  assign n18963 = ( n6019 & ~n6754 ) | ( n6019 & n16413 ) | ( ~n6754 & n16413 ) ;
  assign n18964 = ( n7817 & n18962 ) | ( n7817 & n18963 ) | ( n18962 & n18963 ) ;
  assign n18965 = n9764 & n12594 ;
  assign n18966 = n18965 ^ n14495 ^ 1'b0 ;
  assign n18967 = n4594 ^ n3043 ^ 1'b0 ;
  assign n18968 = n18967 ^ n11556 ^ 1'b0 ;
  assign n18969 = n9054 | n18968 ;
  assign n18970 = n18969 ^ n10162 ^ 1'b0 ;
  assign n18971 = n18193 ^ n1838 ^ 1'b0 ;
  assign n18972 = n2539 & n18971 ;
  assign n18974 = n9394 & ~n17288 ;
  assign n18973 = n17368 ^ n4705 ^ x110 ;
  assign n18975 = n18974 ^ n18973 ^ 1'b0 ;
  assign n18976 = n3832 | n18068 ;
  assign n18977 = n3088 & ~n18976 ;
  assign n18978 = n9401 ^ n822 ^ 1'b0 ;
  assign n18979 = n18978 ^ x119 ^ 1'b0 ;
  assign n18980 = n16163 & ~n18979 ;
  assign n18981 = n2015 & n5079 ;
  assign n18982 = ~n10618 & n17775 ;
  assign n18983 = n18981 & n18982 ;
  assign n18984 = n16103 | n18983 ;
  assign n18986 = n1269 & n16729 ;
  assign n18987 = ~n4100 & n18986 ;
  assign n18985 = ~n12747 & n12983 ;
  assign n18988 = n18987 ^ n18985 ^ 1'b0 ;
  assign n18989 = ~n4057 & n7726 ;
  assign n18990 = n5103 & ~n10326 ;
  assign n18991 = n12346 & ~n18990 ;
  assign n18992 = n12018 & n18991 ;
  assign n18993 = n8648 ^ n478 ^ 1'b0 ;
  assign n18994 = n968 & n4529 ;
  assign n18995 = n6060 | n18994 ;
  assign n18996 = n18995 ^ n7992 ^ 1'b0 ;
  assign n18997 = n4442 ^ n1605 ^ 1'b0 ;
  assign n19001 = n2041 & n6432 ;
  assign n18998 = ( n1289 & ~n3062 ) | ( n1289 & n5869 ) | ( ~n3062 & n5869 ) ;
  assign n18999 = ~n3312 & n6934 ;
  assign n19000 = n18998 & ~n18999 ;
  assign n19002 = n19001 ^ n19000 ^ 1'b0 ;
  assign n19003 = ~n2105 & n13707 ;
  assign n19004 = n15910 ^ n2350 ^ 1'b0 ;
  assign n19005 = n17281 & n19004 ;
  assign n19006 = n3700 & n6717 ;
  assign n19007 = n19006 ^ n1071 ^ 1'b0 ;
  assign n19008 = n4659 & n7924 ;
  assign n19009 = ( n2407 & n8083 ) | ( n2407 & n13063 ) | ( n8083 & n13063 ) ;
  assign n19010 = ( n7697 & n19008 ) | ( n7697 & ~n19009 ) | ( n19008 & ~n19009 ) ;
  assign n19011 = n18089 ^ n14868 ^ n12963 ;
  assign n19012 = n2915 & ~n11014 ;
  assign n19013 = n3388 ^ n1800 ^ 1'b0 ;
  assign n19014 = n14841 & n19013 ;
  assign n19015 = ( n1722 & n3127 ) | ( n1722 & n15994 ) | ( n3127 & n15994 ) ;
  assign n19016 = ~n4590 & n7859 ;
  assign n19017 = n19016 ^ n7208 ^ 1'b0 ;
  assign n19018 = n19017 ^ n1072 ^ 1'b0 ;
  assign n19019 = n3088 & ~n11227 ;
  assign n19020 = n5556 | n19019 ;
  assign n19021 = ~n7627 & n9331 ;
  assign n19022 = n6721 ^ n1865 ^ 1'b0 ;
  assign n19023 = n13573 & ~n19022 ;
  assign n19024 = n11380 ^ n4711 ^ 1'b0 ;
  assign n19025 = n1082 | n19024 ;
  assign n19026 = n12169 ^ n2909 ^ 1'b0 ;
  assign n19027 = n3107 & ~n19026 ;
  assign n19028 = n19027 ^ n10123 ^ 1'b0 ;
  assign n19029 = n19025 | n19028 ;
  assign n19032 = n718 | n878 ;
  assign n19033 = n19032 ^ n3845 ^ 1'b0 ;
  assign n19031 = n1033 & n3007 ;
  assign n19034 = n19033 ^ n19031 ^ 1'b0 ;
  assign n19035 = n19034 ^ n2690 ^ 1'b0 ;
  assign n19030 = n7832 & n12959 ;
  assign n19036 = n19035 ^ n19030 ^ n6895 ;
  assign n19037 = n12734 ^ n9525 ^ 1'b0 ;
  assign n19039 = n9992 ^ n4631 ^ 1'b0 ;
  assign n19038 = n559 & n14076 ;
  assign n19040 = n19039 ^ n19038 ^ 1'b0 ;
  assign n19041 = n4236 & ~n19040 ;
  assign n19044 = ~x64 & n6811 ;
  assign n19045 = ~n3682 & n19044 ;
  assign n19042 = n1430 ^ n663 ^ 1'b0 ;
  assign n19043 = n8579 & ~n19042 ;
  assign n19046 = n19045 ^ n19043 ^ 1'b0 ;
  assign n19047 = ~n14041 & n19046 ;
  assign n19048 = n14595 ^ n3501 ^ 1'b0 ;
  assign n19049 = n8112 & n9942 ;
  assign n19050 = ~n2636 & n11489 ;
  assign n19051 = n19050 ^ n17979 ^ 1'b0 ;
  assign n19052 = n15585 | n19051 ;
  assign n19053 = n16922 ^ n15851 ^ 1'b0 ;
  assign n19054 = n14179 & n19053 ;
  assign n19059 = n4272 | n8701 ;
  assign n19060 = n14071 | n19059 ;
  assign n19055 = x58 | n549 ;
  assign n19056 = n19055 ^ n1548 ^ n1023 ;
  assign n19057 = n19056 ^ n3169 ^ 1'b0 ;
  assign n19058 = n19057 ^ n11737 ^ n2105 ;
  assign n19061 = n19060 ^ n19058 ^ n3924 ;
  assign n19062 = ( n14269 & n14816 ) | ( n14269 & n15381 ) | ( n14816 & n15381 ) ;
  assign n19063 = n3081 & ~n3680 ;
  assign n19064 = n1212 & n19063 ;
  assign n19065 = n4804 ^ n2148 ^ 1'b0 ;
  assign n19066 = ~n10443 & n19065 ;
  assign n19067 = n8588 ^ n8484 ^ n4356 ;
  assign n19068 = n1220 & n4376 ;
  assign n19069 = n19068 ^ n2068 ^ 1'b0 ;
  assign n19070 = ( n19066 & n19067 ) | ( n19066 & n19069 ) | ( n19067 & n19069 ) ;
  assign n19071 = ~n19064 & n19070 ;
  assign n19072 = n19071 ^ n6372 ^ 1'b0 ;
  assign n19077 = n8899 ^ n3729 ^ n1093 ;
  assign n19073 = ~n5949 & n13052 ;
  assign n19074 = ~x146 & n19073 ;
  assign n19075 = n14633 & ~n19074 ;
  assign n19076 = n19075 ^ n10387 ^ 1'b0 ;
  assign n19078 = n19077 ^ n19076 ^ n8901 ;
  assign n19079 = ( x123 & n2005 ) | ( x123 & ~n3556 ) | ( n2005 & ~n3556 ) ;
  assign n19080 = n10763 | n10893 ;
  assign n19081 = n19079 & ~n19080 ;
  assign n19082 = n19081 ^ n15602 ^ 1'b0 ;
  assign n19083 = ~n16185 & n19082 ;
  assign n19085 = ( ~n6215 & n7577 ) | ( ~n6215 & n11411 ) | ( n7577 & n11411 ) ;
  assign n19084 = n6218 & ~n15635 ;
  assign n19086 = n19085 ^ n19084 ^ 1'b0 ;
  assign n19087 = n19086 ^ n9642 ^ 1'b0 ;
  assign n19088 = n14918 & ~n19087 ;
  assign n19089 = n9023 ^ n4826 ^ 1'b0 ;
  assign n19090 = ~n647 & n7239 ;
  assign n19091 = ~n8071 & n19090 ;
  assign n19092 = n3113 & n19091 ;
  assign n19093 = n8805 ^ n6952 ^ n5452 ;
  assign n19094 = n9382 & ~n15305 ;
  assign n19095 = ~n790 & n19094 ;
  assign n19096 = n2061 | n19095 ;
  assign n19097 = n5744 & ~n19096 ;
  assign n19103 = n14750 ^ n13373 ^ 1'b0 ;
  assign n19104 = n1677 & n19103 ;
  assign n19105 = ~n8851 & n19104 ;
  assign n19099 = ( n4009 & n6375 ) | ( n4009 & n10605 ) | ( n6375 & n10605 ) ;
  assign n19100 = n4610 | n19099 ;
  assign n19098 = n7575 & ~n18692 ;
  assign n19101 = n19100 ^ n19098 ^ 1'b0 ;
  assign n19102 = ( n7093 & n11494 ) | ( n7093 & ~n19101 ) | ( n11494 & ~n19101 ) ;
  assign n19106 = n19105 ^ n19102 ^ n7184 ;
  assign n19113 = ( n759 & ~n1261 ) | ( n759 & n6314 ) | ( ~n1261 & n6314 ) ;
  assign n19107 = n10313 ^ n5338 ^ 1'b0 ;
  assign n19108 = n6888 & n19107 ;
  assign n19109 = n19108 ^ n16596 ^ 1'b0 ;
  assign n19110 = n8942 & n19109 ;
  assign n19111 = ~n12717 & n19110 ;
  assign n19112 = n19111 ^ n12382 ^ n9489 ;
  assign n19114 = n19113 ^ n19112 ^ 1'b0 ;
  assign n19115 = n9111 & n19114 ;
  assign n19116 = ( n3229 & n6615 ) | ( n3229 & n11432 ) | ( n6615 & n11432 ) ;
  assign n19117 = n4753 & n19116 ;
  assign n19118 = n2653 & n9934 ;
  assign n19120 = ~n5509 & n5542 ;
  assign n19121 = n19120 ^ n16338 ^ 1'b0 ;
  assign n19119 = n14696 | n16985 ;
  assign n19122 = n19121 ^ n19119 ^ 1'b0 ;
  assign n19123 = n9371 & ~n19122 ;
  assign n19124 = ( n3864 & ~n9860 ) | ( n3864 & n10092 ) | ( ~n9860 & n10092 ) ;
  assign n19125 = n13214 ^ n2469 ^ 1'b0 ;
  assign n19126 = ( n469 & ~n9638 ) | ( n469 & n18629 ) | ( ~n9638 & n18629 ) ;
  assign n19127 = n19126 ^ n17164 ^ 1'b0 ;
  assign n19128 = n5073 & ~n10066 ;
  assign n19129 = ~n10097 & n19128 ;
  assign n19130 = n16578 | n19129 ;
  assign n19131 = n19130 ^ n5992 ^ 1'b0 ;
  assign n19132 = n19131 ^ n1380 ^ 1'b0 ;
  assign n19133 = ~n3904 & n15418 ;
  assign n19134 = n19133 ^ n6550 ^ 1'b0 ;
  assign n19135 = n13756 ^ n11728 ^ n1686 ;
  assign n19137 = n7930 ^ n7096 ^ n5077 ;
  assign n19136 = n6274 & ~n12952 ;
  assign n19138 = n19137 ^ n19136 ^ 1'b0 ;
  assign n19139 = ( n514 & ~n14777 ) | ( n514 & n19138 ) | ( ~n14777 & n19138 ) ;
  assign n19143 = n5022 & n14010 ;
  assign n19140 = n9259 ^ n4009 ^ 1'b0 ;
  assign n19141 = n3992 & ~n19140 ;
  assign n19142 = n19141 ^ n16054 ^ 1'b0 ;
  assign n19144 = n19143 ^ n19142 ^ 1'b0 ;
  assign n19145 = n2253 & ~n12839 ;
  assign n19146 = ~n10738 & n15406 ;
  assign n19147 = n19146 ^ n3899 ^ 1'b0 ;
  assign n19148 = n19147 ^ n600 ^ 1'b0 ;
  assign n19149 = ~n10901 & n19148 ;
  assign n19150 = n15013 ^ n7477 ^ n2055 ;
  assign n19151 = n13920 ^ n2250 ^ 1'b0 ;
  assign n19152 = n19151 ^ n11850 ^ 1'b0 ;
  assign n19153 = n19150 & ~n19152 ;
  assign n19154 = n1917 | n17036 ;
  assign n19155 = n19154 ^ n674 ^ 1'b0 ;
  assign n19156 = n19155 ^ n13982 ^ n12085 ;
  assign n19157 = n19156 ^ n18156 ^ n12350 ;
  assign n19158 = ( n4985 & n6462 ) | ( n4985 & n9694 ) | ( n6462 & n9694 ) ;
  assign n19159 = n4364 & n4793 ;
  assign n19160 = n7440 | n12723 ;
  assign n19161 = n11703 & ~n19160 ;
  assign n19162 = n19161 ^ n11388 ^ n843 ;
  assign n19163 = n10948 ^ n3824 ^ 1'b0 ;
  assign n19164 = n19163 ^ n13014 ^ 1'b0 ;
  assign n19165 = n11097 | n14618 ;
  assign n19166 = n4434 | n19165 ;
  assign n19167 = n7753 & n19166 ;
  assign n19168 = n10779 | n11951 ;
  assign n19169 = ( n751 & n12624 ) | ( n751 & n12819 ) | ( n12624 & n12819 ) ;
  assign n19170 = n19169 ^ n9772 ^ 1'b0 ;
  assign n19171 = ~n4812 & n9241 ;
  assign n19172 = n10339 | n19171 ;
  assign n19173 = n14135 | n19172 ;
  assign n19174 = n14341 ^ n13048 ^ 1'b0 ;
  assign n19175 = ~n15926 & n19174 ;
  assign n19176 = n9858 ^ n7646 ^ 1'b0 ;
  assign n19177 = n8190 & n19176 ;
  assign n19178 = ( x108 & ~n1015 ) | ( x108 & n13157 ) | ( ~n1015 & n13157 ) ;
  assign n19179 = n19178 ^ n11393 ^ 1'b0 ;
  assign n19180 = n12169 & n19179 ;
  assign n19181 = ~n7110 & n19180 ;
  assign n19182 = n19177 & n19181 ;
  assign n19183 = n19182 ^ n14796 ^ 1'b0 ;
  assign n19187 = n14732 ^ n7698 ^ 1'b0 ;
  assign n19186 = ( n5988 & n6693 ) | ( n5988 & ~n11153 ) | ( n6693 & ~n11153 ) ;
  assign n19184 = n1209 & ~n8362 ;
  assign n19185 = n13209 & n19184 ;
  assign n19188 = n19187 ^ n19186 ^ n19185 ;
  assign n19189 = n1175 & ~n19188 ;
  assign n19190 = x106 & ~n11017 ;
  assign n19191 = ( n1000 & ~n2441 ) | ( n1000 & n11291 ) | ( ~n2441 & n11291 ) ;
  assign n19192 = ~n14997 & n19191 ;
  assign n19193 = n19192 ^ n2255 ^ x84 ;
  assign n19194 = ( ~n569 & n11251 ) | ( ~n569 & n18473 ) | ( n11251 & n18473 ) ;
  assign n19195 = ( n3223 & n4261 ) | ( n3223 & ~n6058 ) | ( n4261 & ~n6058 ) ;
  assign n19196 = ~n8058 & n19195 ;
  assign n19197 = n5198 & ~n19196 ;
  assign n19198 = n19197 ^ n8702 ^ 1'b0 ;
  assign n19199 = n16464 ^ n7710 ^ 1'b0 ;
  assign n19200 = n6228 & ~n19199 ;
  assign n19201 = ~n8815 & n19200 ;
  assign n19202 = n19198 & n19201 ;
  assign n19207 = n3456 & n7322 ;
  assign n19208 = n19207 ^ n433 ^ 1'b0 ;
  assign n19209 = n558 & n19208 ;
  assign n19204 = n14940 ^ n8078 ^ 1'b0 ;
  assign n19203 = ~n1450 & n3441 ;
  assign n19205 = n19204 ^ n19203 ^ 1'b0 ;
  assign n19206 = n2413 & ~n19205 ;
  assign n19210 = n19209 ^ n19206 ^ 1'b0 ;
  assign n19211 = n2022 & ~n19210 ;
  assign n19212 = n6506 & n19211 ;
  assign n19213 = n9342 | n19212 ;
  assign n19214 = n19202 & ~n19213 ;
  assign n19215 = n5924 & ~n16767 ;
  assign n19216 = n12323 | n18079 ;
  assign n19217 = n2739 & ~n19216 ;
  assign n19218 = n2548 ^ x179 ^ 1'b0 ;
  assign n19219 = n19218 ^ n6305 ^ 1'b0 ;
  assign n19220 = n8246 & n19219 ;
  assign n19221 = ~n19217 & n19220 ;
  assign n19222 = n13137 & n19221 ;
  assign n19223 = n19222 ^ n12582 ^ 1'b0 ;
  assign n19224 = n12856 & ~n19223 ;
  assign n19225 = n14589 & ~n19224 ;
  assign n19226 = n19225 ^ n7909 ^ 1'b0 ;
  assign n19227 = n19118 & n19226 ;
  assign n19228 = n19227 ^ n3568 ^ 1'b0 ;
  assign n19229 = n369 | n5997 ;
  assign n19230 = n5934 | n19229 ;
  assign n19231 = n19230 ^ n5072 ^ 1'b0 ;
  assign n19232 = n8016 & n19231 ;
  assign n19233 = n3388 & n19232 ;
  assign n19234 = n10601 ^ n6800 ^ 1'b0 ;
  assign n19235 = n13456 ^ n4884 ^ n1124 ;
  assign n19236 = ~n15508 & n19235 ;
  assign n19237 = ~x108 & n1809 ;
  assign n19238 = n5742 | n19237 ;
  assign n19239 = n5800 ^ n3139 ^ n376 ;
  assign n19240 = n5387 & n19239 ;
  assign n19241 = n14945 ^ n13347 ^ 1'b0 ;
  assign n19242 = ~n2673 & n19241 ;
  assign n19243 = n5645 & ~n6388 ;
  assign n19244 = ~x53 & n19243 ;
  assign n19245 = n19244 ^ n10029 ^ n3067 ;
  assign n19247 = n12102 ^ n3405 ^ 1'b0 ;
  assign n19246 = ~n5141 & n14813 ;
  assign n19248 = n19247 ^ n19246 ^ 1'b0 ;
  assign n19249 = n2428 & n15571 ;
  assign n19250 = n4169 | n4241 ;
  assign n19251 = n19250 ^ n2504 ^ 1'b0 ;
  assign n19254 = ~x163 & n15987 ;
  assign n19252 = ( ~x7 & n459 ) | ( ~x7 & n3583 ) | ( n459 & n3583 ) ;
  assign n19253 = n19252 ^ n18742 ^ 1'b0 ;
  assign n19255 = n19254 ^ n19253 ^ n7151 ;
  assign n19256 = n3551 & ~n18026 ;
  assign n19257 = ~n3599 & n19256 ;
  assign n19258 = n3257 | n7912 ;
  assign n19259 = ( ~n13975 & n17519 ) | ( ~n13975 & n19258 ) | ( n17519 & n19258 ) ;
  assign n19260 = n15776 ^ n13981 ^ 1'b0 ;
  assign n19261 = ~n600 & n19260 ;
  assign n19262 = ~n10707 & n19261 ;
  assign n19263 = n19262 ^ n9798 ^ 1'b0 ;
  assign n19264 = n16954 ^ n16140 ^ n770 ;
  assign n19265 = n11465 | n14421 ;
  assign n19266 = n12957 ^ n5473 ^ 1'b0 ;
  assign n19267 = n8811 | n19266 ;
  assign n19271 = ~n4216 & n5452 ;
  assign n19272 = n19271 ^ n3536 ^ 1'b0 ;
  assign n19268 = n399 & ~n1515 ;
  assign n19269 = n19268 ^ n2988 ^ 1'b0 ;
  assign n19270 = n1354 | n19269 ;
  assign n19273 = n19272 ^ n19270 ^ 1'b0 ;
  assign n19274 = ( ~n7517 & n19267 ) | ( ~n7517 & n19273 ) | ( n19267 & n19273 ) ;
  assign n19276 = n5653 & ~n8647 ;
  assign n19275 = n9091 & ~n17120 ;
  assign n19277 = n19276 ^ n19275 ^ 1'b0 ;
  assign n19278 = ( n2279 & n8369 ) | ( n2279 & n11966 ) | ( n8369 & n11966 ) ;
  assign n19279 = n4556 | n19278 ;
  assign n19280 = n11186 | n19279 ;
  assign n19281 = n19280 ^ n14086 ^ 1'b0 ;
  assign n19284 = n7186 & ~n8978 ;
  assign n19285 = n9490 & n19284 ;
  assign n19286 = n19285 ^ n11783 ^ 1'b0 ;
  assign n19287 = n4937 & ~n19286 ;
  assign n19282 = n11067 & n15795 ;
  assign n19283 = n19282 ^ n11741 ^ 1'b0 ;
  assign n19288 = n19287 ^ n19283 ^ 1'b0 ;
  assign n19289 = ~n19281 & n19288 ;
  assign n19290 = n3131 | n8682 ;
  assign n19291 = n4606 & n7316 ;
  assign n19292 = n19291 ^ n6218 ^ 1'b0 ;
  assign n19293 = ( n322 & n1804 ) | ( n322 & ~n19292 ) | ( n1804 & ~n19292 ) ;
  assign n19297 = n5110 ^ x14 ^ 1'b0 ;
  assign n19298 = n7668 & n19297 ;
  assign n19294 = n1528 & ~n4545 ;
  assign n19295 = n19294 ^ n8247 ^ 1'b0 ;
  assign n19296 = n18521 | n19295 ;
  assign n19299 = n19298 ^ n19296 ^ 1'b0 ;
  assign n19300 = n17295 ^ n407 ^ 1'b0 ;
  assign n19301 = n745 & n19300 ;
  assign n19302 = ( n1004 & n19299 ) | ( n1004 & n19301 ) | ( n19299 & n19301 ) ;
  assign n19303 = n6927 ^ n4123 ^ 1'b0 ;
  assign n19307 = ( n1665 & n3523 ) | ( n1665 & n8440 ) | ( n3523 & n8440 ) ;
  assign n19304 = ~n1433 & n18854 ;
  assign n19305 = n19304 ^ n8997 ^ n6930 ;
  assign n19306 = ~n7389 & n19305 ;
  assign n19308 = n19307 ^ n19306 ^ 1'b0 ;
  assign n19309 = ~n363 & n13240 ;
  assign n19310 = n19309 ^ n2096 ^ 1'b0 ;
  assign n19311 = n19310 ^ n5255 ^ 1'b0 ;
  assign n19312 = n19308 | n19311 ;
  assign n19313 = n19303 & ~n19312 ;
  assign n19314 = n2052 | n15666 ;
  assign n19315 = n5143 & n12271 ;
  assign n19316 = ~n19314 & n19315 ;
  assign n19317 = n19316 ^ n11341 ^ 1'b0 ;
  assign n19318 = n4555 ^ x188 ^ 1'b0 ;
  assign n19319 = n9689 | n14371 ;
  assign n19320 = ( ~n6428 & n18284 ) | ( ~n6428 & n18594 ) | ( n18284 & n18594 ) ;
  assign n19321 = n9870 ^ n6574 ^ 1'b0 ;
  assign n19322 = n7071 | n16291 ;
  assign n19323 = n2504 | n19322 ;
  assign n19324 = n5010 ^ n1003 ^ 1'b0 ;
  assign n19325 = n806 & ~n19324 ;
  assign n19326 = ( n1038 & n4585 ) | ( n1038 & ~n19325 ) | ( n4585 & ~n19325 ) ;
  assign n19327 = n8016 & ~n19326 ;
  assign n19328 = ~n19323 & n19327 ;
  assign n19329 = n4718 & ~n4894 ;
  assign n19330 = n4894 & n19329 ;
  assign n19331 = n5139 & ~n19330 ;
  assign n19332 = ~n5139 & n19331 ;
  assign n19333 = x67 & ~n1059 ;
  assign n19334 = ~x67 & n19333 ;
  assign n19335 = n697 & ~n3910 ;
  assign n19336 = n3910 & n19335 ;
  assign n19337 = n5460 & ~n19336 ;
  assign n19338 = n19336 & n19337 ;
  assign n19339 = n19334 & ~n19338 ;
  assign n19340 = n1869 & n19339 ;
  assign n19341 = n19332 & n19340 ;
  assign n19342 = n4089 | n5527 ;
  assign n19343 = n4089 & ~n19342 ;
  assign n19344 = n3421 & ~n19343 ;
  assign n19345 = ~n3421 & n19344 ;
  assign n19346 = n344 & n1930 ;
  assign n19347 = ~n344 & n19346 ;
  assign n19348 = n1142 | n2214 ;
  assign n19349 = n19347 & ~n19348 ;
  assign n19350 = n3469 & n19349 ;
  assign n19351 = n4698 | n8352 ;
  assign n19352 = n8352 & ~n19351 ;
  assign n19353 = ~n2450 & n10937 ;
  assign n19354 = n19352 & n19353 ;
  assign n19355 = n19350 | n19354 ;
  assign n19356 = n19350 & ~n19355 ;
  assign n19357 = n7700 | n19356 ;
  assign n19358 = n19357 ^ n4068 ^ 1'b0 ;
  assign n19359 = ~n19345 & n19358 ;
  assign n19360 = ~n13185 & n19359 ;
  assign n19361 = n19341 & n19360 ;
  assign n19362 = ( x126 & ~n2955 ) | ( x126 & n4394 ) | ( ~n2955 & n4394 ) ;
  assign n19363 = x83 & n19362 ;
  assign n19364 = n19363 ^ n9401 ^ n1761 ;
  assign n19365 = n14790 ^ n11360 ^ n4404 ;
  assign n19366 = n14991 ^ n12305 ^ 1'b0 ;
  assign n19367 = ~n2846 & n5179 ;
  assign n19368 = x215 & ~n3554 ;
  assign n19369 = ( n5634 & n14936 ) | ( n5634 & ~n19368 ) | ( n14936 & ~n19368 ) ;
  assign n19370 = n9377 ^ n4325 ^ n4320 ;
  assign n19371 = n19198 & n19370 ;
  assign n19372 = ~n2176 & n7766 ;
  assign n19373 = ~n3486 & n19372 ;
  assign n19374 = n19373 ^ n14025 ^ 1'b0 ;
  assign n19375 = ( x186 & n7490 ) | ( x186 & ~n13955 ) | ( n7490 & ~n13955 ) ;
  assign n19376 = ( ~n3782 & n11960 ) | ( ~n3782 & n18509 ) | ( n11960 & n18509 ) ;
  assign n19377 = n6694 & n16683 ;
  assign n19378 = ~n19376 & n19377 ;
  assign n19379 = ~n15703 & n18888 ;
  assign n19380 = n19379 ^ n11308 ^ 1'b0 ;
  assign n19381 = n19380 ^ n14609 ^ 1'b0 ;
  assign n19382 = n19381 ^ n10537 ^ n1992 ;
  assign n19383 = n791 | n7109 ;
  assign n19384 = n7270 | n19383 ;
  assign n19385 = n11046 ^ n4073 ^ n3199 ;
  assign n19386 = n3610 | n14057 ;
  assign n19387 = n19386 ^ x33 ^ 1'b0 ;
  assign n19388 = n14687 ^ n10186 ^ n759 ;
  assign n19389 = n2264 | n19388 ;
  assign n19390 = ( ~n1478 & n11374 ) | ( ~n1478 & n14450 ) | ( n11374 & n14450 ) ;
  assign n19391 = n1909 & n11431 ;
  assign n19392 = n19390 & n19391 ;
  assign n19393 = n9544 & n19392 ;
  assign n19394 = n8203 & n13251 ;
  assign n19395 = n19394 ^ n3047 ^ n1524 ;
  assign n19396 = n815 & n13596 ;
  assign n19397 = n4306 ^ n4231 ^ 1'b0 ;
  assign n19398 = n19396 | n19397 ;
  assign n19399 = n15694 ^ n3641 ^ 1'b0 ;
  assign n19400 = n1034 ^ x63 ^ 1'b0 ;
  assign n19401 = n6636 | n8851 ;
  assign n19402 = n12125 & ~n19401 ;
  assign n19403 = n13134 | n17020 ;
  assign n19404 = n14335 & ~n19403 ;
  assign n19405 = n7805 & ~n19404 ;
  assign n19406 = n19405 ^ x59 ^ 1'b0 ;
  assign n19407 = n18899 ^ n9476 ^ 1'b0 ;
  assign n19408 = n4326 ^ n639 ^ 1'b0 ;
  assign n19409 = n19408 ^ n10511 ^ 1'b0 ;
  assign n19410 = ( n10979 & ~n13740 ) | ( n10979 & n19409 ) | ( ~n13740 & n19409 ) ;
  assign n19411 = n7190 ^ n2864 ^ 1'b0 ;
  assign n19413 = n2586 | n6873 ;
  assign n19412 = n8183 & n14000 ;
  assign n19414 = n19413 ^ n19412 ^ 1'b0 ;
  assign n19415 = n18634 & ~n19414 ;
  assign n19416 = ~n19411 & n19415 ;
  assign n19418 = n18284 ^ n7429 ^ 1'b0 ;
  assign n19417 = n7785 & ~n18329 ;
  assign n19419 = n19418 ^ n19417 ^ 1'b0 ;
  assign n19420 = ~n4857 & n11552 ;
  assign n19421 = n19420 ^ n9263 ^ 1'b0 ;
  assign n19422 = n5230 | n13903 ;
  assign n19424 = n7437 | n12853 ;
  assign n19425 = n3664 | n19424 ;
  assign n19423 = ~n7654 & n11345 ;
  assign n19426 = n19425 ^ n19423 ^ 1'b0 ;
  assign n19427 = n3984 & ~n19426 ;
  assign n19428 = n5213 ^ n3957 ^ 1'b0 ;
  assign n19429 = ~n4890 & n15037 ;
  assign n19430 = ( n3783 & ~n9281 ) | ( n3783 & n19429 ) | ( ~n9281 & n19429 ) ;
  assign n19431 = n984 & n16101 ;
  assign n19432 = n19431 ^ n17375 ^ 1'b0 ;
  assign n19433 = n4973 | n13481 ;
  assign n19434 = n19433 ^ n17554 ^ 1'b0 ;
  assign n19435 = ( n1214 & ~n18218 ) | ( n1214 & n19434 ) | ( ~n18218 & n19434 ) ;
  assign n19436 = n617 | n11113 ;
  assign n19440 = ~x49 & n3302 ;
  assign n19437 = n6720 & ~n8323 ;
  assign n19438 = n9983 & n19437 ;
  assign n19439 = n5047 | n19438 ;
  assign n19441 = n19440 ^ n19439 ^ 1'b0 ;
  assign n19442 = ( n7454 & n19436 ) | ( n7454 & n19441 ) | ( n19436 & n19441 ) ;
  assign n19443 = n1706 | n4579 ;
  assign n19444 = n19443 ^ n7303 ^ 1'b0 ;
  assign n19445 = ~n4582 & n19444 ;
  assign n19446 = n8148 ^ n3272 ^ 1'b0 ;
  assign n19447 = n8480 & ~n19446 ;
  assign n19448 = n2504 | n16000 ;
  assign n19449 = n19447 | n19448 ;
  assign n19450 = n13195 ^ n7748 ^ 1'b0 ;
  assign n19451 = ~n575 & n15536 ;
  assign n19452 = ~x0 & n271 ;
  assign n19453 = n19452 ^ n16820 ^ 1'b0 ;
  assign n19454 = n12007 ^ n9752 ^ n9331 ;
  assign n19455 = ( n1489 & ~n16925 ) | ( n1489 & n19454 ) | ( ~n16925 & n19454 ) ;
  assign n19456 = n4342 & ~n7270 ;
  assign n19457 = n567 & ~n19456 ;
  assign n19458 = n19457 ^ n3150 ^ 1'b0 ;
  assign n19459 = ~n3584 & n19458 ;
  assign n19460 = n14214 | n16377 ;
  assign n19461 = n14251 & n17106 ;
  assign n19463 = ~n1467 & n16318 ;
  assign n19462 = n8174 ^ n5253 ^ 1'b0 ;
  assign n19464 = n19463 ^ n19462 ^ 1'b0 ;
  assign n19465 = n11380 ^ n7947 ^ n1281 ;
  assign n19466 = n11246 ^ n9889 ^ 1'b0 ;
  assign n19467 = ~n11947 & n19466 ;
  assign n19470 = n4723 ^ n4386 ^ n2471 ;
  assign n19471 = n535 | n19470 ;
  assign n19468 = n11531 ^ n10055 ^ 1'b0 ;
  assign n19469 = n9227 & ~n19468 ;
  assign n19472 = n19471 ^ n19469 ^ n15282 ;
  assign n19473 = n1124 & n19472 ;
  assign n19474 = n5996 & ~n13469 ;
  assign n19475 = ~n19473 & n19474 ;
  assign n19476 = ~n10625 & n11175 ;
  assign n19477 = n6417 & n8645 ;
  assign n19478 = n12361 ^ n7897 ^ n6790 ;
  assign n19479 = n17989 ^ n17277 ^ 1'b0 ;
  assign n19480 = ~n6029 & n19479 ;
  assign n19481 = ( ~n7533 & n8348 ) | ( ~n7533 & n19480 ) | ( n8348 & n19480 ) ;
  assign n19482 = n15388 ^ n5874 ^ 1'b0 ;
  assign n19483 = n11123 ^ n5350 ^ 1'b0 ;
  assign n19484 = n2501 ^ n1941 ^ 1'b0 ;
  assign n19485 = n6856 & ~n19484 ;
  assign n19486 = ( n9594 & n19058 ) | ( n9594 & n19485 ) | ( n19058 & n19485 ) ;
  assign n19487 = ( ~x241 & n2106 ) | ( ~x241 & n12536 ) | ( n2106 & n12536 ) ;
  assign n19488 = n4611 | n19487 ;
  assign n19489 = n19488 ^ n12546 ^ 1'b0 ;
  assign n19490 = ~n1706 & n8051 ;
  assign n19491 = n2795 & n19490 ;
  assign n19492 = n616 | n19491 ;
  assign n19493 = n5433 ^ n5209 ^ 1'b0 ;
  assign n19494 = n5778 & ~n19493 ;
  assign n19495 = n19494 ^ n15054 ^ 1'b0 ;
  assign n19496 = n3332 & ~n15992 ;
  assign n19497 = n19496 ^ n4419 ^ 1'b0 ;
  assign n19505 = n4165 & ~n6205 ;
  assign n19506 = n19505 ^ n18329 ^ 1'b0 ;
  assign n19502 = n1597 & n5550 ;
  assign n19503 = n19502 ^ n3706 ^ 1'b0 ;
  assign n19498 = n1675 & n8501 ;
  assign n19499 = n19498 ^ n17017 ^ 1'b0 ;
  assign n19500 = n19499 ^ n4172 ^ 1'b0 ;
  assign n19501 = n3961 & n19500 ;
  assign n19504 = n19503 ^ n19501 ^ n1935 ;
  assign n19507 = n19506 ^ n19504 ^ 1'b0 ;
  assign n19508 = n19497 | n19507 ;
  assign n19509 = n1963 ^ n1260 ^ 1'b0 ;
  assign n19510 = n9651 & n19509 ;
  assign n19511 = n15145 ^ n5984 ^ 1'b0 ;
  assign n19512 = n19510 | n19511 ;
  assign n19513 = ~n6822 & n17131 ;
  assign n19514 = n8125 & n8296 ;
  assign n19515 = n3885 | n19514 ;
  assign n19516 = n19515 ^ n8152 ^ 1'b0 ;
  assign n19517 = n2873 & ~n13413 ;
  assign n19518 = ( n7244 & n8959 ) | ( n7244 & n13148 ) | ( n8959 & n13148 ) ;
  assign n19519 = n18475 | n19518 ;
  assign n19520 = n3149 | n19519 ;
  assign n19521 = n16581 & n19520 ;
  assign n19522 = n15395 ^ n10636 ^ 1'b0 ;
  assign n19523 = ~n2741 & n5628 ;
  assign n19524 = n19523 ^ n16391 ^ 1'b0 ;
  assign n19525 = n7656 & ~n19524 ;
  assign n19526 = n19525 ^ n2118 ^ 1'b0 ;
  assign n19527 = n19526 ^ n1768 ^ 1'b0 ;
  assign n19528 = n3126 & n19527 ;
  assign n19529 = n6781 ^ n2436 ^ 1'b0 ;
  assign n19530 = n13255 & n16725 ;
  assign n19531 = n19529 & n19530 ;
  assign n19532 = n19531 ^ n15985 ^ n7217 ;
  assign n19533 = n2261 ^ x67 ^ 1'b0 ;
  assign n19534 = n19533 ^ n1306 ^ 1'b0 ;
  assign n19535 = n3145 & ~n19534 ;
  assign n19536 = n19535 ^ n535 ^ 1'b0 ;
  assign n19537 = n15659 & n18294 ;
  assign n19538 = n19536 & n19537 ;
  assign n19539 = n2754 & ~n9230 ;
  assign n19540 = n19538 & n19539 ;
  assign n19541 = n13525 ^ n12802 ^ 1'b0 ;
  assign n19542 = n2781 | n19541 ;
  assign n19543 = ( n6792 & n11997 ) | ( n6792 & ~n17574 ) | ( n11997 & ~n17574 ) ;
  assign n19544 = x159 & n19543 ;
  assign n19545 = n19544 ^ n6435 ^ 1'b0 ;
  assign n19546 = ~n9968 & n10443 ;
  assign n19547 = ( n1795 & n6025 ) | ( n1795 & ~n14304 ) | ( n6025 & ~n14304 ) ;
  assign n19548 = n19546 | n19547 ;
  assign n19549 = ~n936 & n18870 ;
  assign n19550 = n12578 ^ n6529 ^ 1'b0 ;
  assign n19551 = n19549 & ~n19550 ;
  assign n19552 = n19551 ^ n4600 ^ 1'b0 ;
  assign n19553 = n19548 | n19552 ;
  assign n19554 = n6556 | n14421 ;
  assign n19555 = n19554 ^ n18810 ^ 1'b0 ;
  assign n19556 = n9230 | n19555 ;
  assign n19557 = n2983 ^ n1346 ^ 1'b0 ;
  assign n19558 = n19557 ^ n8572 ^ 1'b0 ;
  assign n19559 = n8989 & n13181 ;
  assign n19560 = n19558 & ~n19559 ;
  assign n19561 = n19560 ^ n10661 ^ 1'b0 ;
  assign n19562 = n8417 ^ n4797 ^ 1'b0 ;
  assign n19563 = n2353 & n7543 ;
  assign n19564 = n4026 & n10026 ;
  assign n19565 = ~n3431 & n16543 ;
  assign n19566 = n19565 ^ n19254 ^ 1'b0 ;
  assign n19567 = ~n13278 & n19566 ;
  assign n19568 = ~n18508 & n19567 ;
  assign n19569 = n8942 | n12743 ;
  assign n19570 = n8417 & ~n12592 ;
  assign n19571 = n5974 ^ n4428 ^ 1'b0 ;
  assign n19572 = n1254 & ~n19571 ;
  assign n19573 = n19572 ^ n17032 ^ 1'b0 ;
  assign n19574 = n851 & n19573 ;
  assign n19575 = ( n5336 & n12268 ) | ( n5336 & ~n12321 ) | ( n12268 & ~n12321 ) ;
  assign n19577 = ~n3403 & n3938 ;
  assign n19578 = ~n3809 & n19577 ;
  assign n19576 = n5491 & ~n8852 ;
  assign n19579 = n19578 ^ n19576 ^ 1'b0 ;
  assign n19580 = n15741 ^ n15121 ^ 1'b0 ;
  assign n19581 = n3138 & ~n19580 ;
  assign n19582 = ~n19579 & n19581 ;
  assign n19583 = n9769 & ~n13744 ;
  assign n19584 = n18337 ^ n482 ^ 1'b0 ;
  assign n19585 = n19583 & ~n19584 ;
  assign n19586 = n2660 | n2974 ;
  assign n19587 = n19586 ^ n4312 ^ 1'b0 ;
  assign n19588 = n19587 ^ n17219 ^ 1'b0 ;
  assign n19589 = n19585 & n19588 ;
  assign n19590 = n17137 ^ n16513 ^ 1'b0 ;
  assign n19591 = n19589 | n19590 ;
  assign n19592 = n3918 & n8477 ;
  assign n19593 = n19592 ^ n4991 ^ 1'b0 ;
  assign n19594 = n17796 ^ n5451 ^ 1'b0 ;
  assign n19595 = n19594 ^ n4274 ^ 1'b0 ;
  assign n19596 = n18030 | n19595 ;
  assign n19597 = n15531 ^ n1705 ^ n1612 ;
  assign n19598 = n19597 ^ n1393 ^ 1'b0 ;
  assign n19599 = n16165 & ~n19598 ;
  assign n19600 = n6352 ^ n2041 ^ 1'b0 ;
  assign n19601 = n8957 ^ n4455 ^ 1'b0 ;
  assign n19602 = ( ~n5870 & n8253 ) | ( ~n5870 & n9413 ) | ( n8253 & n9413 ) ;
  assign n19603 = n6936 & n19602 ;
  assign n19604 = ( n7962 & n19601 ) | ( n7962 & ~n19603 ) | ( n19601 & ~n19603 ) ;
  assign n19605 = n19604 ^ n6846 ^ 1'b0 ;
  assign n19606 = n13179 | n19605 ;
  assign n19607 = ( n2922 & n14448 ) | ( n2922 & ~n18114 ) | ( n14448 & ~n18114 ) ;
  assign n19608 = n15463 ^ n6911 ^ 1'b0 ;
  assign n19609 = ( n3088 & n4184 ) | ( n3088 & n4569 ) | ( n4184 & n4569 ) ;
  assign n19611 = n12140 ^ n1935 ^ 1'b0 ;
  assign n19612 = n12906 & ~n19611 ;
  assign n19610 = n14179 & ~n14790 ;
  assign n19613 = n19612 ^ n19610 ^ 1'b0 ;
  assign n19614 = n13717 ^ n8772 ^ 1'b0 ;
  assign n19615 = n5159 & ~n13742 ;
  assign n19616 = n3573 & n19615 ;
  assign n19617 = n19616 ^ n6601 ^ 1'b0 ;
  assign n19618 = n9762 & n19617 ;
  assign n19619 = n19618 ^ n5519 ^ 1'b0 ;
  assign n19620 = n15583 ^ n2346 ^ 1'b0 ;
  assign n19621 = n10605 ^ n575 ^ 1'b0 ;
  assign n19622 = ( n10657 & n14017 ) | ( n10657 & n19621 ) | ( n14017 & n19621 ) ;
  assign n19625 = n16390 ^ n6834 ^ 1'b0 ;
  assign n19623 = ~n800 & n5934 ;
  assign n19624 = n19623 ^ n14378 ^ 1'b0 ;
  assign n19626 = n19625 ^ n19624 ^ 1'b0 ;
  assign n19627 = ( n14677 & n14983 ) | ( n14677 & n18166 ) | ( n14983 & n18166 ) ;
  assign n19628 = n5264 ^ x237 ^ 1'b0 ;
  assign n19629 = n7547 & n19628 ;
  assign n19630 = ~n3794 & n19121 ;
  assign n19631 = n10863 & n19630 ;
  assign n19632 = n19629 & ~n19631 ;
  assign n19633 = ~n12237 & n19632 ;
  assign n19634 = n8963 | n19633 ;
  assign n19638 = n18915 ^ n7420 ^ 1'b0 ;
  assign n19639 = n4654 | n19638 ;
  assign n19635 = n13169 ^ n5893 ^ 1'b0 ;
  assign n19636 = n1731 ^ n723 ^ 1'b0 ;
  assign n19637 = n19635 & ~n19636 ;
  assign n19640 = n19639 ^ n19637 ^ 1'b0 ;
  assign n19641 = n2739 ^ x218 ^ 1'b0 ;
  assign n19642 = n6967 | n19641 ;
  assign n19643 = n19640 & ~n19642 ;
  assign n19644 = x59 & ~n1137 ;
  assign n19645 = n19644 ^ x111 ^ 1'b0 ;
  assign n19646 = n11872 | n19645 ;
  assign n19647 = n19646 ^ n5829 ^ 1'b0 ;
  assign n19648 = ( n10493 & ~n14505 ) | ( n10493 & n18163 ) | ( ~n14505 & n18163 ) ;
  assign n19649 = n16134 ^ n9933 ^ 1'b0 ;
  assign n19650 = n19649 ^ n9021 ^ 1'b0 ;
  assign n19651 = n19285 ^ n17048 ^ n7411 ;
  assign n19652 = n5084 | n10040 ;
  assign n19653 = ~n8363 & n19652 ;
  assign n19654 = n19653 ^ n8601 ^ 1'b0 ;
  assign n19655 = n9849 ^ n5022 ^ 1'b0 ;
  assign n19656 = ~n2648 & n19655 ;
  assign n19657 = ( n12341 & ~n16826 ) | ( n12341 & n19656 ) | ( ~n16826 & n19656 ) ;
  assign n19658 = ( n756 & ~n3470 ) | ( n756 & n16106 ) | ( ~n3470 & n16106 ) ;
  assign n19659 = n8138 & ~n8214 ;
  assign n19660 = n10325 | n19659 ;
  assign n19661 = n19658 & ~n19660 ;
  assign n19662 = n18417 ^ n1874 ^ 1'b0 ;
  assign n19663 = n14151 ^ x209 ^ 1'b0 ;
  assign n19664 = n8674 & ~n19663 ;
  assign n19665 = n11688 & n19664 ;
  assign n19666 = n15289 & ~n19665 ;
  assign n19667 = n11563 ^ n1314 ^ 1'b0 ;
  assign n19668 = n14093 ^ n2228 ^ 1'b0 ;
  assign n19669 = n6214 ^ n4819 ^ x38 ;
  assign n19670 = n563 & n11684 ;
  assign n19671 = n19670 ^ n11781 ^ 1'b0 ;
  assign n19672 = n19671 ^ n18920 ^ n4207 ;
  assign n19673 = n16660 ^ n4380 ^ 1'b0 ;
  assign n19674 = ~n10169 & n19673 ;
  assign n19675 = n14016 & n19674 ;
  assign n19677 = ( ~n1024 & n1600 ) | ( ~n1024 & n9748 ) | ( n1600 & n9748 ) ;
  assign n19676 = n2877 & n9502 ;
  assign n19678 = n19677 ^ n19676 ^ 1'b0 ;
  assign n19679 = n3554 & ~n5674 ;
  assign n19680 = n19679 ^ n9383 ^ 1'b0 ;
  assign n19681 = n19680 ^ n5668 ^ 1'b0 ;
  assign n19682 = n8122 | n19681 ;
  assign n19683 = n10786 | n19682 ;
  assign n19684 = n6711 ^ n5880 ^ 1'b0 ;
  assign n19685 = n19684 ^ n8570 ^ 1'b0 ;
  assign n19686 = n12123 & ~n19685 ;
  assign n19687 = n19686 ^ n3147 ^ 1'b0 ;
  assign n19689 = ( n2932 & n13608 ) | ( n2932 & ~n14520 ) | ( n13608 & ~n14520 ) ;
  assign n19688 = n6015 ^ n2686 ^ 1'b0 ;
  assign n19690 = n19689 ^ n19688 ^ 1'b0 ;
  assign n19691 = n3108 ^ n1776 ^ 1'b0 ;
  assign n19692 = n8709 & n19691 ;
  assign n19695 = n2670 & ~n15465 ;
  assign n19693 = x18 & n8901 ;
  assign n19694 = n1728 & n19693 ;
  assign n19696 = n19695 ^ n19694 ^ n13644 ;
  assign n19697 = n19696 ^ n13781 ^ 1'b0 ;
  assign n19698 = n10090 & ~n13251 ;
  assign n19699 = ~n11091 & n19698 ;
  assign n19700 = n8117 & n15969 ;
  assign n19701 = ~n16101 & n19700 ;
  assign n19702 = n1651 & ~n5751 ;
  assign n19703 = ( n15294 & n17297 ) | ( n15294 & ~n19702 ) | ( n17297 & ~n19702 ) ;
  assign n19704 = ( ~n2132 & n2180 ) | ( ~n2132 & n10171 ) | ( n2180 & n10171 ) ;
  assign n19705 = n1442 | n19704 ;
  assign n19706 = n15196 | n19705 ;
  assign n19707 = n8163 | n17260 ;
  assign n19708 = n10213 | n19707 ;
  assign n19709 = n19708 ^ n8298 ^ 1'b0 ;
  assign n19710 = n18846 & ~n19709 ;
  assign n19711 = n19038 | n19293 ;
  assign n19712 = n8984 | n19711 ;
  assign n19714 = n13165 ^ n2431 ^ 1'b0 ;
  assign n19715 = n19714 ^ n19503 ^ n11285 ;
  assign n19713 = n9999 ^ n1869 ^ 1'b0 ;
  assign n19716 = n19715 ^ n19713 ^ 1'b0 ;
  assign n19717 = n3479 & ~n19716 ;
  assign n19718 = n19717 ^ n3058 ^ 1'b0 ;
  assign n19719 = n2755 & ~n3568 ;
  assign n19720 = n14696 & n18759 ;
  assign n19724 = ~n5851 & n11261 ;
  assign n19721 = n4286 & ~n10897 ;
  assign n19722 = n19721 ^ n8666 ^ 1'b0 ;
  assign n19723 = n19722 ^ n3100 ^ 1'b0 ;
  assign n19725 = n19724 ^ n19723 ^ 1'b0 ;
  assign n19726 = n14876 ^ n3129 ^ 1'b0 ;
  assign n19727 = x100 & ~n19726 ;
  assign n19728 = n4158 | n12766 ;
  assign n19729 = n6561 ^ n5720 ^ 1'b0 ;
  assign n19731 = n4331 ^ n4031 ^ 1'b0 ;
  assign n19732 = ~n2073 & n19731 ;
  assign n19733 = n19732 ^ n5099 ^ n1022 ;
  assign n19730 = n4323 & ~n4534 ;
  assign n19734 = n19733 ^ n19730 ^ 1'b0 ;
  assign n19735 = n1120 | n15123 ;
  assign n19736 = n8477 | n19735 ;
  assign n19737 = n3910 | n19736 ;
  assign n19738 = ( n8225 & ~n9856 ) | ( n8225 & n9911 ) | ( ~n9856 & n9911 ) ;
  assign n19739 = ( n5726 & n13651 ) | ( n5726 & n15422 ) | ( n13651 & n15422 ) ;
  assign n19740 = ~n8453 & n13239 ;
  assign n19741 = n7305 & n19740 ;
  assign n19742 = ( n1761 & ~n7382 ) | ( n1761 & n8129 ) | ( ~n7382 & n8129 ) ;
  assign n19743 = ~n1056 & n14985 ;
  assign n19744 = ( n3588 & n19742 ) | ( n3588 & n19743 ) | ( n19742 & n19743 ) ;
  assign n19745 = ~n11486 & n17440 ;
  assign n19746 = ~n5960 & n19745 ;
  assign n19747 = n13039 | n13980 ;
  assign n19748 = n6847 ^ n5388 ^ 1'b0 ;
  assign n19749 = n12068 & ~n19748 ;
  assign n19750 = n19749 ^ n7987 ^ 1'b0 ;
  assign n19751 = n14481 ^ n11291 ^ n4264 ;
  assign n19753 = ( ~n5719 & n8094 ) | ( ~n5719 & n8287 ) | ( n8094 & n8287 ) ;
  assign n19754 = n14633 ^ n10579 ^ x106 ;
  assign n19755 = n19754 ^ n7374 ^ 1'b0 ;
  assign n19756 = ~n19753 & n19755 ;
  assign n19752 = n9882 & n14833 ;
  assign n19757 = n19756 ^ n19752 ^ 1'b0 ;
  assign n19758 = n2324 ^ n520 ^ 1'b0 ;
  assign n19759 = ( n3027 & ~n4478 ) | ( n3027 & n19758 ) | ( ~n4478 & n19758 ) ;
  assign n19760 = n19757 | n19759 ;
  assign n19761 = ~n2171 & n9981 ;
  assign n19762 = n1241 & n2449 ;
  assign n19763 = x235 & n10056 ;
  assign n19764 = n7180 | n17042 ;
  assign n19765 = n6354 & ~n19764 ;
  assign n19766 = n19765 ^ n6149 ^ 1'b0 ;
  assign n19767 = n19763 & n19766 ;
  assign n19768 = n9835 | n17016 ;
  assign n19771 = x142 & ~n2951 ;
  assign n19772 = ~n12574 & n19771 ;
  assign n19773 = n19772 ^ n4097 ^ 1'b0 ;
  assign n19774 = n6464 ^ n1140 ^ 1'b0 ;
  assign n19775 = n19774 ^ n2762 ^ 1'b0 ;
  assign n19776 = n19773 | n19775 ;
  assign n19777 = n11703 | n19776 ;
  assign n19778 = n3885 & ~n19777 ;
  assign n19779 = n15734 & ~n19778 ;
  assign n19780 = ~n1687 & n19779 ;
  assign n19769 = n4900 | n7761 ;
  assign n19770 = ~n11309 & n19769 ;
  assign n19781 = n19780 ^ n19770 ^ 1'b0 ;
  assign n19782 = n2133 ^ n905 ^ 1'b0 ;
  assign n19783 = n1162 | n19782 ;
  assign n19784 = n718 | n19783 ;
  assign n19785 = n19784 ^ n3472 ^ 1'b0 ;
  assign n19786 = n3754 | n13937 ;
  assign n19787 = n19785 | n19786 ;
  assign n19788 = n14746 ^ n2608 ^ 1'b0 ;
  assign n19789 = n1665 & ~n5637 ;
  assign n19790 = n19789 ^ n10268 ^ 1'b0 ;
  assign n19791 = n9192 & ~n19790 ;
  assign n19792 = x188 & n6644 ;
  assign n19793 = x0 | n19792 ;
  assign n19794 = ( n11432 & ~n14856 ) | ( n11432 & n19793 ) | ( ~n14856 & n19793 ) ;
  assign n19795 = x226 & n887 ;
  assign n19796 = n19795 ^ n11875 ^ 1'b0 ;
  assign n19800 = n907 | n3316 ;
  assign n19798 = ( ~n3791 & n4775 ) | ( ~n3791 & n17101 ) | ( n4775 & n17101 ) ;
  assign n19799 = n19798 ^ x14 ^ 1'b0 ;
  assign n19801 = n19800 ^ n19799 ^ 1'b0 ;
  assign n19802 = n6660 | n19801 ;
  assign n19797 = n559 | n13135 ;
  assign n19803 = n19802 ^ n19797 ^ 1'b0 ;
  assign n19804 = n7960 & n9722 ;
  assign n19805 = ~n14777 & n19804 ;
  assign n19806 = n19805 ^ n9542 ^ 1'b0 ;
  assign n19807 = n12162 ^ n8629 ^ 1'b0 ;
  assign n19808 = n4148 | n19807 ;
  assign n19809 = n8125 | n19135 ;
  assign n19810 = n2855 & ~n19809 ;
  assign n19811 = ( n6077 & n19808 ) | ( n6077 & n19810 ) | ( n19808 & n19810 ) ;
  assign n19812 = n2543 & n15870 ;
  assign n19813 = n19812 ^ n15609 ^ 1'b0 ;
  assign n19814 = n5043 ^ x29 ^ 1'b0 ;
  assign n19815 = n19814 ^ n5421 ^ 1'b0 ;
  assign n19816 = ~n15162 & n19815 ;
  assign n19817 = n7790 & ~n16486 ;
  assign n19818 = n19817 ^ n6292 ^ 1'b0 ;
  assign n19819 = n9380 ^ n2113 ^ 1'b0 ;
  assign n19820 = n6526 & n19819 ;
  assign n19821 = n19820 ^ n11559 ^ 1'b0 ;
  assign n19822 = n19821 ^ n7617 ^ n2074 ;
  assign n19823 = ( x114 & n18425 ) | ( x114 & n19822 ) | ( n18425 & n19822 ) ;
  assign n19824 = n10479 ^ n5714 ^ 1'b0 ;
  assign n19825 = n19067 | n19824 ;
  assign n19826 = n10122 ^ n3554 ^ 1'b0 ;
  assign n19827 = n18282 & ~n19826 ;
  assign n19828 = ( n7113 & n19825 ) | ( n7113 & ~n19827 ) | ( n19825 & ~n19827 ) ;
  assign n19829 = n19828 ^ n9479 ^ 1'b0 ;
  assign n19830 = ~n9450 & n19829 ;
  assign n19831 = n5801 | n19830 ;
  assign n19835 = n15834 ^ n6979 ^ 1'b0 ;
  assign n19836 = n13330 | n19835 ;
  assign n19832 = n3419 ^ n1703 ^ 1'b0 ;
  assign n19833 = n19832 ^ n13757 ^ 1'b0 ;
  assign n19834 = n19833 ^ n8903 ^ 1'b0 ;
  assign n19837 = n19836 ^ n19834 ^ n3270 ;
  assign n19838 = n19837 ^ n11647 ^ 1'b0 ;
  assign n19839 = n8025 | n19838 ;
  assign n19840 = ~n8689 & n12228 ;
  assign n19841 = n19840 ^ n5901 ^ 1'b0 ;
  assign n19842 = n19841 ^ n7650 ^ 1'b0 ;
  assign n19843 = n11995 | n17221 ;
  assign n19844 = n18734 & ~n19843 ;
  assign n19845 = n6333 ^ n5286 ^ n1194 ;
  assign n19846 = n4000 ^ n3884 ^ 1'b0 ;
  assign n19847 = n19845 & n19846 ;
  assign n19848 = n2521 ^ n2502 ^ 1'b0 ;
  assign n19849 = n19848 ^ n10873 ^ n1829 ;
  assign n19850 = ( n7185 & n19109 ) | ( n7185 & ~n19849 ) | ( n19109 & ~n19849 ) ;
  assign n19851 = n19850 ^ n6871 ^ 1'b0 ;
  assign n19852 = n19847 & n19851 ;
  assign n19853 = n3267 & ~n8851 ;
  assign n19854 = ~n9028 & n19853 ;
  assign n19855 = n8976 ^ n4487 ^ n3628 ;
  assign n19856 = n10469 | n13936 ;
  assign n19857 = n19855 & n19856 ;
  assign n19858 = n15168 ^ n5302 ^ 1'b0 ;
  assign n19859 = n16279 & n19858 ;
  assign n19862 = n3653 ^ n513 ^ 1'b0 ;
  assign n19863 = n2063 & n19862 ;
  assign n19860 = n16169 ^ n10803 ^ n2120 ;
  assign n19861 = n19860 ^ n2445 ^ 1'b0 ;
  assign n19864 = n19863 ^ n19861 ^ n16644 ;
  assign n19865 = n2071 & ~n10885 ;
  assign n19866 = n19865 ^ n8332 ^ 1'b0 ;
  assign n19867 = n5431 ^ n5296 ^ 1'b0 ;
  assign n19868 = n5263 | n19867 ;
  assign n19869 = ( n15080 & ~n19866 ) | ( n15080 & n19868 ) | ( ~n19866 & n19868 ) ;
  assign n19870 = n5330 ^ n4826 ^ 1'b0 ;
  assign n19871 = ~n8017 & n15772 ;
  assign n19872 = ~n486 & n2539 ;
  assign n19873 = n2854 & n4359 ;
  assign n19874 = n19873 ^ n9188 ^ 1'b0 ;
  assign n19875 = n14580 | n19874 ;
  assign n19876 = n19872 & ~n19875 ;
  assign n19877 = n11494 | n15462 ;
  assign n19878 = n19877 ^ n317 ^ 1'b0 ;
  assign n19879 = n5963 | n9872 ;
  assign n19880 = n19879 ^ n13120 ^ 1'b0 ;
  assign n19881 = n19880 ^ n8296 ^ n4907 ;
  assign n19882 = n698 | n14388 ;
  assign n19883 = ~n2134 & n2749 ;
  assign n19884 = n19882 & n19883 ;
  assign n19885 = ~n7466 & n19884 ;
  assign n19886 = n4775 ^ n1832 ^ 1'b0 ;
  assign n19887 = n1521 & n19886 ;
  assign n19888 = n19887 ^ n10716 ^ 1'b0 ;
  assign n19889 = n3468 & ~n19888 ;
  assign n19890 = ( ~n5980 & n6667 ) | ( ~n5980 & n19889 ) | ( n6667 & n19889 ) ;
  assign n19891 = ~n1488 & n3718 ;
  assign n19892 = ~n19890 & n19891 ;
  assign n19893 = n16634 & n19892 ;
  assign n19894 = ( ~n1184 & n1209 ) | ( ~n1184 & n19893 ) | ( n1209 & n19893 ) ;
  assign n19895 = ( n18037 & ~n19885 ) | ( n18037 & n19894 ) | ( ~n19885 & n19894 ) ;
  assign n19896 = n12834 ^ n12158 ^ 1'b0 ;
  assign n19897 = n10289 ^ n8295 ^ 1'b0 ;
  assign n19898 = x28 & n19897 ;
  assign n19899 = n19898 ^ n12150 ^ 1'b0 ;
  assign n19900 = n19899 ^ n19462 ^ 1'b0 ;
  assign n19901 = ( n4038 & n17493 ) | ( n4038 & ~n19603 ) | ( n17493 & ~n19603 ) ;
  assign n19902 = n1543 & n18867 ;
  assign n19903 = n9402 & ~n19902 ;
  assign n19904 = ( n774 & ~n3709 ) | ( n774 & n15194 ) | ( ~n3709 & n15194 ) ;
  assign n19905 = n12546 ^ n4047 ^ 1'b0 ;
  assign n19906 = ( n2739 & n4210 ) | ( n2739 & n19905 ) | ( n4210 & n19905 ) ;
  assign n19907 = n7735 ^ n5726 ^ n4274 ;
  assign n19908 = n19907 ^ n15566 ^ 1'b0 ;
  assign n19909 = n19908 ^ n4915 ^ 1'b0 ;
  assign n19910 = n3133 ^ n1350 ^ 1'b0 ;
  assign n19911 = n19909 & n19910 ;
  assign n19912 = n9036 & ~n16224 ;
  assign n19913 = n2721 | n19912 ;
  assign n19914 = n539 & ~n19913 ;
  assign n19915 = n19914 ^ n10120 ^ 1'b0 ;
  assign n19916 = ~n13059 & n15882 ;
  assign n19917 = n3209 ^ x76 ^ 1'b0 ;
  assign n19918 = x4 & ~n19917 ;
  assign n19919 = n19918 ^ n4846 ^ 1'b0 ;
  assign n19920 = n13017 & ~n19919 ;
  assign n19921 = n5311 | n8226 ;
  assign n19922 = n9470 & ~n19921 ;
  assign n19923 = n19922 ^ n9836 ^ 1'b0 ;
  assign n19924 = n13692 ^ n8278 ^ 1'b0 ;
  assign n19925 = n8936 | n19924 ;
  assign n19926 = n3694 & n9776 ;
  assign n19927 = n19926 ^ n2543 ^ 1'b0 ;
  assign n19928 = n6362 & n10448 ;
  assign n19929 = n19927 & n19928 ;
  assign n19930 = ~n3450 & n11479 ;
  assign n19931 = n19930 ^ n19516 ^ 1'b0 ;
  assign n19932 = ~n2430 & n8978 ;
  assign n19933 = n6881 & ~n19932 ;
  assign n19934 = ~n12110 & n19933 ;
  assign n19935 = ( ~n836 & n15576 ) | ( ~n836 & n17716 ) | ( n15576 & n17716 ) ;
  assign n19937 = n1957 & n9222 ;
  assign n19936 = n4758 & ~n12410 ;
  assign n19938 = n19937 ^ n19936 ^ 1'b0 ;
  assign n19939 = n19938 ^ n1376 ^ 1'b0 ;
  assign n19940 = n6005 ^ n4531 ^ 1'b0 ;
  assign n19944 = n3960 | n6321 ;
  assign n19945 = n560 & n19944 ;
  assign n19946 = ~n4268 & n19945 ;
  assign n19941 = ~n4050 & n16071 ;
  assign n19942 = n19941 ^ n2134 ^ 1'b0 ;
  assign n19943 = n3215 & n19942 ;
  assign n19947 = n19946 ^ n19943 ^ 1'b0 ;
  assign n19948 = n15567 | n19947 ;
  assign n19949 = n19940 & ~n19948 ;
  assign n19950 = n19949 ^ n15079 ^ 1'b0 ;
  assign n19951 = n259 & n4342 ;
  assign n19952 = n19951 ^ n7407 ^ 1'b0 ;
  assign n19953 = ~n1992 & n10146 ;
  assign n19954 = n19953 ^ n19866 ^ 1'b0 ;
  assign n19955 = n13249 | n19954 ;
  assign n19956 = n12619 & ~n19955 ;
  assign n19957 = ~n19952 & n19956 ;
  assign n19958 = n5905 & ~n13556 ;
  assign n19959 = ~n2634 & n13293 ;
  assign n19960 = n19959 ^ n18622 ^ n17298 ;
  assign n19961 = n10653 ^ n7439 ^ 1'b0 ;
  assign n19962 = n3942 & n19961 ;
  assign n19963 = n1843 & n2640 ;
  assign n19964 = n12161 & ~n19963 ;
  assign n19965 = n19962 & n19964 ;
  assign n19966 = ~n13621 & n19965 ;
  assign n19967 = n5893 & ~n9257 ;
  assign n19968 = n1464 & n19967 ;
  assign n19969 = n19968 ^ n3422 ^ 1'b0 ;
  assign n19970 = n8294 | n19969 ;
  assign n19972 = n2277 | n3557 ;
  assign n19973 = n1209 | n19972 ;
  assign n19971 = n19868 ^ n15996 ^ n4007 ;
  assign n19974 = n19973 ^ n19971 ^ 1'b0 ;
  assign n19975 = n12953 | n19974 ;
  assign n19976 = n12066 & ~n19975 ;
  assign n19977 = n11480 ^ n1217 ^ 1'b0 ;
  assign n19978 = n2839 | n19977 ;
  assign n19979 = n4857 ^ n1665 ^ 1'b0 ;
  assign n19980 = n19979 ^ n13227 ^ 1'b0 ;
  assign n19981 = ~n5757 & n7078 ;
  assign n19982 = n19981 ^ n10707 ^ 1'b0 ;
  assign n19983 = n19982 ^ n9307 ^ 1'b0 ;
  assign n19984 = n2830 & n19983 ;
  assign n19985 = n19984 ^ n16502 ^ 1'b0 ;
  assign n19986 = n380 | n4317 ;
  assign n19987 = n6257 ^ n1200 ^ 1'b0 ;
  assign n19988 = n11066 | n19987 ;
  assign n19989 = n8813 ^ n1239 ^ 1'b0 ;
  assign n19990 = n8245 & n19989 ;
  assign n19991 = n19990 ^ n15074 ^ 1'b0 ;
  assign n19992 = n14016 ^ n550 ^ 1'b0 ;
  assign n19993 = n19992 ^ n5820 ^ 1'b0 ;
  assign n19994 = n1610 & n19993 ;
  assign n19995 = n5304 & ~n14329 ;
  assign n19996 = n2224 | n11818 ;
  assign n19997 = ~n3560 & n9157 ;
  assign n19998 = n19997 ^ n3296 ^ 1'b0 ;
  assign n19999 = n19998 ^ n7454 ^ 1'b0 ;
  assign n20000 = n5423 & ~n19999 ;
  assign n20001 = n10550 | n20000 ;
  assign n20002 = n9371 ^ n7724 ^ 1'b0 ;
  assign n20003 = n2124 | n8358 ;
  assign n20004 = n20003 ^ n360 ^ 1'b0 ;
  assign n20005 = n20004 ^ n10097 ^ 1'b0 ;
  assign n20006 = n20002 & ~n20005 ;
  assign n20011 = n6461 ^ n5395 ^ 1'b0 ;
  assign n20007 = n3767 | n18829 ;
  assign n20008 = n790 & n20007 ;
  assign n20009 = n19161 & n20008 ;
  assign n20010 = n20009 ^ n5105 ^ 1'b0 ;
  assign n20012 = n20011 ^ n20010 ^ 1'b0 ;
  assign n20013 = n17256 ^ n5844 ^ n1663 ;
  assign n20014 = n9903 ^ n865 ^ 1'b0 ;
  assign n20015 = n13757 & n20014 ;
  assign n20018 = n7609 ^ n3448 ^ 1'b0 ;
  assign n20019 = n3746 & n20018 ;
  assign n20017 = n2699 & ~n16138 ;
  assign n20020 = n20019 ^ n20017 ^ 1'b0 ;
  assign n20016 = n1213 & ~n16186 ;
  assign n20021 = n20020 ^ n20016 ^ 1'b0 ;
  assign n20022 = n15602 ^ n3759 ^ 1'b0 ;
  assign n20023 = n17875 & ~n20022 ;
  assign n20024 = n6569 & ~n12344 ;
  assign n20026 = n17974 ^ n9763 ^ n3381 ;
  assign n20025 = n7049 & n16739 ;
  assign n20027 = n20026 ^ n20025 ^ 1'b0 ;
  assign n20028 = ~n6636 & n20027 ;
  assign n20029 = n9365 ^ n5850 ^ x199 ;
  assign n20030 = ( n1310 & ~n3354 ) | ( n1310 & n6092 ) | ( ~n3354 & n6092 ) ;
  assign n20031 = n14538 | n20030 ;
  assign n20032 = n20031 ^ n16841 ^ 1'b0 ;
  assign n20033 = n19292 | n20032 ;
  assign n20034 = n2437 & n6465 ;
  assign n20035 = n9311 & ~n20034 ;
  assign n20036 = ~n9467 & n10160 ;
  assign n20037 = n20036 ^ n7127 ^ 1'b0 ;
  assign n20038 = n11436 ^ n1667 ^ 1'b0 ;
  assign n20039 = n20038 ^ n10965 ^ x216 ;
  assign n20040 = n20039 ^ n4734 ^ 1'b0 ;
  assign n20041 = ~n2213 & n3504 ;
  assign n20042 = n4305 | n20041 ;
  assign n20043 = n15986 ^ n2409 ^ n1919 ;
  assign n20044 = n13975 ^ n6206 ^ 1'b0 ;
  assign n20045 = n20044 ^ n13925 ^ 1'b0 ;
  assign n20046 = ~n20043 & n20045 ;
  assign n20047 = ( ~n11379 & n12656 ) | ( ~n11379 & n20046 ) | ( n12656 & n20046 ) ;
  assign n20048 = n19390 ^ n11321 ^ 1'b0 ;
  assign n20049 = n20047 & ~n20048 ;
  assign n20050 = ( n6011 & ~n10408 ) | ( n6011 & n10464 ) | ( ~n10408 & n10464 ) ;
  assign n20051 = n20050 ^ n17516 ^ n5597 ;
  assign n20052 = n5979 ^ n1244 ^ 1'b0 ;
  assign n20053 = n20051 | n20052 ;
  assign n20057 = n7186 ^ x0 ^ 1'b0 ;
  assign n20055 = n6386 ^ n3955 ^ n3716 ;
  assign n20054 = n4910 ^ n2483 ^ 1'b0 ;
  assign n20056 = n20055 ^ n20054 ^ 1'b0 ;
  assign n20058 = n20057 ^ n20056 ^ n17935 ;
  assign n20059 = ~n17081 & n18283 ;
  assign n20060 = n5535 & ~n9300 ;
  assign n20061 = n821 & ~n20060 ;
  assign n20062 = ( n6338 & n11140 ) | ( n6338 & ~n15341 ) | ( n11140 & ~n15341 ) ;
  assign n20063 = n19973 ^ n650 ^ 1'b0 ;
  assign n20064 = n11910 | n20063 ;
  assign n20065 = n14553 ^ n13873 ^ 1'b0 ;
  assign n20066 = n13938 ^ n8170 ^ n773 ;
  assign n20067 = n4287 & n10070 ;
  assign n20068 = n20067 ^ n7253 ^ n3445 ;
  assign n20069 = n5159 ^ n4201 ^ 1'b0 ;
  assign n20070 = n3938 & ~n20069 ;
  assign n20071 = n3773 | n5833 ;
  assign n20072 = ~n8244 & n11774 ;
  assign n20073 = n20072 ^ n5396 ^ 1'b0 ;
  assign n20074 = ~n9579 & n20073 ;
  assign n20075 = n17238 ^ n12959 ^ 1'b0 ;
  assign n20076 = n4812 & ~n20075 ;
  assign n20077 = n20076 ^ n16905 ^ 1'b0 ;
  assign n20078 = n19845 ^ n6681 ^ n5614 ;
  assign n20079 = ( ~n5207 & n9028 ) | ( ~n5207 & n19952 ) | ( n9028 & n19952 ) ;
  assign n20080 = n10311 ^ n7495 ^ 1'b0 ;
  assign n20081 = n1393 & n7215 ;
  assign n20082 = n20081 ^ n10428 ^ 1'b0 ;
  assign n20083 = x103 & ~n20082 ;
  assign n20084 = ~n20080 & n20083 ;
  assign n20085 = n6616 & ~n20084 ;
  assign n20086 = n20085 ^ n903 ^ 1'b0 ;
  assign n20087 = n13768 & n20086 ;
  assign n20088 = ( n3648 & n10172 ) | ( n3648 & n10520 ) | ( n10172 & n10520 ) ;
  assign n20089 = n20088 ^ n10818 ^ 1'b0 ;
  assign n20090 = n17685 | n20089 ;
  assign n20091 = n20090 ^ n5431 ^ 1'b0 ;
  assign n20092 = n15675 & ~n19934 ;
  assign n20093 = ~n9906 & n20092 ;
  assign n20094 = n908 | n6724 ;
  assign n20095 = n4810 | n20094 ;
  assign n20096 = n6775 & n20095 ;
  assign n20097 = n20096 ^ n19673 ^ 1'b0 ;
  assign n20098 = n2142 & ~n20097 ;
  assign n20099 = n20098 ^ n6152 ^ 1'b0 ;
  assign n20100 = n4037 | n10516 ;
  assign n20101 = n20100 ^ n8830 ^ 1'b0 ;
  assign n20102 = n11344 ^ n1369 ^ 1'b0 ;
  assign n20103 = n3342 | n20102 ;
  assign n20104 = n3318 | n14270 ;
  assign n20105 = n20103 & ~n20104 ;
  assign n20106 = n20105 ^ n874 ^ 1'b0 ;
  assign n20107 = n538 & ~n20106 ;
  assign n20108 = n15669 & ~n20107 ;
  assign n20109 = ( n15827 & n20101 ) | ( n15827 & n20108 ) | ( n20101 & n20108 ) ;
  assign n20110 = n6739 ^ n5460 ^ 1'b0 ;
  assign n20111 = ~n15712 & n20110 ;
  assign n20112 = n6066 | n13765 ;
  assign n20113 = ~n8260 & n20112 ;
  assign n20114 = ~n20111 & n20113 ;
  assign n20116 = n13623 ^ n5521 ^ 1'b0 ;
  assign n20117 = ~n642 & n20116 ;
  assign n20118 = n12213 & n20117 ;
  assign n20115 = ~n789 & n3854 ;
  assign n20119 = n20118 ^ n20115 ^ 1'b0 ;
  assign n20120 = n14668 ^ n3281 ^ 1'b0 ;
  assign n20121 = ~n5025 & n8760 ;
  assign n20122 = n5535 & n11791 ;
  assign n20123 = ~n7365 & n7384 ;
  assign n20124 = n8594 ^ n4448 ^ n989 ;
  assign n20129 = ~n6949 & n13574 ;
  assign n20130 = ~n13030 & n20129 ;
  assign n20127 = n5956 ^ n4765 ^ 1'b0 ;
  assign n20128 = ~n13589 & n20127 ;
  assign n20125 = n14233 ^ n9753 ^ 1'b0 ;
  assign n20126 = n14127 | n20125 ;
  assign n20131 = n20130 ^ n20128 ^ n20126 ;
  assign n20132 = n20124 & n20131 ;
  assign n20133 = n20132 ^ n13994 ^ 1'b0 ;
  assign n20134 = n17506 ^ n5519 ^ 1'b0 ;
  assign n20135 = n11244 ^ n755 ^ x4 ;
  assign n20136 = n10593 & ~n12372 ;
  assign n20137 = n20136 ^ n8545 ^ 1'b0 ;
  assign n20138 = n20137 ^ n4170 ^ 1'b0 ;
  assign n20139 = n10935 ^ n3176 ^ 1'b0 ;
  assign n20140 = ~n16415 & n20139 ;
  assign n20141 = n8328 & ~n8698 ;
  assign n20142 = n291 | n20141 ;
  assign n20143 = n20142 ^ n8490 ^ 1'b0 ;
  assign n20144 = n20143 ^ n17697 ^ 1'b0 ;
  assign n20145 = n326 & ~n6565 ;
  assign n20146 = n20145 ^ n6159 ^ 1'b0 ;
  assign n20147 = n12699 ^ n2617 ^ 1'b0 ;
  assign n20148 = n20146 & n20147 ;
  assign n20149 = n1836 | n18125 ;
  assign n20150 = n12198 & ~n20149 ;
  assign n20151 = n11933 ^ n3109 ^ 1'b0 ;
  assign n20152 = n6312 | n19388 ;
  assign n20153 = n15222 ^ n1005 ^ 1'b0 ;
  assign n20154 = n9356 & ~n12218 ;
  assign n20155 = ~n14801 & n20154 ;
  assign n20156 = n2125 & ~n7282 ;
  assign n20157 = n2686 | n20156 ;
  assign n20158 = ( x82 & n13189 ) | ( x82 & ~n16483 ) | ( n13189 & ~n16483 ) ;
  assign n20159 = n20158 ^ n12761 ^ n6307 ;
  assign n20160 = ~n6798 & n20159 ;
  assign n20161 = n17820 ^ n5116 ^ n2183 ;
  assign n20162 = ( ~n3504 & n6019 ) | ( ~n3504 & n20161 ) | ( n6019 & n20161 ) ;
  assign n20165 = n6164 ^ n4902 ^ 1'b0 ;
  assign n20163 = n14132 ^ n9477 ^ n5952 ;
  assign n20164 = n4100 & ~n20163 ;
  assign n20166 = n20165 ^ n20164 ^ 1'b0 ;
  assign n20167 = n20166 ^ x22 ^ 1'b0 ;
  assign n20168 = n1469 & n20167 ;
  assign n20169 = n17059 ^ n10343 ^ 1'b0 ;
  assign n20170 = n12295 ^ n716 ^ 1'b0 ;
  assign n20171 = n20170 ^ n1764 ^ 1'b0 ;
  assign n20172 = n8823 & ~n20171 ;
  assign n20173 = n20172 ^ n2530 ^ 1'b0 ;
  assign n20174 = n2353 & n9688 ;
  assign n20175 = n4216 & n20174 ;
  assign n20176 = n10106 & n10495 ;
  assign n20177 = n17468 & n20176 ;
  assign n20178 = n11140 | n11728 ;
  assign n20179 = ~n11672 & n20178 ;
  assign n20180 = n2186 & ~n4460 ;
  assign n20181 = n16023 & n20180 ;
  assign n20182 = n5932 & n12820 ;
  assign n20183 = n2614 & n20182 ;
  assign n20184 = n6354 | n8115 ;
  assign n20185 = n14807 & ~n20184 ;
  assign n20186 = n8528 | n20185 ;
  assign n20187 = n20186 ^ n17963 ^ 1'b0 ;
  assign n20190 = ( ~n6655 & n9579 ) | ( ~n6655 & n20054 ) | ( n9579 & n20054 ) ;
  assign n20191 = ~n3806 & n6385 ;
  assign n20192 = n5586 & n20191 ;
  assign n20193 = n20192 ^ n17290 ^ 1'b0 ;
  assign n20194 = n20190 & n20193 ;
  assign n20188 = n10548 ^ n6413 ^ 1'b0 ;
  assign n20189 = ~n16891 & n20188 ;
  assign n20195 = n20194 ^ n20189 ^ 1'b0 ;
  assign n20196 = ( x0 & n731 ) | ( x0 & ~n8627 ) | ( n731 & ~n8627 ) ;
  assign n20197 = ~n15978 & n15980 ;
  assign n20198 = n9154 ^ n4895 ^ 1'b0 ;
  assign n20199 = n12526 | n20198 ;
  assign n20200 = n749 & ~n20199 ;
  assign n20201 = n20200 ^ n8417 ^ 1'b0 ;
  assign n20202 = n20201 ^ n12042 ^ n752 ;
  assign n20203 = n3920 & ~n8581 ;
  assign n20204 = n2918 | n7452 ;
  assign n20205 = n20204 ^ n2690 ^ 1'b0 ;
  assign n20206 = n4183 & ~n20205 ;
  assign n20207 = n20203 | n20206 ;
  assign n20208 = n11408 | n20207 ;
  assign n20209 = ~n2057 & n2749 ;
  assign n20210 = n762 & n20209 ;
  assign n20211 = ~n9042 & n12876 ;
  assign n20212 = ~n19943 & n20211 ;
  assign n20213 = n20212 ^ n7021 ^ 1'b0 ;
  assign n20214 = ~n20210 & n20213 ;
  assign n20219 = ( n7399 & n13892 ) | ( n7399 & ~n16170 ) | ( n13892 & ~n16170 ) ;
  assign n20215 = n4872 ^ n1102 ^ 1'b0 ;
  assign n20216 = ~n1894 & n20215 ;
  assign n20217 = n20216 ^ n3587 ^ 1'b0 ;
  assign n20218 = n9653 | n20217 ;
  assign n20220 = n20219 ^ n20218 ^ 1'b0 ;
  assign n20221 = n20214 & ~n20220 ;
  assign n20222 = ~n301 & n18872 ;
  assign n20223 = n20222 ^ n10563 ^ 1'b0 ;
  assign n20224 = n4679 | n20223 ;
  assign n20225 = ( n2513 & ~n4741 ) | ( n2513 & n6715 ) | ( ~n4741 & n6715 ) ;
  assign n20226 = n20225 ^ n8391 ^ 1'b0 ;
  assign n20227 = ( x248 & n1084 ) | ( x248 & ~n8019 ) | ( n1084 & ~n8019 ) ;
  assign n20228 = n11458 & ~n20227 ;
  assign n20229 = n20228 ^ n14564 ^ 1'b0 ;
  assign n20230 = n17259 ^ n10115 ^ n6590 ;
  assign n20231 = n18724 ^ n12554 ^ 1'b0 ;
  assign n20232 = n8930 | n20231 ;
  assign n20233 = n20232 ^ n2906 ^ 1'b0 ;
  assign n20234 = ( n20229 & ~n20230 ) | ( n20229 & n20233 ) | ( ~n20230 & n20233 ) ;
  assign n20235 = n2796 & n3003 ;
  assign n20236 = n14409 ^ n14085 ^ x16 ;
  assign n20237 = ~n14280 & n20236 ;
  assign n20238 = n5760 & ~n14978 ;
  assign n20239 = n20238 ^ n7575 ^ 1'b0 ;
  assign n20240 = n4222 & n20239 ;
  assign n20241 = n6975 & n18974 ;
  assign n20249 = n4795 & ~n11102 ;
  assign n20250 = n20249 ^ n492 ^ 1'b0 ;
  assign n20251 = n11505 & n20250 ;
  assign n20242 = n19209 ^ n831 ^ 1'b0 ;
  assign n20243 = ~n1274 & n20242 ;
  assign n20244 = n4095 | n6354 ;
  assign n20245 = n6523 & ~n20244 ;
  assign n20246 = x71 & n2333 ;
  assign n20247 = n20245 & n20246 ;
  assign n20248 = n20243 & ~n20247 ;
  assign n20252 = n20251 ^ n20248 ^ 1'b0 ;
  assign n20253 = n20241 & n20252 ;
  assign n20254 = ~n11142 & n20253 ;
  assign n20255 = n4783 & n13644 ;
  assign n20256 = ~n1411 & n2603 ;
  assign n20257 = n20256 ^ n7978 ^ 1'b0 ;
  assign n20258 = n20257 ^ n10066 ^ 1'b0 ;
  assign n20259 = n1938 | n20258 ;
  assign n20260 = n20259 ^ x83 ^ 1'b0 ;
  assign n20261 = n20260 ^ n18242 ^ 1'b0 ;
  assign n20262 = n11401 ^ n9084 ^ n853 ;
  assign n20265 = n984 & n3705 ;
  assign n20266 = n20265 ^ n2132 ^ 1'b0 ;
  assign n20263 = ~n4438 & n7101 ;
  assign n20264 = n13712 & ~n20263 ;
  assign n20267 = n20266 ^ n20264 ^ 1'b0 ;
  assign n20268 = n3632 & n17407 ;
  assign n20269 = n1139 ^ x229 ^ 1'b0 ;
  assign n20270 = ( n9526 & n15502 ) | ( n9526 & n20269 ) | ( n15502 & n20269 ) ;
  assign n20271 = n1362 & n7859 ;
  assign n20272 = ~n353 & n20271 ;
  assign n20273 = n12443 ^ n7624 ^ n1044 ;
  assign n20274 = n20273 ^ n17582 ^ 1'b0 ;
  assign n20275 = n20272 | n20274 ;
  assign n20276 = n4537 ^ n2483 ^ 1'b0 ;
  assign n20277 = n7157 & n20276 ;
  assign n20278 = n7109 | n8164 ;
  assign n20279 = n20278 ^ n1546 ^ 1'b0 ;
  assign n20280 = n13608 & ~n20279 ;
  assign n20281 = ~n8093 & n20280 ;
  assign n20282 = n20281 ^ n6241 ^ 1'b0 ;
  assign n20283 = n20282 ^ n10149 ^ n3726 ;
  assign n20284 = n7278 & n20080 ;
  assign n20285 = n2048 ^ n1180 ^ 1'b0 ;
  assign n20286 = n20285 ^ n13196 ^ 1'b0 ;
  assign n20287 = n20284 & n20286 ;
  assign n20288 = ~n19696 & n20287 ;
  assign n20289 = ( x37 & x40 ) | ( x37 & ~n1807 ) | ( x40 & ~n1807 ) ;
  assign n20290 = n15237 ^ n6594 ^ 1'b0 ;
  assign n20291 = n20289 & n20290 ;
  assign n20292 = n8241 ^ n3523 ^ 1'b0 ;
  assign n20293 = ( n6907 & ~n8358 ) | ( n6907 & n14675 ) | ( ~n8358 & n14675 ) ;
  assign n20294 = n20293 ^ n11843 ^ n6599 ;
  assign n20295 = n937 & n20294 ;
  assign n20296 = ~n335 & n5579 ;
  assign n20297 = n1935 & n20296 ;
  assign n20298 = n20297 ^ n20239 ^ n14329 ;
  assign n20299 = n15447 ^ n8075 ^ 1'b0 ;
  assign n20300 = x36 | n1943 ;
  assign n20301 = n20300 ^ n11213 ^ 1'b0 ;
  assign n20302 = n15726 ^ n13923 ^ 1'b0 ;
  assign n20303 = ~n6023 & n9388 ;
  assign n20304 = ~n2937 & n20303 ;
  assign n20305 = n11831 | n13277 ;
  assign n20306 = n20304 & ~n20305 ;
  assign n20307 = ( n4452 & n14177 ) | ( n4452 & ~n20306 ) | ( n14177 & ~n20306 ) ;
  assign n20308 = ( n11249 & ~n19734 ) | ( n11249 & n20307 ) | ( ~n19734 & n20307 ) ;
  assign n20309 = n12746 ^ n6950 ^ 1'b0 ;
  assign n20310 = ~n9314 & n10378 ;
  assign n20311 = n20310 ^ n10473 ^ 1'b0 ;
  assign n20312 = n897 & ~n20311 ;
  assign n20313 = ~n3127 & n20312 ;
  assign n20314 = n8178 & n20313 ;
  assign n20315 = n20314 ^ n961 ^ 1'b0 ;
  assign n20316 = n19880 | n20315 ;
  assign n20317 = n20309 & ~n20316 ;
  assign n20318 = ~n6780 & n7411 ;
  assign n20319 = n9005 & n20318 ;
  assign n20320 = n15434 & ~n20319 ;
  assign n20321 = n2050 & n2732 ;
  assign n20322 = n20321 ^ n12031 ^ 1'b0 ;
  assign n20324 = ~n3403 & n5359 ;
  assign n20325 = ~n725 & n20324 ;
  assign n20323 = ( n2846 & n3904 ) | ( n2846 & ~n7152 ) | ( n3904 & ~n7152 ) ;
  assign n20326 = n20325 ^ n20323 ^ 1'b0 ;
  assign n20328 = n3552 & n12536 ;
  assign n20329 = n4688 | n20328 ;
  assign n20330 = n3924 & ~n20329 ;
  assign n20327 = n5708 ^ n5218 ^ n1233 ;
  assign n20331 = n20330 ^ n20327 ^ n5896 ;
  assign n20332 = n6841 & ~n11577 ;
  assign n20333 = n20332 ^ n5569 ^ 1'b0 ;
  assign n20334 = n15760 & ~n20333 ;
  assign n20335 = n2266 & n20334 ;
  assign n20336 = n6468 ^ n2118 ^ 1'b0 ;
  assign n20337 = ~n20335 & n20336 ;
  assign n20338 = ~n6373 & n13948 ;
  assign n20339 = ~n1559 & n20338 ;
  assign n20340 = n20339 ^ n5655 ^ 1'b0 ;
  assign n20341 = n1648 | n9311 ;
  assign n20348 = n5890 | n15955 ;
  assign n20345 = n10443 | n15670 ;
  assign n20346 = ( n2176 & n2486 ) | ( n2176 & n20345 ) | ( n2486 & n20345 ) ;
  assign n20342 = n1077 | n8225 ;
  assign n20343 = n1053 | n20342 ;
  assign n20344 = n8158 & n20343 ;
  assign n20347 = n20346 ^ n20344 ^ 1'b0 ;
  assign n20349 = n20348 ^ n20347 ^ n17529 ;
  assign n20350 = n19738 ^ n16361 ^ n15039 ;
  assign n20351 = n6316 ^ n2605 ^ 1'b0 ;
  assign n20352 = n1742 | n8253 ;
  assign n20353 = ~n20351 & n20352 ;
  assign n20354 = n20353 ^ x231 ^ 1'b0 ;
  assign n20355 = n20354 ^ n4682 ^ 1'b0 ;
  assign n20356 = ~n12337 & n19473 ;
  assign n20357 = n20356 ^ n13854 ^ 1'b0 ;
  assign n20358 = n8112 | n10226 ;
  assign n20359 = n10256 | n20358 ;
  assign n20360 = ~n14151 & n20359 ;
  assign n20361 = ~n13536 & n20360 ;
  assign n20365 = n9461 | n12384 ;
  assign n20366 = n20365 ^ n2495 ^ 1'b0 ;
  assign n20362 = n9828 ^ n8246 ^ 1'b0 ;
  assign n20363 = n20362 ^ n15387 ^ 1'b0 ;
  assign n20364 = n18298 | n20363 ;
  assign n20367 = n20366 ^ n20364 ^ n2543 ;
  assign n20368 = n2445 ^ n2258 ^ 1'b0 ;
  assign n20369 = ~n3383 & n20368 ;
  assign n20370 = n20369 ^ n2208 ^ n1113 ;
  assign n20371 = ( ~n3152 & n12216 ) | ( ~n3152 & n19204 ) | ( n12216 & n19204 ) ;
  assign n20372 = n5976 & ~n12713 ;
  assign n20377 = n9436 ^ n2230 ^ 1'b0 ;
  assign n20373 = n4831 | n13189 ;
  assign n20374 = x187 & ~n2881 ;
  assign n20375 = ~n10256 & n20374 ;
  assign n20376 = n20373 | n20375 ;
  assign n20378 = n20377 ^ n20376 ^ 1'b0 ;
  assign n20379 = ~n20372 & n20378 ;
  assign n20380 = n20379 ^ n8329 ^ n6491 ;
  assign n20381 = n6611 & ~n18222 ;
  assign n20382 = ~n11369 & n20381 ;
  assign n20383 = n3520 & ~n7057 ;
  assign n20384 = n20382 & n20383 ;
  assign n20385 = ~n17339 & n20384 ;
  assign n20386 = n4212 & n11112 ;
  assign n20387 = n16118 ^ n5489 ^ 1'b0 ;
  assign n20388 = n20386 & ~n20387 ;
  assign n20389 = n16684 ^ n11309 ^ 1'b0 ;
  assign n20390 = n9355 ^ n6501 ^ 1'b0 ;
  assign n20391 = n5780 & n11859 ;
  assign n20392 = n20391 ^ n14719 ^ 1'b0 ;
  assign n20393 = n13679 & ~n20392 ;
  assign n20394 = n17115 ^ n8029 ^ 1'b0 ;
  assign n20395 = n8376 ^ n2577 ^ 1'b0 ;
  assign n20396 = n14342 ^ n4921 ^ n4533 ;
  assign n20397 = ~n20395 & n20396 ;
  assign n20398 = ( n6764 & n9638 ) | ( n6764 & ~n20397 ) | ( n9638 & ~n20397 ) ;
  assign n20399 = ~n2610 & n5061 ;
  assign n20400 = n11215 | n17297 ;
  assign n20401 = n20399 & ~n20400 ;
  assign n20402 = n13214 ^ n9502 ^ 1'b0 ;
  assign n20403 = n13543 | n20402 ;
  assign n20404 = n20403 ^ n19480 ^ 1'b0 ;
  assign n20405 = n6690 & ~n20404 ;
  assign n20410 = n6704 ^ n2108 ^ n702 ;
  assign n20406 = ~n677 & n1499 ;
  assign n20407 = ~n4245 & n20406 ;
  assign n20408 = n9880 & n14891 ;
  assign n20409 = n20407 & n20408 ;
  assign n20411 = n20410 ^ n20409 ^ 1'b0 ;
  assign n20412 = ~n18449 & n20411 ;
  assign n20413 = n20412 ^ n1938 ^ 1'b0 ;
  assign n20414 = n19917 ^ n10994 ^ 1'b0 ;
  assign n20415 = ( n2116 & n2713 ) | ( n2116 & n5228 ) | ( n2713 & n5228 ) ;
  assign n20416 = ~n12863 & n15144 ;
  assign n20417 = n9832 ^ n4001 ^ 1'b0 ;
  assign n20418 = n1034 & n20417 ;
  assign n20419 = n11921 | n17263 ;
  assign n20420 = n20418 | n20419 ;
  assign n20421 = n20420 ^ n7988 ^ 1'b0 ;
  assign n20422 = n16718 & ~n20421 ;
  assign n20423 = n20422 ^ n13050 ^ 1'b0 ;
  assign n20424 = n14306 & n20423 ;
  assign n20425 = n16596 ^ n1407 ^ 1'b0 ;
  assign n20426 = n20425 ^ n14251 ^ x201 ;
  assign n20427 = n20426 ^ n19670 ^ n15239 ;
  assign n20428 = n4544 & ~n20427 ;
  assign n20429 = ~n8143 & n20428 ;
  assign n20430 = n9813 & ~n11703 ;
  assign n20431 = n20430 ^ n10360 ^ 1'b0 ;
  assign n20432 = n5722 & ~n14182 ;
  assign n20433 = n20431 & n20432 ;
  assign n20434 = n5864 & n16546 ;
  assign n20435 = n20433 & n20434 ;
  assign n20436 = n14723 & ~n15158 ;
  assign n20437 = n18695 ^ n15609 ^ 1'b0 ;
  assign n20440 = n12228 ^ n3725 ^ 1'b0 ;
  assign n20438 = n1930 | n6537 ;
  assign n20439 = n13142 | n20438 ;
  assign n20441 = n20440 ^ n20439 ^ 1'b0 ;
  assign n20442 = n18196 & n20441 ;
  assign n20443 = n15277 & n19314 ;
  assign n20444 = n4857 | n20443 ;
  assign n20445 = n20444 ^ n11610 ^ 1'b0 ;
  assign n20447 = n3804 ^ n2338 ^ 1'b0 ;
  assign n20446 = n3382 | n4046 ;
  assign n20448 = n20447 ^ n20446 ^ 1'b0 ;
  assign n20449 = n7054 ^ n2108 ^ 1'b0 ;
  assign n20450 = n2794 | n20449 ;
  assign n20451 = n12255 | n13475 ;
  assign n20452 = n20450 & ~n20451 ;
  assign n20453 = n20452 ^ n15063 ^ 1'b0 ;
  assign n20454 = ~n781 & n11869 ;
  assign n20455 = n20454 ^ n1325 ^ 1'b0 ;
  assign n20456 = n20455 ^ n6865 ^ 1'b0 ;
  assign n20457 = n10365 & n20456 ;
  assign n20458 = ~n5223 & n20457 ;
  assign n20459 = n10178 ^ n5343 ^ 1'b0 ;
  assign n20460 = n16386 ^ n2532 ^ 1'b0 ;
  assign n20461 = n3237 | n8170 ;
  assign n20462 = n10030 & n20308 ;
  assign n20463 = n11532 ^ n7353 ^ 1'b0 ;
  assign n20464 = n13523 ^ n3716 ^ 1'b0 ;
  assign n20465 = ~n10223 & n20464 ;
  assign n20466 = ~n9104 & n20465 ;
  assign n20467 = n2553 & ~n14541 ;
  assign n20468 = ~n781 & n20467 ;
  assign n20469 = n20466 & n20468 ;
  assign n20470 = n2979 | n8472 ;
  assign n20471 = n20470 ^ n18350 ^ 1'b0 ;
  assign n20472 = n8148 ^ n6232 ^ n4244 ;
  assign n20473 = n4375 & ~n20472 ;
  assign n20474 = ~n11074 & n20473 ;
  assign n20475 = n15493 & n20474 ;
  assign n20476 = ~n9842 & n11886 ;
  assign n20477 = ~n20475 & n20476 ;
  assign n20478 = n20477 ^ n616 ^ 1'b0 ;
  assign n20480 = n3350 & ~n7990 ;
  assign n20479 = ~n1007 & n16933 ;
  assign n20481 = n20480 ^ n20479 ^ 1'b0 ;
  assign n20482 = n20481 ^ n6501 ^ 1'b0 ;
  assign n20483 = n1297 & n12530 ;
  assign n20484 = ( n13114 & n20482 ) | ( n13114 & ~n20483 ) | ( n20482 & ~n20483 ) ;
  assign n20485 = n17451 ^ n15341 ^ 1'b0 ;
  assign n20486 = n14181 & n20485 ;
  assign n20487 = n1300 & n15100 ;
  assign n20488 = n20487 ^ n19067 ^ n5025 ;
  assign n20489 = ( n14583 & ~n15950 ) | ( n14583 & n20488 ) | ( ~n15950 & n20488 ) ;
  assign n20490 = n9981 | n12922 ;
  assign n20491 = n20489 & ~n20490 ;
  assign n20492 = n6346 & ~n20491 ;
  assign n20493 = n20492 ^ n14591 ^ 1'b0 ;
  assign n20494 = n20493 ^ n8156 ^ n1510 ;
  assign n20495 = ( n2826 & n5449 ) | ( n2826 & ~n10114 ) | ( n5449 & ~n10114 ) ;
  assign n20496 = ( n5179 & n15095 ) | ( n5179 & n20495 ) | ( n15095 & n20495 ) ;
  assign n20497 = ~n10539 & n20496 ;
  assign n20498 = n7469 ^ n3639 ^ 1'b0 ;
  assign n20499 = n1935 & n20498 ;
  assign n20500 = n20497 & n20499 ;
  assign n20501 = ~n6914 & n20500 ;
  assign n20502 = ~n10550 & n19144 ;
  assign n20503 = n2188 & n6312 ;
  assign n20504 = ( n7185 & n7562 ) | ( n7185 & n20503 ) | ( n7562 & n20503 ) ;
  assign n20505 = n10625 ^ n974 ^ 1'b0 ;
  assign n20506 = n19372 ^ n8662 ^ n6835 ;
  assign n20507 = n17207 ^ n12963 ^ n2799 ;
  assign n20508 = n4555 ^ n2714 ^ 1'b0 ;
  assign n20509 = n20508 ^ n11173 ^ 1'b0 ;
  assign n20510 = n2022 & n20509 ;
  assign n20511 = ~n5046 & n20510 ;
  assign n20512 = n12261 | n20511 ;
  assign n20513 = x209 & n3090 ;
  assign n20514 = n20513 ^ n2395 ^ 1'b0 ;
  assign n20515 = ( n4244 & ~n10484 ) | ( n4244 & n20514 ) | ( ~n10484 & n20514 ) ;
  assign n20516 = ( ~n5415 & n5833 ) | ( ~n5415 & n16110 ) | ( n5833 & n16110 ) ;
  assign n20517 = n20516 ^ n8515 ^ n5987 ;
  assign n20518 = n20515 | n20517 ;
  assign n20519 = n19177 | n20518 ;
  assign n20520 = n8312 ^ n2399 ^ 1'b0 ;
  assign n20521 = ( n13707 & n17666 ) | ( n13707 & n20520 ) | ( n17666 & n20520 ) ;
  assign n20522 = n6450 ^ x102 ^ 1'b0 ;
  assign n20523 = ( n1641 & n4242 ) | ( n1641 & ~n20522 ) | ( n4242 & ~n20522 ) ;
  assign n20524 = n11859 ^ n10668 ^ 1'b0 ;
  assign n20525 = n20524 ^ n15762 ^ 1'b0 ;
  assign n20526 = n4359 & ~n9916 ;
  assign n20527 = n20526 ^ n9724 ^ 1'b0 ;
  assign n20528 = n13085 | n20527 ;
  assign n20529 = n2829 & n5980 ;
  assign n20535 = ~n4160 & n9671 ;
  assign n20536 = n13103 & n20535 ;
  assign n20531 = n10596 ^ n385 ^ 1'b0 ;
  assign n20532 = ~n5042 & n20531 ;
  assign n20533 = n20532 ^ n980 ^ 1'b0 ;
  assign n20530 = n7977 | n20203 ;
  assign n20534 = n20533 ^ n20530 ^ 1'b0 ;
  assign n20537 = n20536 ^ n20534 ^ 1'b0 ;
  assign n20538 = n2922 & n4925 ;
  assign n20539 = ( n2968 & ~n5423 ) | ( n2968 & n20538 ) | ( ~n5423 & n20538 ) ;
  assign n20545 = n5603 ^ n1811 ^ 1'b0 ;
  assign n20544 = ( n2442 & n2630 ) | ( n2442 & n9221 ) | ( n2630 & n9221 ) ;
  assign n20546 = n20545 ^ n20544 ^ 1'b0 ;
  assign n20547 = n12671 & ~n14998 ;
  assign n20548 = ~n7954 & n20547 ;
  assign n20549 = n20548 ^ n274 ^ 1'b0 ;
  assign n20550 = n20546 & ~n20549 ;
  assign n20540 = n1139 & n10322 ;
  assign n20541 = n20540 ^ n11262 ^ 1'b0 ;
  assign n20542 = ( x93 & ~n1493 ) | ( x93 & n20541 ) | ( ~n1493 & n20541 ) ;
  assign n20543 = ~n5294 & n20542 ;
  assign n20551 = n20550 ^ n20543 ^ 1'b0 ;
  assign n20552 = ( n10060 & ~n14809 ) | ( n10060 & n15130 ) | ( ~n14809 & n15130 ) ;
  assign n20553 = n19298 ^ n11537 ^ n3808 ;
  assign n20554 = n8190 & n20553 ;
  assign n20555 = n20554 ^ n1442 ^ 1'b0 ;
  assign n20556 = n3542 & n20555 ;
  assign n20557 = n8708 ^ n8129 ^ 1'b0 ;
  assign n20562 = n1188 | n3072 ;
  assign n20563 = n5807 | n20562 ;
  assign n20558 = n7846 ^ n3112 ^ 1'b0 ;
  assign n20559 = n12375 & n20558 ;
  assign n20560 = ~n1558 & n20559 ;
  assign n20561 = ~n14212 & n20560 ;
  assign n20564 = n20563 ^ n20561 ^ 1'b0 ;
  assign n20565 = n16331 | n20564 ;
  assign n20566 = n3968 & n7559 ;
  assign n20567 = n20566 ^ n17005 ^ 1'b0 ;
  assign n20568 = n6617 | n15951 ;
  assign n20569 = n9888 & ~n20568 ;
  assign n20570 = n4917 ^ n3293 ^ 1'b0 ;
  assign n20571 = n10369 ^ n10223 ^ 1'b0 ;
  assign n20572 = n20570 | n20571 ;
  assign n20574 = n19207 ^ n6262 ^ n3015 ;
  assign n20573 = n8683 & n17829 ;
  assign n20575 = n20574 ^ n20573 ^ 1'b0 ;
  assign n20576 = n1435 & ~n12273 ;
  assign n20577 = n20576 ^ n10579 ^ 1'b0 ;
  assign n20578 = n3074 ^ n2995 ^ 1'b0 ;
  assign n20579 = n19015 ^ n6846 ^ 1'b0 ;
  assign n20580 = ~n706 & n20579 ;
  assign n20581 = ~n2292 & n9044 ;
  assign n20582 = n20581 ^ n20095 ^ n1760 ;
  assign n20583 = n12489 ^ n11239 ^ 1'b0 ;
  assign n20584 = x148 & ~n20583 ;
  assign n20585 = n404 & n2141 ;
  assign n20586 = n20585 ^ n653 ^ 1'b0 ;
  assign n20587 = n20586 ^ n5437 ^ n1998 ;
  assign n20588 = n20584 & n20587 ;
  assign n20589 = n20582 & n20588 ;
  assign n20590 = n16773 ^ n1572 ^ 1'b0 ;
  assign n20591 = ~n3904 & n15679 ;
  assign n20592 = n20591 ^ n10023 ^ 1'b0 ;
  assign n20593 = n17942 & ~n20592 ;
  assign n20594 = n4160 ^ n1011 ^ n838 ;
  assign n20595 = n20594 ^ n8589 ^ n3710 ;
  assign n20596 = n13616 | n20595 ;
  assign n20597 = n4724 & n7915 ;
  assign n20598 = n13742 ^ n12327 ^ n1814 ;
  assign n20599 = x214 & ~n13333 ;
  assign n20600 = n20599 ^ n11393 ^ n10028 ;
  assign n20601 = x57 & ~n1757 ;
  assign n20602 = n20601 ^ n3622 ^ 1'b0 ;
  assign n20603 = n1427 | n4746 ;
  assign n20605 = n4855 & ~n6750 ;
  assign n20604 = n14062 ^ n6776 ^ 1'b0 ;
  assign n20606 = n20605 ^ n20604 ^ 1'b0 ;
  assign n20607 = n20603 & ~n20606 ;
  assign n20608 = n12663 ^ n6690 ^ n4509 ;
  assign n20609 = n16923 & ~n19747 ;
  assign n20610 = n18003 & n20609 ;
  assign n20611 = n14329 ^ n3464 ^ 1'b0 ;
  assign n20612 = n20611 ^ n16259 ^ 1'b0 ;
  assign n20613 = ~n15693 & n20612 ;
  assign n20614 = n961 & ~n968 ;
  assign n20615 = n20614 ^ n3521 ^ 1'b0 ;
  assign n20616 = n1279 & n20615 ;
  assign n20617 = n17462 & n20616 ;
  assign n20618 = n20617 ^ n12131 ^ 1'b0 ;
  assign n20619 = n13264 & ~n20618 ;
  assign n20620 = n20619 ^ n10813 ^ 1'b0 ;
  assign n20621 = n20620 ^ n982 ^ 1'b0 ;
  assign n20622 = ( n1925 & ~n13711 ) | ( n1925 & n18380 ) | ( ~n13711 & n18380 ) ;
  assign n20623 = ~n6520 & n11432 ;
  assign n20624 = n15513 ^ n4751 ^ n616 ;
  assign n20625 = ~n2667 & n5644 ;
  assign n20626 = n1626 & ~n20625 ;
  assign n20627 = n20624 & n20626 ;
  assign n20628 = n20627 ^ n12097 ^ 1'b0 ;
  assign n20629 = n19723 & n20628 ;
  assign n20630 = n17526 ^ n9614 ^ 1'b0 ;
  assign n20631 = n4764 & ~n20630 ;
  assign n20632 = n9885 & n20631 ;
  assign n20633 = n15320 & n20632 ;
  assign n20634 = n16536 ^ n2830 ^ 1'b0 ;
  assign n20635 = n8311 | n15653 ;
  assign n20636 = n5023 & n20635 ;
  assign n20637 = n20634 & n20636 ;
  assign n20638 = n1374 & ~n20637 ;
  assign n20639 = n17424 ^ n14341 ^ n8131 ;
  assign n20640 = n15471 & ~n20639 ;
  assign n20641 = ~n3788 & n10122 ;
  assign n20642 = n20641 ^ n7172 ^ 1'b0 ;
  assign n20643 = n3898 ^ n2966 ^ n509 ;
  assign n20644 = n4448 ^ n552 ^ 1'b0 ;
  assign n20645 = n20644 ^ n7621 ^ n4279 ;
  assign n20646 = n20645 ^ n2914 ^ 1'b0 ;
  assign n20647 = n20643 & ~n20646 ;
  assign n20650 = n13492 ^ n4826 ^ 1'b0 ;
  assign n20651 = n20650 ^ n8370 ^ 1'b0 ;
  assign n20648 = n6079 ^ n560 ^ 1'b0 ;
  assign n20649 = n10923 & ~n20648 ;
  assign n20652 = n20651 ^ n20649 ^ 1'b0 ;
  assign n20653 = n7264 | n14513 ;
  assign n20654 = n9220 & ~n20653 ;
  assign n20655 = n19521 ^ n18835 ^ 1'b0 ;
  assign n20656 = n19891 & ~n20655 ;
  assign n20657 = n1598 | n3894 ;
  assign n20658 = n20657 ^ n13334 ^ 1'b0 ;
  assign n20659 = x227 & ~n20658 ;
  assign n20660 = n20659 ^ x210 ^ 1'b0 ;
  assign n20661 = ~n702 & n9275 ;
  assign n20662 = n20661 ^ n14220 ^ 1'b0 ;
  assign n20663 = n20662 ^ n1192 ^ 1'b0 ;
  assign n20664 = ~n4460 & n11479 ;
  assign n20665 = n20664 ^ x129 ^ 1'b0 ;
  assign n20666 = n6874 ^ n6708 ^ n4142 ;
  assign n20667 = ( ~n2925 & n20665 ) | ( ~n2925 & n20666 ) | ( n20665 & n20666 ) ;
  assign n20668 = n20667 ^ n18340 ^ 1'b0 ;
  assign n20669 = n12600 ^ n3460 ^ 1'b0 ;
  assign n20670 = ( n4062 & n8623 ) | ( n4062 & n12966 ) | ( n8623 & n12966 ) ;
  assign n20671 = n13460 ^ n11072 ^ 1'b0 ;
  assign n20672 = n20671 ^ n17222 ^ 1'b0 ;
  assign n20673 = ( n20496 & ~n20670 ) | ( n20496 & n20672 ) | ( ~n20670 & n20672 ) ;
  assign n20674 = n8433 & n11386 ;
  assign n20675 = n20674 ^ n2176 ^ 1'b0 ;
  assign n20676 = n19440 ^ n14667 ^ n2401 ;
  assign n20677 = ( n16998 & n20675 ) | ( n16998 & n20676 ) | ( n20675 & n20676 ) ;
  assign n20678 = x14 & ~n966 ;
  assign n20679 = ~n3833 & n19467 ;
  assign n20680 = ~n20678 & n20679 ;
  assign n20681 = x104 & n19633 ;
  assign n20682 = n4783 ^ n3841 ^ 1'b0 ;
  assign n20683 = n2129 ^ n1788 ^ 1'b0 ;
  assign n20684 = ~n11837 & n20683 ;
  assign n20685 = n20684 ^ n428 ^ 1'b0 ;
  assign n20686 = n11569 ^ n5785 ^ n2360 ;
  assign n20687 = n20685 & n20686 ;
  assign n20688 = n20687 ^ n10842 ^ 1'b0 ;
  assign n20689 = n20688 ^ n19056 ^ 1'b0 ;
  assign n20690 = n20682 & ~n20689 ;
  assign n20691 = n840 & n2993 ;
  assign n20692 = n5361 & n16928 ;
  assign n20693 = n12365 ^ n5554 ^ 1'b0 ;
  assign n20694 = n2103 & ~n20693 ;
  assign n20695 = n3059 & ~n4216 ;
  assign n20696 = ~n7122 & n20695 ;
  assign n20697 = ~n2033 & n20696 ;
  assign n20698 = n13574 ^ n9666 ^ 1'b0 ;
  assign n20699 = n18758 & ~n20698 ;
  assign n20700 = ~n2272 & n5971 ;
  assign n20701 = n20700 ^ n10787 ^ 1'b0 ;
  assign n20702 = ~n3340 & n6805 ;
  assign n20703 = ~n1137 & n7663 ;
  assign n20704 = n20703 ^ n20520 ^ n7644 ;
  assign n20705 = n2208 | n7474 ;
  assign n20706 = n5626 ^ n5182 ^ 1'b0 ;
  assign n20707 = ( n476 & n14693 ) | ( n476 & ~n20706 ) | ( n14693 & ~n20706 ) ;
  assign n20708 = n20707 ^ x84 ^ 1'b0 ;
  assign n20709 = ~n20705 & n20708 ;
  assign n20710 = ~n3067 & n6447 ;
  assign n20712 = n3275 ^ n2284 ^ 1'b0 ;
  assign n20711 = n2660 | n10720 ;
  assign n20713 = n20712 ^ n20711 ^ 1'b0 ;
  assign n20714 = n9875 & ~n12613 ;
  assign n20715 = n5445 & n20714 ;
  assign n20716 = n18490 ^ n13192 ^ 1'b0 ;
  assign n20717 = n358 & ~n3874 ;
  assign n20721 = n2235 & n5788 ;
  assign n20718 = n1941 & ~n5127 ;
  assign n20719 = ~n2307 & n10090 ;
  assign n20720 = n20718 & n20719 ;
  assign n20722 = n20721 ^ n20720 ^ n1833 ;
  assign n20723 = n7047 ^ n2192 ^ 1'b0 ;
  assign n20724 = n20723 ^ n8666 ^ 1'b0 ;
  assign n20725 = n17665 & ~n20724 ;
  assign n20726 = n13543 | n16546 ;
  assign n20727 = ~n11515 & n20726 ;
  assign n20728 = n20727 ^ n18938 ^ 1'b0 ;
  assign n20732 = ( n9042 & n10632 ) | ( n9042 & ~n18006 ) | ( n10632 & ~n18006 ) ;
  assign n20729 = n860 & n5918 ;
  assign n20730 = n20729 ^ n8351 ^ 1'b0 ;
  assign n20731 = ( n4830 & n18288 ) | ( n4830 & n20730 ) | ( n18288 & n20730 ) ;
  assign n20733 = n20732 ^ n20731 ^ 1'b0 ;
  assign n20734 = n14002 | n20733 ;
  assign n20735 = ~n456 & n3856 ;
  assign n20736 = n20735 ^ n12361 ^ 1'b0 ;
  assign n20737 = n9870 ^ n2365 ^ 1'b0 ;
  assign n20738 = n12045 | n20737 ;
  assign n20739 = n10186 & n15671 ;
  assign n20740 = n20738 & n20739 ;
  assign n20741 = n2746 ^ n2548 ^ n2337 ;
  assign n20742 = ~n2329 & n3396 ;
  assign n20743 = ~n5203 & n20742 ;
  assign n20744 = n20743 ^ n15651 ^ 1'b0 ;
  assign n20745 = n20741 | n20744 ;
  assign n20746 = ( n5398 & n13944 ) | ( n5398 & ~n18375 ) | ( n13944 & ~n18375 ) ;
  assign n20747 = n17202 ^ n13277 ^ n2369 ;
  assign n20749 = n5461 & ~n5674 ;
  assign n20748 = ~n5006 & n15196 ;
  assign n20750 = n20749 ^ n20748 ^ 1'b0 ;
  assign n20751 = ~n6088 & n8545 ;
  assign n20752 = n11310 & n20751 ;
  assign n20753 = n20752 ^ n6204 ^ 1'b0 ;
  assign n20754 = n20753 ^ n6327 ^ 1'b0 ;
  assign n20755 = n1254 & n20754 ;
  assign n20756 = n5467 & n6615 ;
  assign n20757 = n20755 & n20756 ;
  assign n20758 = n20036 ^ n2791 ^ 1'b0 ;
  assign n20759 = n18282 & n20758 ;
  assign n20760 = ( n1833 & n5196 ) | ( n1833 & ~n20759 ) | ( n5196 & ~n20759 ) ;
  assign n20761 = n478 & ~n7068 ;
  assign n20762 = n20761 ^ n1480 ^ 1'b0 ;
  assign n20763 = n13583 & n20762 ;
  assign n20764 = n20763 ^ n12176 ^ 1'b0 ;
  assign n20765 = ~n704 & n18601 ;
  assign n20766 = ~n6364 & n20765 ;
  assign n20767 = ~n2794 & n4881 ;
  assign n20768 = n20767 ^ n8649 ^ 1'b0 ;
  assign n20769 = n20768 ^ n12124 ^ 1'b0 ;
  assign n20770 = ~n6688 & n11208 ;
  assign n20771 = n20770 ^ n9888 ^ 1'b0 ;
  assign n20772 = ~x15 & n20771 ;
  assign n20773 = n20769 & n20772 ;
  assign n20774 = n10008 ^ n7099 ^ 1'b0 ;
  assign n20775 = n5510 & n16581 ;
  assign n20776 = ~n20774 & n20775 ;
  assign n20782 = n6082 ^ n2955 ^ 1'b0 ;
  assign n20783 = n2473 | n20782 ;
  assign n20784 = ( ~n2990 & n8451 ) | ( ~n2990 & n20783 ) | ( n8451 & n20783 ) ;
  assign n20777 = n8106 ^ n4189 ^ n3884 ;
  assign n20778 = n20777 ^ n7673 ^ n4501 ;
  assign n20779 = n20778 ^ n13803 ^ 1'b0 ;
  assign n20780 = n8259 & ~n10568 ;
  assign n20781 = n20779 & n20780 ;
  assign n20785 = n20784 ^ n20781 ^ n8077 ;
  assign n20786 = n3842 & n11145 ;
  assign n20787 = ~n1521 & n18668 ;
  assign n20788 = n12257 ^ n2253 ^ 1'b0 ;
  assign n20789 = n4951 | n10182 ;
  assign n20790 = n3326 | n20789 ;
  assign n20791 = n10043 & n14108 ;
  assign n20792 = n20790 | n20791 ;
  assign n20795 = n3826 & ~n9730 ;
  assign n20796 = n17128 & n20795 ;
  assign n20797 = n552 & n20796 ;
  assign n20793 = ~n10336 & n15020 ;
  assign n20794 = ~n2057 & n20793 ;
  assign n20798 = n20797 ^ n20794 ^ 1'b0 ;
  assign n20799 = n20508 ^ n1446 ^ 1'b0 ;
  assign n20800 = n19641 | n20236 ;
  assign n20801 = n20800 ^ n759 ^ 1'b0 ;
  assign n20802 = n2151 & n20801 ;
  assign n20803 = ~n6600 & n20802 ;
  assign n20804 = n5879 ^ n877 ^ 1'b0 ;
  assign n20805 = n20804 ^ n10518 ^ 1'b0 ;
  assign n20806 = n4772 | n20805 ;
  assign n20807 = n20806 ^ n5637 ^ 1'b0 ;
  assign n20808 = n6391 | n18981 ;
  assign n20809 = n3315 & ~n20808 ;
  assign n20810 = n7522 | n20809 ;
  assign n20811 = ( n11812 & n13562 ) | ( n11812 & n15700 ) | ( n13562 & n15700 ) ;
  assign n20812 = n7184 & n15734 ;
  assign n20813 = n20812 ^ n761 ^ 1'b0 ;
  assign n20814 = n7277 & n11927 ;
  assign n20815 = n20814 ^ n5984 ^ 1'b0 ;
  assign n20816 = n16727 ^ n7908 ^ 1'b0 ;
  assign n20817 = n17178 | n20816 ;
  assign n20818 = n12551 ^ n9222 ^ 1'b0 ;
  assign n20819 = n11175 | n20818 ;
  assign n20820 = n18473 ^ n4765 ^ 1'b0 ;
  assign n20821 = n10859 & n20161 ;
  assign n20822 = n20821 ^ n16587 ^ 1'b0 ;
  assign n20823 = n7060 & ~n18645 ;
  assign n20824 = ~n7007 & n20823 ;
  assign n20825 = n20822 & n20824 ;
  assign n20826 = n20825 ^ n18274 ^ 1'b0 ;
  assign n20827 = n2856 ^ n1952 ^ 1'b0 ;
  assign n20828 = n14341 ^ n8117 ^ 1'b0 ;
  assign n20829 = n13167 | n20422 ;
  assign n20830 = n7521 & n18951 ;
  assign n20831 = n20830 ^ n5319 ^ 1'b0 ;
  assign n20832 = n8410 & n9170 ;
  assign n20833 = n18451 & n20832 ;
  assign n20834 = ~n4037 & n20833 ;
  assign n20835 = n1070 & ~n1717 ;
  assign n20836 = n20835 ^ n18912 ^ 1'b0 ;
  assign n20837 = n3878 & ~n7396 ;
  assign n20838 = n20837 ^ n8229 ^ 1'b0 ;
  assign n20839 = n20838 ^ n4036 ^ 1'b0 ;
  assign n20840 = n15710 & ~n20839 ;
  assign n20841 = n20002 ^ n6601 ^ 1'b0 ;
  assign n20842 = n10144 & n13920 ;
  assign n20843 = n19436 & n20842 ;
  assign n20844 = n20843 ^ n19422 ^ 1'b0 ;
  assign n20845 = ~n5931 & n16889 ;
  assign n20846 = n2168 | n20845 ;
  assign n20847 = n5304 | n20846 ;
  assign n20848 = ( n6371 & n6563 ) | ( n6371 & n20847 ) | ( n6563 & n20847 ) ;
  assign n20849 = n2017 & ~n5025 ;
  assign n20850 = n20849 ^ n5164 ^ 1'b0 ;
  assign n20851 = n1261 & n20850 ;
  assign n20852 = n2713 & n6781 ;
  assign n20853 = n20852 ^ n4023 ^ 1'b0 ;
  assign n20854 = ~n8029 & n20853 ;
  assign n20855 = n20854 ^ n4987 ^ 1'b0 ;
  assign n20856 = n9583 & ~n20855 ;
  assign n20857 = n20851 & n20856 ;
  assign n20858 = n5483 & n17724 ;
  assign n20859 = n14054 ^ n9694 ^ 1'b0 ;
  assign n20860 = n13915 ^ n7713 ^ 1'b0 ;
  assign n20861 = ~n20783 & n20860 ;
  assign n20862 = n16920 ^ n4300 ^ n3523 ;
  assign n20863 = n3917 | n13547 ;
  assign n20864 = n20863 ^ n7089 ^ 1'b0 ;
  assign n20865 = n14143 & n20864 ;
  assign n20866 = ~n4970 & n20865 ;
  assign n20867 = n20866 ^ n14477 ^ 1'b0 ;
  assign n20868 = n5154 ^ n2941 ^ n2523 ;
  assign n20869 = n14536 ^ n5598 ^ 1'b0 ;
  assign n20870 = ~n17940 & n20869 ;
  assign n20871 = ( n13543 & ~n20868 ) | ( n13543 & n20870 ) | ( ~n20868 & n20870 ) ;
  assign n20872 = ~n19091 & n19425 ;
  assign n20873 = n20872 ^ n11053 ^ 1'b0 ;
  assign n20877 = ( ~n5666 & n13752 ) | ( ~n5666 & n20312 ) | ( n13752 & n20312 ) ;
  assign n20874 = n4652 & ~n6314 ;
  assign n20875 = n7926 | n13873 ;
  assign n20876 = n20874 | n20875 ;
  assign n20878 = n20877 ^ n20876 ^ 1'b0 ;
  assign n20879 = n3061 & n5988 ;
  assign n20880 = n15338 ^ n3866 ^ 1'b0 ;
  assign n20881 = n10364 & ~n20880 ;
  assign n20882 = n909 & n13212 ;
  assign n20883 = n20882 ^ n14035 ^ 1'b0 ;
  assign n20884 = n1156 | n20883 ;
  assign n20886 = ~n516 & n18310 ;
  assign n20887 = ~n13617 & n20886 ;
  assign n20888 = n2932 ^ n1803 ^ 1'b0 ;
  assign n20889 = ~n20887 & n20888 ;
  assign n20890 = ( ~n9373 & n12090 ) | ( ~n9373 & n20889 ) | ( n12090 & n20889 ) ;
  assign n20885 = n5528 & n14769 ;
  assign n20891 = n20890 ^ n20885 ^ 1'b0 ;
  assign n20896 = ( ~n7046 & n7587 ) | ( ~n7046 & n9279 ) | ( n7587 & n9279 ) ;
  assign n20892 = n2670 | n13021 ;
  assign n20893 = n20892 ^ n2575 ^ 1'b0 ;
  assign n20894 = n19191 & ~n20893 ;
  assign n20895 = n20894 ^ n16005 ^ 1'b0 ;
  assign n20897 = n20896 ^ n20895 ^ n10694 ;
  assign n20898 = n15406 ^ n7972 ^ 1'b0 ;
  assign n20899 = n12480 ^ n3531 ^ 1'b0 ;
  assign n20900 = n3360 & ~n20899 ;
  assign n20901 = n6751 & ~n20843 ;
  assign n20902 = ~n5060 & n17392 ;
  assign n20903 = n16305 & ~n20902 ;
  assign n20904 = n20903 ^ n10923 ^ 1'b0 ;
  assign n20905 = n11884 | n20904 ;
  assign n20906 = n20905 ^ n5864 ^ 1'b0 ;
  assign n20911 = ~n1974 & n2024 ;
  assign n20912 = n556 & n20911 ;
  assign n20907 = n8924 | n9008 ;
  assign n20908 = n1202 & ~n20907 ;
  assign n20909 = ~n17759 & n20908 ;
  assign n20910 = ~n13328 & n20909 ;
  assign n20913 = n20912 ^ n20910 ^ n18190 ;
  assign n20914 = ( n957 & n5207 ) | ( n957 & ~n7088 ) | ( n5207 & ~n7088 ) ;
  assign n20915 = n20914 ^ n13753 ^ 1'b0 ;
  assign n20916 = ~n1274 & n20915 ;
  assign n20917 = n6613 ^ n1060 ^ 1'b0 ;
  assign n20918 = n706 & ~n20917 ;
  assign n20919 = n6700 & n20918 ;
  assign n20920 = n4527 & n20919 ;
  assign n20921 = n8463 & n8719 ;
  assign n20922 = ( n5566 & n6599 ) | ( n5566 & n18187 ) | ( n6599 & n18187 ) ;
  assign n20923 = ( ~n10310 & n20921 ) | ( ~n10310 & n20922 ) | ( n20921 & n20922 ) ;
  assign n20924 = ~n10723 & n20923 ;
  assign n20925 = n11371 & n13608 ;
  assign n20926 = n20925 ^ n5073 ^ 1'b0 ;
  assign n20927 = n20926 ^ n20833 ^ 1'b0 ;
  assign n20928 = ~n14344 & n20927 ;
  assign n20929 = n3472 | n9096 ;
  assign n20930 = n6622 & n9671 ;
  assign n20934 = n706 & n9298 ;
  assign n20935 = n20934 ^ n434 ^ 1'b0 ;
  assign n20931 = n2528 | n12771 ;
  assign n20932 = n20931 ^ n11741 ^ 1'b0 ;
  assign n20933 = ~n4597 & n20932 ;
  assign n20936 = n20935 ^ n20933 ^ 1'b0 ;
  assign n20939 = ~n5790 & n13543 ;
  assign n20937 = n9798 ^ n4174 ^ 1'b0 ;
  assign n20938 = n4500 & n20937 ;
  assign n20940 = n20939 ^ n20938 ^ 1'b0 ;
  assign n20941 = n14876 ^ n11246 ^ n2352 ;
  assign n20942 = n3148 & ~n20941 ;
  assign n20943 = n19583 ^ x83 ^ 1'b0 ;
  assign n20944 = n20943 ^ n11328 ^ 1'b0 ;
  assign n20945 = n19033 ^ n12001 ^ 1'b0 ;
  assign n20946 = n20945 ^ n18480 ^ n11903 ;
  assign n20947 = n16908 & ~n20946 ;
  assign n20948 = ~n20944 & n20947 ;
  assign n20949 = ~n3997 & n17619 ;
  assign n20950 = n518 & ~n9559 ;
  assign n20951 = n20950 ^ n14329 ^ 1'b0 ;
  assign n20952 = ~n2833 & n14918 ;
  assign n20953 = n17681 & ~n20952 ;
  assign n20954 = n20953 ^ n20131 ^ 1'b0 ;
  assign n20956 = x229 | n1907 ;
  assign n20955 = ~n2232 & n13950 ;
  assign n20957 = n20956 ^ n20955 ^ 1'b0 ;
  assign n20958 = ~n513 & n6290 ;
  assign n20959 = n20957 | n20958 ;
  assign n20960 = n20959 ^ n4991 ^ 1'b0 ;
  assign n20961 = n14329 & n20960 ;
  assign n20962 = n8512 & n20961 ;
  assign n20963 = n12705 & n19451 ;
  assign n20964 = ( ~n8344 & n13090 ) | ( ~n8344 & n18131 ) | ( n13090 & n18131 ) ;
  assign n20965 = n20964 ^ n16296 ^ 1'b0 ;
  assign n20966 = ~n11251 & n20965 ;
  assign n20967 = n20966 ^ n11457 ^ 1'b0 ;
  assign n20968 = n11910 ^ n5560 ^ n5232 ;
  assign n20969 = n9331 | n16482 ;
  assign n20970 = n20969 ^ n1510 ^ 1'b0 ;
  assign n20971 = n20968 | n20970 ;
  assign n20972 = n1058 & ~n4078 ;
  assign n20973 = n2802 & n6509 ;
  assign n20974 = ~n20972 & n20973 ;
  assign n20975 = ~n16964 & n20974 ;
  assign n20976 = ( x248 & n2824 ) | ( x248 & ~n17501 ) | ( n2824 & ~n17501 ) ;
  assign n20977 = n12529 & ~n20976 ;
  assign n20978 = n7495 & n15941 ;
  assign n20979 = n8729 & n13690 ;
  assign n20980 = x161 | n7731 ;
  assign n20981 = n20980 ^ n14784 ^ 1'b0 ;
  assign n20982 = n20979 | n20981 ;
  assign n20983 = n4076 & n9088 ;
  assign n20984 = n20983 ^ n1741 ^ 1'b0 ;
  assign n20985 = n950 & n15193 ;
  assign n20986 = ~n20984 & n20985 ;
  assign n20987 = ~n2897 & n19209 ;
  assign n20988 = n20987 ^ n12616 ^ 1'b0 ;
  assign n20989 = n12440 | n20988 ;
  assign n20990 = n11764 ^ n5504 ^ 1'b0 ;
  assign n20991 = n18231 & n20990 ;
  assign n20992 = n20991 ^ n7180 ^ 1'b0 ;
  assign n20993 = n5155 ^ n3709 ^ 1'b0 ;
  assign n20994 = n20993 ^ n2387 ^ 1'b0 ;
  assign n20995 = ~n15709 & n20994 ;
  assign n20996 = n9752 & ~n20995 ;
  assign n20997 = n20996 ^ n8451 ^ 1'b0 ;
  assign n20998 = x178 & ~n8517 ;
  assign n20999 = n3504 & ~n7564 ;
  assign n21000 = n1518 & n20999 ;
  assign n21001 = n4799 | n21000 ;
  assign n21002 = n21001 ^ n12970 ^ n3755 ;
  assign n21003 = ~n3926 & n10344 ;
  assign n21004 = n12690 ^ n2294 ^ 1'b0 ;
  assign n21005 = n1692 | n7726 ;
  assign n21006 = n21005 ^ n12209 ^ n326 ;
  assign n21007 = ( n733 & ~n7946 ) | ( n733 & n16164 ) | ( ~n7946 & n16164 ) ;
  assign n21008 = n17903 ^ n1605 ^ 1'b0 ;
  assign n21009 = n5154 & n21008 ;
  assign n21010 = n6798 & ~n15193 ;
  assign n21011 = n21010 ^ n20838 ^ 1'b0 ;
  assign n21012 = n9468 ^ n4222 ^ 1'b0 ;
  assign n21013 = n6232 | n21012 ;
  assign n21017 = n714 | n13467 ;
  assign n21014 = n6599 ^ n2656 ^ 1'b0 ;
  assign n21015 = n8214 & n21014 ;
  assign n21016 = n17142 & n21015 ;
  assign n21018 = n21017 ^ n21016 ^ 1'b0 ;
  assign n21019 = ~n3572 & n21018 ;
  assign n21020 = n2627 & n10600 ;
  assign n21021 = ( n5864 & n17654 ) | ( n5864 & ~n21020 ) | ( n17654 & ~n21020 ) ;
  assign n21022 = ~n8708 & n21021 ;
  assign n21023 = n21022 ^ n20431 ^ 1'b0 ;
  assign n21024 = n20386 ^ n11365 ^ n6866 ;
  assign n21025 = n21024 ^ n12500 ^ 1'b0 ;
  assign n21026 = n21023 & n21025 ;
  assign n21027 = ~n18850 & n21026 ;
  assign n21028 = n7326 & ~n10071 ;
  assign n21029 = n8174 ^ n5754 ^ n288 ;
  assign n21030 = n21029 ^ n8994 ^ 1'b0 ;
  assign n21031 = ~n21028 & n21030 ;
  assign n21034 = n12881 ^ n2851 ^ 1'b0 ;
  assign n21032 = n1758 & n3170 ;
  assign n21033 = ~n10369 & n21032 ;
  assign n21035 = n21034 ^ n21033 ^ 1'b0 ;
  assign n21036 = ( n6951 & ~n16668 ) | ( n6951 & n21035 ) | ( ~n16668 & n21035 ) ;
  assign n21037 = ~n15228 & n21036 ;
  assign n21038 = n21037 ^ n10405 ^ 1'b0 ;
  assign n21041 = ( n681 & ~n6772 ) | ( n681 & n7769 ) | ( ~n6772 & n7769 ) ;
  assign n21039 = ~n4751 & n12943 ;
  assign n21040 = ~n5760 & n21039 ;
  assign n21042 = n21041 ^ n21040 ^ n7237 ;
  assign n21043 = n1980 & n3587 ;
  assign n21044 = ~n18028 & n19494 ;
  assign n21045 = ~n3253 & n14262 ;
  assign n21046 = ~n14324 & n21045 ;
  assign n21053 = n1151 & ~n2856 ;
  assign n21054 = ~x216 & n2397 ;
  assign n21055 = ( ~n6213 & n21053 ) | ( ~n6213 & n21054 ) | ( n21053 & n21054 ) ;
  assign n21048 = ~n11262 & n16651 ;
  assign n21049 = n5465 | n8823 ;
  assign n21050 = n21049 ^ n6298 ^ 1'b0 ;
  assign n21051 = n21050 ^ n7897 ^ n1698 ;
  assign n21052 = n21048 | n21051 ;
  assign n21056 = n21055 ^ n21052 ^ 1'b0 ;
  assign n21057 = n2332 & n21056 ;
  assign n21047 = n11190 & ~n20384 ;
  assign n21058 = n21057 ^ n21047 ^ 1'b0 ;
  assign n21059 = n9686 | n21058 ;
  assign n21060 = n9735 ^ n5930 ^ 1'b0 ;
  assign n21061 = n20054 ^ n10352 ^ n2587 ;
  assign n21062 = ( n15609 & ~n15964 ) | ( n15609 & n21061 ) | ( ~n15964 & n21061 ) ;
  assign n21063 = n7080 | n21062 ;
  assign n21064 = n21060 & ~n21063 ;
  assign n21065 = n21064 ^ n13732 ^ n1850 ;
  assign n21066 = n4480 ^ n2257 ^ 1'b0 ;
  assign n21067 = ~n7499 & n21066 ;
  assign n21068 = n12485 ^ n5372 ^ 1'b0 ;
  assign n21069 = n7133 | n21068 ;
  assign n21070 = ( n3091 & ~n21067 ) | ( n3091 & n21069 ) | ( ~n21067 & n21069 ) ;
  assign n21071 = ~n5121 & n7658 ;
  assign n21072 = n21071 ^ n15756 ^ 1'b0 ;
  assign n21073 = n7972 & n21072 ;
  assign n21074 = ~n11874 & n15511 ;
  assign n21075 = n2984 ^ n1139 ^ 1'b0 ;
  assign n21076 = n21075 ^ n11353 ^ n10416 ;
  assign n21077 = n20611 | n21076 ;
  assign n21078 = n7102 | n21077 ;
  assign n21079 = n9838 ^ n4927 ^ x200 ;
  assign n21080 = ( n5575 & ~n6628 ) | ( n5575 & n9658 ) | ( ~n6628 & n9658 ) ;
  assign n21081 = n21079 & ~n21080 ;
  assign n21082 = n10812 ^ n3043 ^ 1'b0 ;
  assign n21083 = x219 & ~n21082 ;
  assign n21084 = n21083 ^ n15089 ^ 1'b0 ;
  assign n21085 = ( n8531 & ~n20686 ) | ( n8531 & n21084 ) | ( ~n20686 & n21084 ) ;
  assign n21086 = ~n20086 & n21085 ;
  assign n21087 = n19025 ^ n10876 ^ n8910 ;
  assign n21089 = ( n645 & n5278 ) | ( n645 & ~n5953 ) | ( n5278 & ~n5953 ) ;
  assign n21088 = n10056 & n10230 ;
  assign n21090 = n21089 ^ n21088 ^ 1'b0 ;
  assign n21091 = ~n1906 & n20899 ;
  assign n21092 = n7101 & n7443 ;
  assign n21093 = n21092 ^ n15181 ^ 1'b0 ;
  assign n21094 = n21091 | n21093 ;
  assign n21095 = n21094 ^ n20868 ^ 1'b0 ;
  assign n21096 = ( n3676 & n4985 ) | ( n3676 & n10464 ) | ( n4985 & n10464 ) ;
  assign n21097 = n6307 & ~n21096 ;
  assign n21098 = n15231 & n21097 ;
  assign n21109 = n4905 & n9607 ;
  assign n21099 = n3877 ^ n3422 ^ 1'b0 ;
  assign n21100 = n21099 ^ n11375 ^ n4346 ;
  assign n21102 = n879 & ~n15264 ;
  assign n21103 = n397 & n21102 ;
  assign n21104 = n21103 ^ n904 ^ 1'b0 ;
  assign n21105 = ~n6613 & n21104 ;
  assign n21101 = n7062 & ~n9332 ;
  assign n21106 = n21105 ^ n21101 ^ 1'b0 ;
  assign n21107 = n21106 ^ n5432 ^ 1'b0 ;
  assign n21108 = n21100 | n21107 ;
  assign n21110 = n21109 ^ n21108 ^ 1'b0 ;
  assign n21111 = n12310 ^ n637 ^ 1'b0 ;
  assign n21112 = ~n12824 & n21111 ;
  assign n21113 = n13892 & n21112 ;
  assign n21114 = ~n17428 & n21113 ;
  assign n21115 = n14481 & n17316 ;
  assign n21116 = ~n12800 & n21115 ;
  assign n21117 = n10312 ^ n1930 ^ 1'b0 ;
  assign n21118 = n19438 & ~n21117 ;
  assign n21119 = ~n5056 & n12209 ;
  assign n21120 = n20864 ^ n11666 ^ 1'b0 ;
  assign n21121 = n11706 & ~n21120 ;
  assign n21122 = n749 | n21121 ;
  assign n21123 = n10092 & ~n15703 ;
  assign n21124 = n21122 & n21123 ;
  assign n21125 = n21119 | n21124 ;
  assign n21126 = n13132 ^ n2190 ^ 1'b0 ;
  assign n21127 = ~n19650 & n21126 ;
  assign n21128 = ~n4616 & n8845 ;
  assign n21129 = n21128 ^ n2047 ^ 1'b0 ;
  assign n21130 = n3059 | n4917 ;
  assign n21131 = n4286 & ~n21130 ;
  assign n21132 = ( n7450 & ~n16757 ) | ( n7450 & n21131 ) | ( ~n16757 & n21131 ) ;
  assign n21136 = ( ~n455 & n3388 ) | ( ~n455 & n11937 ) | ( n3388 & n11937 ) ;
  assign n21133 = n4679 | n15098 ;
  assign n21134 = n565 & n9245 ;
  assign n21135 = ~n21133 & n21134 ;
  assign n21137 = n21136 ^ n21135 ^ n20269 ;
  assign n21138 = n12319 | n21005 ;
  assign n21139 = n19394 & n21138 ;
  assign n21140 = n10451 & ~n21139 ;
  assign n21141 = n15320 ^ n10255 ^ 1'b0 ;
  assign n21142 = ~n3922 & n18882 ;
  assign n21143 = n13952 & n21142 ;
  assign n21144 = ( n3215 & n13957 ) | ( n3215 & ~n16949 ) | ( n13957 & ~n16949 ) ;
  assign n21145 = n15123 ^ n1404 ^ 1'b0 ;
  assign n21146 = x101 & n8767 ;
  assign n21147 = ~n16510 & n21146 ;
  assign n21148 = n12271 & n12906 ;
  assign n21149 = n21148 ^ n4261 ^ 1'b0 ;
  assign n21150 = n21149 ^ n9960 ^ 1'b0 ;
  assign n21151 = n15856 ^ n11006 ^ n4803 ;
  assign n21152 = n21151 ^ n14145 ^ 1'b0 ;
  assign n21153 = n8848 & ~n14994 ;
  assign n21154 = n11594 ^ n3907 ^ 1'b0 ;
  assign n21155 = n18030 ^ n11553 ^ 1'b0 ;
  assign n21156 = n1070 & ~n21155 ;
  assign n21157 = n7214 ^ n5760 ^ 1'b0 ;
  assign n21158 = ~n10709 & n21157 ;
  assign n21159 = n5656 | n13641 ;
  assign n21160 = n21159 ^ n12797 ^ 1'b0 ;
  assign n21161 = n16865 ^ n4956 ^ 1'b0 ;
  assign n21162 = ( ~n7038 & n21160 ) | ( ~n7038 & n21161 ) | ( n21160 & n21161 ) ;
  assign n21163 = ( n1453 & ~n2445 ) | ( n1453 & n11878 ) | ( ~n2445 & n11878 ) ;
  assign n21164 = n7019 | n9530 ;
  assign n21165 = n21164 ^ n10121 ^ 1'b0 ;
  assign n21166 = n21165 ^ n10377 ^ 1'b0 ;
  assign n21167 = n15737 & ~n21166 ;
  assign n21168 = n13232 & n17483 ;
  assign n21169 = ~n20194 & n21168 ;
  assign n21170 = ( n747 & n2483 ) | ( n747 & n15194 ) | ( n2483 & n15194 ) ;
  assign n21171 = n5656 ^ n3982 ^ 1'b0 ;
  assign n21172 = n21170 | n21171 ;
  assign n21173 = n6373 ^ n3135 ^ 1'b0 ;
  assign n21174 = n21173 ^ n11904 ^ 1'b0 ;
  assign n21175 = n6559 ^ n2495 ^ 1'b0 ;
  assign n21176 = n2810 | n21175 ;
  assign n21177 = x30 & n294 ;
  assign n21178 = n21177 ^ n11864 ^ 1'b0 ;
  assign n21179 = ~n10625 & n21178 ;
  assign n21180 = n12429 ^ n9231 ^ 1'b0 ;
  assign n21181 = n7056 & n7660 ;
  assign n21182 = n21181 ^ n13521 ^ 1'b0 ;
  assign n21183 = n21182 ^ n6611 ^ 1'b0 ;
  assign n21184 = n14873 & n21183 ;
  assign n21185 = ( n3926 & ~n10572 ) | ( n3926 & n21184 ) | ( ~n10572 & n21184 ) ;
  assign n21186 = n12922 | n17169 ;
  assign n21187 = n16570 ^ n8865 ^ 1'b0 ;
  assign n21188 = n5549 | n13254 ;
  assign n21189 = n21188 ^ n8319 ^ 1'b0 ;
  assign n21190 = n19499 ^ x85 ^ 1'b0 ;
  assign n21191 = n21190 ^ n9236 ^ n734 ;
  assign n21192 = n2492 | n7768 ;
  assign n21193 = n11133 ^ n4094 ^ 1'b0 ;
  assign n21194 = n21192 | n21193 ;
  assign n21195 = n12069 & n14848 ;
  assign n21196 = n21195 ^ n13891 ^ 1'b0 ;
  assign n21197 = ~n4083 & n16119 ;
  assign n21198 = ~x82 & n21197 ;
  assign n21199 = ~n21196 & n21198 ;
  assign n21200 = n7282 | n13555 ;
  assign n21201 = n17387 & ~n21200 ;
  assign n21202 = n21201 ^ n15381 ^ 1'b0 ;
  assign n21203 = n11974 ^ n2947 ^ 1'b0 ;
  assign n21204 = ~n21202 & n21203 ;
  assign n21205 = n16479 ^ n16194 ^ 1'b0 ;
  assign n21206 = n2393 | n21205 ;
  assign n21207 = n21206 ^ n18147 ^ n9313 ;
  assign n21208 = n1928 | n2726 ;
  assign n21209 = ( ~n3402 & n5246 ) | ( ~n3402 & n10104 ) | ( n5246 & n10104 ) ;
  assign n21210 = n8956 ^ n7044 ^ n2333 ;
  assign n21211 = n21210 ^ n7767 ^ 1'b0 ;
  assign n21212 = n21209 & ~n21211 ;
  assign n21213 = n9103 | n17578 ;
  assign n21214 = n12785 | n21213 ;
  assign n21215 = n5637 & ~n6553 ;
  assign n21216 = n13756 & n21215 ;
  assign n21217 = n5721 | n21216 ;
  assign n21218 = n18303 | n21217 ;
  assign n21219 = ( ~n1763 & n3097 ) | ( ~n1763 & n13781 ) | ( n3097 & n13781 ) ;
  assign n21220 = n6397 ^ n940 ^ 1'b0 ;
  assign n21221 = n12029 ^ n1937 ^ 1'b0 ;
  assign n21222 = n21220 | n21221 ;
  assign n21223 = n21222 ^ n19222 ^ 1'b0 ;
  assign n21224 = n5115 | n16507 ;
  assign n21225 = n5282 | n21224 ;
  assign n21228 = n20210 ^ n5872 ^ 1'b0 ;
  assign n21229 = n2509 & ~n21228 ;
  assign n21230 = ( n11917 & n18831 ) | ( n11917 & ~n21229 ) | ( n18831 & ~n21229 ) ;
  assign n21231 = n21230 ^ n10008 ^ 1'b0 ;
  assign n21226 = n7567 & ~n10231 ;
  assign n21227 = n21226 ^ n911 ^ 1'b0 ;
  assign n21232 = n21231 ^ n21227 ^ 1'b0 ;
  assign n21233 = n19695 ^ n16009 ^ 1'b0 ;
  assign n21234 = n21230 | n21233 ;
  assign n21235 = n13671 & ~n21234 ;
  assign n21236 = ~n1752 & n21235 ;
  assign n21237 = n959 | n3891 ;
  assign n21238 = n6332 & n9869 ;
  assign n21239 = n3116 & ~n9078 ;
  assign n21240 = n21239 ^ x111 ^ 1'b0 ;
  assign n21241 = n9054 | n20987 ;
  assign n21242 = n21241 ^ n16238 ^ 1'b0 ;
  assign n21243 = n21242 ^ n8030 ^ 1'b0 ;
  assign n21244 = n18736 ^ n15028 ^ n2930 ;
  assign n21245 = n11457 ^ n5503 ^ n3852 ;
  assign n21246 = ~n20464 & n21245 ;
  assign n21247 = n10948 & n21246 ;
  assign n21248 = n935 & ~n2203 ;
  assign n21249 = n296 & n21248 ;
  assign n21250 = n21234 ^ n17293 ^ 1'b0 ;
  assign n21251 = ~n365 & n12592 ;
  assign n21252 = ( n5140 & n5571 ) | ( n5140 & ~n18380 ) | ( n5571 & ~n18380 ) ;
  assign n21253 = n21252 ^ n17747 ^ 1'b0 ;
  assign n21254 = n21252 & n21253 ;
  assign n21256 = n5711 | n9451 ;
  assign n21257 = n1515 & ~n21256 ;
  assign n21255 = n12464 | n15305 ;
  assign n21258 = n21257 ^ n21255 ^ 1'b0 ;
  assign n21259 = n21254 & ~n21258 ;
  assign n21260 = n14456 & n21259 ;
  assign n21261 = n2949 & n12529 ;
  assign n21262 = n3698 & n11153 ;
  assign n21263 = n13035 ^ n12869 ^ 1'b0 ;
  assign n21264 = n1217 & n21263 ;
  assign n21265 = n21264 ^ n16910 ^ 1'b0 ;
  assign n21266 = n5864 & ~n21265 ;
  assign n21269 = n5949 ^ n2909 ^ 1'b0 ;
  assign n21270 = n5765 | n21269 ;
  assign n21271 = n21270 ^ n7175 ^ n1541 ;
  assign n21272 = n21271 ^ n7573 ^ 1'b0 ;
  assign n21273 = n18337 & n21272 ;
  assign n21274 = n21273 ^ n3939 ^ 1'b0 ;
  assign n21267 = n4241 & n7672 ;
  assign n21268 = n3315 & n21267 ;
  assign n21275 = n21274 ^ n21268 ^ n4402 ;
  assign n21276 = n8567 ^ n1817 ^ 1'b0 ;
  assign n21277 = ~n3511 & n15242 ;
  assign n21278 = n21277 ^ n20843 ^ 1'b0 ;
  assign n21279 = n21278 ^ n14708 ^ n6597 ;
  assign n21280 = n298 & ~n3903 ;
  assign n21281 = n1140 & ~n19536 ;
  assign n21283 = n9968 ^ n3104 ^ 1'b0 ;
  assign n21282 = n2344 & ~n15321 ;
  assign n21284 = n21283 ^ n21282 ^ 1'b0 ;
  assign n21285 = n21284 ^ n21138 ^ 1'b0 ;
  assign n21286 = n12091 ^ x30 ^ 1'b0 ;
  assign n21287 = n3185 & ~n21286 ;
  assign n21288 = n9269 & n21287 ;
  assign n21289 = n14679 ^ n12820 ^ n3882 ;
  assign n21290 = n8636 & n16192 ;
  assign n21291 = ( n1777 & n9528 ) | ( n1777 & ~n16586 ) | ( n9528 & ~n16586 ) ;
  assign n21292 = n14379 ^ n12763 ^ 1'b0 ;
  assign n21293 = n15383 ^ n11479 ^ 1'b0 ;
  assign n21294 = ( n2943 & n12228 ) | ( n2943 & n21293 ) | ( n12228 & n21293 ) ;
  assign n21295 = n20127 ^ n17192 ^ n10016 ;
  assign n21296 = n6163 ^ n5304 ^ 1'b0 ;
  assign n21297 = n17176 ^ x86 ^ 1'b0 ;
  assign n21298 = n21296 | n21297 ;
  assign n21299 = ~n11873 & n14244 ;
  assign n21300 = n21299 ^ n19155 ^ 1'b0 ;
  assign n21301 = n16953 ^ n889 ^ 1'b0 ;
  assign n21302 = n17755 | n21301 ;
  assign n21303 = n1486 & n7745 ;
  assign n21304 = n9528 ^ n2544 ^ 1'b0 ;
  assign n21305 = ( n4056 & ~n8077 ) | ( n4056 & n11447 ) | ( ~n8077 & n11447 ) ;
  assign n21306 = n16264 | n20134 ;
  assign n21307 = ~n8548 & n9500 ;
  assign n21308 = ~n21202 & n21307 ;
  assign n21309 = n21308 ^ n11694 ^ 1'b0 ;
  assign n21310 = n1922 & n21309 ;
  assign n21311 = n2202 & n21310 ;
  assign n21312 = n15930 ^ n3888 ^ n2645 ;
  assign n21313 = ~n1582 & n17000 ;
  assign n21315 = n9245 ^ n2248 ^ 1'b0 ;
  assign n21316 = n10129 & n21315 ;
  assign n21314 = n6342 & ~n20962 ;
  assign n21317 = n21316 ^ n21314 ^ 1'b0 ;
  assign n21318 = ( n12750 & n15694 ) | ( n12750 & n18593 ) | ( n15694 & n18593 ) ;
  assign n21319 = n8805 ^ n5059 ^ 1'b0 ;
  assign n21320 = n7070 & ~n21319 ;
  assign n21321 = n21320 ^ n5135 ^ 1'b0 ;
  assign n21322 = n8823 ^ n2489 ^ 1'b0 ;
  assign n21323 = n3273 & ~n21322 ;
  assign n21324 = n16900 ^ n3104 ^ 1'b0 ;
  assign n21325 = n3119 & n10222 ;
  assign n21326 = n21324 & n21325 ;
  assign n21327 = ~n1442 & n12371 ;
  assign n21328 = n21327 ^ n6884 ^ 1'b0 ;
  assign n21330 = n20574 ^ n2673 ^ n2130 ;
  assign n21329 = n16966 & n17424 ;
  assign n21331 = n21330 ^ n21329 ^ 1'b0 ;
  assign n21332 = n16924 ^ n2106 ^ 1'b0 ;
  assign n21333 = n6379 ^ n2416 ^ 1'b0 ;
  assign n21334 = n650 & ~n21333 ;
  assign n21335 = n8808 ^ n7469 ^ 1'b0 ;
  assign n21336 = n21334 & ~n21335 ;
  assign n21337 = n5934 & n10168 ;
  assign n21338 = ~n21336 & n21337 ;
  assign n21339 = n4920 & ~n8669 ;
  assign n21340 = n21338 & n21339 ;
  assign n21351 = n10185 ^ n4128 ^ 1'b0 ;
  assign n21350 = n19914 ^ n3210 ^ 1'b0 ;
  assign n21348 = ( n3794 & n4144 ) | ( n3794 & n5422 ) | ( n4144 & n5422 ) ;
  assign n21341 = n9295 ^ n3551 ^ 1'b0 ;
  assign n21342 = n2357 & n5729 ;
  assign n21343 = n3985 & n21342 ;
  assign n21344 = n21343 ^ n3913 ^ 1'b0 ;
  assign n21345 = n2144 | n21344 ;
  assign n21346 = n21341 | n21345 ;
  assign n21347 = ~x83 & n21346 ;
  assign n21349 = n21348 ^ n21347 ^ 1'b0 ;
  assign n21352 = n21351 ^ n21350 ^ n21349 ;
  assign n21353 = n8719 & n9249 ;
  assign n21354 = n2486 | n7490 ;
  assign n21355 = n21354 ^ n17190 ^ 1'b0 ;
  assign n21356 = n3236 & ~n19833 ;
  assign n21357 = n10289 ^ n2997 ^ 1'b0 ;
  assign n21358 = n8370 ^ n5145 ^ 1'b0 ;
  assign n21359 = n21358 ^ n2234 ^ n1665 ;
  assign n21360 = ~n14919 & n17166 ;
  assign n21361 = ~n3249 & n21360 ;
  assign n21362 = ( n5626 & n13635 ) | ( n5626 & ~n17114 ) | ( n13635 & ~n17114 ) ;
  assign n21363 = n21361 | n21362 ;
  assign n21364 = n21363 ^ n11158 ^ 1'b0 ;
  assign n21365 = n16952 & n21364 ;
  assign n21366 = n1736 & ~n8957 ;
  assign n21367 = n21366 ^ n6188 ^ 1'b0 ;
  assign n21368 = n21367 ^ n2637 ^ 1'b0 ;
  assign n21369 = n21365 & ~n21368 ;
  assign n21370 = n17422 ^ n4229 ^ 1'b0 ;
  assign n21371 = n11498 & n21370 ;
  assign n21372 = ~n19656 & n21371 ;
  assign n21373 = n11252 ^ n1312 ^ 1'b0 ;
  assign n21374 = n4560 & ~n21373 ;
  assign n21375 = n21374 ^ n17549 ^ 1'b0 ;
  assign n21376 = n9772 ^ x158 ^ 1'b0 ;
  assign n21377 = n778 | n21376 ;
  assign n21378 = n7786 | n21377 ;
  assign n21379 = n21378 ^ n13793 ^ 1'b0 ;
  assign n21380 = ~n6672 & n15899 ;
  assign n21381 = n17080 & n21380 ;
  assign n21382 = n5099 ^ n4216 ^ 1'b0 ;
  assign n21383 = n21381 | n21382 ;
  assign n21384 = n15054 ^ n5271 ^ 1'b0 ;
  assign n21385 = n15701 ^ n8765 ^ n3043 ;
  assign n21386 = ( n4194 & n10475 ) | ( n4194 & ~n21385 ) | ( n10475 & ~n21385 ) ;
  assign n21387 = ~n5793 & n12802 ;
  assign n21388 = n21387 ^ n12023 ^ 1'b0 ;
  assign n21390 = ~n4191 & n8415 ;
  assign n21391 = n4298 | n21390 ;
  assign n21392 = n21391 ^ n12783 ^ 1'b0 ;
  assign n21389 = n753 | n8554 ;
  assign n21393 = n21392 ^ n21389 ^ n10118 ;
  assign n21394 = ( n3215 & ~n21388 ) | ( n3215 & n21393 ) | ( ~n21388 & n21393 ) ;
  assign n21395 = n8107 ^ n2997 ^ 1'b0 ;
  assign n21396 = n12417 & ~n14913 ;
  assign n21397 = n5209 & ~n21396 ;
  assign n21398 = n21397 ^ n7201 ^ 1'b0 ;
  assign n21399 = ~n723 & n8560 ;
  assign n21400 = n21399 ^ n3016 ^ 1'b0 ;
  assign n21401 = n15869 ^ n7565 ^ 1'b0 ;
  assign n21402 = n1959 & n21401 ;
  assign n21403 = n10694 | n16950 ;
  assign n21404 = n21403 ^ n5963 ^ 1'b0 ;
  assign n21405 = ~n2214 & n13538 ;
  assign n21406 = n11408 & n21405 ;
  assign n21407 = n2108 | n8270 ;
  assign n21408 = n2099 | n7106 ;
  assign n21409 = n21408 ^ n16296 ^ 1'b0 ;
  assign n21410 = n21232 ^ n1079 ^ 1'b0 ;
  assign n21412 = n16305 ^ n1689 ^ 1'b0 ;
  assign n21413 = n6276 & n21412 ;
  assign n21411 = n2430 | n4704 ;
  assign n21414 = n21413 ^ n21411 ^ 1'b0 ;
  assign n21415 = n5778 & n21414 ;
  assign n21417 = n8618 ^ n2224 ^ 1'b0 ;
  assign n21416 = ~n1418 & n13393 ;
  assign n21418 = n21417 ^ n21416 ^ 1'b0 ;
  assign n21419 = n4373 ^ n3976 ^ x40 ;
  assign n21420 = n17985 & n21419 ;
  assign n21421 = ~n1175 & n2991 ;
  assign n21422 = n673 | n20141 ;
  assign n21423 = n7895 ^ n3791 ^ 1'b0 ;
  assign n21424 = n21422 | n21423 ;
  assign n21425 = n11689 | n21424 ;
  assign n21426 = n21425 ^ n473 ^ 1'b0 ;
  assign n21427 = n5177 ^ n2471 ^ 1'b0 ;
  assign n21428 = n1138 & n21427 ;
  assign n21429 = ~n8839 & n21428 ;
  assign n21430 = n21429 ^ n13159 ^ 1'b0 ;
  assign n21431 = n8484 & n21430 ;
  assign n21432 = n21431 ^ n7859 ^ 1'b0 ;
  assign n21433 = n13151 ^ n2553 ^ 1'b0 ;
  assign n21434 = ~n15265 & n21433 ;
  assign n21435 = n4732 | n8090 ;
  assign n21436 = n21434 | n21435 ;
  assign n21437 = n21436 ^ n13383 ^ 1'b0 ;
  assign n21438 = n2966 & ~n17725 ;
  assign n21439 = ~n17595 & n21438 ;
  assign n21440 = ~n7795 & n10333 ;
  assign n21441 = n4954 & n21440 ;
  assign n21442 = n4042 | n8382 ;
  assign n21443 = n16029 ^ n10973 ^ 1'b0 ;
  assign n21444 = n5569 | n20737 ;
  assign n21445 = n2325 | n21444 ;
  assign n21446 = n739 & ~n4993 ;
  assign n21447 = n9942 & ~n21446 ;
  assign n21448 = n20673 & n21447 ;
  assign n21449 = n15147 ^ n11064 ^ 1'b0 ;
  assign n21450 = n19151 & n21449 ;
  assign n21451 = n21450 ^ n3307 ^ 1'b0 ;
  assign n21452 = n14406 ^ n5689 ^ 1'b0 ;
  assign n21453 = n5455 & ~n21452 ;
  assign n21454 = n19532 & n21453 ;
  assign n21455 = n21443 ^ n2305 ^ 1'b0 ;
  assign n21456 = ~n16650 & n20531 ;
  assign n21457 = n21456 ^ n6481 ^ 1'b0 ;
  assign n21458 = ( n2810 & n7091 ) | ( n2810 & ~n21457 ) | ( n7091 & ~n21457 ) ;
  assign n21459 = n7912 & ~n21458 ;
  assign n21463 = n8403 & n11134 ;
  assign n21464 = n21463 ^ n7165 ^ 1'b0 ;
  assign n21460 = n4229 ^ n2054 ^ 1'b0 ;
  assign n21461 = ( n4001 & n11284 ) | ( n4001 & n21460 ) | ( n11284 & n21460 ) ;
  assign n21462 = n10322 | n21461 ;
  assign n21465 = n21464 ^ n21462 ^ n6563 ;
  assign n21467 = n5630 ^ n3207 ^ n677 ;
  assign n21468 = n21467 ^ n5468 ^ 1'b0 ;
  assign n21466 = ~n9221 & n14123 ;
  assign n21469 = n21468 ^ n21466 ^ 1'b0 ;
  assign n21470 = n2588 | n19876 ;
  assign n21471 = n7844 & ~n21470 ;
  assign n21472 = n4800 ^ n3056 ^ n2118 ;
  assign n21473 = n14143 ^ n10280 ^ 1'b0 ;
  assign n21474 = n4764 ^ n1829 ^ 1'b0 ;
  assign n21475 = n4907 | n21474 ;
  assign n21476 = ~n15564 & n21475 ;
  assign n21477 = n3598 & ~n20505 ;
  assign n21478 = n14965 & n21477 ;
  assign n21479 = n17836 ^ n3756 ^ n972 ;
  assign n21480 = x158 | n10040 ;
  assign n21481 = n15118 ^ n4385 ^ n663 ;
  assign n21482 = n5910 | n11030 ;
  assign n21483 = ( n6690 & n21481 ) | ( n6690 & ~n21482 ) | ( n21481 & ~n21482 ) ;
  assign n21484 = n9200 ^ n6643 ^ 1'b0 ;
  assign n21485 = ~n15087 & n21484 ;
  assign n21486 = ( x153 & n4074 ) | ( x153 & n21485 ) | ( n4074 & n21485 ) ;
  assign n21487 = ( n449 & n2548 ) | ( n449 & ~n9851 ) | ( n2548 & ~n9851 ) ;
  assign n21488 = n10593 & ~n21487 ;
  assign n21489 = n21488 ^ n11061 ^ 1'b0 ;
  assign n21490 = ( n7703 & n11721 ) | ( n7703 & ~n17517 ) | ( n11721 & ~n17517 ) ;
  assign n21491 = n12609 ^ n7813 ^ 1'b0 ;
  assign n21492 = n21491 ^ n14461 ^ 1'b0 ;
  assign n21493 = n21490 & ~n21492 ;
  assign n21494 = n10636 ^ n7914 ^ 1'b0 ;
  assign n21495 = n21493 | n21494 ;
  assign n21496 = ( n7047 & n9075 ) | ( n7047 & n21495 ) | ( n9075 & n21495 ) ;
  assign n21497 = n1768 & n18336 ;
  assign n21498 = n8938 & n21497 ;
  assign n21499 = n7519 & ~n21498 ;
  assign n21500 = n8953 & n14325 ;
  assign n21501 = n3749 | n7308 ;
  assign n21502 = n13053 ^ n3126 ^ 1'b0 ;
  assign n21503 = n18116 ^ n17532 ^ n8997 ;
  assign n21508 = n8131 | n19820 ;
  assign n21504 = ( n918 & n1486 ) | ( n918 & ~n3597 ) | ( n1486 & ~n3597 ) ;
  assign n21505 = n2228 & ~n2751 ;
  assign n21506 = ~n21504 & n21505 ;
  assign n21507 = x22 & ~n21506 ;
  assign n21509 = n21508 ^ n21507 ^ 1'b0 ;
  assign n21510 = ~n9465 & n21509 ;
  assign n21511 = n21510 ^ n14777 ^ 1'b0 ;
  assign n21512 = n18589 & ~n21511 ;
  assign n21513 = ( n3093 & n8529 ) | ( n3093 & ~n8690 ) | ( n8529 & ~n8690 ) ;
  assign n21514 = n5507 & n20864 ;
  assign n21515 = n21514 ^ n15307 ^ 1'b0 ;
  assign n21516 = ( n10522 & ~n12064 ) | ( n10522 & n21515 ) | ( ~n12064 & n21515 ) ;
  assign n21517 = n21516 ^ n14660 ^ 1'b0 ;
  assign n21518 = n1307 & ~n18398 ;
  assign n21519 = n21518 ^ n5037 ^ 1'b0 ;
  assign n21520 = n4677 & n18874 ;
  assign n21521 = n21520 ^ n12864 ^ 1'b0 ;
  assign n21522 = n10569 & n21521 ;
  assign n21523 = n5695 | n6047 ;
  assign n21524 = n6972 & n21523 ;
  assign n21525 = n8957 ^ n6312 ^ 1'b0 ;
  assign n21526 = n21524 & ~n21525 ;
  assign n21527 = n21526 ^ n10032 ^ n4076 ;
  assign n21528 = ~n12009 & n21527 ;
  assign n21529 = ( n11056 & n21372 ) | ( n11056 & n21528 ) | ( n21372 & n21528 ) ;
  assign n21530 = n20755 ^ n1873 ^ 1'b0 ;
  assign n21532 = n13943 ^ n7499 ^ 1'b0 ;
  assign n21533 = n5215 & n21532 ;
  assign n21531 = n19276 ^ n1653 ^ 1'b0 ;
  assign n21534 = n21533 ^ n21531 ^ n647 ;
  assign n21537 = n10226 & ~n15915 ;
  assign n21535 = ~n3761 & n19715 ;
  assign n21536 = n21535 ^ n3610 ^ 1'b0 ;
  assign n21538 = n21537 ^ n21536 ^ 1'b0 ;
  assign n21539 = n8800 ^ n3555 ^ 1'b0 ;
  assign n21540 = n11093 | n21539 ;
  assign n21541 = n11466 | n13988 ;
  assign n21542 = n13988 & ~n21541 ;
  assign n21543 = n3404 & n21542 ;
  assign n21544 = ~n11039 & n21543 ;
  assign n21545 = n11039 & n21544 ;
  assign n21546 = ~n11215 & n21545 ;
  assign n21547 = ~n21540 & n21546 ;
  assign n21548 = n8830 ^ n5663 ^ n3027 ;
  assign n21549 = n12877 ^ n10183 ^ 1'b0 ;
  assign n21550 = n21548 & n21549 ;
  assign n21551 = n650 ^ x60 ^ 1'b0 ;
  assign n21552 = n21550 | n21551 ;
  assign n21553 = n21552 ^ n5428 ^ 1'b0 ;
  assign n21555 = n4108 ^ n1155 ^ 1'b0 ;
  assign n21556 = ~n5730 & n21555 ;
  assign n21554 = n2958 & ~n15551 ;
  assign n21557 = n21556 ^ n21554 ^ n9011 ;
  assign n21558 = n21557 ^ n10585 ^ 1'b0 ;
  assign n21559 = n12905 ^ x61 ^ 1'b0 ;
  assign n21560 = ( ~n1000 & n5515 ) | ( ~n1000 & n7371 ) | ( n5515 & n7371 ) ;
  assign n21561 = n8643 ^ n4189 ^ 1'b0 ;
  assign n21562 = n21560 & n21561 ;
  assign n21563 = n21562 ^ n14673 ^ n1871 ;
  assign n21564 = ( ~n1455 & n3362 ) | ( ~n1455 & n4203 ) | ( n3362 & n4203 ) ;
  assign n21565 = ( n17405 & ~n17488 ) | ( n17405 & n21564 ) | ( ~n17488 & n21564 ) ;
  assign n21566 = n17991 & n21565 ;
  assign n21567 = n21566 ^ n20146 ^ 1'b0 ;
  assign n21568 = n18087 ^ n12822 ^ 1'b0 ;
  assign n21569 = ~n12097 & n21568 ;
  assign n21570 = n9652 ^ n814 ^ 1'b0 ;
  assign n21571 = ~n18613 & n21570 ;
  assign n21572 = ~n1553 & n2966 ;
  assign n21573 = n21572 ^ n12671 ^ n11448 ;
  assign n21574 = ~n17616 & n20357 ;
  assign n21575 = n21574 ^ n5139 ^ 1'b0 ;
  assign n21576 = n21573 & ~n21575 ;
  assign n21577 = n21576 ^ n5399 ^ 1'b0 ;
  assign n21578 = n4389 & n5162 ;
  assign n21579 = n9913 ^ n6745 ^ 1'b0 ;
  assign n21580 = n18910 ^ n10578 ^ 1'b0 ;
  assign n21581 = ~n21579 & n21580 ;
  assign n21582 = x62 & n21581 ;
  assign n21583 = n21582 ^ n1256 ^ 1'b0 ;
  assign n21584 = n21583 ^ n18600 ^ 1'b0 ;
  assign n21585 = n8729 | n21584 ;
  assign n21586 = n1889 & n21585 ;
  assign n21587 = n455 | n17525 ;
  assign n21591 = n4907 ^ n2307 ^ n1500 ;
  assign n21592 = ( ~n1457 & n2376 ) | ( ~n1457 & n21591 ) | ( n2376 & n21591 ) ;
  assign n21588 = n11448 ^ n4981 ^ 1'b0 ;
  assign n21589 = ~n3534 & n21588 ;
  assign n21590 = ( ~n13220 & n17728 ) | ( ~n13220 & n21589 ) | ( n17728 & n21589 ) ;
  assign n21593 = n21592 ^ n21590 ^ 1'b0 ;
  assign n21594 = n860 & ~n13278 ;
  assign n21595 = n21594 ^ n18738 ^ 1'b0 ;
  assign n21596 = ~n4184 & n17655 ;
  assign n21597 = n21596 ^ n2827 ^ 1'b0 ;
  assign n21598 = ~n3273 & n4126 ;
  assign n21599 = n8567 ^ n7726 ^ 1'b0 ;
  assign n21600 = n4907 & n6432 ;
  assign n21601 = n16684 & ~n21600 ;
  assign n21602 = n9934 ^ n9428 ^ 1'b0 ;
  assign n21603 = n7049 & n21602 ;
  assign n21604 = n21603 ^ n19510 ^ 1'b0 ;
  assign n21605 = ~n5954 & n21604 ;
  assign n21606 = n12864 ^ n8648 ^ 1'b0 ;
  assign n21607 = n21606 ^ n12121 ^ n9993 ;
  assign n21608 = n15395 ^ n8340 ^ n5598 ;
  assign n21609 = n21608 ^ n5786 ^ 1'b0 ;
  assign n21610 = ( n4081 & n12651 ) | ( n4081 & ~n21609 ) | ( n12651 & ~n21609 ) ;
  assign n21611 = n17948 ^ n16560 ^ n1528 ;
  assign n21612 = ( ~x84 & n2618 ) | ( ~x84 & n21611 ) | ( n2618 & n21611 ) ;
  assign n21613 = n2725 & ~n3198 ;
  assign n21614 = ~n12131 & n21613 ;
  assign n21615 = n7206 | n8945 ;
  assign n21616 = n21615 ^ n4078 ^ 1'b0 ;
  assign n21617 = n12746 | n21616 ;
  assign n21618 = n13297 | n21617 ;
  assign n21619 = n10547 ^ n1899 ^ 1'b0 ;
  assign n21620 = n8548 | n21619 ;
  assign n21621 = n21620 ^ n18675 ^ 1'b0 ;
  assign n21622 = n16711 ^ n6372 ^ 1'b0 ;
  assign n21623 = ~n20805 & n21622 ;
  assign n21624 = n20304 | n21607 ;
  assign n21625 = n9286 ^ x183 ^ 1'b0 ;
  assign n21626 = n18544 ^ x15 ^ 1'b0 ;
  assign n21627 = n21626 ^ n884 ^ 1'b0 ;
  assign n21628 = ~n940 & n10223 ;
  assign n21629 = n21628 ^ n3776 ^ 1'b0 ;
  assign n21630 = ( ~n776 & n12218 ) | ( ~n776 & n21629 ) | ( n12218 & n21629 ) ;
  assign n21631 = n19254 | n21630 ;
  assign n21632 = n21627 & ~n21631 ;
  assign n21633 = n16237 ^ n749 ^ 1'b0 ;
  assign n21634 = n11518 & n21633 ;
  assign n21635 = n21634 ^ n15489 ^ 1'b0 ;
  assign n21636 = n8783 | n15483 ;
  assign n21637 = n5853 & n13775 ;
  assign n21638 = ~n10742 & n21637 ;
  assign n21639 = ( ~n315 & n21636 ) | ( ~n315 & n21638 ) | ( n21636 & n21638 ) ;
  assign n21640 = n6235 & ~n16826 ;
  assign n21641 = n21640 ^ x13 ^ 1'b0 ;
  assign n21642 = n2378 & ~n2538 ;
  assign n21643 = n21642 ^ n18434 ^ 1'b0 ;
  assign n21644 = n21643 ^ x108 ^ 1'b0 ;
  assign n21646 = n9761 ^ n2382 ^ 1'b0 ;
  assign n21645 = ~n6606 & n18581 ;
  assign n21647 = n21646 ^ n21645 ^ 1'b0 ;
  assign n21648 = n18935 ^ n7380 ^ 1'b0 ;
  assign n21649 = n18429 & ~n21648 ;
  assign n21650 = n10378 & n21649 ;
  assign n21651 = ~n16764 & n21650 ;
  assign n21652 = n5864 & n16018 ;
  assign n21653 = n14192 ^ n3104 ^ 1'b0 ;
  assign n21654 = n21652 & n21653 ;
  assign n21655 = ~n5326 & n12705 ;
  assign n21656 = n21654 & n21655 ;
  assign n21657 = n7587 & n21656 ;
  assign n21658 = n4985 & n21657 ;
  assign n21659 = n4338 & ~n8688 ;
  assign n21660 = n21659 ^ n17380 ^ n1998 ;
  assign n21661 = ( n3570 & n5733 ) | ( n3570 & n9091 ) | ( n5733 & n9091 ) ;
  assign n21662 = n4287 & ~n8960 ;
  assign n21663 = n14784 ^ n9713 ^ 1'b0 ;
  assign n21664 = n519 & ~n21663 ;
  assign n21665 = n12828 | n16562 ;
  assign n21666 = n14452 & ~n21665 ;
  assign n21667 = n19706 ^ n9127 ^ n8051 ;
  assign n21668 = n2277 | n13635 ;
  assign n21669 = n15593 & ~n21668 ;
  assign n21670 = n6811 ^ n5108 ^ 1'b0 ;
  assign n21671 = ~n4361 & n21670 ;
  assign n21672 = n16572 & n21671 ;
  assign n21673 = n21672 ^ n9263 ^ 1'b0 ;
  assign n21674 = n634 | n6338 ;
  assign n21675 = n21674 ^ n9575 ^ 1'b0 ;
  assign n21676 = ~n2581 & n18650 ;
  assign n21677 = ~n21675 & n21676 ;
  assign n21678 = ( n3959 & n5626 ) | ( n3959 & n21677 ) | ( n5626 & n21677 ) ;
  assign n21679 = n349 ^ x85 ^ 1'b0 ;
  assign n21680 = n4569 | n21679 ;
  assign n21681 = n13458 & n21680 ;
  assign n21682 = n21681 ^ n9364 ^ 1'b0 ;
  assign n21683 = n1360 & n21682 ;
  assign n21687 = ~n2869 & n7021 ;
  assign n21688 = n4995 & ~n21687 ;
  assign n21689 = n21688 ^ n7122 ^ 1'b0 ;
  assign n21684 = n4218 & ~n13495 ;
  assign n21685 = n11798 & n21684 ;
  assign n21686 = n15043 & ~n21685 ;
  assign n21690 = n21689 ^ n21686 ^ 1'b0 ;
  assign n21691 = n13356 & ~n19364 ;
  assign n21692 = ~n3333 & n21691 ;
  assign n21693 = ~n4610 & n17820 ;
  assign n21694 = n21693 ^ n10755 ^ 1'b0 ;
  assign n21695 = ( x164 & n4150 ) | ( x164 & ~n8472 ) | ( n4150 & ~n8472 ) ;
  assign n21696 = n377 | n10768 ;
  assign n21697 = n21696 ^ n4157 ^ 1'b0 ;
  assign n21698 = n21697 ^ n14481 ^ 1'b0 ;
  assign n21699 = n21695 & ~n21698 ;
  assign n21700 = n5874 ^ n3790 ^ 1'b0 ;
  assign n21701 = n3822 & n15490 ;
  assign n21702 = ~n6821 & n21701 ;
  assign n21703 = n7928 | n21702 ;
  assign n21704 = ~n2823 & n6435 ;
  assign n21705 = n21704 ^ n6655 ^ 1'b0 ;
  assign n21706 = n21705 ^ n15255 ^ n2178 ;
  assign n21722 = n2437 & n7016 ;
  assign n21723 = ~n7016 & n21722 ;
  assign n21724 = n5693 | n20809 ;
  assign n21725 = n20809 & ~n21724 ;
  assign n21726 = n2059 | n11312 ;
  assign n21727 = ~n21725 & n21726 ;
  assign n21728 = n21723 & n21727 ;
  assign n21729 = n18997 | n21728 ;
  assign n21707 = n9297 ^ n3547 ^ n506 ;
  assign n21708 = ( n4524 & ~n5918 ) | ( n4524 & n21707 ) | ( ~n5918 & n21707 ) ;
  assign n21709 = n18387 | n21708 ;
  assign n21714 = n4582 & n5354 ;
  assign n21710 = n15646 ^ n1855 ^ 1'b0 ;
  assign n21711 = n2896 | n21710 ;
  assign n21712 = x101 & ~n21711 ;
  assign n21713 = n21712 ^ n1499 ^ 1'b0 ;
  assign n21715 = n21714 ^ n21713 ^ 1'b0 ;
  assign n21716 = n4641 & n21715 ;
  assign n21717 = ~n21709 & n21716 ;
  assign n21718 = ~n3376 & n8892 ;
  assign n21719 = n21717 | n21718 ;
  assign n21720 = n21717 & ~n21719 ;
  assign n21721 = n8411 | n21720 ;
  assign n21730 = n21729 ^ n21721 ^ 1'b0 ;
  assign n21731 = ~n3036 & n3225 ;
  assign n21732 = n2826 & n21731 ;
  assign n21733 = ( ~n1435 & n12133 ) | ( ~n1435 & n21732 ) | ( n12133 & n21732 ) ;
  assign n21734 = n6134 & n6737 ;
  assign n21735 = n21733 | n21734 ;
  assign n21736 = n16725 | n21735 ;
  assign n21737 = n7643 & n16630 ;
  assign n21738 = n6671 ^ n5255 ^ 1'b0 ;
  assign n21739 = ~n6762 & n21738 ;
  assign n21740 = ( n1622 & ~n2782 ) | ( n1622 & n8001 ) | ( ~n2782 & n8001 ) ;
  assign n21741 = n21739 & n21740 ;
  assign n21742 = ~n21737 & n21741 ;
  assign n21743 = n14592 ^ n8549 ^ 1'b0 ;
  assign n21744 = n7297 & ~n21743 ;
  assign n21745 = n21744 ^ n3911 ^ 1'b0 ;
  assign n21746 = n2590 & n10886 ;
  assign n21747 = n8966 & n21746 ;
  assign n21748 = ~n9170 & n21747 ;
  assign n21749 = ~n917 & n16119 ;
  assign n21750 = n9445 ^ n4574 ^ 1'b0 ;
  assign n21751 = n21749 & n21750 ;
  assign n21752 = n12048 & n21751 ;
  assign n21753 = ~n4450 & n16644 ;
  assign n21754 = n14122 ^ n6397 ^ 1'b0 ;
  assign n21755 = ~n17290 & n21754 ;
  assign n21756 = ( n8129 & n13609 ) | ( n8129 & n21755 ) | ( n13609 & n21755 ) ;
  assign n21757 = ~n2029 & n21756 ;
  assign n21758 = n21757 ^ n6352 ^ 1'b0 ;
  assign n21759 = n21753 | n21758 ;
  assign n21760 = ~n2480 & n9562 ;
  assign n21761 = ~n1110 & n21760 ;
  assign n21762 = n21761 ^ n6100 ^ 1'b0 ;
  assign n21763 = n14547 ^ n4773 ^ 1'b0 ;
  assign n21764 = ~n3278 & n10895 ;
  assign n21765 = n21764 ^ n15694 ^ 1'b0 ;
  assign n21766 = n21763 & ~n21765 ;
  assign n21767 = ( ~n1130 & n5339 ) | ( ~n1130 & n18418 ) | ( n5339 & n18418 ) ;
  assign n21768 = ~n3943 & n13909 ;
  assign n21769 = n940 | n10928 ;
  assign n21770 = n2336 | n21769 ;
  assign n21771 = n13544 ^ n3785 ^ 1'b0 ;
  assign n21772 = n7647 | n21771 ;
  assign n21773 = n21770 | n21772 ;
  assign n21774 = ~n21768 & n21773 ;
  assign n21775 = n21774 ^ n1263 ^ 1'b0 ;
  assign n21776 = ( ~n369 & n21767 ) | ( ~n369 & n21775 ) | ( n21767 & n21775 ) ;
  assign n21777 = n12900 ^ n7532 ^ 1'b0 ;
  assign n21778 = ~n6267 & n10521 ;
  assign n21779 = n21777 & n21778 ;
  assign n21782 = ~n13468 & n18727 ;
  assign n21783 = ~x110 & n21782 ;
  assign n21780 = ~n7172 & n11538 ;
  assign n21781 = n21780 ^ n16664 ^ 1'b0 ;
  assign n21784 = n21783 ^ n21781 ^ 1'b0 ;
  assign n21785 = n21784 ^ n13407 ^ n11966 ;
  assign n21786 = n21785 ^ n8594 ^ 1'b0 ;
  assign n21787 = n9606 ^ n8978 ^ 1'b0 ;
  assign n21788 = n20582 & n21787 ;
  assign n21789 = n21788 ^ n13657 ^ n12140 ;
  assign n21790 = n10222 & n15391 ;
  assign n21791 = n21790 ^ n19857 ^ 1'b0 ;
  assign n21792 = n13739 ^ n8803 ^ n3034 ;
  assign n21793 = n2399 & ~n3997 ;
  assign n21794 = n21793 ^ n13292 ^ 1'b0 ;
  assign n21795 = n5314 ^ n4509 ^ 1'b0 ;
  assign n21796 = n14473 ^ n9117 ^ n345 ;
  assign n21797 = n6098 & ~n21796 ;
  assign n21798 = n512 | n6186 ;
  assign n21799 = n21798 ^ n3694 ^ 1'b0 ;
  assign n21800 = n7726 & n21799 ;
  assign n21801 = ( n582 & n5885 ) | ( n582 & ~n15696 ) | ( n5885 & ~n15696 ) ;
  assign n21802 = n718 | n21801 ;
  assign n21803 = n4286 & ~n21802 ;
  assign n21804 = n7536 & ~n17313 ;
  assign n21805 = n21804 ^ n9001 ^ 1'b0 ;
  assign n21806 = n706 | n12537 ;
  assign n21807 = n17862 ^ n10955 ^ 1'b0 ;
  assign n21808 = ~n5354 & n9059 ;
  assign n21809 = n21808 ^ n21777 ^ 1'b0 ;
  assign n21810 = ~n673 & n12818 ;
  assign n21811 = n3854 & ~n19754 ;
  assign n21812 = n21810 & n21811 ;
  assign n21813 = ( n3958 & ~n16642 ) | ( n3958 & n19583 ) | ( ~n16642 & n19583 ) ;
  assign n21814 = ~n9352 & n9379 ;
  assign n21815 = n21814 ^ n3009 ^ 1'b0 ;
  assign n21816 = ( n12853 & n13527 ) | ( n12853 & n21815 ) | ( n13527 & n21815 ) ;
  assign n21817 = n21816 ^ x37 ^ 1'b0 ;
  assign n21818 = ( n6638 & ~n6808 ) | ( n6638 & n21817 ) | ( ~n6808 & n21817 ) ;
  assign n21819 = n1616 | n12609 ;
  assign n21820 = n21819 ^ n13930 ^ 1'b0 ;
  assign n21821 = n11718 ^ n1266 ^ 1'b0 ;
  assign n21822 = n3903 | n21821 ;
  assign n21823 = n2830 & ~n19559 ;
  assign n21824 = n21822 & n21823 ;
  assign n21825 = n2264 & n15747 ;
  assign n21826 = n21825 ^ n2516 ^ 1'b0 ;
  assign n21827 = ~n7293 & n17716 ;
  assign n21828 = n9178 & n13571 ;
  assign n21829 = n19517 ^ n989 ^ 1'b0 ;
  assign n21830 = n2266 | n13316 ;
  assign n21831 = n12020 & ~n21830 ;
  assign n21832 = x191 & n21831 ;
  assign n21833 = ~n5233 & n21832 ;
  assign n21834 = ~n8095 & n21833 ;
  assign n21835 = n16891 & ~n21834 ;
  assign n21836 = ~n13780 & n20624 ;
  assign n21837 = n21836 ^ n10316 ^ 1'b0 ;
  assign n21838 = n3055 & n3467 ;
  assign n21839 = n6975 & n15056 ;
  assign n21840 = ~n6344 & n21839 ;
  assign n21841 = ( n14115 & n21838 ) | ( n14115 & ~n21840 ) | ( n21838 & ~n21840 ) ;
  assign n21842 = n11509 ^ n9374 ^ 1'b0 ;
  assign n21843 = n19939 ^ n7915 ^ 1'b0 ;
  assign n21844 = n6093 & n21843 ;
  assign n21845 = n6081 ^ n1033 ^ 1'b0 ;
  assign n21846 = n14122 | n21845 ;
  assign n21847 = ( ~n1806 & n6158 ) | ( ~n1806 & n21846 ) | ( n6158 & n21846 ) ;
  assign n21848 = n11348 ^ n756 ^ 1'b0 ;
  assign n21852 = n4395 & n8839 ;
  assign n21853 = n21852 ^ n11328 ^ 1'b0 ;
  assign n21849 = ~n5295 & n6084 ;
  assign n21850 = n3374 & n21849 ;
  assign n21851 = n21850 ^ n11672 ^ n2910 ;
  assign n21854 = n21853 ^ n21851 ^ 1'b0 ;
  assign n21855 = x159 & n21854 ;
  assign n21856 = n10685 & n17905 ;
  assign n21857 = n16967 | n17792 ;
  assign n21858 = n20268 | n21857 ;
  assign n21859 = n15295 ^ n10521 ^ 1'b0 ;
  assign n21860 = n21859 ^ n10621 ^ n4762 ;
  assign n21861 = n1472 | n2404 ;
  assign n21862 = n4376 | n21861 ;
  assign n21863 = n8649 | n21862 ;
  assign n21864 = n3202 | n16825 ;
  assign n21865 = n657 | n21864 ;
  assign n21866 = n19177 & n21865 ;
  assign n21867 = n17761 & n21866 ;
  assign n21868 = n3340 & n8829 ;
  assign n21869 = ( n2651 & n14023 ) | ( n2651 & n21868 ) | ( n14023 & n21868 ) ;
  assign n21870 = n21869 ^ n20667 ^ 1'b0 ;
  assign n21871 = n8620 ^ n6692 ^ 1'b0 ;
  assign n21872 = n18993 & ~n21871 ;
  assign n21873 = n11013 & ~n16738 ;
  assign n21874 = n11461 & ~n21873 ;
  assign n21875 = n2036 & ~n3380 ;
  assign n21876 = n8226 | n21875 ;
  assign n21877 = n8060 | n21876 ;
  assign n21878 = ( ~n15158 & n21874 ) | ( ~n15158 & n21877 ) | ( n21874 & n21877 ) ;
  assign n21879 = ~n867 & n1643 ;
  assign n21880 = n12717 & ~n21879 ;
  assign n21881 = ~n17377 & n21880 ;
  assign n21882 = n21878 & n21881 ;
  assign n21883 = n6359 & ~n12642 ;
  assign n21884 = ~n16766 & n21883 ;
  assign n21885 = n17560 ^ n961 ^ 1'b0 ;
  assign n21886 = n17631 | n21885 ;
  assign n21887 = ~n1663 & n10385 ;
  assign n21888 = n21887 ^ n10612 ^ 1'b0 ;
  assign n21889 = n8780 & n17598 ;
  assign n21890 = n12241 & n21889 ;
  assign n21891 = n11802 ^ n2684 ^ 1'b0 ;
  assign n21892 = n549 | n21891 ;
  assign n21893 = n19566 ^ n14093 ^ n5331 ;
  assign n21894 = n3641 | n15330 ;
  assign n21895 = n17772 | n21894 ;
  assign n21896 = n5945 & n21895 ;
  assign n21897 = ~n8370 & n18846 ;
  assign n21899 = n12009 ^ n10122 ^ 1'b0 ;
  assign n21898 = n9854 ^ n7768 ^ n732 ;
  assign n21900 = n21899 ^ n21898 ^ n17733 ;
  assign n21901 = n2732 | n4298 ;
  assign n21902 = n21901 ^ n1488 ^ 1'b0 ;
  assign n21903 = n10595 & n21902 ;
  assign n21906 = n12485 ^ n1897 ^ 1'b0 ;
  assign n21907 = x237 & n21906 ;
  assign n21904 = n20603 ^ n4902 ^ 1'b0 ;
  assign n21905 = n6736 | n21904 ;
  assign n21908 = n21907 ^ n21905 ^ n7844 ;
  assign n21909 = n2500 ^ n2057 ^ 1'b0 ;
  assign n21910 = n271 & ~n21909 ;
  assign n21911 = ( x11 & n1952 ) | ( x11 & ~n21910 ) | ( n1952 & ~n21910 ) ;
  assign n21912 = ( ~n4242 & n4423 ) | ( ~n4242 & n21911 ) | ( n4423 & n21911 ) ;
  assign n21913 = n14339 & ~n21912 ;
  assign n21914 = n9862 ^ n4595 ^ n2965 ;
  assign n21915 = ( ~n4772 & n6200 ) | ( ~n4772 & n6526 ) | ( n6200 & n6526 ) ;
  assign n21916 = ( n9379 & ~n17889 ) | ( n9379 & n21915 ) | ( ~n17889 & n21915 ) ;
  assign n21917 = n21916 ^ n3483 ^ n1687 ;
  assign n21918 = n13466 | n16194 ;
  assign n21919 = n5843 | n21918 ;
  assign n21920 = n20853 ^ n20056 ^ 1'b0 ;
  assign n21921 = n3750 & n15105 ;
  assign n21922 = n21921 ^ n6223 ^ 1'b0 ;
  assign n21923 = n21922 ^ n11737 ^ 1'b0 ;
  assign n21924 = n5765 ^ n4333 ^ 1'b0 ;
  assign n21925 = n15952 ^ n10011 ^ n3638 ;
  assign n21927 = n12001 ^ n1101 ^ 1'b0 ;
  assign n21928 = n985 | n21927 ;
  assign n21926 = n6683 & ~n10529 ;
  assign n21929 = n21928 ^ n21926 ^ 1'b0 ;
  assign n21934 = n11667 ^ n6975 ^ 1'b0 ;
  assign n21930 = ( n3119 & n5588 ) | ( n3119 & ~n15938 ) | ( n5588 & ~n15938 ) ;
  assign n21931 = n21930 ^ n2106 ^ 1'b0 ;
  assign n21932 = n21931 ^ n13192 ^ 1'b0 ;
  assign n21933 = ~n4766 & n21932 ;
  assign n21935 = n21934 ^ n21933 ^ 1'b0 ;
  assign n21936 = n7571 ^ n4674 ^ 1'b0 ;
  assign n21937 = n14258 | n21936 ;
  assign n21938 = n13556 ^ n2957 ^ 1'b0 ;
  assign n21939 = n15829 ^ n5230 ^ 1'b0 ;
  assign n21940 = n10214 ^ n4094 ^ 1'b0 ;
  assign n21941 = n21940 ^ n1192 ^ 1'b0 ;
  assign n21942 = n3322 & n8404 ;
  assign n21943 = ~n1483 & n21942 ;
  assign n21944 = n9752 ^ n9619 ^ 1'b0 ;
  assign n21945 = n9259 & n21944 ;
  assign n21946 = n21945 ^ n3797 ^ 1'b0 ;
  assign n21947 = n12767 ^ n1528 ^ 1'b0 ;
  assign n21948 = n21947 ^ n13384 ^ 1'b0 ;
  assign n21949 = ~n1223 & n9108 ;
  assign n21950 = n4497 ^ x234 ^ 1'b0 ;
  assign n21951 = ( n3492 & ~n5816 ) | ( n3492 & n9351 ) | ( ~n5816 & n9351 ) ;
  assign n21952 = ~n5656 & n21951 ;
  assign n21953 = ( n7145 & n21950 ) | ( n7145 & ~n21952 ) | ( n21950 & ~n21952 ) ;
  assign n21954 = ~n13623 & n21953 ;
  assign n21955 = ~n21949 & n21954 ;
  assign n21956 = n1453 | n11799 ;
  assign n21957 = n21956 ^ n5121 ^ 1'b0 ;
  assign n21958 = n20536 ^ n13742 ^ 1'b0 ;
  assign n21959 = ~n685 & n21958 ;
  assign n21964 = n21021 ^ n320 ^ 1'b0 ;
  assign n21965 = n21964 ^ n9201 ^ x247 ;
  assign n21966 = n19339 & n21965 ;
  assign n21967 = ~n19339 & n21966 ;
  assign n21960 = ~n639 & n4718 ;
  assign n21961 = n639 & n21960 ;
  assign n21962 = n3922 | n21961 ;
  assign n21963 = n3922 & ~n21962 ;
  assign n21968 = n21967 ^ n21963 ^ n18915 ;
  assign n21969 = n16373 & n17730 ;
  assign n21970 = ~n16373 & n21969 ;
  assign n21971 = n21968 & ~n21970 ;
  assign n21972 = ~n21959 & n21971 ;
  assign n21973 = n14294 ^ n6720 ^ 1'b0 ;
  assign n21974 = n5923 & n21973 ;
  assign n21975 = n14339 ^ n10378 ^ 1'b0 ;
  assign n21976 = ~n5216 & n11975 ;
  assign n21977 = n21976 ^ n18545 ^ n9960 ;
  assign n21978 = n21977 ^ n11607 ^ 1'b0 ;
  assign n21979 = x84 & ~n21978 ;
  assign n21980 = n21979 ^ n1499 ^ 1'b0 ;
  assign n21981 = n12923 ^ n11531 ^ n4328 ;
  assign n21982 = n21981 ^ n9432 ^ 1'b0 ;
  assign n21983 = n19116 & ~n21982 ;
  assign n21984 = ( ~n4595 & n7439 ) | ( ~n4595 & n19748 ) | ( n7439 & n19748 ) ;
  assign n21985 = ~n9605 & n17442 ;
  assign n21986 = n20584 ^ n16691 ^ 1'b0 ;
  assign n21987 = n3734 ^ n3237 ^ 1'b0 ;
  assign n21988 = ~n5263 & n21987 ;
  assign n21989 = n13384 ^ n10422 ^ 1'b0 ;
  assign n21990 = n21988 & n21989 ;
  assign n21991 = n14624 | n21990 ;
  assign n21992 = n21009 & n21991 ;
  assign n21993 = ~n369 & n6196 ;
  assign n21994 = n9763 & n16968 ;
  assign n21995 = ~n21993 & n21994 ;
  assign n21996 = ( n14150 & n15705 ) | ( n14150 & ~n21995 ) | ( n15705 & ~n21995 ) ;
  assign n21997 = ( n6310 & ~n10293 ) | ( n6310 & n21996 ) | ( ~n10293 & n21996 ) ;
  assign n21998 = n15689 | n21458 ;
  assign n21999 = n21998 ^ n13992 ^ 1'b0 ;
  assign n22000 = n4797 & n21999 ;
  assign n22001 = ~n8509 & n22000 ;
  assign n22002 = ~n2592 & n11821 ;
  assign n22003 = n2428 & ~n16058 ;
  assign n22004 = n22002 & n22003 ;
  assign n22005 = n4150 | n6464 ;
  assign n22006 = n3835 | n22005 ;
  assign n22008 = n12864 ^ n4775 ^ 1'b0 ;
  assign n22009 = n13887 & n22008 ;
  assign n22007 = ~n4562 & n14207 ;
  assign n22010 = n22009 ^ n22007 ^ 1'b0 ;
  assign n22011 = n7573 ^ n7102 ^ 1'b0 ;
  assign n22012 = ~n14566 & n18871 ;
  assign n22013 = n13917 ^ n8602 ^ 1'b0 ;
  assign n22014 = n1407 & n22013 ;
  assign n22015 = n16021 ^ x212 ^ 1'b0 ;
  assign n22016 = n4716 ^ n4620 ^ 1'b0 ;
  assign n22017 = n22016 ^ n21928 ^ 1'b0 ;
  assign n22018 = n8041 | n22017 ;
  assign n22019 = n22018 ^ n9986 ^ 1'b0 ;
  assign n22020 = n2217 | n17485 ;
  assign n22021 = ( n9077 & n17495 ) | ( n9077 & n22020 ) | ( n17495 & n22020 ) ;
  assign n22022 = ~n918 & n3856 ;
  assign n22023 = n3927 | n22022 ;
  assign n22025 = n10753 ^ n729 ^ 1'b0 ;
  assign n22026 = n11066 | n22025 ;
  assign n22027 = n22026 ^ n14052 ^ 1'b0 ;
  assign n22024 = n1476 & ~n12745 ;
  assign n22028 = n22027 ^ n22024 ^ 1'b0 ;
  assign n22029 = n14762 ^ n10036 ^ 1'b0 ;
  assign n22030 = n16631 & n22029 ;
  assign n22031 = n3586 & ~n6329 ;
  assign n22032 = n7081 | n9432 ;
  assign n22033 = n22032 ^ n5140 ^ 1'b0 ;
  assign n22034 = n6910 & ~n22033 ;
  assign n22035 = ~n10432 & n22034 ;
  assign n22036 = n22031 & ~n22035 ;
  assign n22037 = n22036 ^ n1477 ^ 1'b0 ;
  assign n22038 = n22037 ^ n10518 ^ 1'b0 ;
  assign n22039 = ~n740 & n22038 ;
  assign n22040 = n7830 ^ n7748 ^ 1'b0 ;
  assign n22041 = n22040 ^ n18551 ^ n3320 ;
  assign n22042 = ( n5124 & n5525 ) | ( n5124 & ~n6384 ) | ( n5525 & ~n6384 ) ;
  assign n22043 = n22042 ^ n3866 ^ 1'b0 ;
  assign n22044 = n11657 ^ n984 ^ 1'b0 ;
  assign n22045 = ~n2916 & n3394 ;
  assign n22046 = n22045 ^ n12385 ^ 1'b0 ;
  assign n22047 = ( ~n4631 & n5084 ) | ( ~n4631 & n11316 ) | ( n5084 & n11316 ) ;
  assign n22048 = ( x116 & ~n3880 ) | ( x116 & n22047 ) | ( ~n3880 & n22047 ) ;
  assign n22049 = n22048 ^ n10709 ^ 1'b0 ;
  assign n22050 = n10825 | n22049 ;
  assign n22051 = ~n4124 & n13081 ;
  assign n22052 = n22051 ^ n9767 ^ 1'b0 ;
  assign n22053 = n1767 & n22052 ;
  assign n22054 = n5020 & ~n18346 ;
  assign n22055 = n22054 ^ n6531 ^ 1'b0 ;
  assign n22056 = n13277 | n22055 ;
  assign n22057 = n10066 | n22056 ;
  assign n22062 = n3161 ^ n2896 ^ n2261 ;
  assign n22061 = n2957 & ~n9998 ;
  assign n22063 = n22062 ^ n22061 ^ 1'b0 ;
  assign n22064 = n22063 ^ n17358 ^ 1'b0 ;
  assign n22058 = x51 & n14856 ;
  assign n22059 = n2914 & n22058 ;
  assign n22060 = n2488 & ~n22059 ;
  assign n22065 = n22064 ^ n22060 ^ 1'b0 ;
  assign n22074 = n5912 & n7709 ;
  assign n22066 = x148 & ~n4824 ;
  assign n22067 = n3160 | n4655 ;
  assign n22068 = ~n1823 & n22067 ;
  assign n22069 = n5757 ^ n2224 ^ 1'b0 ;
  assign n22070 = ~n10501 & n22069 ;
  assign n22071 = n1548 & n22070 ;
  assign n22072 = ( n22066 & n22068 ) | ( n22066 & n22071 ) | ( n22068 & n22071 ) ;
  assign n22073 = n22072 ^ n3687 ^ 1'b0 ;
  assign n22075 = n22074 ^ n22073 ^ n20288 ;
  assign n22076 = n1694 & n10043 ;
  assign n22077 = n9263 ^ n327 ^ 1'b0 ;
  assign n22078 = n8236 & n22077 ;
  assign n22079 = n7273 & ~n22078 ;
  assign n22080 = ( ~n1110 & n6240 ) | ( ~n1110 & n8675 ) | ( n6240 & n8675 ) ;
  assign n22081 = ~n22079 & n22080 ;
  assign n22082 = n10694 & ~n22081 ;
  assign n22083 = n22082 ^ n19180 ^ 1'b0 ;
  assign n22084 = ~n376 & n1106 ;
  assign n22085 = n7984 ^ n2628 ^ 1'b0 ;
  assign n22086 = n22084 | n22085 ;
  assign n22087 = ~n535 & n18053 ;
  assign n22088 = n22087 ^ n6271 ^ 1'b0 ;
  assign n22089 = n22088 ^ n2164 ^ 1'b0 ;
  assign n22090 = ( ~x75 & n2078 ) | ( ~x75 & n6369 ) | ( n2078 & n6369 ) ;
  assign n22091 = n2077 | n6400 ;
  assign n22092 = n22091 ^ n1024 ^ 1'b0 ;
  assign n22093 = n2687 & n18119 ;
  assign n22094 = ~n17544 & n22093 ;
  assign n22095 = n14852 & n20723 ;
  assign n22096 = n22095 ^ n9554 ^ 1'b0 ;
  assign n22097 = n22096 ^ n5324 ^ 1'b0 ;
  assign n22098 = ~n20438 & n22097 ;
  assign n22099 = n22094 & n22098 ;
  assign n22100 = n22092 | n22099 ;
  assign n22101 = n22090 & ~n22100 ;
  assign n22102 = ( ~n1903 & n7960 ) | ( ~n1903 & n16129 ) | ( n7960 & n16129 ) ;
  assign n22103 = n13063 | n22102 ;
  assign n22104 = n22103 ^ n8090 ^ 1'b0 ;
  assign n22105 = n4994 ^ n875 ^ 1'b0 ;
  assign n22106 = n11322 | n20976 ;
  assign n22107 = n22106 ^ n13231 ^ 1'b0 ;
  assign n22108 = n1030 & ~n9979 ;
  assign n22109 = n22108 ^ n13843 ^ 1'b0 ;
  assign n22110 = n22109 ^ n12281 ^ n5250 ;
  assign n22111 = n18850 & ~n22110 ;
  assign n22112 = n3411 & n10793 ;
  assign n22113 = n13367 & n22112 ;
  assign n22114 = n15141 ^ n4317 ^ n3551 ;
  assign n22115 = n22114 ^ n1876 ^ 1'b0 ;
  assign n22116 = n10045 | n22115 ;
  assign n22117 = n9912 & n14068 ;
  assign n22118 = ~n9514 & n10946 ;
  assign n22119 = n6019 & n22118 ;
  assign n22120 = ~n19911 & n20537 ;
  assign n22121 = n12526 ^ n2513 ^ 1'b0 ;
  assign n22122 = n2707 & ~n22121 ;
  assign n22123 = n2048 & ~n10296 ;
  assign n22124 = n17916 & n22123 ;
  assign n22125 = n22122 & n22124 ;
  assign n22126 = n8932 | n15294 ;
  assign n22127 = n8708 ^ n1777 ^ 1'b0 ;
  assign n22128 = n22126 & n22127 ;
  assign n22129 = n22128 ^ n10691 ^ 1'b0 ;
  assign n22130 = n10850 & n18598 ;
  assign n22131 = ( ~n301 & n3150 ) | ( ~n301 & n8527 ) | ( n3150 & n8527 ) ;
  assign n22133 = n9188 ^ n6088 ^ n5736 ;
  assign n22132 = n4173 | n13802 ;
  assign n22134 = n22133 ^ n22132 ^ 1'b0 ;
  assign n22135 = n319 | n10215 ;
  assign n22136 = n22134 & ~n22135 ;
  assign n22137 = n21334 ^ n1509 ^ 1'b0 ;
  assign n22139 = n7231 & n11537 ;
  assign n22138 = n4731 & ~n4967 ;
  assign n22140 = n22139 ^ n22138 ^ n8623 ;
  assign n22141 = ( n6429 & n17645 ) | ( n6429 & n22140 ) | ( n17645 & n22140 ) ;
  assign n22142 = n8126 ^ n6596 ^ n3685 ;
  assign n22143 = ( n2721 & n6493 ) | ( n2721 & n22142 ) | ( n6493 & n22142 ) ;
  assign n22144 = n22143 ^ n15604 ^ 1'b0 ;
  assign n22145 = n8548 & n14178 ;
  assign n22146 = n9394 & ~n18200 ;
  assign n22147 = x14 & ~n6119 ;
  assign n22148 = ~x30 & n22147 ;
  assign n22149 = ~x153 & n10653 ;
  assign n22150 = n22149 ^ n5155 ^ 1'b0 ;
  assign n22151 = n14366 ^ n2743 ^ 1'b0 ;
  assign n22152 = n14059 & n22151 ;
  assign n22153 = ~n19968 & n22152 ;
  assign n22154 = ~n22150 & n22153 ;
  assign n22155 = ~n10882 & n13806 ;
  assign n22156 = n13520 ^ n2258 ^ 1'b0 ;
  assign n22157 = n20486 ^ n7809 ^ 1'b0 ;
  assign n22158 = n17638 | n22157 ;
  assign n22159 = ~n729 & n9832 ;
  assign n22160 = n22159 ^ n489 ^ 1'b0 ;
  assign n22161 = n22160 ^ n13584 ^ 1'b0 ;
  assign n22162 = n5780 ^ n1804 ^ 1'b0 ;
  assign n22163 = n12654 ^ n12580 ^ n11274 ;
  assign n22164 = n12061 ^ n4300 ^ n805 ;
  assign n22165 = ~n22163 & n22164 ;
  assign n22166 = ( n13320 & ~n17102 ) | ( n13320 & n18020 ) | ( ~n17102 & n18020 ) ;
  assign n22171 = ~n7962 & n10580 ;
  assign n22172 = n22171 ^ n12158 ^ 1'b0 ;
  assign n22167 = n5927 & ~n11864 ;
  assign n22168 = n14169 & n22167 ;
  assign n22169 = ~n22167 & n22168 ;
  assign n22170 = n22169 ^ n288 ^ 1'b0 ;
  assign n22173 = n22172 ^ n22170 ^ n11718 ;
  assign n22174 = n22173 ^ n10532 ^ 1'b0 ;
  assign n22175 = n7267 ^ n3050 ^ n1407 ;
  assign n22176 = n19121 & n22175 ;
  assign n22177 = n4580 & n22176 ;
  assign n22178 = n4042 | n10125 ;
  assign n22179 = n22177 & ~n22178 ;
  assign n22180 = n1961 & ~n6057 ;
  assign n22181 = x91 & ~n690 ;
  assign n22182 = n22181 ^ n692 ^ 1'b0 ;
  assign n22183 = n22067 ^ n7404 ^ 1'b0 ;
  assign n22184 = n10983 & n22183 ;
  assign n22185 = n4423 & n7017 ;
  assign n22186 = n22185 ^ n12562 ^ 1'b0 ;
  assign n22188 = n3821 ^ n948 ^ 1'b0 ;
  assign n22187 = ~n283 & n8789 ;
  assign n22189 = n22188 ^ n22187 ^ 1'b0 ;
  assign n22190 = n8639 & n22189 ;
  assign n22191 = ~n22186 & n22190 ;
  assign n22192 = n20932 & ~n22191 ;
  assign n22193 = ~n22184 & n22192 ;
  assign n22194 = ( n1489 & n16477 ) | ( n1489 & n18336 ) | ( n16477 & n18336 ) ;
  assign n22195 = ~n7264 & n20019 ;
  assign n22196 = n22195 ^ n6021 ^ 1'b0 ;
  assign n22197 = n22194 & n22196 ;
  assign n22198 = n5985 & n12495 ;
  assign n22199 = ~n18403 & n22198 ;
  assign n22200 = n10736 & ~n12694 ;
  assign n22201 = n22200 ^ n4775 ^ 1'b0 ;
  assign n22202 = n13740 & ~n22201 ;
  assign n22206 = n6018 ^ n5034 ^ x39 ;
  assign n22203 = n1913 & ~n4306 ;
  assign n22204 = ~n817 & n22203 ;
  assign n22205 = n12413 & n22204 ;
  assign n22207 = n22206 ^ n22205 ^ n18603 ;
  assign n22208 = ~n12741 & n18013 ;
  assign n22209 = n11351 ^ n2054 ^ 1'b0 ;
  assign n22210 = n1218 & ~n22209 ;
  assign n22211 = n12131 & n22210 ;
  assign n22212 = ~n13391 & n22211 ;
  assign n22213 = n1524 | n7040 ;
  assign n22214 = n1733 | n16094 ;
  assign n22215 = ~n4065 & n22214 ;
  assign n22216 = n9870 & ~n22215 ;
  assign n22217 = n22216 ^ n342 ^ 1'b0 ;
  assign n22218 = ~n349 & n17585 ;
  assign n22220 = n4657 & ~n11306 ;
  assign n22219 = n11446 ^ n11328 ^ n9684 ;
  assign n22221 = n22220 ^ n22219 ^ 1'b0 ;
  assign n22222 = n6091 ^ n1021 ^ 1'b0 ;
  assign n22223 = n1524 & n22222 ;
  assign n22224 = n11716 ^ n10438 ^ 1'b0 ;
  assign n22225 = n2428 & ~n22224 ;
  assign n22226 = n16207 ^ n11042 ^ 1'b0 ;
  assign n22227 = ( n7429 & n13992 ) | ( n7429 & ~n18783 ) | ( n13992 & ~n18783 ) ;
  assign n22228 = n22227 ^ n9172 ^ 1'b0 ;
  assign n22229 = n749 | n15670 ;
  assign n22230 = n739 & ~n19193 ;
  assign n22231 = n22230 ^ n19137 ^ 1'b0 ;
  assign n22232 = n8826 & n21158 ;
  assign n22233 = n5597 ^ n2306 ^ 1'b0 ;
  assign n22234 = n7398 & n22233 ;
  assign n22235 = n22234 ^ n6345 ^ n6299 ;
  assign n22236 = n11886 & n14635 ;
  assign n22237 = ~n12189 & n22236 ;
  assign n22238 = n17704 ^ n12376 ^ n9329 ;
  assign n22239 = n17982 | n22238 ;
  assign n22240 = n22239 ^ n9276 ^ 1'b0 ;
  assign n22241 = x131 & ~n11228 ;
  assign n22242 = n3662 & n22241 ;
  assign n22243 = n22242 ^ n7822 ^ 1'b0 ;
  assign n22249 = n459 & ~n10221 ;
  assign n22250 = n10221 & n22249 ;
  assign n22251 = n672 & ~n22250 ;
  assign n22252 = ~n672 & n22251 ;
  assign n22253 = n1989 & n22252 ;
  assign n22244 = ~n322 & n6700 ;
  assign n22245 = n22244 ^ n5387 ^ 1'b0 ;
  assign n22246 = n12536 ^ n1830 ^ 1'b0 ;
  assign n22247 = n1086 & ~n22246 ;
  assign n22248 = n22245 & n22247 ;
  assign n22254 = n22253 ^ n22248 ^ 1'b0 ;
  assign n22255 = n15747 & n22254 ;
  assign n22256 = n13945 ^ n9668 ^ n2542 ;
  assign n22257 = n1239 & n22256 ;
  assign n22258 = n21683 & n22257 ;
  assign n22259 = n1203 & ~n4460 ;
  assign n22260 = n6599 | n10532 ;
  assign n22261 = n22260 ^ n9317 ^ 1'b0 ;
  assign n22262 = n22261 ^ n21910 ^ n6402 ;
  assign n22263 = n2641 | n14740 ;
  assign n22264 = n20692 ^ n2670 ^ 1'b0 ;
  assign n22265 = n10187 | n22264 ;
  assign n22266 = ~n7004 & n9208 ;
  assign n22269 = n1866 ^ n959 ^ 1'b0 ;
  assign n22267 = ~n7788 & n14881 ;
  assign n22268 = n22267 ^ n6674 ^ 1'b0 ;
  assign n22270 = n22269 ^ n22268 ^ n2146 ;
  assign n22271 = n19866 ^ n4087 ^ 1'b0 ;
  assign n22272 = n10897 | n12947 ;
  assign n22273 = n12207 ^ n5920 ^ 1'b0 ;
  assign n22274 = ~n6934 & n22273 ;
  assign n22275 = ~n15671 & n22274 ;
  assign n22276 = n9944 & ~n10268 ;
  assign n22277 = ~n18129 & n22276 ;
  assign n22278 = n22277 ^ n5893 ^ 1'b0 ;
  assign n22279 = n6214 | n12823 ;
  assign n22280 = n6234 & ~n22279 ;
  assign n22281 = n1993 & n22280 ;
  assign n22282 = n12199 | n22281 ;
  assign n22283 = n22282 ^ n2924 ^ 1'b0 ;
  assign n22284 = n5029 | n6215 ;
  assign n22285 = n18169 | n22284 ;
  assign n22286 = n22159 ^ n10548 ^ n5826 ;
  assign n22287 = n22286 ^ n19121 ^ n4939 ;
  assign n22288 = n22285 & n22287 ;
  assign n22289 = ( ~n4479 & n17663 ) | ( ~n4479 & n18270 ) | ( n17663 & n18270 ) ;
  assign n22290 = ( n2282 & ~n4953 ) | ( n2282 & n8585 ) | ( ~n4953 & n8585 ) ;
  assign n22291 = x170 & n22290 ;
  assign n22292 = ~n22289 & n22291 ;
  assign n22293 = n18398 ^ n15657 ^ n13889 ;
  assign n22294 = n4891 & n14468 ;
  assign n22295 = ~n1622 & n22294 ;
  assign n22296 = n20382 | n22295 ;
  assign n22297 = n22296 ^ n9820 ^ 1'b0 ;
  assign n22298 = n4826 | n12950 ;
  assign n22299 = n8698 | n22298 ;
  assign n22300 = n13716 | n21290 ;
  assign n22301 = n3965 & ~n16747 ;
  assign n22302 = n11466 ^ n4354 ^ 1'b0 ;
  assign n22303 = n15119 & n22302 ;
  assign n22304 = n8200 ^ n4469 ^ n4458 ;
  assign n22307 = ~x170 & n8941 ;
  assign n22308 = n22307 ^ n1228 ^ 1'b0 ;
  assign n22309 = n18246 & n22308 ;
  assign n22305 = n19907 ^ n2477 ^ 1'b0 ;
  assign n22306 = n7308 & ~n22305 ;
  assign n22310 = n22309 ^ n22306 ^ n6874 ;
  assign n22311 = n13764 | n18276 ;
  assign n22312 = n6336 ^ n2460 ^ 1'b0 ;
  assign n22313 = ~n11642 & n22312 ;
  assign n22314 = n22313 ^ n6310 ^ 1'b0 ;
  assign n22315 = n22314 ^ n4831 ^ 1'b0 ;
  assign n22316 = n3388 | n7172 ;
  assign n22317 = n22316 ^ n5124 ^ x68 ;
  assign n22318 = n22317 ^ n5004 ^ 1'b0 ;
  assign n22319 = n1758 & n22318 ;
  assign n22320 = n7282 ^ n2696 ^ 1'b0 ;
  assign n22321 = n1153 | n5013 ;
  assign n22322 = n9154 & ~n22321 ;
  assign n22323 = n2763 & n21272 ;
  assign n22324 = n22323 ^ n11175 ^ 1'b0 ;
  assign n22325 = n13641 ^ n9671 ^ n8598 ;
  assign n22326 = n9490 ^ n3696 ^ 1'b0 ;
  assign n22327 = n3097 & n22326 ;
  assign n22328 = n22327 ^ n10361 ^ 1'b0 ;
  assign n22329 = n22325 | n22328 ;
  assign n22330 = n11694 & ~n22329 ;
  assign n22331 = n22330 ^ n5601 ^ 1'b0 ;
  assign n22332 = ~n7975 & n12494 ;
  assign n22333 = n8695 & n22332 ;
  assign n22334 = n22333 ^ n19659 ^ n19456 ;
  assign n22335 = ~n1655 & n11917 ;
  assign n22336 = n11999 | n22335 ;
  assign n22337 = n9471 & ~n11333 ;
  assign n22338 = n1489 & n22337 ;
  assign n22340 = n6572 | n14517 ;
  assign n22341 = n3380 & n12228 ;
  assign n22342 = n10091 & n22341 ;
  assign n22343 = n22340 & n22342 ;
  assign n22339 = x161 & ~n7409 ;
  assign n22344 = n22343 ^ n22339 ^ 1'b0 ;
  assign n22345 = n6723 & n18272 ;
  assign n22346 = n22345 ^ n17544 ^ 1'b0 ;
  assign n22347 = n5288 ^ n308 ^ 1'b0 ;
  assign n22348 = n13333 & n22347 ;
  assign n22349 = n22348 ^ n12672 ^ n8763 ;
  assign n22350 = ~n8908 & n11585 ;
  assign n22353 = x179 & ~n10751 ;
  assign n22354 = n5739 & n22353 ;
  assign n22351 = n3567 ^ n896 ^ 1'b0 ;
  assign n22352 = n10089 | n22351 ;
  assign n22355 = n22354 ^ n22352 ^ 1'b0 ;
  assign n22356 = n17369 ^ n1462 ^ 1'b0 ;
  assign n22357 = n8202 & n15966 ;
  assign n22358 = ~n6385 & n22357 ;
  assign n22359 = n5154 & ~n13360 ;
  assign n22360 = n22359 ^ n9676 ^ 1'b0 ;
  assign n22361 = n20482 & ~n22360 ;
  assign n22362 = n22361 ^ n2191 ^ 1'b0 ;
  assign n22363 = ( n8159 & n10252 ) | ( n8159 & ~n22362 ) | ( n10252 & ~n22362 ) ;
  assign n22364 = x223 | n366 ;
  assign n22365 = n19137 ^ n6923 ^ 1'b0 ;
  assign n22366 = n6412 & n22365 ;
  assign n22369 = n4471 & ~n13746 ;
  assign n22370 = n11123 & n22369 ;
  assign n22367 = n4684 | n16203 ;
  assign n22368 = n8275 & ~n22367 ;
  assign n22371 = n22370 ^ n22368 ^ 1'b0 ;
  assign n22372 = n22366 & ~n22371 ;
  assign n22373 = ( ~n4084 & n16129 ) | ( ~n4084 & n19891 ) | ( n16129 & n19891 ) ;
  assign n22374 = n7590 ^ n2033 ^ 1'b0 ;
  assign n22375 = n22374 ^ n14449 ^ 1'b0 ;
  assign n22376 = ( n6508 & ~n22373 ) | ( n6508 & n22375 ) | ( ~n22373 & n22375 ) ;
  assign n22378 = n18829 ^ n15936 ^ 1'b0 ;
  assign n22379 = n1900 | n22378 ;
  assign n22377 = n9352 | n15946 ;
  assign n22380 = n22379 ^ n22377 ^ 1'b0 ;
  assign n22381 = n2706 & n22380 ;
  assign n22382 = n2006 & ~n15992 ;
  assign n22383 = n22382 ^ n2332 ^ 1'b0 ;
  assign n22384 = ~n6704 & n12522 ;
  assign n22385 = n13159 & n22384 ;
  assign n22386 = ~n7569 & n19575 ;
  assign n22387 = n4312 | n8842 ;
  assign n22388 = ( n13391 & n15415 ) | ( n13391 & n22273 ) | ( n15415 & n22273 ) ;
  assign n22390 = n18725 ^ n4818 ^ 1'b0 ;
  assign n22391 = n22390 ^ n7928 ^ n5776 ;
  assign n22389 = n12640 & n12647 ;
  assign n22392 = n22391 ^ n22389 ^ 1'b0 ;
  assign n22393 = n15928 | n22392 ;
  assign n22397 = n6987 & n7217 ;
  assign n22398 = n14738 & n22397 ;
  assign n22394 = n7317 ^ n2746 ^ 1'b0 ;
  assign n22395 = n22394 ^ n7370 ^ 1'b0 ;
  assign n22396 = n3097 & n22395 ;
  assign n22399 = n22398 ^ n22396 ^ 1'b0 ;
  assign n22400 = n5912 ^ n2725 ^ 1'b0 ;
  assign n22401 = n9987 ^ n397 ^ 1'b0 ;
  assign n22402 = ( n1989 & n22400 ) | ( n1989 & n22401 ) | ( n22400 & n22401 ) ;
  assign n22403 = n289 & n17728 ;
  assign n22404 = ~n9569 & n22403 ;
  assign n22405 = n6929 & ~n10851 ;
  assign n22406 = n22405 ^ n12310 ^ 1'b0 ;
  assign n22407 = n16261 ^ n7856 ^ n7778 ;
  assign n22408 = n3025 | n3843 ;
  assign n22409 = n22408 ^ n12639 ^ 1'b0 ;
  assign n22410 = ~n7097 & n22409 ;
  assign n22411 = ~n4953 & n22410 ;
  assign n22412 = ~n22407 & n22411 ;
  assign n22413 = n22412 ^ n16723 ^ n10742 ;
  assign n22414 = ~n1003 & n18835 ;
  assign n22415 = ( n10336 & ~n22314 ) | ( n10336 & n22414 ) | ( ~n22314 & n22414 ) ;
  assign n22416 = ~n10176 & n22415 ;
  assign n22417 = n22416 ^ n19804 ^ 1'b0 ;
  assign n22418 = ~n5724 & n22417 ;
  assign n22419 = n2366 & n7554 ;
  assign n22420 = n1830 | n18338 ;
  assign n22421 = n22419 | n22420 ;
  assign n22422 = n11516 ^ n10396 ^ 1'b0 ;
  assign n22423 = n13552 ^ n4535 ^ n1776 ;
  assign n22424 = n9780 & n22423 ;
  assign n22425 = n9154 & n22424 ;
  assign n22426 = n1648 | n7847 ;
  assign n22427 = ~n11350 & n12201 ;
  assign n22428 = n21091 & n22427 ;
  assign n22429 = n5546 & ~n22070 ;
  assign n22430 = n22429 ^ n2983 ^ 1'b0 ;
  assign n22431 = n21516 & n22430 ;
  assign n22432 = ~n5778 & n21523 ;
  assign n22433 = ~n3402 & n22432 ;
  assign n22434 = ( n3737 & ~n6392 ) | ( n3737 & n9496 ) | ( ~n6392 & n9496 ) ;
  assign n22435 = n22434 ^ n3123 ^ 1'b0 ;
  assign n22436 = n22433 | n22435 ;
  assign n22438 = n1924 & n6764 ;
  assign n22437 = ~n3025 & n8577 ;
  assign n22439 = n22438 ^ n22437 ^ 1'b0 ;
  assign n22440 = n3681 & ~n22439 ;
  assign n22441 = n17051 & n22440 ;
  assign n22443 = n9540 ^ n555 ^ 1'b0 ;
  assign n22442 = n6409 ^ n2773 ^ 1'b0 ;
  assign n22444 = n22443 ^ n22442 ^ n14236 ;
  assign n22445 = n11115 ^ n1700 ^ 1'b0 ;
  assign n22446 = n22445 ^ n21539 ^ n6874 ;
  assign n22447 = n9200 & n11605 ;
  assign n22448 = n17089 ^ n15985 ^ 1'b0 ;
  assign n22449 = n22447 | n22448 ;
  assign n22450 = n19845 ^ n3880 ^ n1284 ;
  assign n22451 = n17758 ^ n7139 ^ 1'b0 ;
  assign n22452 = n6368 & ~n22451 ;
  assign n22453 = n21117 | n22452 ;
  assign n22454 = ( ~n5389 & n16845 ) | ( ~n5389 & n22453 ) | ( n16845 & n22453 ) ;
  assign n22455 = n6847 | n10979 ;
  assign n22456 = n6188 & n15165 ;
  assign n22457 = n22455 & n22456 ;
  assign n22458 = n7001 ^ n4258 ^ 1'b0 ;
  assign n22459 = n6114 & ~n22458 ;
  assign n22460 = ~n2406 & n3369 ;
  assign n22461 = n22460 ^ n14965 ^ 1'b0 ;
  assign n22462 = n11663 & ~n22461 ;
  assign n22463 = n6035 & n22462 ;
  assign n22464 = n18323 ^ n1038 ^ 1'b0 ;
  assign n22465 = ~n785 & n22464 ;
  assign n22466 = n13407 & n21023 ;
  assign n22467 = n22466 ^ n5003 ^ 1'b0 ;
  assign n22468 = n1382 ^ n393 ^ 1'b0 ;
  assign n22469 = n15901 ^ n15198 ^ n1127 ;
  assign n22470 = ~n22468 & n22469 ;
  assign n22471 = ~n6338 & n11133 ;
  assign n22472 = n4910 | n9865 ;
  assign n22473 = n22472 ^ n10796 ^ 1'b0 ;
  assign n22474 = ~n1797 & n22473 ;
  assign n22475 = n2347 & n22474 ;
  assign n22476 = ( ~n755 & n10709 ) | ( ~n755 & n22475 ) | ( n10709 & n22475 ) ;
  assign n22477 = n1780 & n21716 ;
  assign n22478 = ~n15509 & n22477 ;
  assign n22479 = n22478 ^ n20602 ^ n10227 ;
  assign n22480 = n21446 ^ n14776 ^ 1'b0 ;
  assign n22481 = n14629 & ~n22480 ;
  assign n22482 = n21186 ^ n19308 ^ n4019 ;
  assign n22483 = ( n5013 & n5243 ) | ( n5013 & n11772 ) | ( n5243 & n11772 ) ;
  assign n22484 = n6138 ^ n2475 ^ 1'b0 ;
  assign n22485 = n15785 ^ n12548 ^ 1'b0 ;
  assign n22486 = n20359 & ~n22485 ;
  assign n22487 = ( n4354 & n14123 ) | ( n4354 & n20983 ) | ( n14123 & n20983 ) ;
  assign n22488 = n22486 & ~n22487 ;
  assign n22489 = n22488 ^ n3023 ^ 1'b0 ;
  assign n22490 = n1401 | n2795 ;
  assign n22491 = n636 & n22490 ;
  assign n22492 = ~n18655 & n22491 ;
  assign n22493 = n22492 ^ n10279 ^ 1'b0 ;
  assign n22494 = ( ~n3694 & n20041 ) | ( ~n3694 & n21270 ) | ( n20041 & n21270 ) ;
  assign n22495 = ~n7391 & n7675 ;
  assign n22496 = n22495 ^ n8893 ^ 1'b0 ;
  assign n22497 = ( ~n1021 & n7953 ) | ( ~n1021 & n18998 ) | ( n7953 & n18998 ) ;
  assign n22498 = n22497 ^ n20732 ^ 1'b0 ;
  assign n22499 = n16169 & n22498 ;
  assign n22500 = ~n10532 & n13727 ;
  assign n22501 = ~n14316 & n22500 ;
  assign n22506 = n19716 ^ n9714 ^ 1'b0 ;
  assign n22503 = n5121 & ~n11833 ;
  assign n22502 = ~n3481 & n5414 ;
  assign n22504 = n22503 ^ n22502 ^ 1'b0 ;
  assign n22505 = n11413 | n22504 ;
  assign n22507 = n22506 ^ n22505 ^ 1'b0 ;
  assign n22508 = ~n22501 & n22507 ;
  assign n22509 = n22508 ^ n15517 ^ 1'b0 ;
  assign n22510 = n17942 ^ n14603 ^ 1'b0 ;
  assign n22511 = n22510 ^ n16659 ^ n8276 ;
  assign n22512 = n4817 | n7421 ;
  assign n22513 = ~n11129 & n11333 ;
  assign n22514 = n22513 ^ n18335 ^ n5090 ;
  assign n22515 = ( n948 & n17809 ) | ( n948 & ~n22514 ) | ( n17809 & ~n22514 ) ;
  assign n22516 = ( n4970 & n11114 ) | ( n4970 & n12836 ) | ( n11114 & n12836 ) ;
  assign n22517 = n22516 ^ n6141 ^ 1'b0 ;
  assign n22518 = ( n5946 & ~n6838 ) | ( n5946 & n22517 ) | ( ~n6838 & n22517 ) ;
  assign n22519 = n4858 | n9921 ;
  assign n22520 = n12167 ^ n1255 ^ 1'b0 ;
  assign n22521 = n8905 | n22520 ;
  assign n22522 = n9555 ^ n1991 ^ 1'b0 ;
  assign n22523 = n6516 ^ n1613 ^ 1'b0 ;
  assign n22524 = n13079 | n22523 ;
  assign n22525 = n10313 ^ n9537 ^ 1'b0 ;
  assign n22526 = n18465 & n22525 ;
  assign n22527 = n19002 & n22526 ;
  assign n22528 = n20181 ^ n4211 ^ 1'b0 ;
  assign n22529 = n1310 | n6934 ;
  assign n22530 = n4872 & ~n9472 ;
  assign n22531 = ~n22529 & n22530 ;
  assign n22532 = n10447 | n18926 ;
  assign n22533 = n3933 | n22532 ;
  assign n22534 = n22533 ^ n8253 ^ 1'b0 ;
  assign n22535 = n18722 ^ x158 ^ 1'b0 ;
  assign n22536 = n18803 & ~n22535 ;
  assign n22538 = n1761 | n13115 ;
  assign n22537 = n2327 & ~n20551 ;
  assign n22539 = n22538 ^ n22537 ^ 1'b0 ;
  assign n22540 = n10046 & n19180 ;
  assign n22541 = ( n286 & n16949 ) | ( n286 & ~n17565 ) | ( n16949 & ~n17565 ) ;
  assign n22542 = ( n6831 & n9192 ) | ( n6831 & n11865 ) | ( n9192 & n11865 ) ;
  assign n22543 = ~n8705 & n8752 ;
  assign n22544 = n2563 & n22543 ;
  assign n22545 = n14677 ^ n13521 ^ 1'b0 ;
  assign n22546 = n4764 & n22545 ;
  assign n22547 = ~n4918 & n22546 ;
  assign n22548 = n2479 & n12472 ;
  assign n22549 = n22434 ^ n6668 ^ 1'b0 ;
  assign n22550 = n22549 ^ n19430 ^ 1'b0 ;
  assign n22551 = n14865 ^ n7787 ^ 1'b0 ;
  assign n22552 = n8850 | n22551 ;
  assign n22553 = n20219 ^ n7690 ^ 1'b0 ;
  assign n22554 = n14924 & ~n22553 ;
  assign n22555 = ~n604 & n15179 ;
  assign n22556 = n10973 | n22555 ;
  assign n22557 = n8831 | n19398 ;
  assign n22558 = ~n6597 & n18934 ;
  assign n22559 = n12373 ^ n7540 ^ 1'b0 ;
  assign n22560 = n22559 ^ n19442 ^ 1'b0 ;
  assign n22561 = n3518 & ~n7406 ;
  assign n22562 = n20330 & n22561 ;
  assign n22563 = ~n5523 & n10045 ;
  assign n22564 = ( n2991 & n6944 ) | ( n2991 & n22563 ) | ( n6944 & n22563 ) ;
  assign n22565 = n9890 & ~n22564 ;
  assign n22566 = n1515 & n22565 ;
  assign n22567 = ( n1038 & ~n2610 ) | ( n1038 & n5581 ) | ( ~n2610 & n5581 ) ;
  assign n22568 = ~n4528 & n18616 ;
  assign n22569 = n18987 ^ n6526 ^ 1'b0 ;
  assign n22570 = ( n22567 & ~n22568 ) | ( n22567 & n22569 ) | ( ~n22568 & n22569 ) ;
  assign n22571 = ( n2405 & ~n22566 ) | ( n2405 & n22570 ) | ( ~n22566 & n22570 ) ;
  assign n22572 = n12189 ^ n9345 ^ n8893 ;
  assign n22573 = n22572 ^ n21526 ^ 1'b0 ;
  assign n22574 = n22573 ^ n5765 ^ 1'b0 ;
  assign n22575 = n2988 & ~n22574 ;
  assign n22576 = ~n22571 & n22575 ;
  assign n22577 = n20196 ^ n16363 ^ n9561 ;
  assign n22578 = ( n2843 & n18371 ) | ( n2843 & ~n18692 ) | ( n18371 & ~n18692 ) ;
  assign n22579 = n7447 & n14486 ;
  assign n22580 = n289 & ~n1347 ;
  assign n22581 = n8294 | n10865 ;
  assign n22582 = n17654 ^ n2084 ^ 1'b0 ;
  assign n22583 = ~n8458 & n22582 ;
  assign n22584 = n758 | n22583 ;
  assign n22585 = n277 & n10425 ;
  assign n22586 = n22585 ^ n6842 ^ 1'b0 ;
  assign n22587 = ~n19018 & n22586 ;
  assign n22588 = ~n3998 & n22587 ;
  assign n22589 = n21746 ^ n8421 ^ 1'b0 ;
  assign n22590 = ~n13513 & n22589 ;
  assign n22591 = n14845 ^ n1458 ^ 1'b0 ;
  assign n22592 = ~n719 & n4911 ;
  assign n22593 = ~n3978 & n22592 ;
  assign n22594 = n21785 ^ n5814 ^ 1'b0 ;
  assign n22595 = ~n22593 & n22594 ;
  assign n22596 = n20791 & n22595 ;
  assign n22597 = n5805 ^ n4676 ^ 1'b0 ;
  assign n22598 = ~n12051 & n22597 ;
  assign n22599 = n22598 ^ n15717 ^ 1'b0 ;
  assign n22600 = n7488 | n22599 ;
  assign n22601 = n22600 ^ n6646 ^ 1'b0 ;
  assign n22602 = n3468 ^ n2775 ^ 1'b0 ;
  assign n22605 = ( n1173 & n6694 ) | ( n1173 & n7807 ) | ( n6694 & n7807 ) ;
  assign n22603 = n14644 & ~n16861 ;
  assign n22604 = ~n5599 & n22603 ;
  assign n22606 = n22605 ^ n22604 ^ n12514 ;
  assign n22607 = n20080 ^ n9094 ^ 1'b0 ;
  assign n22608 = n22606 & n22607 ;
  assign n22609 = n3299 | n19658 ;
  assign n22610 = n5866 & ~n22609 ;
  assign n22611 = n9358 & ~n22610 ;
  assign n22612 = n22611 ^ n2437 ^ 1'b0 ;
  assign n22613 = n20107 ^ n14310 ^ 1'b0 ;
  assign n22614 = n7719 & ~n13661 ;
  assign n22615 = ( n1298 & n4722 ) | ( n1298 & ~n21556 ) | ( n4722 & ~n21556 ) ;
  assign n22616 = n2246 & n2306 ;
  assign n22617 = n22616 ^ n469 ^ 1'b0 ;
  assign n22618 = n10455 & ~n22617 ;
  assign n22619 = n1733 & n2973 ;
  assign n22620 = ~n2915 & n3118 ;
  assign n22621 = n9339 & n22620 ;
  assign n22622 = n22619 | n22621 ;
  assign n22623 = n3480 & ~n12275 ;
  assign n22624 = n22623 ^ n6432 ^ 1'b0 ;
  assign n22625 = ( n3568 & n5672 ) | ( n3568 & n7723 ) | ( n5672 & n7723 ) ;
  assign n22626 = n22625 ^ n13167 ^ 1'b0 ;
  assign n22627 = ( n5748 & n20983 ) | ( n5748 & n22626 ) | ( n20983 & n22626 ) ;
  assign n22628 = n3094 & ~n6325 ;
  assign n22629 = x36 | n4320 ;
  assign n22630 = ( n2169 & n22628 ) | ( n2169 & ~n22629 ) | ( n22628 & ~n22629 ) ;
  assign n22631 = n6522 & n22630 ;
  assign n22632 = n15595 & ~n20086 ;
  assign n22633 = ~n5865 & n22632 ;
  assign n22634 = n9496 ^ n5400 ^ 1'b0 ;
  assign n22635 = ( n2534 & ~n7857 ) | ( n2534 & n11802 ) | ( ~n7857 & n11802 ) ;
  assign n22636 = n18807 & ~n22635 ;
  assign n22637 = n6100 & n15338 ;
  assign n22638 = n22637 ^ n11959 ^ 1'b0 ;
  assign n22639 = n10300 & ~n10512 ;
  assign n22640 = ~n8169 & n22639 ;
  assign n22641 = ~n12503 & n22640 ;
  assign n22642 = n984 & n6788 ;
  assign n22643 = n3850 & n22642 ;
  assign n22644 = n6938 & ~n22643 ;
  assign n22645 = n22644 ^ n2786 ^ 1'b0 ;
  assign n22646 = ( ~n5244 & n5482 ) | ( ~n5244 & n5853 ) | ( n5482 & n5853 ) ;
  assign n22647 = ( n1242 & n4287 ) | ( n1242 & n22646 ) | ( n4287 & n22646 ) ;
  assign n22648 = n6145 ^ n546 ^ 1'b0 ;
  assign n22649 = ~n22647 & n22648 ;
  assign n22650 = ( n15773 & n22645 ) | ( n15773 & n22649 ) | ( n22645 & n22649 ) ;
  assign n22651 = n15986 ^ n12282 ^ 1'b0 ;
  assign n22652 = ( n2100 & n3882 ) | ( n2100 & n22651 ) | ( n3882 & n22651 ) ;
  assign n22654 = n8164 ^ n1837 ^ 1'b0 ;
  assign n22655 = ~n1105 & n22654 ;
  assign n22653 = n1595 & n4722 ;
  assign n22656 = n22655 ^ n22653 ^ 1'b0 ;
  assign n22658 = n4547 ^ n275 ^ 1'b0 ;
  assign n22659 = ~n1758 & n9986 ;
  assign n22660 = ~n15585 & n22659 ;
  assign n22661 = n22658 & n22660 ;
  assign n22657 = n3927 | n20340 ;
  assign n22662 = n22661 ^ n22657 ^ 1'b0 ;
  assign n22663 = ~n6045 & n13448 ;
  assign n22664 = n13655 & n22663 ;
  assign n22665 = n2002 ^ x185 ^ 1'b0 ;
  assign n22666 = ~n22664 & n22665 ;
  assign n22667 = ~n886 & n6467 ;
  assign n22668 = ~n7853 & n22667 ;
  assign n22669 = ( n1132 & n5068 ) | ( n1132 & ~n5798 ) | ( n5068 & ~n5798 ) ;
  assign n22670 = n22669 ^ n17181 ^ 1'b0 ;
  assign n22671 = n22668 | n22670 ;
  assign n22672 = ( n20455 & n22666 ) | ( n20455 & ~n22671 ) | ( n22666 & ~n22671 ) ;
  assign n22673 = n2421 ^ n2302 ^ 1'b0 ;
  assign n22674 = n3980 & n22673 ;
  assign n22675 = ~n19442 & n22674 ;
  assign n22676 = n22675 ^ n11666 ^ 1'b0 ;
  assign n22677 = n8696 ^ n4172 ^ 1'b0 ;
  assign n22678 = n22677 ^ n14335 ^ n8906 ;
  assign n22679 = ( n19237 & n20155 ) | ( n19237 & n22678 ) | ( n20155 & n22678 ) ;
  assign n22680 = n7701 ^ n5216 ^ 1'b0 ;
  assign n22681 = n11064 ^ x199 ^ 1'b0 ;
  assign n22682 = n17666 & ~n22681 ;
  assign n22683 = ( n4975 & n8381 ) | ( n4975 & n22682 ) | ( n8381 & n22682 ) ;
  assign n22684 = n11421 ^ n6479 ^ 1'b0 ;
  assign n22685 = n4458 & ~n11585 ;
  assign n22686 = n22685 ^ x91 ^ 1'b0 ;
  assign n22687 = n12177 ^ n1760 ^ 1'b0 ;
  assign n22688 = n21915 & ~n22687 ;
  assign n22689 = n16830 & ~n22688 ;
  assign n22690 = n9401 & n22689 ;
  assign n22691 = n10261 & n12444 ;
  assign n22692 = n8245 ^ n7974 ^ 1'b0 ;
  assign n22693 = n1486 & n22692 ;
  assign n22694 = ( n9399 & n22691 ) | ( n9399 & n22693 ) | ( n22691 & n22693 ) ;
  assign n22695 = ~n15630 & n22694 ;
  assign n22696 = n5754 & ~n6961 ;
  assign n22697 = n16885 & ~n22696 ;
  assign n22698 = n22697 ^ n1935 ^ 1'b0 ;
  assign n22699 = n5043 & ~n22083 ;
  assign n22700 = n22699 ^ n20800 ^ 1'b0 ;
  assign n22701 = n432 & ~n16542 ;
  assign n22702 = ( n2907 & ~n10774 ) | ( n2907 & n18793 ) | ( ~n10774 & n18793 ) ;
  assign n22703 = n2044 & ~n7609 ;
  assign n22704 = n4104 ^ n1895 ^ x184 ;
  assign n22705 = n7126 ^ n4666 ^ 1'b0 ;
  assign n22706 = n14998 | n22705 ;
  assign n22707 = n22704 | n22706 ;
  assign n22708 = ~n4947 & n17544 ;
  assign n22709 = ~n8048 & n22708 ;
  assign n22710 = ~n16810 & n18643 ;
  assign n22711 = n22709 & n22710 ;
  assign n22712 = n9231 & n19116 ;
  assign n22713 = ~n5366 & n22712 ;
  assign n22714 = n21481 | n22713 ;
  assign n22715 = n5744 ^ n4216 ^ 1'b0 ;
  assign n22716 = n1467 & n11471 ;
  assign n22717 = n22715 & ~n22716 ;
  assign n22718 = n22717 ^ n16617 ^ 1'b0 ;
  assign n22720 = ( n367 & n1496 ) | ( n367 & n6309 ) | ( n1496 & n6309 ) ;
  assign n22719 = n13010 ^ n7670 ^ 1'b0 ;
  assign n22721 = n22720 ^ n22719 ^ 1'b0 ;
  assign n22722 = ~n2392 & n20624 ;
  assign n22723 = n22722 ^ n3776 ^ x70 ;
  assign n22724 = n16521 ^ n13592 ^ 1'b0 ;
  assign n22725 = n7097 & ~n10557 ;
  assign n22726 = n22724 & n22725 ;
  assign n22727 = ~n877 & n10865 ;
  assign n22728 = n22727 ^ n20637 ^ 1'b0 ;
  assign n22729 = n3782 ^ n3592 ^ n2093 ;
  assign n22730 = ( n10826 & ~n13079 ) | ( n10826 & n22729 ) | ( ~n13079 & n22729 ) ;
  assign n22731 = n8084 | n10534 ;
  assign n22732 = n4060 & ~n22731 ;
  assign n22733 = n20411 ^ n18257 ^ 1'b0 ;
  assign n22734 = n21118 & ~n22733 ;
  assign n22735 = n16341 & n22734 ;
  assign n22736 = n11810 & ~n22735 ;
  assign n22737 = n20787 ^ n14241 ^ 1'b0 ;
  assign n22738 = x118 & n9252 ;
  assign n22739 = ( n7876 & n16307 ) | ( n7876 & ~n22738 ) | ( n16307 & ~n22738 ) ;
  assign n22740 = n3487 & ~n7029 ;
  assign n22741 = n2457 & n22740 ;
  assign n22742 = n1996 & n6198 ;
  assign n22743 = ~n15535 & n19121 ;
  assign n22744 = n22743 ^ n14985 ^ 1'b0 ;
  assign n22745 = ~n22742 & n22744 ;
  assign n22746 = n22745 ^ n7338 ^ 1'b0 ;
  assign n22747 = n22746 ^ n6906 ^ 1'b0 ;
  assign n22748 = ~n22741 & n22747 ;
  assign n22749 = ( n6461 & n9788 ) | ( n6461 & ~n15268 ) | ( n9788 & ~n15268 ) ;
  assign n22750 = n5229 & n18176 ;
  assign n22751 = n22749 & n22750 ;
  assign n22752 = n22751 ^ n2819 ^ 1'b0 ;
  assign n22753 = ( n1499 & ~n2191 ) | ( n1499 & n8141 ) | ( ~n2191 & n8141 ) ;
  assign n22754 = n22753 ^ n18058 ^ 1'b0 ;
  assign n22755 = n10584 | n22754 ;
  assign n22756 = ~n4347 & n9911 ;
  assign n22757 = ~n4880 & n19312 ;
  assign n22758 = n5420 & n19787 ;
  assign n22759 = n22758 ^ n20157 ^ 1'b0 ;
  assign n22760 = n21388 ^ n11920 ^ 1'b0 ;
  assign n22761 = ( n1376 & ~n22759 ) | ( n1376 & n22760 ) | ( ~n22759 & n22760 ) ;
  assign n22762 = n9358 ^ n7844 ^ 1'b0 ;
  assign n22763 = n853 & n4196 ;
  assign n22764 = n393 & n22763 ;
  assign n22765 = n7492 | n22764 ;
  assign n22766 = n22765 ^ n6151 ^ 1'b0 ;
  assign n22767 = n853 & ~n22766 ;
  assign n22768 = n22767 ^ n1457 ^ 1'b0 ;
  assign n22769 = n12835 | n22768 ;
  assign n22770 = n20219 ^ n4931 ^ n4636 ;
  assign n22771 = n489 & n3700 ;
  assign n22772 = ~n1328 & n22771 ;
  assign n22773 = n6663 & ~n22772 ;
  assign n22774 = n10274 & n22773 ;
  assign n22775 = n6484 ^ n5476 ^ 1'b0 ;
  assign n22776 = n11959 | n22775 ;
  assign n22777 = n22193 ^ n7167 ^ 1'b0 ;
  assign n22778 = n2574 ^ x56 ^ 1'b0 ;
  assign n22779 = ( n3536 & ~n6192 ) | ( n3536 & n22778 ) | ( ~n6192 & n22778 ) ;
  assign n22780 = n22779 ^ n4460 ^ n1353 ;
  assign n22781 = n9222 & ~n22780 ;
  assign n22782 = n1996 | n6943 ;
  assign n22783 = n22781 | n22782 ;
  assign n22784 = n6136 | n12564 ;
  assign n22785 = ~n3154 & n9711 ;
  assign n22786 = n283 | n2617 ;
  assign n22787 = n15971 | n22786 ;
  assign n22788 = n22787 ^ n9780 ^ 1'b0 ;
  assign n22789 = ~n22785 & n22788 ;
  assign n22790 = ~n1821 & n22789 ;
  assign n22791 = n5725 & n22790 ;
  assign n22792 = n22791 ^ n3692 ^ 1'b0 ;
  assign n22793 = n22784 | n22792 ;
  assign n22794 = n369 | n13787 ;
  assign n22795 = n6700 | n22794 ;
  assign n22796 = n5493 & ~n19030 ;
  assign n22797 = ~n22795 & n22796 ;
  assign n22798 = x170 & n14922 ;
  assign n22799 = n17557 & n22798 ;
  assign n22800 = n14776 ^ n14696 ^ n10811 ;
  assign n22801 = ~n15988 & n18147 ;
  assign n22802 = ~n22800 & n22801 ;
  assign n22803 = n20643 ^ n1629 ^ 1'b0 ;
  assign n22804 = n22803 ^ n20013 ^ n5241 ;
  assign n22805 = n936 & n21634 ;
  assign n22806 = n22805 ^ n17778 ^ 1'b0 ;
  assign n22807 = ( n7110 & n21682 ) | ( n7110 & ~n22806 ) | ( n21682 & ~n22806 ) ;
  assign n22808 = n17282 ^ n16429 ^ 1'b0 ;
  assign n22809 = n4259 | n13248 ;
  assign n22810 = n22809 ^ n20034 ^ 1'b0 ;
  assign n22811 = n5790 | n8844 ;
  assign n22812 = n22811 ^ n15388 ^ 1'b0 ;
  assign n22813 = n17120 ^ x186 ^ 1'b0 ;
  assign n22814 = ~n4686 & n22813 ;
  assign n22815 = n9028 ^ n749 ^ 1'b0 ;
  assign n22816 = n22814 & ~n22815 ;
  assign n22817 = x242 & n22816 ;
  assign n22818 = ~n787 & n22817 ;
  assign n22819 = n22818 ^ n6941 ^ 1'b0 ;
  assign n22820 = n9846 ^ n8345 ^ 1'b0 ;
  assign n22821 = n22604 ^ n8317 ^ n1930 ;
  assign n22822 = n14135 ^ n3688 ^ 1'b0 ;
  assign n22823 = ~n17991 & n22822 ;
  assign n22824 = ( n2452 & n14179 ) | ( n2452 & n15793 ) | ( n14179 & n15793 ) ;
  assign n22825 = n8274 | n22824 ;
  assign n22826 = n22825 ^ n10063 ^ 1'b0 ;
  assign n22827 = n8721 & n10777 ;
  assign n22828 = n22827 ^ n2718 ^ 1'b0 ;
  assign n22829 = n4518 | n22828 ;
  assign n22830 = n4848 & ~n22829 ;
  assign n22833 = ~n529 & n7303 ;
  assign n22831 = n6488 | n10557 ;
  assign n22832 = n22831 ^ n9959 ^ 1'b0 ;
  assign n22834 = n22833 ^ n22832 ^ n6206 ;
  assign n22835 = n6365 & ~n6772 ;
  assign n22836 = n22835 ^ n11872 ^ 1'b0 ;
  assign n22837 = ~n16129 & n22836 ;
  assign n22838 = n5931 ^ n3321 ^ 1'b0 ;
  assign n22839 = n7879 | n18940 ;
  assign n22840 = n22838 | n22839 ;
  assign n22841 = n18339 & n22840 ;
  assign n22842 = ~n14989 & n22841 ;
  assign n22843 = n1478 & ~n12772 ;
  assign n22844 = n2930 & ~n7841 ;
  assign n22845 = n3166 | n22844 ;
  assign n22846 = n4865 & ~n17110 ;
  assign n22847 = n8968 & n22846 ;
  assign n22848 = n9222 & ~n12728 ;
  assign n22849 = ~n20252 & n22848 ;
  assign n22851 = n8419 ^ n8152 ^ 1'b0 ;
  assign n22852 = x204 & ~n22851 ;
  assign n22850 = n5793 | n20741 ;
  assign n22853 = n22852 ^ n22850 ^ 1'b0 ;
  assign n22854 = n22853 ^ n17154 ^ 1'b0 ;
  assign n22855 = n11281 ^ n4333 ^ 1'b0 ;
  assign n22856 = n7400 ^ n7001 ^ 1'b0 ;
  assign n22857 = ~n22855 & n22856 ;
  assign n22858 = n3111 & n7743 ;
  assign n22859 = ~n12154 & n22858 ;
  assign n22860 = n3326 & n22859 ;
  assign n22861 = n22860 ^ n5157 ^ 1'b0 ;
  assign n22862 = n3095 & ~n6599 ;
  assign n22863 = n7165 & n22862 ;
  assign n22865 = n3077 & n10595 ;
  assign n22864 = n1386 & n5748 ;
  assign n22866 = n22865 ^ n22864 ^ n3958 ;
  assign n22869 = n16371 ^ n9583 ^ 1'b0 ;
  assign n22870 = n22869 ^ n20648 ^ 1'b0 ;
  assign n22867 = n9215 & ~n9848 ;
  assign n22868 = ~n1965 & n22867 ;
  assign n22871 = n22870 ^ n22868 ^ n12990 ;
  assign n22872 = n3743 ^ n557 ^ 1'b0 ;
  assign n22873 = ~n6713 & n22872 ;
  assign n22874 = ~n3324 & n22873 ;
  assign n22875 = n22874 ^ n20166 ^ 1'b0 ;
  assign n22876 = n8731 ^ x22 ^ 1'b0 ;
  assign n22877 = n10222 & ~n22876 ;
  assign n22880 = n2941 ^ n886 ^ 1'b0 ;
  assign n22881 = ~n8054 & n22880 ;
  assign n22878 = n2324 | n11367 ;
  assign n22879 = n8416 | n22878 ;
  assign n22882 = n22881 ^ n22879 ^ 1'b0 ;
  assign n22883 = ( n3542 & n12253 ) | ( n3542 & n15756 ) | ( n12253 & n15756 ) ;
  assign n22884 = n593 | n2592 ;
  assign n22885 = n16073 | n22884 ;
  assign n22886 = n2846 | n22885 ;
  assign n22887 = n22883 & n22886 ;
  assign n22888 = ~n1843 & n4923 ;
  assign n22889 = ~n906 & n22888 ;
  assign n22890 = ~n15284 & n22889 ;
  assign n22891 = ~n7597 & n22890 ;
  assign n22894 = x81 & n8346 ;
  assign n22893 = n5112 | n6472 ;
  assign n22895 = n22894 ^ n22893 ^ 1'b0 ;
  assign n22892 = x185 & ~n11196 ;
  assign n22896 = n22895 ^ n22892 ^ 1'b0 ;
  assign n22897 = ( n3263 & n10143 ) | ( n3263 & ~n17122 ) | ( n10143 & ~n17122 ) ;
  assign n22898 = n13754 & n22897 ;
  assign n22899 = n22898 ^ n4718 ^ 1'b0 ;
  assign n22900 = n1439 & ~n22899 ;
  assign n22901 = n4966 & ~n12002 ;
  assign n22902 = ( n3638 & n12223 ) | ( n3638 & n22901 ) | ( n12223 & n22901 ) ;
  assign n22903 = n22902 ^ n7572 ^ 1'b0 ;
  assign n22904 = ~x170 & n22903 ;
  assign n22905 = n20868 ^ n8484 ^ 1'b0 ;
  assign n22906 = ~n1822 & n2799 ;
  assign n22907 = ( n874 & n5164 ) | ( n874 & n22906 ) | ( n5164 & n22906 ) ;
  assign n22908 = n524 & n22907 ;
  assign n22909 = n22908 ^ n2834 ^ 1'b0 ;
  assign n22910 = n12573 ^ n6573 ^ 1'b0 ;
  assign n22911 = n7323 & ~n22910 ;
  assign n22912 = ( n22803 & n22909 ) | ( n22803 & n22911 ) | ( n22909 & n22911 ) ;
  assign n22913 = n9691 & n13978 ;
  assign n22914 = n22913 ^ n13458 ^ 1'b0 ;
  assign n22915 = n22914 ^ n1315 ^ 1'b0 ;
  assign n22916 = x193 & ~n18762 ;
  assign n22917 = ~n15362 & n22916 ;
  assign n22918 = ~n4421 & n6646 ;
  assign n22919 = ~n14119 & n22918 ;
  assign n22920 = ~n653 & n14338 ;
  assign n22921 = n22920 ^ n9200 ^ 1'b0 ;
  assign n22922 = ~n3827 & n17771 ;
  assign n22925 = n3804 ^ n354 ^ 1'b0 ;
  assign n22926 = ~n9969 & n22925 ;
  assign n22927 = n6319 | n22926 ;
  assign n22923 = x91 | n19295 ;
  assign n22924 = n6966 & ~n22923 ;
  assign n22928 = n22927 ^ n22924 ^ x229 ;
  assign n22929 = n4831 & ~n12386 ;
  assign n22930 = ~n5092 & n22929 ;
  assign n22931 = ~n292 & n12261 ;
  assign n22932 = n22930 & n22931 ;
  assign n22933 = n11472 & n22932 ;
  assign n22934 = n3755 & ~n22933 ;
  assign n22935 = n3822 & n6021 ;
  assign n22936 = n22935 ^ n10226 ^ 1'b0 ;
  assign n22937 = n3415 & ~n22936 ;
  assign n22938 = n14935 ^ n9709 ^ 1'b0 ;
  assign n22939 = n17769 & n22938 ;
  assign n22940 = n5861 ^ n681 ^ 1'b0 ;
  assign n22941 = n22940 ^ n18188 ^ n7015 ;
  assign n22942 = n4907 & ~n12633 ;
  assign n22943 = ~n14110 & n22942 ;
  assign n22946 = n7894 ^ n7598 ^ 1'b0 ;
  assign n22947 = n22150 & n22946 ;
  assign n22944 = n4842 & ~n8395 ;
  assign n22945 = ~n12908 & n22944 ;
  assign n22948 = n22947 ^ n22945 ^ n21502 ;
  assign n22949 = n15985 ^ n6907 ^ 1'b0 ;
  assign n22950 = n20197 & n22949 ;
  assign n22951 = n12419 ^ n6838 ^ 1'b0 ;
  assign n22952 = n5448 & n22951 ;
  assign n22953 = n22952 ^ n824 ^ 1'b0 ;
  assign n22954 = n1571 | n9247 ;
  assign n22955 = n22954 ^ n11836 ^ 1'b0 ;
  assign n22956 = n12909 | n13924 ;
  assign n22957 = n22956 ^ n5544 ^ 1'b0 ;
  assign n22958 = ~n1558 & n22957 ;
  assign n22959 = ( n4171 & ~n18942 ) | ( n4171 & n22958 ) | ( ~n18942 & n22958 ) ;
  assign n22960 = n2054 & n2664 ;
  assign n22961 = n22960 ^ n1661 ^ 1'b0 ;
  assign n22962 = n18069 ^ n15666 ^ 1'b0 ;
  assign n22963 = n22961 | n22962 ;
  assign n22964 = n22959 & ~n22963 ;
  assign n22965 = n4793 & ~n4872 ;
  assign n22966 = ~n5549 & n22965 ;
  assign n22967 = ~n19470 & n22966 ;
  assign n22968 = ~n18914 & n22967 ;
  assign n22969 = ( ~n1365 & n8769 ) | ( ~n1365 & n10794 ) | ( n8769 & n10794 ) ;
  assign n22970 = ~n2651 & n16883 ;
  assign n22971 = n22970 ^ n498 ^ 1'b0 ;
  assign n22972 = ~n1291 & n22971 ;
  assign n22973 = ( n3307 & n22969 ) | ( n3307 & n22972 ) | ( n22969 & n22972 ) ;
  assign n22974 = n4995 & ~n22973 ;
  assign n22975 = n14371 ^ n8226 ^ 1'b0 ;
  assign n22976 = ~n371 & n22975 ;
  assign n22977 = n22976 ^ n14233 ^ 1'b0 ;
  assign n22978 = n1181 | n7311 ;
  assign n22979 = n445 & ~n20730 ;
  assign n22980 = n22978 & n22979 ;
  assign n22981 = n22980 ^ n11519 ^ n10400 ;
  assign n22982 = n15158 ^ n2480 ^ 1'b0 ;
  assign n22983 = n14134 ^ n11345 ^ 1'b0 ;
  assign n22984 = n12097 | n17568 ;
  assign n22985 = n438 & n2447 ;
  assign n22986 = n13343 | n22985 ;
  assign n22987 = n22986 ^ n1097 ^ 1'b0 ;
  assign n22988 = n22987 ^ n2259 ^ n1575 ;
  assign n22989 = n12624 & ~n22988 ;
  assign n22990 = n22989 ^ n20671 ^ 1'b0 ;
  assign n22991 = n5989 | n6512 ;
  assign n22992 = n22991 ^ n16987 ^ 1'b0 ;
  assign n22993 = ~n7178 & n22992 ;
  assign n22994 = n5304 ^ n3668 ^ 1'b0 ;
  assign n22995 = n22994 ^ n8384 ^ 1'b0 ;
  assign n22996 = ( n3425 & n16830 ) | ( n3425 & n20889 ) | ( n16830 & n20889 ) ;
  assign n22997 = n22996 ^ n5054 ^ n4803 ;
  assign n22998 = n20643 ^ n9183 ^ 1'b0 ;
  assign n22999 = n16415 ^ n6618 ^ 1'b0 ;
  assign n23004 = ( n772 & n1397 ) | ( n772 & ~n20431 ) | ( n1397 & ~n20431 ) ;
  assign n23000 = ~n2630 & n7905 ;
  assign n23001 = n10806 & n23000 ;
  assign n23002 = n15994 & ~n23001 ;
  assign n23003 = n17971 & n23002 ;
  assign n23005 = n23004 ^ n23003 ^ 1'b0 ;
  assign n23006 = ( n4643 & ~n22999 ) | ( n4643 & n23005 ) | ( ~n22999 & n23005 ) ;
  assign n23007 = ( n585 & n12427 ) | ( n585 & ~n15632 ) | ( n12427 & ~n15632 ) ;
  assign n23008 = n21075 ^ n12812 ^ 1'b0 ;
  assign n23009 = ~n23007 & n23008 ;
  assign n23010 = n1033 | n16891 ;
  assign n23011 = n18832 | n23010 ;
  assign n23012 = n7569 & n23011 ;
  assign n23013 = n10830 ^ n9518 ^ n305 ;
  assign n23014 = n1871 & n23013 ;
  assign n23015 = n23014 ^ n17953 ^ 1'b0 ;
  assign n23016 = ( n3321 & n7128 ) | ( n3321 & n10216 ) | ( n7128 & n10216 ) ;
  assign n23017 = ( n7833 & n11640 ) | ( n7833 & n23016 ) | ( n11640 & n23016 ) ;
  assign n23018 = n11263 & n21615 ;
  assign n23019 = ~n4434 & n23018 ;
  assign n23020 = n20260 & ~n23019 ;
  assign n23021 = n3249 & n12755 ;
  assign n23022 = n12776 & n23021 ;
  assign n23023 = ~x65 & n20420 ;
  assign n23024 = n5590 | n20036 ;
  assign n23025 = ( n17313 & ~n23023 ) | ( n17313 & n23024 ) | ( ~n23023 & n23024 ) ;
  assign n23026 = n1377 & ~n4508 ;
  assign n23027 = n789 & n23026 ;
  assign n23028 = n23027 ^ n15986 ^ 1'b0 ;
  assign n23029 = n1524 & n3672 ;
  assign n23030 = ~n793 & n3611 ;
  assign n23031 = n4438 & n23030 ;
  assign n23032 = n23031 ^ n20325 ^ n3627 ;
  assign n23033 = n23029 & ~n23032 ;
  assign n23034 = n16138 ^ n351 ^ 1'b0 ;
  assign n23035 = ~n16569 & n23034 ;
  assign n23036 = n1603 ^ n614 ^ 1'b0 ;
  assign n23037 = x0 | n23036 ;
  assign n23038 = n12236 | n23037 ;
  assign n23039 = n23035 | n23038 ;
  assign n23040 = n7258 & n23039 ;
  assign n23041 = n23040 ^ n21930 ^ 1'b0 ;
  assign n23042 = n13052 ^ n1955 ^ 1'b0 ;
  assign n23043 = ~n23041 & n23042 ;
  assign n23044 = n23043 ^ n10749 ^ n3415 ;
  assign n23045 = x36 & n558 ;
  assign n23046 = ~n10056 & n23045 ;
  assign n23047 = n23046 ^ n16224 ^ 1'b0 ;
  assign n23048 = n8834 & n8898 ;
  assign n23049 = n23048 ^ n19002 ^ 1'b0 ;
  assign n23050 = n10214 & n14339 ;
  assign n23051 = n23050 ^ n13643 ^ 1'b0 ;
  assign n23052 = n3135 | n21351 ;
  assign n23053 = n23051 & ~n23052 ;
  assign n23054 = ~n2131 & n10675 ;
  assign n23055 = n1733 & n23054 ;
  assign n23056 = n3067 & ~n18603 ;
  assign n23057 = n23055 & n23056 ;
  assign n23058 = ( ~n3490 & n21231 ) | ( ~n3490 & n23057 ) | ( n21231 & n23057 ) ;
  assign n23059 = n9691 ^ n1296 ^ 1'b0 ;
  assign n23060 = n23059 ^ n9437 ^ n6686 ;
  assign n23061 = ( ~n593 & n22741 ) | ( ~n593 & n23060 ) | ( n22741 & n23060 ) ;
  assign n23062 = n5656 | n10193 ;
  assign n23063 = n23033 & n23062 ;
  assign n23065 = n4644 & ~n12922 ;
  assign n23066 = n23065 ^ n7487 ^ 1'b0 ;
  assign n23067 = n20533 ^ n15009 ^ 1'b0 ;
  assign n23068 = n23066 & n23067 ;
  assign n23064 = n577 & ~n6607 ;
  assign n23069 = n23068 ^ n23064 ^ 1'b0 ;
  assign n23070 = n8523 ^ n5947 ^ 1'b0 ;
  assign n23071 = n18406 & ~n23070 ;
  assign n23072 = n3814 & n11913 ;
  assign n23073 = n3018 ^ n2537 ^ 1'b0 ;
  assign n23074 = x58 & n23073 ;
  assign n23075 = n23074 ^ n5085 ^ 1'b0 ;
  assign n23076 = n23072 | n23075 ;
  assign n23077 = n23076 ^ n12823 ^ 1'b0 ;
  assign n23078 = n23071 & n23077 ;
  assign n23079 = n19572 ^ n16307 ^ n10626 ;
  assign n23080 = n8570 | n9314 ;
  assign n23081 = n23080 ^ n1281 ^ 1'b0 ;
  assign n23082 = n23081 ^ n17181 ^ n9830 ;
  assign n23083 = n2078 & n5312 ;
  assign n23084 = ~n1377 & n23083 ;
  assign n23085 = n6690 ^ n4232 ^ 1'b0 ;
  assign n23086 = n3406 & ~n8535 ;
  assign n23087 = n23086 ^ n9456 ^ 1'b0 ;
  assign n23088 = n12929 & n23087 ;
  assign n23089 = n12456 ^ n395 ^ 1'b0 ;
  assign n23090 = n23088 & ~n23089 ;
  assign n23091 = n17433 & ~n22509 ;
  assign n23093 = n3421 & n5453 ;
  assign n23094 = ~n5592 & n23093 ;
  assign n23095 = n4253 & n23094 ;
  assign n23096 = n23095 ^ n20644 ^ 1'b0 ;
  assign n23092 = n462 & n3129 ;
  assign n23097 = n23096 ^ n23092 ^ 1'b0 ;
  assign n23098 = ~n7194 & n10661 ;
  assign n23099 = ~n12932 & n23098 ;
  assign n23100 = x15 | n11810 ;
  assign n23101 = n4144 | n23100 ;
  assign n23102 = ( ~x17 & n13448 ) | ( ~x17 & n21636 ) | ( n13448 & n21636 ) ;
  assign n23103 = n23102 ^ n14020 ^ 1'b0 ;
  assign n23104 = n23101 & ~n23103 ;
  assign n23105 = n5136 ^ n970 ^ 1'b0 ;
  assign n23106 = ~n3779 & n3986 ;
  assign n23107 = ( n6215 & n16126 ) | ( n6215 & n23106 ) | ( n16126 & n23106 ) ;
  assign n23108 = n23107 ^ n10255 ^ 1'b0 ;
  assign n23110 = n7870 & n9086 ;
  assign n23111 = ( ~n5724 & n12177 ) | ( ~n5724 & n23110 ) | ( n12177 & n23110 ) ;
  assign n23109 = n6341 | n10171 ;
  assign n23112 = n23111 ^ n23109 ^ 1'b0 ;
  assign n23113 = n6885 ^ n1382 ^ 1'b0 ;
  assign n23114 = n12548 & n23113 ;
  assign n23115 = n7925 & ~n15670 ;
  assign n23116 = n10141 ^ n4323 ^ 1'b0 ;
  assign n23117 = n23115 | n23116 ;
  assign n23118 = n16516 ^ n2675 ^ 1'b0 ;
  assign n23119 = n22286 ^ n15747 ^ n14394 ;
  assign n23120 = ~n9914 & n15115 ;
  assign n23121 = n23120 ^ n3138 ^ n2941 ;
  assign n23122 = ~n3189 & n4057 ;
  assign n23136 = ~n337 & n488 ;
  assign n23137 = ~n488 & n23136 ;
  assign n23138 = ~n4624 & n23137 ;
  assign n23123 = n3920 & ~n5013 ;
  assign n23124 = ~n3920 & n23123 ;
  assign n23125 = n661 & ~n23124 ;
  assign n23126 = n918 & n2399 ;
  assign n23127 = ~n918 & n23126 ;
  assign n23128 = n6238 & ~n23127 ;
  assign n23129 = n23127 & n23128 ;
  assign n23130 = n8500 | n19872 ;
  assign n23131 = n23130 ^ n16235 ^ 1'b0 ;
  assign n23132 = n8595 & n10845 ;
  assign n23133 = ~n23131 & n23132 ;
  assign n23134 = ( x69 & ~n23129 ) | ( x69 & n23133 ) | ( ~n23129 & n23133 ) ;
  assign n23135 = ~n23125 & n23134 ;
  assign n23139 = n23138 ^ n23135 ^ 1'b0 ;
  assign n23140 = ~n9269 & n13671 ;
  assign n23141 = ~n20060 & n23140 ;
  assign n23142 = n14697 ^ n10063 ^ n947 ;
  assign n23143 = n23142 ^ n5209 ^ 1'b0 ;
  assign n23144 = n4284 & ~n23143 ;
  assign n23145 = n3770 | n15312 ;
  assign n23146 = n23145 ^ n4840 ^ n998 ;
  assign n23147 = n14603 ^ n13574 ^ 1'b0 ;
  assign n23148 = n23147 ^ n10702 ^ 1'b0 ;
  assign n23149 = ( n23144 & n23146 ) | ( n23144 & ~n23148 ) | ( n23146 & ~n23148 ) ;
  assign n23150 = ~n773 & n19763 ;
  assign n23151 = n6385 & n10424 ;
  assign n23152 = ( ~n1082 & n4953 ) | ( ~n1082 & n21241 ) | ( n4953 & n21241 ) ;
  assign n23153 = ~n4275 & n23152 ;
  assign n23154 = n12201 ^ n7690 ^ 1'b0 ;
  assign n23155 = n13308 | n23154 ;
  assign n23156 = n23155 ^ n11950 ^ n3293 ;
  assign n23157 = n23153 & ~n23156 ;
  assign n23158 = n13698 ^ n12980 ^ 1'b0 ;
  assign n23159 = n23060 | n23158 ;
  assign n23160 = n1763 | n21359 ;
  assign n23161 = n23160 ^ n2543 ^ 1'b0 ;
  assign n23162 = n23161 ^ n9252 ^ 1'b0 ;
  assign n23163 = ~n1946 & n23162 ;
  assign n23164 = n8228 ^ n1965 ^ 1'b0 ;
  assign n23165 = n7220 & n23164 ;
  assign n23166 = n5052 ^ n2259 ^ n1415 ;
  assign n23167 = n6793 & n21173 ;
  assign n23168 = ~n21993 & n23167 ;
  assign n23169 = ( ~n9296 & n23166 ) | ( ~n9296 & n23168 ) | ( n23166 & n23168 ) ;
  assign n23170 = n15222 ^ n7990 ^ n3808 ;
  assign n23172 = n5589 ^ n5102 ^ 1'b0 ;
  assign n23171 = ~n1139 & n19799 ;
  assign n23173 = n23172 ^ n23171 ^ 1'b0 ;
  assign n23174 = n15296 ^ n7774 ^ 1'b0 ;
  assign n23175 = n23173 | n23174 ;
  assign n23176 = ~n4293 & n9638 ;
  assign n23177 = n3123 | n23176 ;
  assign n23178 = n23177 ^ n6602 ^ 1'b0 ;
  assign n23179 = n13536 & ~n23178 ;
  assign n23180 = n22830 ^ n3129 ^ n1600 ;
  assign n23181 = n7070 & n18271 ;
  assign n23182 = ~n12776 & n23181 ;
  assign n23183 = ( n8102 & n16862 ) | ( n8102 & n23182 ) | ( n16862 & n23182 ) ;
  assign n23184 = n22939 ^ n10736 ^ 1'b0 ;
  assign n23185 = n12678 | n23184 ;
  assign n23186 = n12170 ^ n4137 ^ 1'b0 ;
  assign n23187 = n23186 ^ n256 ^ 1'b0 ;
  assign n23188 = n15870 & n23187 ;
  assign n23189 = n23188 ^ n12002 ^ 1'b0 ;
  assign n23190 = n538 & ~n23189 ;
  assign n23192 = ~n1388 & n2970 ;
  assign n23191 = n1246 & ~n9983 ;
  assign n23193 = n23192 ^ n23191 ^ 1'b0 ;
  assign n23194 = n4563 & n22886 ;
  assign n23195 = n22317 | n23194 ;
  assign n23196 = n23195 ^ n16420 ^ 1'b0 ;
  assign n23197 = n8067 ^ n3003 ^ n1665 ;
  assign n23198 = n2314 ^ n347 ^ x16 ;
  assign n23199 = ( n22564 & n23197 ) | ( n22564 & n23198 ) | ( n23197 & n23198 ) ;
  assign n23200 = n17230 ^ n16310 ^ 1'b0 ;
  assign n23201 = n23199 | n23200 ;
  assign n23203 = n4065 | n12016 ;
  assign n23202 = n6736 ^ n5987 ^ n1055 ;
  assign n23204 = n23203 ^ n23202 ^ 1'b0 ;
  assign n23205 = n10081 & ~n23204 ;
  assign n23206 = n19525 ^ n17782 ^ 1'b0 ;
  assign n23207 = n7559 & n23206 ;
  assign n23208 = ~n686 & n8867 ;
  assign n23209 = n2619 & n23208 ;
  assign n23210 = n5350 | n23209 ;
  assign n23211 = n23210 ^ n6698 ^ 1'b0 ;
  assign n23212 = n23207 | n23211 ;
  assign n23213 = n11718 ^ n10397 ^ n3435 ;
  assign n23214 = ~n15350 & n23213 ;
  assign n23215 = n20420 | n23214 ;
  assign n23216 = n3495 & n23215 ;
  assign n23217 = n21863 & n23216 ;
  assign n23218 = n21921 ^ n12105 ^ 1'b0 ;
  assign n23219 = ~n8783 & n21105 ;
  assign n23220 = n10173 ^ n1272 ^ 1'b0 ;
  assign n23221 = n1724 | n14119 ;
  assign n23222 = ( n2116 & n6294 ) | ( n2116 & ~n23221 ) | ( n6294 & ~n23221 ) ;
  assign n23223 = ( ~n9831 & n9925 ) | ( ~n9831 & n23222 ) | ( n9925 & n23222 ) ;
  assign n23224 = n5947 ^ n3207 ^ 1'b0 ;
  assign n23225 = n2939 & ~n23224 ;
  assign n23226 = n5049 & n13265 ;
  assign n23227 = n6121 ^ n1736 ^ 1'b0 ;
  assign n23228 = n23226 | n23227 ;
  assign n23229 = n1535 ^ n1121 ^ 1'b0 ;
  assign n23230 = n23229 ^ n2709 ^ n2225 ;
  assign n23231 = n12444 & ~n23230 ;
  assign n23232 = ~n4050 & n23231 ;
  assign n23233 = n1088 & n3175 ;
  assign n23234 = n23233 ^ n759 ^ 1'b0 ;
  assign n23235 = n23234 ^ n21480 ^ 1'b0 ;
  assign n23236 = n23232 | n23235 ;
  assign n23237 = n11083 | n17453 ;
  assign n23238 = n23237 ^ n3263 ^ 1'b0 ;
  assign n23239 = n5013 | n15054 ;
  assign n23240 = n14551 ^ n1953 ^ 1'b0 ;
  assign n23241 = ~n2448 & n23240 ;
  assign n23242 = n23239 & n23241 ;
  assign n23243 = n577 & n14595 ;
  assign n23244 = n23243 ^ n13520 ^ 1'b0 ;
  assign n23245 = n16245 | n23244 ;
  assign n23246 = ( n19874 & n23242 ) | ( n19874 & n23245 ) | ( n23242 & n23245 ) ;
  assign n23247 = ( n907 & ~n4770 ) | ( n907 & n12464 ) | ( ~n4770 & n12464 ) ;
  assign n23248 = n13698 & ~n16861 ;
  assign n23249 = n4180 & n23248 ;
  assign n23250 = n17046 | n18893 ;
  assign n23251 = n7559 & ~n11706 ;
  assign n23255 = n3693 & ~n6422 ;
  assign n23252 = n8411 ^ n504 ^ 1'b0 ;
  assign n23253 = n7788 | n23252 ;
  assign n23254 = n13454 & n23253 ;
  assign n23256 = n23255 ^ n23254 ^ 1'b0 ;
  assign n23257 = n23256 ^ n20330 ^ n14256 ;
  assign n23258 = n19432 ^ n12236 ^ 1'b0 ;
  assign n23259 = n6388 | n8370 ;
  assign n23260 = n23259 ^ n8351 ^ 1'b0 ;
  assign n23261 = ~n15244 & n23260 ;
  assign n23262 = n23261 ^ n11517 ^ 1'b0 ;
  assign n23264 = n1633 | n3009 ;
  assign n23265 = n12475 & ~n23264 ;
  assign n23263 = n4950 & n5714 ;
  assign n23266 = n23265 ^ n23263 ^ 1'b0 ;
  assign n23267 = ( ~x41 & n575 ) | ( ~x41 & n3172 ) | ( n575 & n3172 ) ;
  assign n23268 = ( n3642 & ~n10689 ) | ( n3642 & n17030 ) | ( ~n10689 & n17030 ) ;
  assign n23269 = ~n16261 & n20522 ;
  assign n23270 = n7344 ^ n7323 ^ 1'b0 ;
  assign n23271 = n10104 & ~n23270 ;
  assign n23274 = n18151 ^ n13927 ^ n3434 ;
  assign n23272 = n2995 | n17602 ;
  assign n23273 = n7307 & n23272 ;
  assign n23275 = n23274 ^ n23273 ^ 1'b0 ;
  assign n23280 = n5905 | n7161 ;
  assign n23281 = n5129 & n23280 ;
  assign n23282 = n23281 ^ n1347 ^ 1'b0 ;
  assign n23276 = n3058 & ~n8690 ;
  assign n23277 = n553 | n23276 ;
  assign n23278 = n14769 & n23277 ;
  assign n23279 = ~n10218 & n23278 ;
  assign n23283 = n23282 ^ n23279 ^ 1'b0 ;
  assign n23284 = n6889 | n13896 ;
  assign n23285 = n10521 ^ n3530 ^ 1'b0 ;
  assign n23286 = n2141 & ~n23285 ;
  assign n23287 = n23286 ^ n17758 ^ 1'b0 ;
  assign n23291 = ~n3921 & n4030 ;
  assign n23292 = n23291 ^ n1209 ^ 1'b0 ;
  assign n23293 = n14583 | n23292 ;
  assign n23288 = n18839 ^ n12858 ^ 1'b0 ;
  assign n23289 = n4905 & n23288 ;
  assign n23290 = ~n21035 & n23289 ;
  assign n23294 = n23293 ^ n23290 ^ 1'b0 ;
  assign n23295 = n5315 & ~n23294 ;
  assign n23296 = ~n2202 & n4565 ;
  assign n23297 = ~n17424 & n23296 ;
  assign n23298 = n10234 & ~n23297 ;
  assign n23299 = n23298 ^ n14848 ^ 1'b0 ;
  assign n23300 = n17588 & ~n21461 ;
  assign n23301 = ~n15200 & n23300 ;
  assign n23302 = n3777 | n6645 ;
  assign n23303 = n18881 ^ n7230 ^ 1'b0 ;
  assign n23304 = ~n12405 & n16325 ;
  assign n23305 = ~n1570 & n9056 ;
  assign n23306 = n10826 & ~n23305 ;
  assign n23307 = n23306 ^ n8776 ^ 1'b0 ;
  assign n23308 = n11007 & ~n23307 ;
  assign n23309 = ~n3776 & n23308 ;
  assign n23310 = n2237 ^ n1483 ^ 1'b0 ;
  assign n23311 = ~n3160 & n23310 ;
  assign n23312 = n12515 & n21895 ;
  assign n23313 = ~n23311 & n23312 ;
  assign n23314 = ~n4590 & n8101 ;
  assign n23315 = n7783 & ~n14073 ;
  assign n23316 = n23315 ^ n6728 ^ 1'b0 ;
  assign n23317 = n8774 & n23316 ;
  assign n23318 = n23317 ^ n18337 ^ 1'b0 ;
  assign n23319 = ( n4184 & ~n5203 ) | ( n4184 & n23318 ) | ( ~n5203 & n23318 ) ;
  assign n23320 = n7399 | n8610 ;
  assign n23321 = n9139 ^ n1635 ^ 1'b0 ;
  assign n23322 = n13506 | n23321 ;
  assign n23323 = n23322 ^ n14675 ^ 1'b0 ;
  assign n23324 = n12074 ^ n11656 ^ 1'b0 ;
  assign n23325 = n16729 & ~n23324 ;
  assign n23326 = n23325 ^ n18780 ^ 1'b0 ;
  assign n23327 = ( n7530 & n10504 ) | ( n7530 & ~n23326 ) | ( n10504 & ~n23326 ) ;
  assign n23328 = ~n1703 & n15168 ;
  assign n23329 = n23328 ^ n4827 ^ 1'b0 ;
  assign n23330 = ~n790 & n14008 ;
  assign n23331 = n7777 & n23330 ;
  assign n23332 = n9913 ^ n6694 ^ 1'b0 ;
  assign n23333 = n11123 & n13090 ;
  assign n23334 = ~n23332 & n23333 ;
  assign n23335 = ~n1308 & n6386 ;
  assign n23336 = n2106 & n23335 ;
  assign n23337 = n23336 ^ n16110 ^ n7381 ;
  assign n23338 = n23337 ^ n13009 ^ n1091 ;
  assign n23339 = n23334 | n23338 ;
  assign n23340 = n9586 & ~n23339 ;
  assign n23343 = n3150 | n15051 ;
  assign n23341 = n2131 | n7686 ;
  assign n23342 = n7636 & ~n23341 ;
  assign n23344 = n23343 ^ n23342 ^ 1'b0 ;
  assign n23345 = n14719 & ~n22453 ;
  assign n23346 = ( n9675 & n11425 ) | ( n9675 & n12130 ) | ( n11425 & n12130 ) ;
  assign n23347 = n1856 | n10035 ;
  assign n23348 = n16505 ^ n4312 ^ n2488 ;
  assign n23349 = n12494 ^ n7007 ^ n5102 ;
  assign n23350 = ~n7871 & n23349 ;
  assign n23355 = n2206 & n5972 ;
  assign n23356 = ~n9638 & n23355 ;
  assign n23351 = n5244 & n19579 ;
  assign n23352 = n8370 & n23351 ;
  assign n23353 = n18475 & ~n23352 ;
  assign n23354 = ~n10600 & n23353 ;
  assign n23357 = n23356 ^ n23354 ^ 1'b0 ;
  assign n23358 = n7376 | n13708 ;
  assign n23359 = n11432 & ~n23358 ;
  assign n23360 = n4898 ^ n1314 ^ 1'b0 ;
  assign n23361 = n16464 ^ n5468 ^ 1'b0 ;
  assign n23362 = n23360 | n23361 ;
  assign n23366 = n1140 & n5154 ;
  assign n23364 = n1532 | n18622 ;
  assign n23365 = n9103 & ~n23364 ;
  assign n23367 = n23366 ^ n23365 ^ 1'b0 ;
  assign n23363 = n21067 ^ n7506 ^ 1'b0 ;
  assign n23368 = n23367 ^ n23363 ^ n4284 ;
  assign n23369 = n23362 & ~n23368 ;
  assign n23370 = n11490 | n12176 ;
  assign n23371 = n18643 & ~n23370 ;
  assign n23372 = n12923 ^ n3716 ^ 1'b0 ;
  assign n23373 = n12399 | n23372 ;
  assign n23374 = ( n6105 & n18357 ) | ( n6105 & n23373 ) | ( n18357 & n23373 ) ;
  assign n23375 = n10140 ^ n9559 ^ 1'b0 ;
  assign n23376 = n21079 & n23375 ;
  assign n23377 = x228 & n11408 ;
  assign n23378 = n23377 ^ n20509 ^ 1'b0 ;
  assign n23379 = n22210 ^ n21406 ^ 1'b0 ;
  assign n23380 = n1666 | n6844 ;
  assign n23381 = n4552 & n23380 ;
  assign n23382 = ~n16770 & n23381 ;
  assign n23383 = n9800 & ~n20778 ;
  assign n23384 = n1902 & n23383 ;
  assign n23385 = n2346 & ~n23384 ;
  assign n23386 = n9949 ^ n5632 ^ 1'b0 ;
  assign n23387 = n18561 ^ n12201 ^ 1'b0 ;
  assign n23389 = n418 | n3573 ;
  assign n23390 = n5980 | n23389 ;
  assign n23391 = n23390 ^ n5321 ^ 1'b0 ;
  assign n23388 = ~n2406 & n20603 ;
  assign n23392 = n23391 ^ n23388 ^ 1'b0 ;
  assign n23393 = n23392 ^ n18645 ^ 1'b0 ;
  assign n23394 = n10411 ^ n7199 ^ 1'b0 ;
  assign n23395 = n20958 | n23394 ;
  assign n23396 = n15956 ^ x140 ^ 1'b0 ;
  assign n23397 = n18156 | n18762 ;
  assign n23398 = n23396 & ~n23397 ;
  assign n23404 = n1340 & ~n4652 ;
  assign n23405 = n23404 ^ n1302 ^ 1'b0 ;
  assign n23406 = ( ~n2216 & n18381 ) | ( ~n2216 & n23405 ) | ( n18381 & n23405 ) ;
  assign n23407 = ~n11887 & n23406 ;
  assign n23401 = ~n7607 & n20795 ;
  assign n23399 = n12128 ^ n5975 ^ 1'b0 ;
  assign n23400 = n20054 & n23399 ;
  assign n23402 = n23401 ^ n23400 ^ n9546 ;
  assign n23403 = n23402 ^ n15440 ^ n10867 ;
  assign n23408 = n23407 ^ n23403 ^ 1'b0 ;
  assign n23409 = n9309 & ~n22476 ;
  assign n23410 = ~n23408 & n23409 ;
  assign n23411 = n6398 ^ n1177 ^ 1'b0 ;
  assign n23412 = n2969 | n5431 ;
  assign n23413 = n23412 ^ n13302 ^ n13044 ;
  assign n23414 = ~n3520 & n5958 ;
  assign n23415 = n6193 & ~n23414 ;
  assign n23416 = ( n9930 & n23413 ) | ( n9930 & ~n23415 ) | ( n23413 & ~n23415 ) ;
  assign n23417 = ( n1486 & n10378 ) | ( n1486 & ~n19249 ) | ( n10378 & ~n19249 ) ;
  assign n23418 = n666 & n6569 ;
  assign n23419 = n19638 & n23418 ;
  assign n23420 = ( n743 & n16862 ) | ( n743 & n23207 ) | ( n16862 & n23207 ) ;
  assign n23421 = n4140 | n6025 ;
  assign n23422 = n23421 ^ n972 ^ 1'b0 ;
  assign n23423 = n9133 & ~n18636 ;
  assign n23424 = n23422 & n23423 ;
  assign n23425 = n16439 | n21515 ;
  assign n23426 = n21082 & ~n23425 ;
  assign n23427 = ( n3218 & n5720 ) | ( n3218 & ~n23426 ) | ( n5720 & ~n23426 ) ;
  assign n23429 = ~n2727 & n3149 ;
  assign n23428 = n6373 ^ n2534 ^ 1'b0 ;
  assign n23430 = n23429 ^ n23428 ^ x118 ;
  assign n23431 = n1879 & ~n8207 ;
  assign n23432 = n23431 ^ n10525 ^ 1'b0 ;
  assign n23433 = n3289 & n23432 ;
  assign n23434 = ~n19178 & n23433 ;
  assign n23435 = n4792 & ~n9247 ;
  assign n23436 = n23435 ^ n3817 ^ 1'b0 ;
  assign n23437 = n365 | n8264 ;
  assign n23438 = n23437 ^ n20908 ^ 1'b0 ;
  assign n23439 = ( x7 & n23436 ) | ( x7 & n23438 ) | ( n23436 & n23438 ) ;
  assign n23440 = ( x2 & ~n4168 ) | ( x2 & n16885 ) | ( ~n4168 & n16885 ) ;
  assign n23441 = n23440 ^ n16757 ^ 1'b0 ;
  assign n23442 = n304 | n8919 ;
  assign n23443 = ~n2361 & n5479 ;
  assign n23444 = n23442 & n23443 ;
  assign n23445 = n8793 ^ n2276 ^ 1'b0 ;
  assign n23446 = n8947 & ~n23445 ;
  assign n23447 = ~n2649 & n11879 ;
  assign n23448 = ~n4136 & n21569 ;
  assign n23449 = n13549 ^ n2903 ^ 1'b0 ;
  assign n23450 = ~n10066 & n23449 ;
  assign n23451 = n14481 & ~n20026 ;
  assign n23452 = x41 & n1752 ;
  assign n23453 = n4652 | n23452 ;
  assign n23454 = n23453 ^ n7033 ^ 1'b0 ;
  assign n23455 = n2277 & ~n9735 ;
  assign n23456 = n23436 ^ n9663 ^ 1'b0 ;
  assign n23457 = n13956 & n21388 ;
  assign n23458 = n23457 ^ n11484 ^ 1'b0 ;
  assign n23461 = n2814 ^ n1103 ^ 1'b0 ;
  assign n23462 = n23461 ^ n18485 ^ 1'b0 ;
  assign n23460 = n13848 ^ n10117 ^ n2542 ;
  assign n23459 = n13732 & ~n17358 ;
  assign n23463 = n23462 ^ n23460 ^ n23459 ;
  assign n23464 = n2871 & n9403 ;
  assign n23465 = n23464 ^ n8235 ^ 1'b0 ;
  assign n23466 = ~n7063 & n23465 ;
  assign n23467 = n6553 & n23466 ;
  assign n23468 = n23463 & n23467 ;
  assign n23469 = n23468 ^ n3335 ^ 1'b0 ;
  assign n23470 = n18163 | n20987 ;
  assign n23471 = n23470 ^ n11628 ^ 1'b0 ;
  assign n23472 = n21270 ^ n8458 ^ 1'b0 ;
  assign n23473 = n1147 & n21869 ;
  assign n23474 = n23473 ^ n22516 ^ 1'b0 ;
  assign n23475 = n23474 ^ n20694 ^ 1'b0 ;
  assign n23476 = n9415 & ~n12184 ;
  assign n23477 = n23476 ^ n11548 ^ 1'b0 ;
  assign n23478 = n12145 ^ n1180 ^ 1'b0 ;
  assign n23479 = n22985 & ~n23478 ;
  assign n23480 = ~n9816 & n23479 ;
  assign n23481 = n23480 ^ n9428 ^ 1'b0 ;
  assign n23482 = n2078 & ~n23481 ;
  assign n23483 = n4792 & ~n20422 ;
  assign n23484 = n13738 ^ n5685 ^ 1'b0 ;
  assign n23485 = n4144 & ~n6792 ;
  assign n23486 = n23484 & n23485 ;
  assign n23487 = n13955 | n23486 ;
  assign n23496 = n14451 ^ n4846 ^ n2800 ;
  assign n23488 = n4395 & ~n4819 ;
  assign n23489 = n23488 ^ n8413 ^ n400 ;
  assign n23490 = n4168 & ~n23489 ;
  assign n23491 = n3140 ^ n1392 ^ 1'b0 ;
  assign n23492 = x176 & ~n23491 ;
  assign n23493 = n10763 ^ n5782 ^ 1'b0 ;
  assign n23494 = ( n19310 & ~n23492 ) | ( n19310 & n23493 ) | ( ~n23492 & n23493 ) ;
  assign n23495 = ( n2653 & ~n23490 ) | ( n2653 & n23494 ) | ( ~n23490 & n23494 ) ;
  assign n23497 = n23496 ^ n23495 ^ n486 ;
  assign n23498 = n5094 | n9200 ;
  assign n23499 = n4086 | n23498 ;
  assign n23500 = n22966 & ~n23499 ;
  assign n23501 = x171 & ~n23500 ;
  assign n23502 = n23501 ^ n3523 ^ 1'b0 ;
  assign n23503 = n23502 ^ n19097 ^ n15876 ;
  assign n23504 = ( n675 & ~n3543 ) | ( n675 & n3933 ) | ( ~n3543 & n3933 ) ;
  assign n23505 = n3338 & ~n6278 ;
  assign n23506 = n23505 ^ n1435 ^ 1'b0 ;
  assign n23507 = n21158 ^ n18050 ^ 1'b0 ;
  assign n23508 = n23506 | n23507 ;
  assign n23509 = n5767 ^ n4769 ^ 1'b0 ;
  assign n23512 = n1705 & ~n3898 ;
  assign n23510 = n16712 ^ n4373 ^ x132 ;
  assign n23511 = n23510 ^ n4139 ^ 1'b0 ;
  assign n23513 = n23512 ^ n23511 ^ n21452 ;
  assign n23514 = ( n4772 & n19083 ) | ( n4772 & ~n20878 ) | ( n19083 & ~n20878 ) ;
  assign n23515 = n23514 ^ n7942 ^ 1'b0 ;
  assign n23516 = n3714 & n13393 ;
  assign n23517 = ( ~n2483 & n9472 ) | ( ~n2483 & n23516 ) | ( n9472 & n23516 ) ;
  assign n23518 = n7943 & n9453 ;
  assign n23519 = n5045 | n15806 ;
  assign n23520 = n8716 | n23519 ;
  assign n23521 = n23520 ^ n428 ^ 1'b0 ;
  assign n23522 = n17032 & ~n23521 ;
  assign n23523 = n23518 & n23522 ;
  assign n23524 = n8516 & n23523 ;
  assign n23525 = n10469 ^ n8185 ^ 1'b0 ;
  assign n23526 = ~n4846 & n23525 ;
  assign n23527 = n5022 ^ n873 ^ 1'b0 ;
  assign n23528 = ~n8148 & n23527 ;
  assign n23529 = n23528 ^ n1863 ^ 1'b0 ;
  assign n23530 = n23529 ^ n13186 ^ n8120 ;
  assign n23531 = ( n12568 & ~n14274 ) | ( n12568 & n22983 ) | ( ~n14274 & n22983 ) ;
  assign n23532 = n300 & n10421 ;
  assign n23533 = ( n15353 & n16547 ) | ( n15353 & ~n23532 ) | ( n16547 & ~n23532 ) ;
  assign n23534 = n8276 ^ n2322 ^ 1'b0 ;
  assign n23535 = n14130 ^ n10059 ^ 1'b0 ;
  assign n23536 = ( ~n12417 & n17336 ) | ( ~n12417 & n23535 ) | ( n17336 & n23535 ) ;
  assign n23537 = ( x182 & ~n1486 ) | ( x182 & n21581 ) | ( ~n1486 & n21581 ) ;
  assign n23538 = n7475 ^ n2271 ^ 1'b0 ;
  assign n23539 = n2226 & n23538 ;
  assign n23540 = n5050 ^ n2103 ^ 1'b0 ;
  assign n23541 = n5370 | n23540 ;
  assign n23542 = n23541 ^ n16134 ^ 1'b0 ;
  assign n23543 = ~n14007 & n23542 ;
  assign n23544 = n13334 & ~n17493 ;
  assign n23545 = n23544 ^ n5508 ^ 1'b0 ;
  assign n23547 = n599 & ~n4290 ;
  assign n23546 = n23352 ^ n8398 ^ 1'b0 ;
  assign n23548 = n23547 ^ n23546 ^ 1'b0 ;
  assign n23549 = n10649 ^ n3951 ^ 1'b0 ;
  assign n23550 = n23548 | n23549 ;
  assign n23551 = n21977 ^ n18454 ^ 1'b0 ;
  assign n23552 = n7873 | n9557 ;
  assign n23553 = n23552 ^ n15564 ^ 1'b0 ;
  assign n23554 = n23551 & n23553 ;
  assign n23555 = n23554 ^ n22914 ^ n15351 ;
  assign n23556 = n18518 ^ n449 ^ 1'b0 ;
  assign n23557 = n729 | n14264 ;
  assign n23558 = ~n617 & n23557 ;
  assign n23559 = n8256 ^ n2291 ^ 1'b0 ;
  assign n23560 = n11226 & n23559 ;
  assign n23561 = n4073 & n23560 ;
  assign n23562 = n2109 | n5127 ;
  assign n23563 = n23562 ^ n9113 ^ n1302 ;
  assign n23564 = x229 & n4260 ;
  assign n23565 = n23564 ^ n14657 ^ n374 ;
  assign n23566 = n3375 | n23565 ;
  assign n23567 = n23566 ^ n8820 ^ 1'b0 ;
  assign n23568 = ~n3299 & n14511 ;
  assign n23569 = n22361 & ~n22941 ;
  assign n23570 = ~n23568 & n23569 ;
  assign n23571 = n6138 | n9320 ;
  assign n23572 = n15614 ^ n4286 ^ 1'b0 ;
  assign n23573 = ~n14805 & n22244 ;
  assign n23574 = n23573 ^ n18288 ^ n5824 ;
  assign n23575 = n23444 ^ n16823 ^ n10166 ;
  assign n23576 = n12674 & n20995 ;
  assign n23577 = ~n3542 & n13978 ;
  assign n23578 = n22674 ^ n8776 ^ 1'b0 ;
  assign n23579 = ~x114 & n23578 ;
  assign n23580 = n17016 ^ n15589 ^ 1'b0 ;
  assign n23581 = n23579 & n23580 ;
  assign n23583 = n3652 & n13837 ;
  assign n23582 = n8829 & ~n9613 ;
  assign n23584 = n23583 ^ n23582 ^ 1'b0 ;
  assign n23585 = n6312 & ~n9879 ;
  assign n23586 = n23585 ^ n7925 ^ 1'b0 ;
  assign n23587 = n14698 & n23586 ;
  assign n23588 = n1404 & n23587 ;
  assign n23589 = n2961 & n3088 ;
  assign n23590 = n23588 & n23589 ;
  assign n23591 = n2549 | n3588 ;
  assign n23594 = n3203 & ~n8170 ;
  assign n23595 = ~n22873 & n23594 ;
  assign n23592 = ~n2272 & n2998 ;
  assign n23593 = ~n6405 & n23592 ;
  assign n23596 = n23595 ^ n23593 ^ 1'b0 ;
  assign n23597 = n952 | n15541 ;
  assign n23598 = n18387 & ~n23597 ;
  assign n23599 = n11291 & ~n13508 ;
  assign n23600 = n20124 ^ n15881 ^ 1'b0 ;
  assign n23601 = n23600 ^ n15229 ^ 1'b0 ;
  assign n23602 = n1829 | n19400 ;
  assign n23603 = n23602 ^ n23411 ^ 1'b0 ;
  assign n23604 = n11568 & n19390 ;
  assign n23605 = n11696 ^ n993 ^ 1'b0 ;
  assign n23606 = n1786 & n23605 ;
  assign n23607 = x236 & ~n20755 ;
  assign n23608 = n23606 & n23607 ;
  assign n23609 = n21257 ^ n7482 ^ 1'b0 ;
  assign n23610 = n10752 ^ n7327 ^ 1'b0 ;
  assign n23616 = n8049 | n14648 ;
  assign n23617 = n1340 | n23616 ;
  assign n23618 = n23617 ^ n9750 ^ 1'b0 ;
  assign n23619 = n6470 | n23618 ;
  assign n23611 = n1935 & ~n5289 ;
  assign n23612 = n23611 ^ n8731 ^ 1'b0 ;
  assign n23613 = n17170 & n23612 ;
  assign n23614 = n23613 ^ n4560 ^ 1'b0 ;
  assign n23615 = n13704 & ~n23614 ;
  assign n23620 = n23619 ^ n23615 ^ 1'b0 ;
  assign n23621 = n531 & ~n1882 ;
  assign n23622 = ~n2800 & n11444 ;
  assign n23623 = n17459 & ~n23622 ;
  assign n23624 = n12937 ^ n10738 ^ 1'b0 ;
  assign n23625 = n23624 ^ n19845 ^ n4714 ;
  assign n23626 = n13781 ^ n12207 ^ n9520 ;
  assign n23627 = n23626 ^ n5230 ^ 1'b0 ;
  assign n23628 = ~n13585 & n23627 ;
  assign n23629 = n19033 ^ n9150 ^ 1'b0 ;
  assign n23630 = n8572 & n23629 ;
  assign n23631 = n4518 | n6172 ;
  assign n23632 = n23631 ^ n10181 ^ 1'b0 ;
  assign n23633 = n6421 ^ x161 ^ 1'b0 ;
  assign n23634 = n3678 | n23633 ;
  assign n23635 = n23632 & ~n23634 ;
  assign n23636 = ~n5327 & n14012 ;
  assign n23640 = n21431 ^ n7760 ^ 1'b0 ;
  assign n23637 = n7595 ^ n5331 ^ 1'b0 ;
  assign n23638 = n3279 & ~n23637 ;
  assign n23639 = ~n17712 & n23638 ;
  assign n23641 = n23640 ^ n23639 ^ 1'b0 ;
  assign n23642 = ( n5224 & n10168 ) | ( n5224 & n12712 ) | ( n10168 & n12712 ) ;
  assign n23644 = ( n4867 & ~n7083 ) | ( n4867 & n7869 ) | ( ~n7083 & n7869 ) ;
  assign n23643 = n880 | n1055 ;
  assign n23645 = n23644 ^ n23643 ^ 1'b0 ;
  assign n23646 = n23642 | n23645 ;
  assign n23647 = n4812 & n9121 ;
  assign n23648 = n1724 | n23647 ;
  assign n23649 = n23648 ^ n10624 ^ 1'b0 ;
  assign n23650 = ( n5327 & n17314 ) | ( n5327 & ~n21353 ) | ( n17314 & ~n21353 ) ;
  assign n23651 = n7500 | n11666 ;
  assign n23652 = n23651 ^ n1922 ^ 1'b0 ;
  assign n23653 = n2617 | n7764 ;
  assign n23654 = ~n10309 & n14041 ;
  assign n23655 = ~n23653 & n23654 ;
  assign n23656 = x62 & n5507 ;
  assign n23657 = ~n8055 & n20956 ;
  assign n23658 = ~n22881 & n23657 ;
  assign n23659 = n19325 & n23658 ;
  assign n23660 = n12612 ^ n1663 ^ 1'b0 ;
  assign n23661 = n6455 & n6854 ;
  assign n23662 = n23661 ^ n14367 ^ n3381 ;
  assign n23663 = n15924 & ~n23662 ;
  assign n23666 = n8565 ^ n5722 ^ 1'b0 ;
  assign n23667 = ~n21822 & n23666 ;
  assign n23664 = n7768 & ~n8470 ;
  assign n23665 = n23664 ^ n8737 ^ 1'b0 ;
  assign n23668 = n23667 ^ n23665 ^ n18990 ;
  assign n23669 = n5725 | n6537 ;
  assign n23670 = ~n10026 & n23669 ;
  assign n23671 = ~n13780 & n23166 ;
  assign n23672 = n23670 & n23671 ;
  assign n23673 = ~n15188 & n20553 ;
  assign n23674 = n23673 ^ n18258 ^ 1'b0 ;
  assign n23675 = n2514 | n15946 ;
  assign n23676 = n21621 & ~n23675 ;
  assign n23677 = n13811 ^ n10130 ^ n5304 ;
  assign n23678 = n9156 ^ n6992 ^ n6788 ;
  assign n23679 = ( n15182 & ~n23677 ) | ( n15182 & n23678 ) | ( ~n23677 & n23678 ) ;
  assign n23680 = n4450 ^ n2755 ^ 1'b0 ;
  assign n23681 = ~n12019 & n23680 ;
  assign n23682 = n593 | n17288 ;
  assign n23683 = n23681 | n23682 ;
  assign n23684 = n650 | n22207 ;
  assign n23685 = n18924 ^ n8944 ^ n4624 ;
  assign n23686 = n7453 & n17884 ;
  assign n23687 = ~n23685 & n23686 ;
  assign n23688 = n14396 ^ n6750 ^ n1978 ;
  assign n23689 = ~n11690 & n23688 ;
  assign n23690 = ( n8898 & ~n10326 ) | ( n8898 & n13837 ) | ( ~n10326 & n13837 ) ;
  assign n23691 = n2711 & ~n17795 ;
  assign n23692 = n23691 ^ n17250 ^ 1'b0 ;
  assign n23693 = n23690 | n23692 ;
  assign n23694 = n18317 ^ n11400 ^ 1'b0 ;
  assign n23695 = n3171 | n10055 ;
  assign n23696 = n23695 ^ n2243 ^ 1'b0 ;
  assign n23697 = n3625 & ~n15153 ;
  assign n23698 = n1645 | n11291 ;
  assign n23699 = ( n6623 & ~n8884 ) | ( n6623 & n10621 ) | ( ~n8884 & n10621 ) ;
  assign n23703 = n3939 ^ x161 ^ 1'b0 ;
  assign n23704 = n6970 & ~n23703 ;
  assign n23700 = n14310 ^ n8783 ^ 1'b0 ;
  assign n23701 = n15642 | n23700 ;
  assign n23702 = n21268 & ~n23701 ;
  assign n23705 = n23704 ^ n23702 ^ 1'b0 ;
  assign n23706 = n23699 & ~n23705 ;
  assign n23707 = ~n23698 & n23706 ;
  assign n23708 = n23707 ^ n17921 ^ 1'b0 ;
  assign n23709 = x132 & n4606 ;
  assign n23710 = ~n6085 & n23709 ;
  assign n23711 = n23710 ^ n1230 ^ 1'b0 ;
  assign n23712 = n11488 & ~n23711 ;
  assign n23713 = n410 | n4440 ;
  assign n23714 = n15020 ^ n1671 ^ n553 ;
  assign n23715 = ~n7809 & n23714 ;
  assign n23716 = ~n13889 & n23715 ;
  assign n23717 = ( n7476 & ~n8106 ) | ( n7476 & n23716 ) | ( ~n8106 & n23716 ) ;
  assign n23718 = n1098 | n2174 ;
  assign n23719 = n1098 & ~n23718 ;
  assign n23720 = n7052 & ~n23719 ;
  assign n23721 = ~n7052 & n23720 ;
  assign n23722 = n1569 & ~n23721 ;
  assign n23723 = n23721 & n23722 ;
  assign n23724 = n8783 | n23723 ;
  assign n23725 = n1010 & ~n3501 ;
  assign n23726 = ~n1010 & n23725 ;
  assign n23727 = ~n4945 & n6921 ;
  assign n23728 = ~n6921 & n23727 ;
  assign n23729 = n23726 | n23728 ;
  assign n23730 = n23724 | n23729 ;
  assign n23731 = n1058 | n7866 ;
  assign n23732 = n10881 & ~n23731 ;
  assign n23733 = n23732 ^ n1702 ^ 1'b0 ;
  assign n23735 = n6510 & ~n13870 ;
  assign n23736 = n23735 ^ n11854 ^ 1'b0 ;
  assign n23734 = n13634 & n14988 ;
  assign n23737 = n23736 ^ n23734 ^ 1'b0 ;
  assign n23738 = n3958 & n18922 ;
  assign n23739 = n495 & ~n5581 ;
  assign n23740 = n8550 ^ x139 ^ 1'b0 ;
  assign n23741 = n23739 | n23740 ;
  assign n23742 = n4759 | n23741 ;
  assign n23743 = n4759 & ~n23742 ;
  assign n23745 = ~n3175 & n12908 ;
  assign n23746 = n23745 ^ n3272 ^ 1'b0 ;
  assign n23744 = ~n2649 & n19286 ;
  assign n23747 = n23746 ^ n23744 ^ 1'b0 ;
  assign n23748 = n23747 ^ n5997 ^ 1'b0 ;
  assign n23749 = ( n14955 & n18707 ) | ( n14955 & ~n23748 ) | ( n18707 & ~n23748 ) ;
  assign n23750 = n8852 ^ n8220 ^ 1'b0 ;
  assign n23751 = ~n1811 & n23750 ;
  assign n23752 = ~n8618 & n23751 ;
  assign n23753 = n2389 | n21621 ;
  assign n23754 = n23753 ^ n17430 ^ 1'b0 ;
  assign n23755 = n10186 ^ n6134 ^ 1'b0 ;
  assign n23756 = x46 | n4026 ;
  assign n23757 = n12713 & ~n23756 ;
  assign n23758 = n23755 & n23757 ;
  assign n23759 = n19411 ^ n2014 ^ 1'b0 ;
  assign n23760 = ( n11302 & ~n11857 ) | ( n11302 & n12527 ) | ( ~n11857 & n12527 ) ;
  assign n23761 = ~n13167 & n23760 ;
  assign n23762 = n16758 ^ n5639 ^ 1'b0 ;
  assign n23763 = n15159 & n23762 ;
  assign n23766 = n2726 & n7137 ;
  assign n23767 = n23766 ^ n2818 ^ 1'b0 ;
  assign n23764 = n10637 & ~n12133 ;
  assign n23765 = n16727 | n23764 ;
  assign n23768 = n23767 ^ n23765 ^ 1'b0 ;
  assign n23769 = n5266 | n7831 ;
  assign n23770 = n2882 | n23769 ;
  assign n23771 = n2463 | n23770 ;
  assign n23773 = n1025 & n20984 ;
  assign n23772 = ~n1353 & n4284 ;
  assign n23774 = n23773 ^ n23772 ^ 1'b0 ;
  assign n23775 = n3675 | n11349 ;
  assign n23776 = n6146 | n23775 ;
  assign n23777 = n23776 ^ n6177 ^ 1'b0 ;
  assign n23780 = n3236 ^ n3121 ^ 1'b0 ;
  assign n23781 = n7321 & n23780 ;
  assign n23782 = n23781 ^ n2756 ^ 1'b0 ;
  assign n23778 = n12399 | n13902 ;
  assign n23779 = n23778 ^ n13759 ^ 1'b0 ;
  assign n23783 = n23782 ^ n23779 ^ n5034 ;
  assign n23784 = ~n15572 & n16413 ;
  assign n23785 = n9588 ^ n1988 ^ 1'b0 ;
  assign n23786 = n3597 & ~n23785 ;
  assign n23787 = n23784 & n23786 ;
  assign n23788 = n3756 & n5958 ;
  assign n23789 = n9895 & n23788 ;
  assign n23790 = n13722 & n23789 ;
  assign n23791 = n4235 & ~n11421 ;
  assign n23792 = ~n9331 & n23791 ;
  assign n23793 = n5238 & n16933 ;
  assign n23794 = n19800 & ~n23793 ;
  assign n23795 = n20720 ^ n15343 ^ 1'b0 ;
  assign n23796 = n392 & n23795 ;
  assign n23797 = n20870 ^ n11375 ^ 1'b0 ;
  assign n23798 = n601 | n8134 ;
  assign n23799 = n21931 & n23798 ;
  assign n23800 = n23799 ^ n22140 ^ 1'b0 ;
  assign n23801 = n23700 ^ n21746 ^ 1'b0 ;
  assign n23802 = n6081 & ~n23801 ;
  assign n23803 = n18734 & n23802 ;
  assign n23804 = n4571 & ~n9914 ;
  assign n23805 = ~x14 & n23804 ;
  assign n23806 = n11884 ^ n4774 ^ 1'b0 ;
  assign n23807 = n23805 | n23806 ;
  assign n23808 = n11918 ^ n6696 ^ 1'b0 ;
  assign n23809 = n4284 & ~n23808 ;
  assign n23810 = n5773 & n7473 ;
  assign n23811 = n8093 ^ n4196 ^ 1'b0 ;
  assign n23812 = n4245 & n23811 ;
  assign n23813 = n2203 | n5857 ;
  assign n23814 = n23813 ^ n3169 ^ 1'b0 ;
  assign n23815 = ( ~n22261 & n23812 ) | ( ~n22261 & n23814 ) | ( n23812 & n23814 ) ;
  assign n23816 = n13135 ^ n6047 ^ 1'b0 ;
  assign n23817 = n20622 & ~n23816 ;
  assign n23818 = ( ~x119 & n867 ) | ( ~x119 & n7253 ) | ( n867 & n7253 ) ;
  assign n23819 = n19734 ^ n13280 ^ 1'b0 ;
  assign n23820 = n2181 & n3891 ;
  assign n23822 = n5037 ^ x28 ^ 1'b0 ;
  assign n23821 = n1307 & ~n12184 ;
  assign n23823 = n23822 ^ n23821 ^ 1'b0 ;
  assign n23825 = n444 | n6409 ;
  assign n23826 = n23825 ^ n9562 ^ 1'b0 ;
  assign n23824 = n15455 | n21230 ;
  assign n23827 = n23826 ^ n23824 ^ 1'b0 ;
  assign n23828 = ~x109 & n1275 ;
  assign n23829 = n3901 | n23828 ;
  assign n23830 = ( n11131 & n17532 ) | ( n11131 & n23829 ) | ( n17532 & n23829 ) ;
  assign n23831 = ~n5812 & n20572 ;
  assign n23832 = n15409 & n23831 ;
  assign n23833 = n6758 & n8085 ;
  assign n23834 = n23833 ^ n11272 ^ 1'b0 ;
  assign n23835 = n17085 & n23834 ;
  assign n23836 = n23835 ^ n10194 ^ 1'b0 ;
  assign n23837 = n514 | n16823 ;
  assign n23838 = n5519 & ~n23837 ;
  assign n23839 = ( ~n2462 & n13990 ) | ( ~n2462 & n22163 ) | ( n13990 & n22163 ) ;
  assign n23840 = n17042 ^ n14928 ^ 1'b0 ;
  assign n23841 = ~n605 & n23590 ;
  assign n23842 = ~n15933 & n21486 ;
  assign n23843 = ~n14102 & n23842 ;
  assign n23844 = ~n5163 & n12970 ;
  assign n23845 = ~n1177 & n17182 ;
  assign n23846 = n1328 & n23845 ;
  assign n23847 = n19011 ^ n4821 ^ 1'b0 ;
  assign n23848 = n23041 ^ n460 ^ 1'b0 ;
  assign n23849 = ~n21761 & n23848 ;
  assign n23850 = n15983 ^ n1259 ^ 1'b0 ;
  assign n23851 = n6591 | n13246 ;
  assign n23852 = n8541 & n23851 ;
  assign n23853 = n23852 ^ n19694 ^ 1'b0 ;
  assign n23854 = n9976 & n10563 ;
  assign n23856 = ~n6572 & n7306 ;
  assign n23857 = ~x244 & n23856 ;
  assign n23855 = n20755 ^ n646 ^ 1'b0 ;
  assign n23858 = n23857 ^ n23855 ^ n18864 ;
  assign n23859 = n5375 | n6460 ;
  assign n23860 = n23859 ^ n1912 ^ 1'b0 ;
  assign n23861 = ~n8220 & n23860 ;
  assign n23862 = n23861 ^ n8912 ^ 1'b0 ;
  assign n23863 = n17066 & ~n20883 ;
  assign n23864 = n23863 ^ n4489 ^ 1'b0 ;
  assign n23865 = n18620 ^ n10813 ^ n8270 ;
  assign n23866 = n23865 ^ n11375 ^ n6127 ;
  assign n23867 = n1775 & n23866 ;
  assign n23868 = ~n5637 & n23867 ;
  assign n23869 = n1641 ^ n1293 ^ 1'b0 ;
  assign n23870 = n9314 | n13977 ;
  assign n23871 = n23869 | n23870 ;
  assign n23872 = n2156 | n8101 ;
  assign n23873 = n23872 ^ n5596 ^ n5347 ;
  assign n23874 = n12685 ^ n7392 ^ n6009 ;
  assign n23875 = ( n2561 & n9035 ) | ( n2561 & n21284 ) | ( n9035 & n21284 ) ;
  assign n23876 = n10117 & n23875 ;
  assign n23877 = n23876 ^ n4435 ^ 1'b0 ;
  assign n23878 = ~n535 & n23877 ;
  assign n23879 = n23878 ^ n5172 ^ 1'b0 ;
  assign n23880 = ~n3570 & n3769 ;
  assign n23881 = n3833 | n20089 ;
  assign n23882 = n23880 & ~n23881 ;
  assign n23883 = ~n4580 & n11222 ;
  assign n23884 = n23883 ^ n9165 ^ n6001 ;
  assign n23886 = n3047 & n12008 ;
  assign n23885 = n269 & n14935 ;
  assign n23887 = n23886 ^ n23885 ^ n13990 ;
  assign n23888 = n3278 & ~n5321 ;
  assign n23889 = n23888 ^ n7466 ^ 1'b0 ;
  assign n23892 = n11087 ^ n7356 ^ n693 ;
  assign n23893 = n23892 ^ n22194 ^ 1'b0 ;
  assign n23894 = n9932 | n23893 ;
  assign n23890 = x236 | n16221 ;
  assign n23891 = n3973 | n23890 ;
  assign n23895 = n23894 ^ n23891 ^ 1'b0 ;
  assign n23896 = ~n1777 & n5907 ;
  assign n23897 = n10671 ^ n6323 ^ 1'b0 ;
  assign n23898 = ~n19518 & n23897 ;
  assign n23899 = n23896 & ~n23898 ;
  assign n23900 = n13896 ^ n7697 ^ 1'b0 ;
  assign n23901 = n4026 ^ n1406 ^ 1'b0 ;
  assign n23902 = n23901 ^ n12208 ^ n3809 ;
  assign n23903 = n1082 | n23902 ;
  assign n23904 = n23903 ^ n14374 ^ 1'b0 ;
  assign n23905 = n3658 | n10966 ;
  assign n23906 = n22998 ^ n4575 ^ 1'b0 ;
  assign n23907 = n18131 ^ n6808 ^ 1'b0 ;
  assign n23908 = n16540 ^ n15236 ^ 1'b0 ;
  assign n23909 = n20440 & n23908 ;
  assign n23910 = n8310 & n16712 ;
  assign n23911 = ~n8310 & n23910 ;
  assign n23912 = n2026 ^ n942 ^ 1'b0 ;
  assign n23913 = n23912 ^ n785 ^ 1'b0 ;
  assign n23914 = ~n17967 & n23913 ;
  assign n23915 = ( n1667 & n4456 ) | ( n1667 & n9699 ) | ( n4456 & n9699 ) ;
  assign n23916 = ( ~n5038 & n11464 ) | ( ~n5038 & n23915 ) | ( n11464 & n23915 ) ;
  assign n23917 = n8310 & ~n19089 ;
  assign n23918 = n23917 ^ n9824 ^ 1'b0 ;
  assign n23920 = n17524 ^ n5666 ^ 1'b0 ;
  assign n23919 = n1432 & n21392 ;
  assign n23921 = n23920 ^ n23919 ^ 1'b0 ;
  assign n23922 = ( ~n2098 & n2781 ) | ( ~n2098 & n10455 ) | ( n2781 & n10455 ) ;
  assign n23923 = n23922 ^ n19205 ^ n7672 ;
  assign n23924 = n15633 ^ n2224 ^ n1496 ;
  assign n23925 = n4525 | n10464 ;
  assign n23926 = n6729 & ~n23925 ;
  assign n23927 = n3533 & ~n23926 ;
  assign n23928 = ~n12495 & n23927 ;
  assign n23929 = n15983 ^ x192 ^ 1'b0 ;
  assign n23930 = n23928 | n23929 ;
  assign n23931 = n8411 & ~n16490 ;
  assign n23932 = ~n18974 & n23931 ;
  assign n23933 = n18348 & ~n23932 ;
  assign n23934 = n23733 & ~n23933 ;
  assign n23935 = n14245 ^ n1179 ^ 1'b0 ;
  assign n23936 = n21592 ^ n9559 ^ 1'b0 ;
  assign n23937 = ( n4511 & n12810 ) | ( n4511 & n23936 ) | ( n12810 & n23936 ) ;
  assign n23938 = ~n2613 & n23937 ;
  assign n23939 = x157 & ~n6349 ;
  assign n23940 = ~n1311 & n23939 ;
  assign n23941 = ~n23603 & n23940 ;
  assign n23942 = n273 & ~n8029 ;
  assign n23943 = n23942 ^ n14387 ^ n3749 ;
  assign n23944 = n10982 & ~n20496 ;
  assign n23945 = n23944 ^ n9656 ^ n6027 ;
  assign n23948 = n15869 | n18124 ;
  assign n23947 = n6220 & n15197 ;
  assign n23946 = n3384 & n12798 ;
  assign n23949 = n23948 ^ n23947 ^ n23946 ;
  assign n23950 = n10023 | n23949 ;
  assign n23951 = n3409 & ~n23950 ;
  assign n23952 = ~n2885 & n17371 ;
  assign n23953 = ~n9697 & n23952 ;
  assign n23954 = n10903 ^ n5173 ^ 1'b0 ;
  assign n23955 = n23954 ^ n13309 ^ 1'b0 ;
  assign n23956 = n5634 | n23955 ;
  assign n23957 = n4618 & n5053 ;
  assign n23958 = x159 & n5650 ;
  assign n23959 = ~n23592 & n23958 ;
  assign n23960 = ~n21713 & n23959 ;
  assign n23961 = ~n2008 & n11328 ;
  assign n23962 = n23961 ^ n11882 ^ 1'b0 ;
  assign n23963 = n11287 & ~n23962 ;
  assign n23964 = n23960 & n23963 ;
  assign n23965 = ( x5 & ~n1669 ) | ( x5 & n2831 ) | ( ~n1669 & n2831 ) ;
  assign n23972 = ( n2392 & ~n3504 ) | ( n2392 & n12916 ) | ( ~n3504 & n12916 ) ;
  assign n23973 = n13140 | n13174 ;
  assign n23974 = n23972 & ~n23973 ;
  assign n23966 = n18791 ^ n16816 ^ 1'b0 ;
  assign n23967 = n1525 & ~n3958 ;
  assign n23968 = n23967 ^ n1406 ^ 1'b0 ;
  assign n23969 = n23968 ^ n10766 ^ 1'b0 ;
  assign n23970 = ( n6253 & n16550 ) | ( n6253 & ~n23969 ) | ( n16550 & ~n23969 ) ;
  assign n23971 = n23966 & ~n23970 ;
  assign n23975 = n23974 ^ n23971 ^ n14926 ;
  assign n23976 = n2829 & n7971 ;
  assign n23977 = ~n15637 & n23976 ;
  assign n23978 = ( n14256 & n19026 ) | ( n14256 & ~n23428 ) | ( n19026 & ~n23428 ) ;
  assign n23979 = n14078 | n23978 ;
  assign n23980 = n18536 ^ n17595 ^ n3880 ;
  assign n23981 = n1899 & ~n10447 ;
  assign n23982 = n1887 & n21358 ;
  assign n23983 = n11504 & n23982 ;
  assign n23984 = n23983 ^ n17272 ^ 1'b0 ;
  assign n23985 = ~n23981 & n23984 ;
  assign n23986 = ( ~n2228 & n6849 ) | ( ~n2228 & n8427 ) | ( n6849 & n8427 ) ;
  assign n23987 = n19623 ^ n1023 ^ 1'b0 ;
  assign n23988 = n15575 & ~n23987 ;
  assign n23989 = n23988 ^ n4757 ^ 1'b0 ;
  assign n23990 = n15221 ^ n5864 ^ 1'b0 ;
  assign n23991 = n2048 & ~n23990 ;
  assign n23992 = n23991 ^ n5375 ^ 1'b0 ;
  assign n23993 = x11 & n1129 ;
  assign n23994 = n11694 & n23993 ;
  assign n23995 = n23994 ^ n21945 ^ 1'b0 ;
  assign n23996 = n622 & n3533 ;
  assign n23997 = n23996 ^ n6927 ^ 1'b0 ;
  assign n23998 = n2360 & n5722 ;
  assign n23999 = n23998 ^ n516 ^ 1'b0 ;
  assign n24000 = n18299 | n23999 ;
  assign n24001 = n9077 ^ n7190 ^ 1'b0 ;
  assign n24002 = n24001 ^ n21139 ^ n14036 ;
  assign n24003 = n8167 & n18378 ;
  assign n24004 = ~n2698 & n13945 ;
  assign n24005 = ~n13928 & n20945 ;
  assign n24006 = n13013 ^ n12978 ^ 1'b0 ;
  assign n24007 = n12002 & ~n24006 ;
  assign n24008 = ~n4340 & n24007 ;
  assign n24009 = n24008 ^ n17523 ^ 1'b0 ;
  assign n24010 = n24009 ^ n10589 ^ 1'b0 ;
  assign n24011 = ( n11072 & n14796 ) | ( n11072 & n18973 ) | ( n14796 & n18973 ) ;
  assign n24012 = ~n10525 & n12237 ;
  assign n24013 = n15093 & n24012 ;
  assign n24014 = n2611 & n20726 ;
  assign n24015 = n4094 & n24014 ;
  assign n24016 = ~n1380 & n16851 ;
  assign n24018 = n6206 & n13391 ;
  assign n24017 = ~n10244 & n18715 ;
  assign n24019 = n24018 ^ n24017 ^ 1'b0 ;
  assign n24020 = n5538 & n24019 ;
  assign n24021 = n1471 & n10790 ;
  assign n24022 = ~n10213 & n24021 ;
  assign n24023 = ( n1742 & ~n17342 ) | ( n1742 & n24022 ) | ( ~n17342 & n24022 ) ;
  assign n24024 = ~n1213 & n22033 ;
  assign n24025 = n18616 ^ n7149 ^ 1'b0 ;
  assign n24026 = n24024 | n24025 ;
  assign n24027 = ~n407 & n7454 ;
  assign n24028 = n6790 ^ n1517 ^ 1'b0 ;
  assign n24029 = n24028 ^ n14815 ^ n7567 ;
  assign n24030 = n2524 ^ n2186 ^ 1'b0 ;
  assign n24031 = ( n1598 & n14246 ) | ( n1598 & n24030 ) | ( n14246 & n24030 ) ;
  assign n24032 = n6330 ^ n5408 ^ 1'b0 ;
  assign n24033 = ( n14219 & n24031 ) | ( n14219 & n24032 ) | ( n24031 & n24032 ) ;
  assign n24034 = n5541 & ~n21326 ;
  assign n24035 = n397 | n4642 ;
  assign n24036 = n24035 ^ n23317 ^ 1'b0 ;
  assign n24041 = n7157 ^ n5790 ^ 1'b0 ;
  assign n24042 = n3825 & ~n24041 ;
  assign n24040 = ~n2061 & n4279 ;
  assign n24043 = n24042 ^ n24040 ^ 1'b0 ;
  assign n24039 = ( n4104 & n8848 ) | ( n4104 & ~n9263 ) | ( n8848 & ~n9263 ) ;
  assign n24037 = n11212 ^ n543 ^ 1'b0 ;
  assign n24038 = n14017 & ~n24037 ;
  assign n24044 = n24043 ^ n24039 ^ n24038 ;
  assign n24045 = n23518 ^ n11672 ^ 1'b0 ;
  assign n24046 = n8197 & ~n24045 ;
  assign n24047 = n24046 ^ n15937 ^ n6409 ;
  assign n24048 = ( n9941 & ~n10490 ) | ( n9941 & n11665 ) | ( ~n10490 & n11665 ) ;
  assign n24049 = ( n2774 & n10963 ) | ( n2774 & n24048 ) | ( n10963 & n24048 ) ;
  assign n24050 = x165 | n24049 ;
  assign n24051 = ~n9180 & n20777 ;
  assign n24052 = n20536 & n24051 ;
  assign n24053 = n17420 | n24052 ;
  assign n24054 = n24053 ^ n10614 ^ 1'b0 ;
  assign n24055 = n16405 ^ n3815 ^ 1'b0 ;
  assign n24056 = n24054 & ~n24055 ;
  assign n24057 = n4699 & n24056 ;
  assign n24058 = n16502 | n23440 ;
  assign n24059 = ( n4080 & n12310 ) | ( n4080 & n24058 ) | ( n12310 & n24058 ) ;
  assign n24060 = ( n4153 & ~n7615 ) | ( n4153 & n20285 ) | ( ~n7615 & n20285 ) ;
  assign n24061 = n24060 ^ n4330 ^ 1'b0 ;
  assign n24062 = n6600 ^ n2454 ^ 1'b0 ;
  assign n24063 = n19380 & ~n24062 ;
  assign n24064 = n24063 ^ n10326 ^ 1'b0 ;
  assign n24065 = ~n20043 & n24064 ;
  assign n24066 = n4247 & ~n15049 ;
  assign n24067 = ( n15656 & n21494 ) | ( n15656 & ~n24066 ) | ( n21494 & ~n24066 ) ;
  assign n24068 = n13063 ^ n7867 ^ 1'b0 ;
  assign n24069 = n24067 | n24068 ;
  assign n24070 = n4931 & n17708 ;
  assign n24071 = n4595 & ~n16203 ;
  assign n24072 = n7844 & n24071 ;
  assign n24073 = n7700 & n24072 ;
  assign n24075 = n3508 & n20987 ;
  assign n24076 = n10688 & n24075 ;
  assign n24074 = n294 & n9196 ;
  assign n24077 = n24076 ^ n24074 ^ 1'b0 ;
  assign n24078 = n9369 & ~n16384 ;
  assign n24079 = n24078 ^ n17259 ^ 1'b0 ;
  assign n24085 = n1801 | n3043 ;
  assign n24080 = n6606 | n20055 ;
  assign n24081 = n24080 ^ n18725 ^ n887 ;
  assign n24082 = n24081 ^ n7473 ^ 1'b0 ;
  assign n24083 = n9298 & ~n24082 ;
  assign n24084 = n24083 ^ n16619 ^ n1228 ;
  assign n24086 = n24085 ^ n24084 ^ 1'b0 ;
  assign n24087 = n6350 | n24086 ;
  assign n24088 = n24079 & ~n24087 ;
  assign n24089 = n12359 & n24088 ;
  assign n24090 = n10144 | n24089 ;
  assign n24091 = n2192 | n5114 ;
  assign n24092 = n24091 ^ n2127 ^ 1'b0 ;
  assign n24093 = n24092 ^ n17288 ^ 1'b0 ;
  assign n24094 = n4376 & n12897 ;
  assign n24095 = n24094 ^ n11421 ^ 1'b0 ;
  assign n24096 = ~n8022 & n16375 ;
  assign n24097 = n24096 ^ n8977 ^ 1'b0 ;
  assign n24098 = n24097 ^ n9489 ^ 1'b0 ;
  assign n24099 = ( n15901 & ~n24095 ) | ( n15901 & n24098 ) | ( ~n24095 & n24098 ) ;
  assign n24100 = n2443 & n7743 ;
  assign n24101 = n24100 ^ n14080 ^ 1'b0 ;
  assign n24102 = ( n6151 & n23901 ) | ( n6151 & n24101 ) | ( n23901 & n24101 ) ;
  assign n24103 = n17731 & ~n24102 ;
  assign n24104 = n24103 ^ n2577 ^ 1'b0 ;
  assign n24105 = n2095 | n6953 ;
  assign n24106 = n14417 ^ n8425 ^ 1'b0 ;
  assign n24107 = n7554 & ~n24106 ;
  assign n24108 = n18047 ^ n5522 ^ 1'b0 ;
  assign n24109 = n966 | n21272 ;
  assign n24110 = n698 | n5334 ;
  assign n24111 = n2755 | n24110 ;
  assign n24112 = n24111 ^ n20485 ^ 1'b0 ;
  assign n24113 = n1872 & n4045 ;
  assign n24114 = n24113 ^ n3895 ^ 1'b0 ;
  assign n24115 = n24114 ^ n11039 ^ n8425 ;
  assign n24116 = n277 & n15141 ;
  assign n24117 = n4832 | n24116 ;
  assign n24118 = n3652 & n8071 ;
  assign n24119 = n7338 & n24118 ;
  assign n24120 = n8441 ^ n4744 ^ 1'b0 ;
  assign n24121 = n14595 ^ n6259 ^ 1'b0 ;
  assign n24122 = ( ~n24119 & n24120 ) | ( ~n24119 & n24121 ) | ( n24120 & n24121 ) ;
  assign n24123 = n17900 ^ n8261 ^ n7571 ;
  assign n24124 = n4732 ^ n4363 ^ 1'b0 ;
  assign n24125 = ~n707 & n24124 ;
  assign n24126 = ( n2124 & n9403 ) | ( n2124 & n18070 ) | ( n9403 & n18070 ) ;
  assign n24127 = ( n919 & n15601 ) | ( n919 & n24126 ) | ( n15601 & n24126 ) ;
  assign n24128 = x178 | n5962 ;
  assign n24129 = n13580 ^ n7448 ^ n1833 ;
  assign n24130 = n24128 & ~n24129 ;
  assign n24131 = n24130 ^ n4738 ^ 1'b0 ;
  assign n24132 = n21172 & ~n24131 ;
  assign n24133 = ( ~x152 & n1336 ) | ( ~x152 & n1372 ) | ( n1336 & n1372 ) ;
  assign n24136 = n2991 | n5423 ;
  assign n24137 = n9236 | n24136 ;
  assign n24134 = n5773 & ~n20997 ;
  assign n24135 = n937 & n24134 ;
  assign n24138 = n24137 ^ n24135 ^ 1'b0 ;
  assign n24139 = n327 & n5676 ;
  assign n24140 = n2214 | n8906 ;
  assign n24141 = n24140 ^ n21930 ^ 1'b0 ;
  assign n24142 = n6371 | n8665 ;
  assign n24143 = n16684 ^ n16507 ^ n16390 ;
  assign n24144 = n11763 & ~n24143 ;
  assign n24145 = n21229 ^ n7369 ^ 1'b0 ;
  assign n24146 = n24145 ^ n8662 ^ 1'b0 ;
  assign n24147 = ( n3000 & ~n5328 ) | ( n3000 & n10359 ) | ( ~n5328 & n10359 ) ;
  assign n24148 = n12837 & n24147 ;
  assign n24149 = ( n14571 & n23142 ) | ( n14571 & ~n24148 ) | ( n23142 & ~n24148 ) ;
  assign n24151 = n20480 ^ n6641 ^ 1'b0 ;
  assign n24150 = n8171 & ~n10639 ;
  assign n24152 = n24151 ^ n24150 ^ 1'b0 ;
  assign n24153 = n8740 & ~n24152 ;
  assign n24154 = ~n1894 & n24153 ;
  assign n24155 = n1005 & n24154 ;
  assign n24156 = n4409 ^ n1254 ^ 1'b0 ;
  assign n24157 = ~n16194 & n24156 ;
  assign n24158 = n8747 & n24157 ;
  assign n24159 = ~n24155 & n24158 ;
  assign n24160 = n10172 ^ n8137 ^ 1'b0 ;
  assign n24161 = n16094 ^ n7604 ^ 1'b0 ;
  assign n24162 = n16255 ^ n13780 ^ 1'b0 ;
  assign n24163 = ~n420 & n24162 ;
  assign n24164 = ~n10145 & n19572 ;
  assign n24165 = n14719 ^ n2041 ^ 1'b0 ;
  assign n24166 = n15496 | n24165 ;
  assign n24167 = n24166 ^ n15957 ^ 1'b0 ;
  assign n24168 = n15365 ^ n8250 ^ 1'b0 ;
  assign n24169 = n13608 ^ n3222 ^ 1'b0 ;
  assign n24170 = n2102 & n24169 ;
  assign n24171 = n24170 ^ n8174 ^ 1'b0 ;
  assign n24172 = n13122 & ~n14242 ;
  assign n24173 = n24172 ^ n5988 ^ 1'b0 ;
  assign n24174 = ( n7015 & ~n8394 ) | ( n7015 & n16163 ) | ( ~n8394 & n16163 ) ;
  assign n24175 = ( ~x71 & n16595 ) | ( ~x71 & n24174 ) | ( n16595 & n24174 ) ;
  assign n24176 = n1886 & ~n18371 ;
  assign n24177 = n14051 ^ n13606 ^ 1'b0 ;
  assign n24178 = n24177 ^ n6188 ^ 1'b0 ;
  assign n24179 = ( ~n24120 & n24176 ) | ( ~n24120 & n24178 ) | ( n24176 & n24178 ) ;
  assign n24180 = n12910 ^ n12202 ^ 1'b0 ;
  assign n24181 = n12780 & ~n24180 ;
  assign n24182 = n24181 ^ n10876 ^ x24 ;
  assign n24183 = n2836 & n3883 ;
  assign n24184 = n24183 ^ x254 ^ 1'b0 ;
  assign n24185 = n8233 & n24184 ;
  assign n24186 = n11074 & n24185 ;
  assign n24187 = n23885 & n24186 ;
  assign n24188 = n23420 ^ n1998 ^ 1'b0 ;
  assign n24189 = n11122 & ~n17343 ;
  assign n24190 = n18874 & n24189 ;
  assign n24191 = ( n7538 & n12947 ) | ( n7538 & ~n14909 ) | ( n12947 & ~n14909 ) ;
  assign n24192 = n8026 & ~n24191 ;
  assign n24193 = n24192 ^ n20260 ^ 1'b0 ;
  assign n24194 = n1038 | n24193 ;
  assign n24195 = n24194 ^ n17982 ^ 1'b0 ;
  assign n24196 = n429 | n4169 ;
  assign n24197 = n6029 ^ n2051 ^ 1'b0 ;
  assign n24198 = ~n24196 & n24197 ;
  assign n24199 = n6709 ^ n1469 ^ 1'b0 ;
  assign n24200 = n24198 & n24199 ;
  assign n24201 = n24200 ^ n11046 ^ 1'b0 ;
  assign n24202 = n2345 | n14515 ;
  assign n24203 = n3160 | n5667 ;
  assign n24204 = n24203 ^ n7649 ^ 1'b0 ;
  assign n24205 = n3112 | n24204 ;
  assign n24206 = n24205 ^ n1239 ^ 1'b0 ;
  assign n24207 = n9237 & n17500 ;
  assign n24208 = n11999 & ~n22110 ;
  assign n24209 = n10311 ^ n5874 ^ 1'b0 ;
  assign n24210 = ~n17060 & n24209 ;
  assign n24211 = n2709 & n10160 ;
  assign n24212 = n24211 ^ n22599 ^ 1'b0 ;
  assign n24213 = n19285 | n24212 ;
  assign n24214 = n24213 ^ n5772 ^ 1'b0 ;
  assign n24215 = ( n19876 & n24210 ) | ( n19876 & n24214 ) | ( n24210 & n24214 ) ;
  assign n24216 = n18521 & n24215 ;
  assign n24217 = ( n3456 & n7488 ) | ( n3456 & n9862 ) | ( n7488 & n9862 ) ;
  assign n24218 = n1197 & n24217 ;
  assign n24219 = n283 & n24218 ;
  assign n24220 = ( n989 & ~n12997 ) | ( n989 & n13704 ) | ( ~n12997 & n13704 ) ;
  assign n24221 = ( n9645 & n10665 ) | ( n9645 & ~n10682 ) | ( n10665 & ~n10682 ) ;
  assign n24222 = n24221 ^ n11377 ^ 1'b0 ;
  assign n24223 = n24220 & n24222 ;
  assign n24224 = n24223 ^ n18879 ^ 1'b0 ;
  assign n24225 = n24219 | n24224 ;
  assign n24226 = n18575 ^ n10056 ^ 1'b0 ;
  assign n24227 = ~n4066 & n24226 ;
  assign n24228 = n13956 & ~n19694 ;
  assign n24229 = n7088 & n24228 ;
  assign n24230 = ~n24227 & n24229 ;
  assign n24231 = n13188 & n24013 ;
  assign n24232 = ( n2133 & n15950 ) | ( n2133 & ~n16106 ) | ( n15950 & ~n16106 ) ;
  assign n24234 = n23337 ^ n892 ^ 1'b0 ;
  assign n24233 = n18091 & ~n18116 ;
  assign n24235 = n24234 ^ n24233 ^ 1'b0 ;
  assign n24236 = n19042 ^ n1190 ^ 1'b0 ;
  assign n24237 = ~n1782 & n21981 ;
  assign n24238 = n24237 ^ n11080 ^ 1'b0 ;
  assign n24239 = n24217 ^ n16271 ^ n2382 ;
  assign n24240 = n15002 | n23031 ;
  assign n24241 = n1819 | n11642 ;
  assign n24242 = n24241 ^ n5039 ^ 1'b0 ;
  assign n24243 = n2194 & n16711 ;
  assign n24244 = n24243 ^ n3721 ^ 1'b0 ;
  assign n24245 = n10886 & ~n24244 ;
  assign n24246 = n24245 ^ n3261 ^ 1'b0 ;
  assign n24247 = ( ~n7000 & n24242 ) | ( ~n7000 & n24246 ) | ( n24242 & n24246 ) ;
  assign n24248 = n24247 ^ n2786 ^ 1'b0 ;
  assign n24249 = ~n16848 & n24248 ;
  assign n24250 = n16134 ^ n6896 ^ 1'b0 ;
  assign n24251 = n24079 | n24250 ;
  assign n24252 = n1761 | n16491 ;
  assign n24253 = n24252 ^ n4741 ^ n4359 ;
  assign n24255 = ( n2447 & n5992 ) | ( n2447 & n12021 ) | ( n5992 & n12021 ) ;
  assign n24254 = n16005 & n20439 ;
  assign n24256 = n24255 ^ n24254 ^ 1'b0 ;
  assign n24257 = ( n2692 & ~n12125 ) | ( n2692 & n24256 ) | ( ~n12125 & n24256 ) ;
  assign n24258 = n1023 | n22605 ;
  assign n24259 = n24258 ^ n17794 ^ 1'b0 ;
  assign n24260 = ~n14030 & n24259 ;
  assign n24264 = ~n8901 & n12922 ;
  assign n24261 = n8250 ^ n5754 ^ 1'b0 ;
  assign n24262 = n10081 & n24261 ;
  assign n24263 = n24262 ^ n13777 ^ 1'b0 ;
  assign n24265 = n24264 ^ n24263 ^ n2519 ;
  assign n24266 = n21827 & n24265 ;
  assign n24267 = n17771 ^ n17232 ^ n851 ;
  assign n24268 = ( n14669 & n20965 ) | ( n14669 & ~n24267 ) | ( n20965 & ~n24267 ) ;
  assign n24269 = n12020 ^ n3645 ^ 1'b0 ;
  assign n24270 = n24269 ^ n3530 ^ 1'b0 ;
  assign n24271 = n24270 ^ n8386 ^ 1'b0 ;
  assign n24272 = ( n315 & ~n4442 ) | ( n315 & n4977 ) | ( ~n4442 & n4977 ) ;
  assign n24273 = n12965 | n24272 ;
  assign n24274 = ( n3989 & n24271 ) | ( n3989 & n24273 ) | ( n24271 & n24273 ) ;
  assign n24275 = n11244 ^ x73 ^ 1'b0 ;
  assign n24276 = ( n5581 & n10473 ) | ( n5581 & ~n12167 ) | ( n10473 & ~n12167 ) ;
  assign n24277 = n6766 ^ n1700 ^ 1'b0 ;
  assign n24278 = n24277 ^ n21654 ^ 1'b0 ;
  assign n24279 = ~n24276 & n24278 ;
  assign n24280 = ~n24275 & n24279 ;
  assign n24281 = n14979 & ~n18060 ;
  assign n24282 = n19402 ^ n2661 ^ 1'b0 ;
  assign n24283 = n24281 & n24282 ;
  assign n24284 = n7695 ^ n2002 ^ 1'b0 ;
  assign n24288 = n9435 | n21487 ;
  assign n24289 = n17099 & ~n24288 ;
  assign n24290 = n6719 | n7311 ;
  assign n24291 = n7655 & ~n24290 ;
  assign n24292 = n24289 & ~n24291 ;
  assign n24285 = n9713 ^ n369 ^ 1'b0 ;
  assign n24286 = n6729 | n24285 ;
  assign n24287 = n11524 | n24286 ;
  assign n24293 = n24292 ^ n24287 ^ 1'b0 ;
  assign n24294 = n1192 ^ n390 ^ 1'b0 ;
  assign n24295 = n3255 & ~n24294 ;
  assign n24296 = n7495 & ~n7710 ;
  assign n24297 = ~n24295 & n24296 ;
  assign n24298 = ( x64 & n1172 ) | ( x64 & n16286 ) | ( n1172 & n16286 ) ;
  assign n24299 = n13057 | n24298 ;
  assign n24300 = n5610 & n9611 ;
  assign n24301 = n3120 & ~n8696 ;
  assign n24302 = n787 & n24301 ;
  assign n24303 = n24302 ^ n17157 ^ n10526 ;
  assign n24304 = n6095 & ~n10636 ;
  assign n24305 = n10779 & n24304 ;
  assign n24306 = n19033 ^ n536 ^ 1'b0 ;
  assign n24307 = ~n1097 & n12818 ;
  assign n24308 = n24307 ^ n17631 ^ 1'b0 ;
  assign n24309 = n6694 ^ n1612 ^ 1'b0 ;
  assign n24310 = n23255 & ~n24309 ;
  assign n24311 = ~n3716 & n24310 ;
  assign n24312 = n24311 ^ n9198 ^ 1'b0 ;
  assign n24313 = ~n2741 & n24312 ;
  assign n24314 = n3797 & n8474 ;
  assign n24315 = n17032 & n24314 ;
  assign n24316 = ~n16639 & n24315 ;
  assign n24317 = ~n13311 & n22659 ;
  assign n24318 = ~n5006 & n19097 ;
  assign n24319 = n24318 ^ n24214 ^ 1'b0 ;
  assign n24320 = n535 & n21548 ;
  assign n24321 = n14441 ^ n2636 ^ 1'b0 ;
  assign n24322 = ~n1786 & n24321 ;
  assign n24323 = n5884 ^ n4879 ^ 1'b0 ;
  assign n24324 = n19579 & n24323 ;
  assign n24325 = n24324 ^ n21229 ^ n9774 ;
  assign n24326 = n18078 ^ n1467 ^ 1'b0 ;
  assign n24327 = n13742 ^ n9065 ^ n987 ;
  assign n24328 = n24327 ^ n686 ^ n580 ;
  assign n24329 = n24328 ^ n20868 ^ n8038 ;
  assign n24330 = n22628 ^ n22453 ^ 1'b0 ;
  assign n24331 = n3141 | n8146 ;
  assign n24332 = n11389 & ~n24331 ;
  assign n24333 = n24332 ^ n22392 ^ 1'b0 ;
  assign n24334 = n3979 | n4981 ;
  assign n24335 = n24334 ^ n351 ^ 1'b0 ;
  assign n24336 = n20731 & n23998 ;
  assign n24337 = ( x224 & n5954 ) | ( x224 & n7358 ) | ( n5954 & n7358 ) ;
  assign n24338 = ~n3145 & n24337 ;
  assign n24339 = n1806 & n4778 ;
  assign n24340 = n4676 ^ n957 ^ 1'b0 ;
  assign n24341 = n24340 ^ n12689 ^ n369 ;
  assign n24342 = ( n5313 & n24339 ) | ( n5313 & n24341 ) | ( n24339 & n24341 ) ;
  assign n24343 = ~n4666 & n24342 ;
  assign n24344 = n9957 | n24343 ;
  assign n24345 = n23560 | n24344 ;
  assign n24346 = n19850 ^ n18329 ^ 1'b0 ;
  assign n24347 = n10212 ^ n3141 ^ 1'b0 ;
  assign n24348 = n6112 & ~n7298 ;
  assign n24349 = n24348 ^ n23317 ^ 1'b0 ;
  assign n24350 = n24347 | n24349 ;
  assign n24351 = n24350 ^ n913 ^ 1'b0 ;
  assign n24352 = ( n15786 & n21150 ) | ( n15786 & ~n22160 ) | ( n21150 & ~n22160 ) ;
  assign n24353 = n8200 ^ n449 ^ 1'b0 ;
  assign n24354 = ~n9767 & n24353 ;
  assign n24355 = n9715 & n14340 ;
  assign n24356 = ( x236 & n24354 ) | ( x236 & ~n24355 ) | ( n24354 & ~n24355 ) ;
  assign n24357 = n6912 | n10650 ;
  assign n24358 = n14166 & ~n24357 ;
  assign n24359 = n24358 ^ n4917 ^ 1'b0 ;
  assign n24360 = ~n13587 & n21154 ;
  assign n24361 = ~n2201 & n24360 ;
  assign n24362 = n8029 | n11935 ;
  assign n24363 = n24362 ^ n10198 ^ 1'b0 ;
  assign n24364 = n10649 & ~n13931 ;
  assign n24365 = n24364 ^ n4312 ^ 1'b0 ;
  assign n24366 = n2151 & ~n4915 ;
  assign n24367 = n15039 & n24366 ;
  assign n24369 = ~n2113 & n7986 ;
  assign n24370 = n24369 ^ n17491 ^ 1'b0 ;
  assign n24368 = n17897 & ~n18853 ;
  assign n24371 = n24370 ^ n24368 ^ 1'b0 ;
  assign n24376 = ~n6882 & n19868 ;
  assign n24372 = n10068 | n13705 ;
  assign n24373 = n14367 & ~n24372 ;
  assign n24374 = n24373 ^ n12594 ^ n8756 ;
  assign n24375 = n17256 | n24374 ;
  assign n24377 = n24376 ^ n24375 ^ 1'b0 ;
  assign n24378 = n12405 & n12600 ;
  assign n24379 = ( n4797 & ~n9093 ) | ( n4797 & n13154 ) | ( ~n9093 & n13154 ) ;
  assign n24380 = n24379 ^ n12590 ^ 1'b0 ;
  assign n24381 = ~n2054 & n3154 ;
  assign n24382 = n3635 | n11765 ;
  assign n24383 = n24382 ^ n8711 ^ 1'b0 ;
  assign n24384 = n5760 & n24383 ;
  assign n24385 = n24384 ^ n15969 ^ n10973 ;
  assign n24386 = ~n2217 & n8548 ;
  assign n24387 = n884 | n17137 ;
  assign n24388 = n24387 ^ n21949 ^ 1'b0 ;
  assign n24389 = ~n2342 & n14631 ;
  assign n24390 = n21882 & n24389 ;
  assign n24391 = n12257 ^ n1742 ^ 1'b0 ;
  assign n24392 = n3765 & ~n24391 ;
  assign n24393 = ~n9355 & n24392 ;
  assign n24394 = ~n16305 & n24393 ;
  assign n24395 = n15857 & ~n24394 ;
  assign n24396 = n7953 & n15432 ;
  assign n24397 = n6694 | n11585 ;
  assign n24398 = n20950 ^ n17956 ^ 1'b0 ;
  assign n24399 = n12069 & n24398 ;
  assign n24400 = n5213 & n24399 ;
  assign n24401 = n1881 & n8399 ;
  assign n24402 = n13215 ^ n8800 ^ 1'b0 ;
  assign n24403 = ( n6673 & ~n16757 ) | ( n6673 & n17027 ) | ( ~n16757 & n17027 ) ;
  assign n24404 = n24403 ^ n12350 ^ 1'b0 ;
  assign n24405 = ( n3039 & n11134 ) | ( n3039 & ~n17371 ) | ( n11134 & ~n17371 ) ;
  assign n24406 = n2819 | n19695 ;
  assign n24407 = n10232 & n18844 ;
  assign n24408 = n6969 | n18473 ;
  assign n24409 = n24408 ^ n11413 ^ 1'b0 ;
  assign n24410 = n19295 ^ n14876 ^ 1'b0 ;
  assign n24411 = n13617 ^ n5261 ^ 1'b0 ;
  assign n24412 = n10881 ^ n1166 ^ 1'b0 ;
  assign n24413 = ~n3972 & n14016 ;
  assign n24414 = n2751 | n5384 ;
  assign n24415 = n24414 ^ n6371 ^ 1'b0 ;
  assign n24416 = n5198 | n24415 ;
  assign n24417 = n24416 ^ n23584 ^ 1'b0 ;
  assign n24418 = n1115 | n15378 ;
  assign n24419 = n24418 ^ n10816 ^ 1'b0 ;
  assign n24420 = n24419 ^ n14320 ^ 1'b0 ;
  assign n24421 = n1544 & n24420 ;
  assign n24422 = n24421 ^ n12557 ^ 1'b0 ;
  assign n24423 = n4331 & ~n24422 ;
  assign n24424 = n8949 ^ n2501 ^ n878 ;
  assign n24425 = n10230 & n24424 ;
  assign n24426 = n557 & n24425 ;
  assign n24427 = ( n8783 & n15874 ) | ( n8783 & n24426 ) | ( n15874 & n24426 ) ;
  assign n24428 = n8769 ^ n7986 ^ 1'b0 ;
  assign n24429 = n6193 & ~n11175 ;
  assign n24430 = ~n21241 & n24429 ;
  assign n24431 = n14341 ^ n2930 ^ 1'b0 ;
  assign n24432 = ~n11799 & n17104 ;
  assign n24433 = n2495 & n24432 ;
  assign n24434 = n24433 ^ n16845 ^ 1'b0 ;
  assign n24438 = n472 & n2963 ;
  assign n24439 = n5613 & n24438 ;
  assign n24440 = n18622 & ~n24439 ;
  assign n24441 = n8049 & n24440 ;
  assign n24435 = n6030 & n16415 ;
  assign n24436 = n24435 ^ n12372 ^ 1'b0 ;
  assign n24437 = n19670 & n24436 ;
  assign n24442 = n24441 ^ n24437 ^ 1'b0 ;
  assign n24443 = n21626 & n24442 ;
  assign n24444 = n24443 ^ n3540 ^ 1'b0 ;
  assign n24445 = ~n11866 & n12419 ;
  assign n24446 = n24445 ^ n22511 ^ 1'b0 ;
  assign n24447 = ~n24444 & n24446 ;
  assign n24448 = n16773 ^ n16450 ^ n1010 ;
  assign n24449 = ( n12498 & ~n18591 ) | ( n12498 & n24072 ) | ( ~n18591 & n24072 ) ;
  assign n24450 = n24337 ^ n22042 ^ 1'b0 ;
  assign n24451 = n24450 ^ n15063 ^ n826 ;
  assign n24452 = n23366 & n24451 ;
  assign n24453 = n9196 ^ n6362 ^ 1'b0 ;
  assign n24454 = ~n5739 & n24453 ;
  assign n24457 = n5603 & ~n10205 ;
  assign n24458 = n24457 ^ n6369 ^ 1'b0 ;
  assign n24455 = n7965 ^ n2847 ^ 1'b0 ;
  assign n24456 = n9831 | n24455 ;
  assign n24459 = n24458 ^ n24456 ^ 1'b0 ;
  assign n24460 = n24454 & n24459 ;
  assign n24461 = n12837 ^ n1850 ^ 1'b0 ;
  assign n24462 = ~n5605 & n6327 ;
  assign n24463 = ( n3734 & n8049 ) | ( n3734 & ~n24462 ) | ( n8049 & ~n24462 ) ;
  assign n24465 = n1011 ^ n791 ^ 1'b0 ;
  assign n24464 = n7909 & n9091 ;
  assign n24466 = n24465 ^ n24464 ^ 1'b0 ;
  assign n24467 = n11499 | n12929 ;
  assign n24468 = n24467 ^ n19743 ^ 1'b0 ;
  assign n24469 = n5809 | n24468 ;
  assign n24470 = n21753 & ~n24469 ;
  assign n24471 = n12961 ^ n10168 ^ n4015 ;
  assign n24472 = n24471 ^ n22770 ^ n10205 ;
  assign n24473 = n21133 & n24472 ;
  assign n24474 = ( n3701 & ~n4170 ) | ( n3701 & n12078 ) | ( ~n4170 & n12078 ) ;
  assign n24475 = n24474 ^ n10664 ^ 1'b0 ;
  assign n24476 = ~n4503 & n12483 ;
  assign n24477 = ( n22094 & n24475 ) | ( n22094 & n24476 ) | ( n24475 & n24476 ) ;
  assign n24481 = n10861 ^ n7437 ^ 1'b0 ;
  assign n24482 = n9954 & ~n24481 ;
  assign n24478 = n4694 ^ n1356 ^ 1'b0 ;
  assign n24479 = n21012 | n24478 ;
  assign n24480 = n14830 | n24479 ;
  assign n24483 = n24482 ^ n24480 ^ 1'b0 ;
  assign n24484 = n5549 & ~n8181 ;
  assign n24485 = n24484 ^ n7773 ^ 1'b0 ;
  assign n24486 = n8640 | n24485 ;
  assign n24487 = n24483 | n24486 ;
  assign n24488 = n6616 ^ n4937 ^ 1'b0 ;
  assign n24489 = ~n8619 & n24488 ;
  assign n24490 = n24489 ^ n11014 ^ n700 ;
  assign n24491 = n7599 & n9694 ;
  assign n24492 = n24491 ^ n11532 ^ 1'b0 ;
  assign n24493 = n9892 & ~n17634 ;
  assign n24494 = n14441 & n24493 ;
  assign n24495 = n22610 ^ n13651 ^ n2836 ;
  assign n24496 = n7632 ^ n5170 ^ 1'b0 ;
  assign n24497 = n4293 & n24496 ;
  assign n24498 = n10406 & n12437 ;
  assign n24499 = ~n3035 & n8455 ;
  assign n24500 = n24498 & n24499 ;
  assign n24503 = n3187 ^ n2359 ^ 1'b0 ;
  assign n24504 = n12897 & n24503 ;
  assign n24505 = ~n8637 & n17993 ;
  assign n24506 = ~n24504 & n24505 ;
  assign n24501 = n7071 | n14967 ;
  assign n24502 = n24501 ^ n10578 ^ 1'b0 ;
  assign n24507 = n24506 ^ n24502 ^ n17180 ;
  assign n24508 = ~n12579 & n18459 ;
  assign n24509 = n24508 ^ n22317 ^ 1'b0 ;
  assign n24510 = ~n3596 & n6232 ;
  assign n24511 = n2253 | n24510 ;
  assign n24512 = n24511 ^ n5008 ^ 1'b0 ;
  assign n24513 = n12330 & n24512 ;
  assign n24514 = n24513 ^ n2040 ^ 1'b0 ;
  assign n24515 = n17510 ^ n7693 ^ 1'b0 ;
  assign n24516 = n20108 & n24515 ;
  assign n24517 = n19587 ^ n258 ^ 1'b0 ;
  assign n24518 = ~n3645 & n24517 ;
  assign n24520 = ( ~n2628 & n10810 ) | ( ~n2628 & n14623 ) | ( n10810 & n14623 ) ;
  assign n24519 = ~n21229 & n23609 ;
  assign n24521 = n24520 ^ n24519 ^ 1'b0 ;
  assign n24522 = n2644 & n22406 ;
  assign n24523 = n3141 ^ n2860 ^ n1713 ;
  assign n24524 = n24523 ^ n3291 ^ 1'b0 ;
  assign n24525 = n8316 | n16884 ;
  assign n24526 = n24524 | n24525 ;
  assign n24527 = n24526 ^ n17903 ^ 1'b0 ;
  assign n24528 = n15366 & ~n24527 ;
  assign n24529 = n5903 ^ x126 ^ 1'b0 ;
  assign n24530 = n7897 & ~n24529 ;
  assign n24531 = n4799 & n5920 ;
  assign n24532 = n24531 ^ n18169 ^ 1'b0 ;
  assign n24533 = n24532 ^ n16176 ^ n9873 ;
  assign n24534 = n24436 ^ n3513 ^ 1'b0 ;
  assign n24535 = n18950 & ~n24534 ;
  assign n24536 = n959 & n8167 ;
  assign n24537 = n24536 ^ n7029 ^ 1'b0 ;
  assign n24538 = ~n1443 & n18176 ;
  assign n24539 = ~n24537 & n24538 ;
  assign n24540 = n24539 ^ n16091 ^ 1'b0 ;
  assign n24541 = n5511 & ~n24540 ;
  assign n24542 = n3540 & n4509 ;
  assign n24543 = n11974 | n20731 ;
  assign n24544 = ~n13416 & n15085 ;
  assign n24545 = ( n24542 & n24543 ) | ( n24542 & ~n24544 ) | ( n24543 & ~n24544 ) ;
  assign n24546 = n21739 ^ n3274 ^ 1'b0 ;
  assign n24547 = n19922 | n24546 ;
  assign n24548 = n24547 ^ n4426 ^ 1'b0 ;
  assign n24549 = n24548 ^ n4200 ^ n1930 ;
  assign n24550 = n12531 & n24549 ;
  assign n24551 = n22966 ^ n16119 ^ n15425 ;
  assign n24552 = ~n983 & n12021 ;
  assign n24553 = n714 & n24552 ;
  assign n24554 = ( ~n16489 & n24551 ) | ( ~n16489 & n24553 ) | ( n24551 & n24553 ) ;
  assign n24555 = ~n444 & n1999 ;
  assign n24556 = ~n5778 & n24555 ;
  assign n24557 = n24556 ^ n20843 ^ 1'b0 ;
  assign n24558 = n1254 | n1430 ;
  assign n24559 = n24558 ^ n12452 ^ 1'b0 ;
  assign n24560 = ( n4081 & ~n4405 ) | ( n4081 & n24559 ) | ( ~n4405 & n24559 ) ;
  assign n24561 = n24560 ^ n5768 ^ 1'b0 ;
  assign n24562 = n2763 & ~n8402 ;
  assign n24563 = n24562 ^ n8715 ^ 1'b0 ;
  assign n24564 = n21708 & ~n24563 ;
  assign n24565 = n3493 & n24564 ;
  assign n24566 = n22927 & ~n24565 ;
  assign n24567 = n24561 & n24566 ;
  assign n24568 = n10097 & ~n11845 ;
  assign n24569 = x34 & n10440 ;
  assign n24570 = n10488 ^ n5138 ^ 1'b0 ;
  assign n24571 = ~n547 & n24570 ;
  assign n24572 = n12601 & n24571 ;
  assign n24573 = ( n4597 & n10013 ) | ( n4597 & n10683 ) | ( n10013 & n10683 ) ;
  assign n24575 = n10394 & ~n14743 ;
  assign n24576 = n24575 ^ n14144 ^ 1'b0 ;
  assign n24574 = n13775 & ~n14796 ;
  assign n24577 = n24576 ^ n24574 ^ 1'b0 ;
  assign n24578 = n20476 ^ n4256 ^ 1'b0 ;
  assign n24579 = n20355 ^ x65 ^ 1'b0 ;
  assign n24580 = ( n11169 & n14095 ) | ( n11169 & n22983 ) | ( n14095 & n22983 ) ;
  assign n24581 = n2395 & n24580 ;
  assign n24582 = n1855 & ~n19326 ;
  assign n24583 = n24582 ^ n21832 ^ 1'b0 ;
  assign n24584 = n19993 ^ n1368 ^ 1'b0 ;
  assign n24585 = n17266 & ~n24584 ;
  assign n24586 = n15316 | n22310 ;
  assign n24587 = ~n3433 & n23461 ;
  assign n24588 = n2449 & n24587 ;
  assign n24589 = n12325 & n24588 ;
  assign n24590 = n23696 ^ n22040 ^ n13817 ;
  assign n24591 = n23957 & ~n24590 ;
  assign n24592 = n17655 ^ n634 ^ 1'b0 ;
  assign n24593 = ~n3056 & n6715 ;
  assign n24594 = ~n1124 & n24593 ;
  assign n24595 = n15188 ^ n4266 ^ 1'b0 ;
  assign n24596 = n12201 & n15723 ;
  assign n24597 = n24596 ^ n11447 ^ 1'b0 ;
  assign n24600 = n17866 ^ n5782 ^ n2924 ;
  assign n24598 = n1255 & n21284 ;
  assign n24599 = ~n1700 & n24598 ;
  assign n24601 = n24600 ^ n24599 ^ n6667 ;
  assign n24602 = n24561 ^ n14258 ^ 1'b0 ;
  assign n24603 = n20658 | n24602 ;
  assign n24604 = n3283 & ~n24603 ;
  assign n24605 = n14245 ^ n11397 ^ 1'b0 ;
  assign n24606 = ( n3600 & n4765 ) | ( n3600 & n24605 ) | ( n4765 & n24605 ) ;
  assign n24607 = n24606 ^ n23918 ^ 1'b0 ;
  assign n24608 = n5243 | n24607 ;
  assign n24613 = n9096 ^ n7391 ^ n5832 ;
  assign n24614 = ~n6126 & n24613 ;
  assign n24609 = n7867 ^ n3632 ^ n2260 ;
  assign n24610 = n5192 & ~n24609 ;
  assign n24611 = n546 & ~n24610 ;
  assign n24612 = n9860 & ~n24611 ;
  assign n24615 = n24614 ^ n24612 ^ n2281 ;
  assign n24620 = n904 & ~n18622 ;
  assign n24616 = n2611 & n8016 ;
  assign n24617 = n24616 ^ n4642 ^ n4518 ;
  assign n24618 = n358 & n24617 ;
  assign n24619 = n14219 & ~n24618 ;
  assign n24621 = n24620 ^ n24619 ^ 1'b0 ;
  assign n24622 = ( n6705 & ~n13673 ) | ( n6705 & n15161 ) | ( ~n13673 & n15161 ) ;
  assign n24624 = n10872 ^ n8825 ^ 1'b0 ;
  assign n24625 = n15295 | n24624 ;
  assign n24623 = n21838 ^ n9350 ^ 1'b0 ;
  assign n24626 = n24625 ^ n24623 ^ n7830 ;
  assign n24630 = n11596 | n21616 ;
  assign n24631 = n2797 & ~n24630 ;
  assign n24627 = n6628 & n19143 ;
  assign n24628 = n24627 ^ n4920 ^ 1'b0 ;
  assign n24629 = n18394 & ~n24628 ;
  assign n24632 = n24631 ^ n24629 ^ 1'b0 ;
  assign n24634 = n22870 ^ n9302 ^ n8655 ;
  assign n24633 = n6047 & n21090 ;
  assign n24635 = n24634 ^ n24633 ^ 1'b0 ;
  assign n24636 = n11268 ^ n3270 ^ 1'b0 ;
  assign n24637 = n24635 & n24636 ;
  assign n24638 = n24637 ^ n9047 ^ 1'b0 ;
  assign n24639 = n3272 & n7049 ;
  assign n24640 = n9919 & n24639 ;
  assign n24641 = ~n12415 & n21510 ;
  assign n24642 = n7380 & ~n12087 ;
  assign n24643 = x182 & ~n5384 ;
  assign n24644 = ~n5100 & n14310 ;
  assign n24645 = n21370 & n24644 ;
  assign n24646 = n433 & n14784 ;
  assign n24647 = ~n23696 & n24646 ;
  assign n24648 = n24647 ^ n1800 ^ 1'b0 ;
  assign n24649 = n3601 ^ n2116 ^ 1'b0 ;
  assign n24650 = ( n444 & ~n3534 ) | ( n444 & n24649 ) | ( ~n3534 & n24649 ) ;
  assign n24651 = ( ~n16905 & n24454 ) | ( ~n16905 & n24650 ) | ( n24454 & n24650 ) ;
  assign n24652 = n21504 & n21644 ;
  assign n24653 = n4358 & n24652 ;
  assign n24654 = n1499 & ~n5635 ;
  assign n24655 = n24654 ^ n3998 ^ 1'b0 ;
  assign n24656 = n8702 & n12755 ;
  assign n24657 = ~n7824 & n24656 ;
  assign n24658 = ( n5369 & ~n16950 ) | ( n5369 & n24657 ) | ( ~n16950 & n24657 ) ;
  assign n24659 = n17507 | n24658 ;
  assign n24660 = n6724 & ~n24659 ;
  assign n24661 = n12091 ^ n10813 ^ 1'b0 ;
  assign n24662 = n18495 & n21570 ;
  assign n24663 = n24661 & n24662 ;
  assign n24664 = n6045 | n7405 ;
  assign n24666 = ( n1147 & n1692 ) | ( n1147 & ~n6132 ) | ( n1692 & ~n6132 ) ;
  assign n24667 = ~n20263 & n24666 ;
  assign n24668 = ~n14100 & n24667 ;
  assign n24665 = n11878 & ~n18898 ;
  assign n24669 = n24668 ^ n24665 ^ 1'b0 ;
  assign n24670 = ~n13234 & n24669 ;
  assign n24671 = n24670 ^ n6372 ^ 1'b0 ;
  assign n24672 = n2580 ^ n634 ^ 1'b0 ;
  assign n24673 = ~n4099 & n24672 ;
  assign n24674 = n24673 ^ n11593 ^ 1'b0 ;
  assign n24675 = n3307 | n24674 ;
  assign n24676 = n13944 & n24675 ;
  assign n24677 = n6977 | n20651 ;
  assign n24678 = n6977 & ~n24677 ;
  assign n24679 = n24678 ^ n9375 ^ 1'b0 ;
  assign n24680 = n1328 & ~n24679 ;
  assign n24681 = n4759 | n22856 ;
  assign n24682 = n14216 ^ n5498 ^ n4934 ;
  assign n24683 = n2405 | n7418 ;
  assign n24684 = n18555 ^ n3835 ^ 1'b0 ;
  assign n24685 = n3681 & ~n6142 ;
  assign n24686 = n24685 ^ n9824 ^ 1'b0 ;
  assign n24687 = n18812 & ~n24686 ;
  assign n24688 = n4973 ^ n2358 ^ 1'b0 ;
  assign n24689 = ( n2754 & n11457 ) | ( n2754 & n24688 ) | ( n11457 & n24688 ) ;
  assign n24690 = n21109 ^ n9077 ^ 1'b0 ;
  assign n24691 = n24689 & n24690 ;
  assign n24692 = ~n2728 & n8459 ;
  assign n24693 = n14945 & ~n24692 ;
  assign n24694 = n7402 ^ n967 ^ 1'b0 ;
  assign n24695 = n11765 ^ n6204 ^ 1'b0 ;
  assign n24696 = n12881 & n24695 ;
  assign n24697 = n15914 & n24492 ;
  assign n24698 = n12762 & ~n20693 ;
  assign n24699 = n677 & ~n24698 ;
  assign n24700 = n17740 & n24699 ;
  assign n24701 = n13201 ^ n10366 ^ 1'b0 ;
  assign n24702 = x25 & n18691 ;
  assign n24703 = n1972 | n14075 ;
  assign n24704 = n19919 & ~n24703 ;
  assign n24705 = n3087 & n7172 ;
  assign n24706 = n24705 ^ n16233 ^ 1'b0 ;
  assign n24709 = n6682 ^ n5255 ^ 1'b0 ;
  assign n24707 = ~n11943 & n19230 ;
  assign n24708 = n7809 | n24707 ;
  assign n24710 = n24709 ^ n24708 ^ 1'b0 ;
  assign n24711 = n7693 | n15607 ;
  assign n24712 = n3915 | n11043 ;
  assign n24713 = ( ~n8032 & n24711 ) | ( ~n8032 & n24712 ) | ( n24711 & n24712 ) ;
  assign n24714 = n11914 ^ n11431 ^ n5943 ;
  assign n24715 = n24714 ^ n13726 ^ 1'b0 ;
  assign n24716 = n13415 ^ n1330 ^ 1'b0 ;
  assign n24717 = ~n14399 & n24716 ;
  assign n24718 = n5312 & ~n23411 ;
  assign n24719 = n24718 ^ n12592 ^ 1'b0 ;
  assign n24720 = n17306 ^ n9341 ^ n2342 ;
  assign n24721 = n24720 ^ n18668 ^ 1'b0 ;
  assign n24722 = n10093 & ~n24721 ;
  assign n24723 = ( n1202 & n6253 ) | ( n1202 & n23480 ) | ( n6253 & n23480 ) ;
  assign n24724 = n9835 ^ n1255 ^ 1'b0 ;
  assign n24725 = n7928 ^ n6325 ^ 1'b0 ;
  assign n24726 = ~n1442 & n15758 ;
  assign n24727 = n24725 & n24726 ;
  assign n24728 = n24727 ^ n12607 ^ 1'b0 ;
  assign n24729 = ( n813 & ~n8592 ) | ( n813 & n11531 ) | ( ~n8592 & n11531 ) ;
  assign n24730 = n24729 ^ n6813 ^ 1'b0 ;
  assign n24731 = ~n1007 & n11904 ;
  assign n24732 = n24731 ^ n23442 ^ 1'b0 ;
  assign n24733 = n11174 & ~n16211 ;
  assign n24734 = n24733 ^ n11784 ^ 1'b0 ;
  assign n24735 = ( n7263 & n18567 ) | ( n7263 & ~n24734 ) | ( n18567 & ~n24734 ) ;
  assign n24737 = n1524 & ~n14010 ;
  assign n24736 = n12517 & n22578 ;
  assign n24738 = n24737 ^ n24736 ^ 1'b0 ;
  assign n24743 = n1982 | n4175 ;
  assign n24742 = n6193 | n7509 ;
  assign n24744 = n24743 ^ n24742 ^ 1'b0 ;
  assign n24739 = n3027 & n4570 ;
  assign n24740 = ( ~n8062 & n12060 ) | ( ~n8062 & n24739 ) | ( n12060 & n24739 ) ;
  assign n24741 = n2956 & n24740 ;
  assign n24745 = n24744 ^ n24741 ^ 1'b0 ;
  assign n24746 = n10312 ^ n4719 ^ 1'b0 ;
  assign n24747 = x221 & ~n24746 ;
  assign n24748 = n24747 ^ n11845 ^ 1'b0 ;
  assign n24749 = n24748 ^ n8891 ^ 1'b0 ;
  assign n24750 = n22985 ^ n20150 ^ n2722 ;
  assign n24751 = n5947 & ~n18509 ;
  assign n24752 = n18562 ^ n17672 ^ 1'b0 ;
  assign n24753 = n3523 | n7306 ;
  assign n24754 = n3422 & ~n24753 ;
  assign n24755 = n24754 ^ n2868 ^ 1'b0 ;
  assign n24756 = n9882 ^ n7615 ^ 1'b0 ;
  assign n24757 = ~n10374 & n24756 ;
  assign n24758 = n12850 & ~n24757 ;
  assign n24759 = n5994 ^ n4444 ^ x94 ;
  assign n24760 = n9899 ^ n7146 ^ 1'b0 ;
  assign n24761 = n20598 ^ n17506 ^ 1'b0 ;
  assign n24762 = n2543 | n23416 ;
  assign n24763 = n3253 & ~n24762 ;
  assign n24764 = n379 | n5716 ;
  assign n24765 = n24764 ^ n21012 ^ 1'b0 ;
  assign n24766 = n12802 & ~n24765 ;
  assign n24767 = n24766 ^ n18020 ^ 1'b0 ;
  assign n24768 = n3296 & ~n7716 ;
  assign n24769 = ( ~n20128 & n22055 ) | ( ~n20128 & n22668 ) | ( n22055 & n22668 ) ;
  assign n24770 = n15969 ^ n824 ^ 1'b0 ;
  assign n24774 = ~n1530 & n4748 ;
  assign n24775 = n24774 ^ n12906 ^ 1'b0 ;
  assign n24771 = n16900 & ~n16958 ;
  assign n24772 = n24771 ^ n15806 ^ 1'b0 ;
  assign n24773 = ~n11747 & n24772 ;
  assign n24776 = n24775 ^ n24773 ^ 1'b0 ;
  assign n24777 = n15998 ^ n374 ^ 1'b0 ;
  assign n24778 = n690 | n24777 ;
  assign n24779 = n10586 ^ n323 ^ 1'b0 ;
  assign n24780 = n24779 ^ n18600 ^ n7444 ;
  assign n24781 = ( n14206 & n24778 ) | ( n14206 & n24780 ) | ( n24778 & n24780 ) ;
  assign n24782 = n22361 ^ n10820 ^ n6544 ;
  assign n24783 = n1551 ^ n1550 ^ n1034 ;
  assign n24784 = n24783 ^ n329 ^ 1'b0 ;
  assign n24785 = n4029 & n24784 ;
  assign n24786 = n4306 ^ n3947 ^ n1811 ;
  assign n24787 = n10365 & n24786 ;
  assign n24788 = n12627 ^ n6128 ^ 1'b0 ;
  assign n24789 = ~n5851 & n14390 ;
  assign n24790 = n24789 ^ n3422 ^ 1'b0 ;
  assign n24791 = ( n6342 & n17128 ) | ( n6342 & n24790 ) | ( n17128 & n24790 ) ;
  assign n24792 = ( n6899 & ~n9614 ) | ( n6899 & n24791 ) | ( ~n9614 & n24791 ) ;
  assign n24793 = ~n7677 & n16625 ;
  assign n24794 = n8446 & n9948 ;
  assign n24795 = ( n6155 & n24793 ) | ( n6155 & ~n24794 ) | ( n24793 & ~n24794 ) ;
  assign n24796 = n439 | n20287 ;
  assign n24797 = n1473 & ~n3027 ;
  assign n24798 = ~n5319 & n8167 ;
  assign n24799 = ~n24797 & n24798 ;
  assign n24800 = n23869 & ~n24799 ;
  assign n24801 = ~n22719 & n24800 ;
  assign n24802 = n21761 ^ n16826 ^ 1'b0 ;
  assign n24803 = ~n18829 & n24802 ;
  assign n24804 = n24803 ^ n15233 ^ n8348 ;
  assign n24805 = n2965 | n18231 ;
  assign n24809 = ~n4283 & n18661 ;
  assign n24806 = n7723 ^ x190 ^ 1'b0 ;
  assign n24807 = n10420 & n24806 ;
  assign n24808 = n13441 & n24807 ;
  assign n24810 = n24809 ^ n24808 ^ 1'b0 ;
  assign n24811 = n22982 ^ n557 ^ 1'b0 ;
  assign n24812 = n3264 | n11407 ;
  assign n24813 = n16165 | n24812 ;
  assign n24814 = x33 & n12653 ;
  assign n24815 = n24814 ^ n13353 ^ 1'b0 ;
  assign n24816 = ~n2950 & n18280 ;
  assign n24817 = n14502 ^ n9001 ^ n4269 ;
  assign n24818 = n24817 ^ n9566 ^ 1'b0 ;
  assign n24819 = n4366 & ~n24818 ;
  assign n24820 = n15027 ^ n10123 ^ 1'b0 ;
  assign n24821 = n5865 & ~n13249 ;
  assign n24822 = n24820 & ~n24821 ;
  assign n24823 = n3287 | n7538 ;
  assign n24824 = n1476 | n24823 ;
  assign n24825 = n12341 | n24824 ;
  assign n24826 = ~n1965 & n12900 ;
  assign n24827 = n4457 & n5003 ;
  assign n24828 = n24827 ^ n12635 ^ 1'b0 ;
  assign n24829 = n24828 ^ n13946 ^ 1'b0 ;
  assign n24830 = n24829 ^ n21428 ^ 1'b0 ;
  assign n24831 = n24531 ^ n5421 ^ 1'b0 ;
  assign n24832 = n14732 ^ n11995 ^ 1'b0 ;
  assign n24833 = n4137 & n24832 ;
  assign n24834 = n24833 ^ n11631 ^ n1760 ;
  assign n24835 = n12390 ^ n4633 ^ 1'b0 ;
  assign n24836 = n24835 ^ n3658 ^ 1'b0 ;
  assign n24837 = n24836 ^ n2692 ^ n845 ;
  assign n24838 = ( ~n4808 & n9023 ) | ( ~n4808 & n24837 ) | ( n9023 & n24837 ) ;
  assign n24839 = n14634 & ~n16157 ;
  assign n24840 = n791 & ~n11729 ;
  assign n24841 = n24840 ^ n10066 ^ 1'b0 ;
  assign n24842 = n21044 ^ n4585 ^ 1'b0 ;
  assign n24843 = ( n1151 & n3164 ) | ( n1151 & n3720 ) | ( n3164 & n3720 ) ;
  assign n24844 = n19135 & n24843 ;
  assign n24845 = n24844 ^ n2918 ^ 1'b0 ;
  assign n24846 = n2871 & n7908 ;
  assign n24847 = ( n1070 & n8951 ) | ( n1070 & n20480 ) | ( n8951 & n20480 ) ;
  assign n24848 = n10646 ^ n6434 ^ 1'b0 ;
  assign n24849 = ~n24847 & n24848 ;
  assign n24850 = ~n4290 & n24849 ;
  assign n24851 = n9045 & n16075 ;
  assign n24852 = n9569 & ~n20598 ;
  assign n24853 = n24852 ^ n21222 ^ 1'b0 ;
  assign n24854 = n24095 ^ n340 ^ 1'b0 ;
  assign n24855 = n10475 & ~n24854 ;
  assign n24856 = n4831 | n24855 ;
  assign n24857 = ~n3888 & n7695 ;
  assign n24858 = n24857 ^ n3504 ^ 1'b0 ;
  assign n24859 = ~n6001 & n24858 ;
  assign n24860 = ( ~n3090 & n4852 ) | ( ~n3090 & n24859 ) | ( n4852 & n24859 ) ;
  assign n24861 = n3087 | n24860 ;
  assign n24862 = n8114 | n24861 ;
  assign n24863 = n2532 & ~n24862 ;
  assign n24865 = n15444 ^ n15087 ^ n6701 ;
  assign n24866 = n24865 ^ n9058 ^ n6669 ;
  assign n24864 = x247 & n3230 ;
  assign n24867 = n24866 ^ n24864 ^ 1'b0 ;
  assign n24868 = n11986 | n22564 ;
  assign n24869 = n9155 & ~n24868 ;
  assign n24870 = n7731 ^ n3198 ^ 1'b0 ;
  assign n24871 = n19245 & n24870 ;
  assign n24872 = x74 & ~n2347 ;
  assign n24873 = n3090 & n24872 ;
  assign n24874 = n24873 ^ n11302 ^ 1'b0 ;
  assign n24875 = n10032 ^ n4046 ^ 1'b0 ;
  assign n24876 = ~n6167 & n24875 ;
  assign n24877 = n8069 & n9111 ;
  assign n24878 = ( ~n3777 & n10757 ) | ( ~n3777 & n11640 ) | ( n10757 & n11640 ) ;
  assign n24879 = n6964 ^ n1273 ^ 1'b0 ;
  assign n24880 = n14194 & ~n24879 ;
  assign n24881 = n24880 ^ n8959 ^ 1'b0 ;
  assign n24882 = ~n8014 & n24881 ;
  assign n24883 = n10908 & n24882 ;
  assign n24884 = n24883 ^ n2916 ^ 1'b0 ;
  assign n24885 = n24884 ^ n9432 ^ 1'b0 ;
  assign n24886 = n19263 & n20536 ;
  assign n24887 = n15045 ^ n4218 ^ 1'b0 ;
  assign n24888 = ~n8662 & n24887 ;
  assign n24889 = ( n9126 & ~n21746 ) | ( n9126 & n24888 ) | ( ~n21746 & n24888 ) ;
  assign n24890 = ( n2473 & n6234 ) | ( n2473 & ~n20968 ) | ( n6234 & ~n20968 ) ;
  assign n24891 = n8978 & n24890 ;
  assign n24892 = n24889 & n24891 ;
  assign n24893 = n4610 | n7278 ;
  assign n24894 = n24892 & ~n24893 ;
  assign n24895 = n17245 & n23043 ;
  assign n24896 = n24895 ^ n14325 ^ 1'b0 ;
  assign n24897 = ~n1005 & n16144 ;
  assign n24898 = ~n1868 & n24897 ;
  assign n24899 = ( n1584 & ~n5127 ) | ( n1584 & n14395 ) | ( ~n5127 & n14395 ) ;
  assign n24901 = n3088 & n3499 ;
  assign n24902 = n24901 ^ n13468 ^ 1'b0 ;
  assign n24900 = n439 | n8719 ;
  assign n24903 = n24902 ^ n24900 ^ n16758 ;
  assign n24904 = n22048 ^ n4593 ^ 1'b0 ;
  assign n24905 = n15063 & n24904 ;
  assign n24906 = ( n7194 & n16316 ) | ( n7194 & n21173 ) | ( n16316 & n21173 ) ;
  assign n24907 = n24906 ^ n18650 ^ 1'b0 ;
  assign n24908 = n24905 & ~n24907 ;
  assign n24909 = n5272 & n13157 ;
  assign n24910 = n4073 & ~n9684 ;
  assign n24911 = ~n7070 & n24910 ;
  assign n24912 = ( n7847 & n24909 ) | ( n7847 & n24911 ) | ( n24909 & n24911 ) ;
  assign n24913 = n20545 ^ n3504 ^ x101 ;
  assign n24914 = ( ~n7029 & n8317 ) | ( ~n7029 & n24913 ) | ( n8317 & n24913 ) ;
  assign n24915 = ~n10188 & n24914 ;
  assign n24916 = ~x238 & n24915 ;
  assign n24917 = n24916 ^ n14738 ^ 1'b0 ;
  assign n24919 = n677 | n9714 ;
  assign n24918 = n7481 | n15856 ;
  assign n24920 = n24919 ^ n24918 ^ n15262 ;
  assign n24921 = n8549 ^ n3556 ^ 1'b0 ;
  assign n24922 = ~n9775 & n24921 ;
  assign n24923 = n10854 & n24922 ;
  assign n24924 = n24923 ^ n6979 ^ 1'b0 ;
  assign n24925 = n399 | n5081 ;
  assign n24926 = n24925 ^ n13448 ^ 1'b0 ;
  assign n24928 = n3134 & ~n9316 ;
  assign n24929 = n24928 ^ n7196 ^ 1'b0 ;
  assign n24930 = n851 & n24929 ;
  assign n24931 = ( n2504 & ~n9316 ) | ( n2504 & n24930 ) | ( ~n9316 & n24930 ) ;
  assign n24927 = n3067 & ~n11039 ;
  assign n24932 = n24931 ^ n24927 ^ n21445 ;
  assign n24933 = n24926 & n24932 ;
  assign n24934 = ~n5719 & n24933 ;
  assign n24935 = ( ~n2378 & n14051 ) | ( ~n2378 & n16093 ) | ( n14051 & n16093 ) ;
  assign n24936 = x149 & n1783 ;
  assign n24937 = n1681 & n24936 ;
  assign n24940 = n3505 & ~n19629 ;
  assign n24938 = ~n8944 & n19638 ;
  assign n24939 = ~n23039 & n24938 ;
  assign n24941 = n24940 ^ n24939 ^ n7398 ;
  assign n24942 = n7277 & n20288 ;
  assign n24943 = ( n24937 & n24941 ) | ( n24937 & ~n24942 ) | ( n24941 & ~n24942 ) ;
  assign n24944 = n1636 | n5699 ;
  assign n24945 = n11596 | n24944 ;
  assign n24946 = n4524 & ~n13314 ;
  assign n24947 = n24946 ^ n16396 ^ 1'b0 ;
  assign n24948 = n24945 & ~n24947 ;
  assign n24949 = ( n3313 & n4018 ) | ( n3313 & n17095 ) | ( n4018 & n17095 ) ;
  assign n24950 = n22162 & n24949 ;
  assign n24951 = n23536 ^ n12429 ^ n548 ;
  assign n24952 = n8398 ^ n5149 ^ 1'b0 ;
  assign n24953 = n6030 & ~n7200 ;
  assign n24954 = n17336 & ~n24953 ;
  assign n24955 = ~n24952 & n24954 ;
  assign n24956 = ( n15546 & n15765 ) | ( n15546 & n18622 ) | ( n15765 & n18622 ) ;
  assign n24958 = n9431 ^ n3278 ^ 1'b0 ;
  assign n24957 = n5515 | n18434 ;
  assign n24959 = n24958 ^ n24957 ^ 1'b0 ;
  assign n24960 = n24275 ^ n3459 ^ 1'b0 ;
  assign n24961 = n9401 | n24960 ;
  assign n24962 = n12976 ^ n2359 ^ 1'b0 ;
  assign n24963 = n4830 & ~n24962 ;
  assign n24964 = n24963 ^ n16029 ^ 1'b0 ;
  assign n24965 = ~n17274 & n24964 ;
  assign n24966 = n6523 & ~n7255 ;
  assign n24967 = n363 | n6170 ;
  assign n24968 = ~n19048 & n24967 ;
  assign n24969 = n24966 & n24968 ;
  assign n24974 = n342 & n9513 ;
  assign n24975 = n24974 ^ n7303 ^ 1'b0 ;
  assign n24970 = n1049 | n19276 ;
  assign n24971 = n24970 ^ n5379 ^ 1'b0 ;
  assign n24972 = ( n5163 & ~n11425 ) | ( n5163 & n24971 ) | ( ~n11425 & n24971 ) ;
  assign n24973 = n24972 ^ n14343 ^ n7312 ;
  assign n24976 = n24975 ^ n24973 ^ n6873 ;
  assign n24977 = n20251 & ~n24976 ;
  assign n24978 = n19606 | n24977 ;
  assign n24979 = n10696 | n24978 ;
  assign n24980 = n24979 ^ n9483 ^ 1'b0 ;
  assign n24981 = n11261 & n13585 ;
  assign n24982 = n23413 & ~n24981 ;
  assign n24983 = ~n14973 & n23533 ;
  assign n24984 = ~n7624 & n11929 ;
  assign n24985 = n1415 & n24984 ;
  assign n24986 = n24985 ^ n24602 ^ n679 ;
  assign n24987 = n4818 & n24986 ;
  assign n24988 = n24987 ^ n11053 ^ 1'b0 ;
  assign n24989 = n23402 ^ n17170 ^ 1'b0 ;
  assign n24990 = n8178 | n24989 ;
  assign n24991 = ( n6147 & n11947 ) | ( n6147 & ~n24990 ) | ( n11947 & ~n24990 ) ;
  assign n24992 = n6463 ^ n5314 ^ 1'b0 ;
  assign n24993 = ( n4447 & ~n15986 ) | ( n4447 & n24992 ) | ( ~n15986 & n24992 ) ;
  assign n24994 = n8320 & n13494 ;
  assign n24995 = n24994 ^ n18980 ^ n7925 ;
  assign n24996 = ( n7527 & n12350 ) | ( n7527 & n24995 ) | ( n12350 & n24995 ) ;
  assign n24997 = n20572 & ~n24610 ;
  assign n24998 = n9484 ^ n1525 ^ 1'b0 ;
  assign n24999 = n24997 & ~n24998 ;
  assign n25000 = n3246 | n15806 ;
  assign n25001 = n24721 | n25000 ;
  assign n25002 = ~n11127 & n18796 ;
  assign n25003 = ~x110 & n25002 ;
  assign n25004 = n25003 ^ n22423 ^ n2870 ;
  assign n25008 = n4578 | n6694 ;
  assign n25009 = n5387 | n25008 ;
  assign n25005 = n13281 ^ x244 ^ 1'b0 ;
  assign n25006 = n25005 ^ n14517 ^ 1'b0 ;
  assign n25007 = n5453 & ~n25006 ;
  assign n25010 = n25009 ^ n25007 ^ 1'b0 ;
  assign n25011 = ~n5133 & n25010 ;
  assign n25012 = ( ~n2924 & n4881 ) | ( ~n2924 & n22067 ) | ( n4881 & n22067 ) ;
  assign n25013 = ~n3898 & n25012 ;
  assign n25014 = n15062 ^ n14324 ^ n2991 ;
  assign n25015 = n11908 | n25014 ;
  assign n25016 = n25015 ^ n10771 ^ 1'b0 ;
  assign n25017 = ( n8884 & n17043 ) | ( n8884 & n19810 ) | ( n17043 & n19810 ) ;
  assign n25018 = ~n1180 & n10961 ;
  assign n25019 = n4323 & n25018 ;
  assign n25020 = ~n1569 & n25019 ;
  assign n25021 = n25020 ^ n12366 ^ n5502 ;
  assign n25022 = n13676 ^ n1904 ^ 1'b0 ;
  assign n25023 = ~n11534 & n25022 ;
  assign n25024 = n9795 | n25023 ;
  assign n25025 = n11564 ^ x186 ^ 1'b0 ;
  assign n25026 = n25025 ^ n14965 ^ 1'b0 ;
  assign n25027 = n1553 & ~n25026 ;
  assign n25029 = n9755 ^ n2202 ^ 1'b0 ;
  assign n25028 = ( n10464 & n11569 ) | ( n10464 & n24217 ) | ( n11569 & n24217 ) ;
  assign n25030 = n25029 ^ n25028 ^ n4677 ;
  assign n25031 = ~n8516 & n15689 ;
  assign n25032 = n18798 & ~n21609 ;
  assign n25033 = n18622 & n25032 ;
  assign n25034 = n22945 ^ n4797 ^ 1'b0 ;
  assign n25035 = n1619 & ~n25034 ;
  assign n25036 = n25035 ^ n2789 ^ 1'b0 ;
  assign n25037 = n13988 ^ n6363 ^ 1'b0 ;
  assign n25038 = ~n11763 & n25037 ;
  assign n25039 = n7230 | n15869 ;
  assign n25040 = ~n5616 & n25039 ;
  assign n25041 = ~n25038 & n25040 ;
  assign n25042 = n24902 ^ n7359 ^ 1'b0 ;
  assign n25043 = n10052 | n24825 ;
  assign n25044 = n8368 & n9550 ;
  assign n25045 = n25044 ^ n3908 ^ 1'b0 ;
  assign n25046 = n19191 & n25045 ;
  assign n25047 = ~n9367 & n20030 ;
  assign n25048 = ~n10593 & n25047 ;
  assign n25049 = n10408 & ~n25048 ;
  assign n25050 = n25046 & n25049 ;
  assign n25051 = n1284 & ~n7997 ;
  assign n25052 = ~n5896 & n25051 ;
  assign n25053 = n12983 & ~n25052 ;
  assign n25054 = ~n21330 & n25053 ;
  assign n25055 = n12557 | n12642 ;
  assign n25056 = n2437 | n25055 ;
  assign n25057 = n25056 ^ n17579 ^ n14589 ;
  assign n25058 = n3473 ^ n2449 ^ 1'b0 ;
  assign n25059 = ~n11509 & n25058 ;
  assign n25060 = n21177 ^ n14493 ^ 1'b0 ;
  assign n25061 = n3088 & ~n25060 ;
  assign n25062 = ~n3398 & n25061 ;
  assign n25063 = ~n25059 & n25062 ;
  assign n25064 = n13756 | n18238 ;
  assign n25071 = n16351 ^ n9101 ^ n2281 ;
  assign n25066 = n10392 ^ n8152 ^ 1'b0 ;
  assign n25065 = n18294 & ~n21082 ;
  assign n25067 = n25066 ^ n25065 ^ 1'b0 ;
  assign n25068 = n5814 & ~n6644 ;
  assign n25069 = n25067 & n25068 ;
  assign n25070 = n5876 & ~n25069 ;
  assign n25072 = n25071 ^ n25070 ^ 1'b0 ;
  assign n25073 = ( n1884 & ~n10387 ) | ( n1884 & n10421 ) | ( ~n10387 & n10421 ) ;
  assign n25074 = n20823 ^ n20269 ^ 1'b0 ;
  assign n25075 = n6063 & n25074 ;
  assign n25076 = ~n11822 & n25075 ;
  assign n25077 = ~n8858 & n9592 ;
  assign n25078 = n1861 & ~n12950 ;
  assign n25079 = ~n7764 & n25078 ;
  assign n25080 = n11168 | n25079 ;
  assign n25081 = x189 | n25080 ;
  assign n25082 = ( ~n271 & n606 ) | ( ~n271 & n14833 ) | ( n606 & n14833 ) ;
  assign n25083 = n25082 ^ n2824 ^ 1'b0 ;
  assign n25084 = n19872 | n25083 ;
  assign n25085 = n18736 | n22724 ;
  assign n25086 = n3166 | n25085 ;
  assign n25087 = n21365 ^ n6139 ^ n6010 ;
  assign n25098 = n5517 | n10150 ;
  assign n25088 = n3734 ^ n509 ^ 1'b0 ;
  assign n25089 = n3911 & ~n25088 ;
  assign n25090 = n3647 | n7149 ;
  assign n25091 = n25090 ^ n593 ^ 1'b0 ;
  assign n25092 = n25089 & ~n25091 ;
  assign n25093 = ~n5230 & n25092 ;
  assign n25094 = n25093 ^ n19624 ^ n13687 ;
  assign n25095 = n14212 ^ n13769 ^ 1'b0 ;
  assign n25096 = n25094 & ~n25095 ;
  assign n25097 = ~n9796 & n25096 ;
  assign n25099 = n25098 ^ n25097 ^ 1'b0 ;
  assign n25100 = n25099 ^ n8523 ^ n3231 ;
  assign n25101 = n7435 | n12456 ;
  assign n25102 = n9196 | n25101 ;
  assign n25103 = n8378 ^ n4995 ^ 1'b0 ;
  assign n25104 = ~n16927 & n25103 ;
  assign n25105 = n20030 & n25104 ;
  assign n25108 = n10956 ^ n3447 ^ 1'b0 ;
  assign n25106 = n1947 & n8159 ;
  assign n25107 = ~n13404 & n25106 ;
  assign n25109 = n25108 ^ n25107 ^ 1'b0 ;
  assign n25110 = n14507 & n25109 ;
  assign n25111 = ~n25105 & n25110 ;
  assign n25112 = n921 & ~n25111 ;
  assign n25113 = n25112 ^ n7925 ^ 1'b0 ;
  assign n25114 = ( n6608 & n10956 ) | ( n6608 & n24466 ) | ( n10956 & n24466 ) ;
  assign n25115 = n19363 ^ n6371 ^ n5834 ;
  assign n25116 = n25115 ^ n6047 ^ 1'b0 ;
  assign n25117 = n4290 & n6005 ;
  assign n25118 = n25117 ^ n20127 ^ 1'b0 ;
  assign n25119 = n15578 ^ n1433 ^ n1160 ;
  assign n25120 = n5850 ^ n2135 ^ 1'b0 ;
  assign n25121 = n11422 & n23282 ;
  assign n25122 = n25120 & n25121 ;
  assign n25123 = n8465 ^ n5243 ^ 1'b0 ;
  assign n25124 = n25123 ^ n9115 ^ n817 ;
  assign n25125 = ~n4584 & n25124 ;
  assign n25126 = n5017 & n10256 ;
  assign n25127 = ~n6964 & n25126 ;
  assign n25128 = n5463 ^ n1903 ^ n674 ;
  assign n25129 = n3697 ^ n1941 ^ 1'b0 ;
  assign n25130 = n25129 ^ n14214 ^ 1'b0 ;
  assign n25131 = n353 & n4140 ;
  assign n25132 = n20582 | n25131 ;
  assign n25133 = x103 & n10333 ;
  assign n25134 = n25133 ^ n13768 ^ 1'b0 ;
  assign n25135 = ( n8117 & n12185 ) | ( n8117 & ~n25134 ) | ( n12185 & ~n25134 ) ;
  assign n25136 = n6865 ^ n441 ^ 1'b0 ;
  assign n25137 = ~n1521 & n25136 ;
  assign n25138 = n7766 & n25137 ;
  assign n25139 = ~n25135 & n25138 ;
  assign n25140 = n9355 & ~n12136 ;
  assign n25142 = n10141 | n18911 ;
  assign n25141 = ~n10534 & n14424 ;
  assign n25143 = n25142 ^ n25141 ^ 1'b0 ;
  assign n25144 = n25143 ^ n8416 ^ 1'b0 ;
  assign n25145 = n3404 & n25144 ;
  assign n25146 = n7690 ^ n5680 ^ n1635 ;
  assign n25147 = n11486 & n25146 ;
  assign n25148 = n9851 ^ n5451 ^ 1'b0 ;
  assign n25149 = ~n1909 & n25148 ;
  assign n25150 = n19506 ^ n16960 ^ 1'b0 ;
  assign n25151 = n25150 ^ n2192 ^ 1'b0 ;
  assign n25152 = n7254 & n25151 ;
  assign n25153 = n1343 | n6297 ;
  assign n25154 = n25125 ^ n11930 ^ n3485 ;
  assign n25155 = ~n9365 & n22348 ;
  assign n25156 = n25155 ^ n21815 ^ 1'b0 ;
  assign n25157 = n802 | n6871 ;
  assign n25158 = n25156 & ~n25157 ;
  assign n25159 = ~n2442 & n15696 ;
  assign n25160 = ~n5517 & n13555 ;
  assign n25161 = n15566 & n25160 ;
  assign n25162 = n25161 ^ n19695 ^ 1'b0 ;
  assign n25163 = n25159 & n25162 ;
  assign n25166 = n20325 ^ n14273 ^ 1'b0 ;
  assign n25167 = n8078 | n25166 ;
  assign n25164 = ( n10055 & ~n18004 ) | ( n10055 & n22611 ) | ( ~n18004 & n22611 ) ;
  assign n25165 = n25164 ^ n17854 ^ 1'b0 ;
  assign n25168 = n25167 ^ n25165 ^ 1'b0 ;
  assign n25169 = x65 & ~n25168 ;
  assign n25170 = n23161 ^ n7650 ^ n2022 ;
  assign n25171 = n1337 & ~n8913 ;
  assign n25172 = n13637 & ~n25171 ;
  assign n25173 = n25172 ^ n24039 ^ 1'b0 ;
  assign n25174 = x169 & n25173 ;
  assign n25175 = n25174 ^ n7327 ^ 1'b0 ;
  assign n25176 = n13921 & ~n25175 ;
  assign n25177 = n25176 ^ n10093 ^ 1'b0 ;
  assign n25178 = n17954 & ~n25177 ;
  assign n25179 = n25170 & n25178 ;
  assign n25180 = n1213 | n5927 ;
  assign n25181 = n25180 ^ n7185 ^ 1'b0 ;
  assign n25182 = ( n13195 & ~n22869 ) | ( n13195 & n25181 ) | ( ~n22869 & n25181 ) ;
  assign n25183 = n12846 ^ n1610 ^ 1'b0 ;
  assign n25184 = n9982 ^ n5042 ^ 1'b0 ;
  assign n25185 = n25183 & ~n25184 ;
  assign n25186 = ~n6698 & n22628 ;
  assign n25187 = ( n1932 & n13373 ) | ( n1932 & ~n25186 ) | ( n13373 & ~n25186 ) ;
  assign n25188 = n12348 ^ n1900 ^ 1'b0 ;
  assign n25189 = n10264 & ~n25188 ;
  assign n25190 = n1270 & n25189 ;
  assign n25191 = ~n25187 & n25190 ;
  assign n25192 = n1033 & n17122 ;
  assign n25193 = n25192 ^ n6801 ^ 1'b0 ;
  assign n25194 = n25193 ^ n11218 ^ n1619 ;
  assign n25195 = n4892 | n25194 ;
  assign n25196 = n2058 & n3720 ;
  assign n25197 = ~n11007 & n25196 ;
  assign n25198 = ~n7306 & n25197 ;
  assign n25199 = ( n1239 & n6384 ) | ( n1239 & n9883 ) | ( n6384 & n9883 ) ;
  assign n25200 = n25199 ^ n22593 ^ 1'b0 ;
  assign n25201 = n10673 & n25200 ;
  assign n25202 = n5905 ^ n2186 ^ 1'b0 ;
  assign n25203 = n25202 ^ n23573 ^ 1'b0 ;
  assign n25204 = n2739 | n25203 ;
  assign n25205 = n25204 ^ n2556 ^ 1'b0 ;
  assign n25206 = n25205 ^ n5975 ^ 1'b0 ;
  assign n25207 = n24150 & n25206 ;
  assign n25208 = ( n4081 & n6360 ) | ( n4081 & n14046 ) | ( n6360 & n14046 ) ;
  assign n25209 = n8101 ^ n3551 ^ 1'b0 ;
  assign n25210 = ( n3024 & n3421 ) | ( n3024 & n13343 ) | ( n3421 & n13343 ) ;
  assign n25211 = n17875 ^ n11713 ^ n2752 ;
  assign n25212 = n781 | n20517 ;
  assign n25213 = n25211 & ~n25212 ;
  assign n25214 = n25213 ^ n12420 ^ 1'b0 ;
  assign n25215 = n25210 & ~n25214 ;
  assign n25216 = n6884 | n25215 ;
  assign n25217 = n940 | n4330 ;
  assign n25218 = n25217 ^ n8163 ^ 1'b0 ;
  assign n25219 = n25218 ^ n10632 ^ 1'b0 ;
  assign n25220 = n818 | n8756 ;
  assign n25221 = n271 | n25220 ;
  assign n25222 = ~n1339 & n25221 ;
  assign n25223 = n18874 & n25222 ;
  assign n25224 = n17157 & n25223 ;
  assign n25225 = n9640 | n25224 ;
  assign n25226 = n25219 & ~n25225 ;
  assign n25227 = ~n8026 & n10316 ;
  assign n25228 = ~n4428 & n25227 ;
  assign n25229 = n25228 ^ n5876 ^ 1'b0 ;
  assign n25230 = ~n12696 & n22317 ;
  assign n25231 = ~n3422 & n25230 ;
  assign n25232 = ( n2475 & n3381 ) | ( n2475 & ~n5917 ) | ( n3381 & ~n5917 ) ;
  assign n25233 = n21449 & n25232 ;
  assign n25234 = ( n1284 & n16904 ) | ( n1284 & ~n24836 ) | ( n16904 & ~n24836 ) ;
  assign n25235 = ~n5639 & n22860 ;
  assign n25236 = n25235 ^ n21338 ^ n14000 ;
  assign n25237 = n15121 ^ n1049 ^ 1'b0 ;
  assign n25238 = ~n1364 & n25237 ;
  assign n25239 = n24376 ^ n2680 ^ 1'b0 ;
  assign n25240 = n25238 & ~n25239 ;
  assign n25241 = ~n14592 & n19317 ;
  assign n25242 = n25241 ^ n12519 ^ 1'b0 ;
  assign n25243 = n6403 | n9342 ;
  assign n25244 = n25243 ^ n12573 ^ 1'b0 ;
  assign n25245 = n25244 ^ n11370 ^ 1'b0 ;
  assign n25246 = n12554 ^ n10736 ^ 1'b0 ;
  assign n25247 = n24926 ^ n22018 ^ n2916 ;
  assign n25248 = ~n5895 & n8500 ;
  assign n25249 = n16128 ^ n10915 ^ 1'b0 ;
  assign n25250 = ~n4029 & n25249 ;
  assign n25251 = n306 & ~n8803 ;
  assign n25252 = ~n25250 & n25251 ;
  assign n25253 = n25252 ^ n7301 ^ 1'b0 ;
  assign n25254 = ~n7424 & n25253 ;
  assign n25255 = ( n1187 & n2569 ) | ( n1187 & n13359 ) | ( n2569 & n13359 ) ;
  assign n25256 = n11204 | n23001 ;
  assign n25257 = n21903 ^ n12153 ^ 1'b0 ;
  assign n25258 = n3253 | n3255 ;
  assign n25259 = n13565 ^ n7270 ^ 1'b0 ;
  assign n25260 = n14084 & n25259 ;
  assign n25261 = ~n18915 & n25260 ;
  assign n25262 = n25261 ^ x65 ^ 1'b0 ;
  assign n25263 = n5263 | n18910 ;
  assign n25264 = n25263 ^ n12008 ^ n2939 ;
  assign n25265 = n18089 ^ n3586 ^ 1'b0 ;
  assign n25266 = n3597 & n25265 ;
  assign n25267 = n18827 ^ n6739 ^ 1'b0 ;
  assign n25268 = n10322 & ~n25267 ;
  assign n25269 = n5243 | n9603 ;
  assign n25270 = n25269 ^ n21829 ^ n579 ;
  assign n25271 = ~n9030 & n11593 ;
  assign n25272 = n24381 & ~n25271 ;
  assign n25273 = n25272 ^ n8612 ^ 1'b0 ;
  assign n25274 = n14798 ^ n8673 ^ n6851 ;
  assign n25275 = n11591 & n25274 ;
  assign n25276 = n3325 & ~n25275 ;
  assign n25277 = n15219 & n25276 ;
  assign n25278 = n25277 ^ n19364 ^ 1'b0 ;
  assign n25279 = ~n18299 & n25278 ;
  assign n25280 = n23623 & n25279 ;
  assign n25281 = n6783 ^ n2173 ^ 1'b0 ;
  assign n25282 = n14595 & ~n25281 ;
  assign n25284 = n20382 ^ n6139 ^ x155 ;
  assign n25283 = n8488 | n10250 ;
  assign n25285 = n25284 ^ n25283 ^ 1'b0 ;
  assign n25286 = ~n3363 & n7910 ;
  assign n25287 = n5411 & n25286 ;
  assign n25288 = n8632 ^ n2428 ^ 1'b0 ;
  assign n25289 = ~n16567 & n25288 ;
  assign n25290 = n6257 ^ x95 ^ 1'b0 ;
  assign n25291 = ~n7194 & n25290 ;
  assign n25292 = n25291 ^ n19411 ^ n18429 ;
  assign n25293 = n25289 & ~n25292 ;
  assign n25294 = n9840 ^ n1458 ^ 1'b0 ;
  assign n25295 = n25294 ^ n17055 ^ 1'b0 ;
  assign n25296 = n16261 | n25295 ;
  assign n25297 = n1107 & ~n10718 ;
  assign n25298 = n25297 ^ n13748 ^ 1'b0 ;
  assign n25299 = n9639 ^ n4604 ^ 1'b0 ;
  assign n25300 = n25298 & n25299 ;
  assign n25301 = n25296 & ~n25300 ;
  assign n25302 = ( n441 & n2756 ) | ( n441 & ~n6605 ) | ( n2756 & ~n6605 ) ;
  assign n25303 = ( n10995 & ~n13780 ) | ( n10995 & n25302 ) | ( ~n13780 & n25302 ) ;
  assign n25304 = n8117 & n25303 ;
  assign n25305 = n7778 ^ n5956 ^ 1'b0 ;
  assign n25306 = ~n25304 & n25305 ;
  assign n25307 = n3176 & n25306 ;
  assign n25308 = ~n10724 & n25307 ;
  assign n25309 = n1829 | n6445 ;
  assign n25310 = n1504 | n25309 ;
  assign n25311 = n25310 ^ n1926 ^ 1'b0 ;
  assign n25312 = n15601 & n25311 ;
  assign n25316 = n4932 ^ n780 ^ 1'b0 ;
  assign n25317 = n10796 & n25316 ;
  assign n25318 = ~n2952 & n25317 ;
  assign n25313 = ~n7281 & n15098 ;
  assign n25314 = n16047 & n25313 ;
  assign n25315 = ( ~n11937 & n24150 ) | ( ~n11937 & n25314 ) | ( n24150 & n25314 ) ;
  assign n25319 = n25318 ^ n25315 ^ n11342 ;
  assign n25320 = n19572 ^ n17935 ^ n6128 ;
  assign n25321 = n22173 ^ n9978 ^ 1'b0 ;
  assign n25322 = n5649 & ~n7532 ;
  assign n25323 = n1288 & n1744 ;
  assign n25324 = n25323 ^ n13774 ^ 1'b0 ;
  assign n25325 = n17733 | n22680 ;
  assign n25326 = ~n13411 & n14214 ;
  assign n25327 = n5213 & n25326 ;
  assign n25328 = n25327 ^ n12329 ^ 1'b0 ;
  assign n25329 = n16855 ^ n806 ^ 1'b0 ;
  assign n25330 = n18468 & n25329 ;
  assign n25331 = n21928 ^ n7270 ^ 1'b0 ;
  assign n25332 = n6215 | n25331 ;
  assign n25333 = ( n3193 & ~n25330 ) | ( n3193 & n25332 ) | ( ~n25330 & n25332 ) ;
  assign n25334 = n20623 ^ n5638 ^ 1'b0 ;
  assign n25335 = n19336 ^ n4780 ^ 1'b0 ;
  assign n25336 = ( n4284 & ~n18803 ) | ( n4284 & n25335 ) | ( ~n18803 & n25335 ) ;
  assign n25337 = n17293 | n25167 ;
  assign n25338 = n25336 & ~n25337 ;
  assign n25339 = ( n3995 & n18315 ) | ( n3995 & ~n25338 ) | ( n18315 & ~n25338 ) ;
  assign n25340 = ( n2101 & n2794 ) | ( n2101 & ~n11595 ) | ( n2794 & ~n11595 ) ;
  assign n25341 = n3910 & ~n25340 ;
  assign n25342 = n502 & ~n10314 ;
  assign n25343 = n6529 ^ n1800 ^ n1407 ;
  assign n25344 = n17980 ^ n9942 ^ n1846 ;
  assign n25345 = ( n13829 & n25343 ) | ( n13829 & n25344 ) | ( n25343 & n25344 ) ;
  assign n25346 = ~n3919 & n17442 ;
  assign n25347 = n439 & n25346 ;
  assign n25348 = ( ~n11090 & n11201 ) | ( ~n11090 & n12366 ) | ( n11201 & n12366 ) ;
  assign n25350 = n4560 & ~n8209 ;
  assign n25351 = n16359 & n25350 ;
  assign n25352 = n3019 | n25351 ;
  assign n25353 = n18948 & ~n25352 ;
  assign n25349 = ~n11350 & n12734 ;
  assign n25354 = n25353 ^ n25349 ^ 1'b0 ;
  assign n25355 = n8343 & n12402 ;
  assign n25356 = n960 & n9224 ;
  assign n25357 = n11641 & n25356 ;
  assign n25358 = n25357 ^ n15486 ^ n1932 ;
  assign n25359 = n25355 | n25358 ;
  assign n25360 = n18719 ^ n9610 ^ 1'b0 ;
  assign n25361 = n25360 ^ n2074 ^ 1'b0 ;
  assign n25362 = n21379 & ~n25361 ;
  assign n25363 = ~n4349 & n6945 ;
  assign n25364 = n17772 & n25363 ;
  assign n25365 = n25364 ^ n5013 ^ 1'b0 ;
  assign n25366 = x128 & n5896 ;
  assign n25367 = n16985 & n25366 ;
  assign n25368 = n21761 ^ n9196 ^ n3469 ;
  assign n25369 = ( n1332 & n3702 ) | ( n1332 & ~n4354 ) | ( n3702 & ~n4354 ) ;
  assign n25370 = ( n7844 & n25368 ) | ( n7844 & n25369 ) | ( n25368 & n25369 ) ;
  assign n25371 = n7688 | n25370 ;
  assign n25372 = ( n23269 & n25367 ) | ( n23269 & ~n25371 ) | ( n25367 & ~n25371 ) ;
  assign n25373 = n582 & ~n23091 ;
  assign n25374 = n3543 & ~n11039 ;
  assign n25375 = n1203 & ~n25374 ;
  assign n25376 = n25375 ^ n3288 ^ 1'b0 ;
  assign n25377 = ~n7578 & n19680 ;
  assign n25378 = n25377 ^ n1458 ^ 1'b0 ;
  assign n25379 = n1246 | n18373 ;
  assign n25380 = n1651 & n18141 ;
  assign n25381 = n25379 & n25380 ;
  assign n25382 = n25381 ^ n14181 ^ n4836 ;
  assign n25383 = n6874 | n14796 ;
  assign n25384 = n3183 | n25383 ;
  assign n25385 = n13725 | n15010 ;
  assign n25386 = n12662 & ~n25385 ;
  assign n25387 = ( n15682 & n25384 ) | ( n15682 & n25386 ) | ( n25384 & n25386 ) ;
  assign n25388 = ( n8515 & ~n21434 ) | ( n8515 & n25387 ) | ( ~n21434 & n25387 ) ;
  assign n25389 = ~n4912 & n8878 ;
  assign n25390 = n25389 ^ n5710 ^ 1'b0 ;
  assign n25391 = n25390 ^ n10234 ^ 1'b0 ;
  assign n25392 = x48 & ~n25391 ;
  assign n25393 = n9816 & ~n13528 ;
  assign n25394 = n16814 & ~n25393 ;
  assign n25395 = n11069 & ~n11380 ;
  assign n25396 = n19285 ^ n9286 ^ 1'b0 ;
  assign n25397 = ( n2539 & n2890 ) | ( n2539 & ~n25396 ) | ( n2890 & ~n25396 ) ;
  assign n25398 = n2357 & n12877 ;
  assign n25399 = ~n12877 & n25398 ;
  assign n25400 = n25399 ^ n4460 ^ n4286 ;
  assign n25401 = n20061 ^ n9268 ^ 1'b0 ;
  assign n25402 = ~n25400 & n25401 ;
  assign n25403 = n15649 ^ n13036 ^ n3502 ;
  assign n25404 = n7209 & n8762 ;
  assign n25405 = n25403 & n25404 ;
  assign n25406 = n3821 ^ n1038 ^ n838 ;
  assign n25407 = n15030 | n25406 ;
  assign n25408 = n25407 ^ n274 ^ 1'b0 ;
  assign n25409 = ~n4340 & n11226 ;
  assign n25410 = n25409 ^ n9734 ^ 1'b0 ;
  assign n25411 = ( n5537 & n24483 ) | ( n5537 & n25410 ) | ( n24483 & n25410 ) ;
  assign n25412 = n7919 ^ n4309 ^ 1'b0 ;
  assign n25413 = n21392 ^ n7962 ^ 1'b0 ;
  assign n25414 = ( n3468 & n25412 ) | ( n3468 & ~n25413 ) | ( n25412 & ~n25413 ) ;
  assign n25415 = n19548 ^ n10941 ^ 1'b0 ;
  assign n25416 = n16192 & ~n25415 ;
  assign n25417 = n16477 & ~n17680 ;
  assign n25418 = n23756 & n25417 ;
  assign n25419 = n21764 ^ n10690 ^ 1'b0 ;
  assign n25422 = n1036 & ~n15876 ;
  assign n25420 = ( n3116 & n16292 ) | ( n3116 & n21868 ) | ( n16292 & n21868 ) ;
  assign n25421 = n21931 & ~n25420 ;
  assign n25423 = n25422 ^ n25421 ^ 1'b0 ;
  assign n25424 = ~n3048 & n4775 ;
  assign n25425 = n21993 ^ n10157 ^ 1'b0 ;
  assign n25426 = n8113 ^ n4726 ^ 1'b0 ;
  assign n25427 = ~n2547 & n25426 ;
  assign n25428 = n14951 & n25427 ;
  assign n25429 = ( n24050 & n25425 ) | ( n24050 & ~n25428 ) | ( n25425 & ~n25428 ) ;
  assign n25430 = n13523 ^ n13264 ^ 1'b0 ;
  assign n25431 = n19503 ^ n3021 ^ 1'b0 ;
  assign n25432 = n25431 ^ n13780 ^ 1'b0 ;
  assign n25433 = n2522 & ~n25432 ;
  assign n25434 = n7976 & ~n17529 ;
  assign n25435 = n25434 ^ n20467 ^ 1'b0 ;
  assign n25436 = ~n12090 & n25435 ;
  assign n25437 = n5295 | n25436 ;
  assign n25438 = n5131 & ~n6309 ;
  assign n25439 = n14502 & n25438 ;
  assign n25440 = n5389 & ~n7916 ;
  assign n25441 = n7370 | n25440 ;
  assign n25442 = n3899 | n25441 ;
  assign n25443 = n25439 & n25442 ;
  assign n25444 = n25443 ^ n15519 ^ 1'b0 ;
  assign n25445 = n16780 ^ n11675 ^ 1'b0 ;
  assign n25446 = n10417 | n25445 ;
  assign n25447 = n25446 ^ n18895 ^ n8293 ;
  assign n25448 = x165 | n3156 ;
  assign n25449 = n25448 ^ n571 ^ 1'b0 ;
  assign n25450 = n25449 ^ n6327 ^ 1'b0 ;
  assign n25451 = ( n4278 & n8549 ) | ( n4278 & ~n25450 ) | ( n8549 & ~n25450 ) ;
  assign n25452 = n8083 ^ x155 ^ 1'b0 ;
  assign n25453 = n25451 & ~n25452 ;
  assign n25455 = n17267 ^ n17204 ^ n1571 ;
  assign n25454 = n351 | n15413 ;
  assign n25456 = n25455 ^ n25454 ^ 1'b0 ;
  assign n25457 = n25456 ^ n16735 ^ 1'b0 ;
  assign n25458 = n4719 & ~n13859 ;
  assign n25459 = n25458 ^ n1703 ^ 1'b0 ;
  assign n25460 = n3332 ^ n978 ^ 1'b0 ;
  assign n25461 = n23912 | n25460 ;
  assign n25462 = n25461 ^ n8959 ^ 1'b0 ;
  assign n25463 = n13753 | n23495 ;
  assign n25464 = n25463 ^ n5384 ^ 1'b0 ;
  assign n25468 = n2281 ^ n1147 ^ 1'b0 ;
  assign n25469 = ~n4366 & n25468 ;
  assign n25470 = ~n6728 & n25469 ;
  assign n25471 = ~n7102 & n25470 ;
  assign n25465 = ~n13103 & n15555 ;
  assign n25466 = ~n17735 & n25465 ;
  assign n25467 = n13165 & n25466 ;
  assign n25472 = n25471 ^ n25467 ^ 1'b0 ;
  assign n25473 = n20300 & n25472 ;
  assign n25474 = n18477 & ~n25473 ;
  assign n25475 = ~n13752 & n14083 ;
  assign n25476 = n25475 ^ n9997 ^ 1'b0 ;
  assign n25477 = n25476 ^ n24860 ^ n10464 ;
  assign n25478 = n7396 & n11317 ;
  assign n25479 = ~x167 & n25478 ;
  assign n25480 = n20386 | n25479 ;
  assign n25481 = n25480 ^ n6196 ^ 1'b0 ;
  assign n25482 = n4926 | n23218 ;
  assign n25485 = n11929 ^ n7653 ^ 1'b0 ;
  assign n25486 = n17953 & n25485 ;
  assign n25483 = n18665 ^ n1473 ^ 1'b0 ;
  assign n25484 = n6548 | n25483 ;
  assign n25487 = n25486 ^ n25484 ^ 1'b0 ;
  assign n25492 = n11401 ^ n2504 ^ 1'b0 ;
  assign n25493 = n4711 & ~n25492 ;
  assign n25494 = n8447 ^ n6177 ^ n5255 ;
  assign n25495 = n11761 ^ n512 ^ 1'b0 ;
  assign n25496 = n25494 | n25495 ;
  assign n25497 = n25493 & ~n25496 ;
  assign n25498 = ( ~n9242 & n23276 ) | ( ~n9242 & n25497 ) | ( n23276 & n25497 ) ;
  assign n25488 = n7077 ^ n7070 ^ n616 ;
  assign n25489 = ~n768 & n13757 ;
  assign n25490 = n25489 ^ n5518 ^ 1'b0 ;
  assign n25491 = ~n25488 & n25490 ;
  assign n25499 = n25498 ^ n25491 ^ 1'b0 ;
  assign n25500 = n19449 & n21932 ;
  assign n25501 = ~n12024 & n25500 ;
  assign n25502 = n15387 & n22709 ;
  assign n25503 = n25502 ^ n6163 ^ 1'b0 ;
  assign n25510 = n4395 ^ n908 ^ 1'b0 ;
  assign n25504 = x76 & n5922 ;
  assign n25505 = n25504 ^ n7980 ^ 1'b0 ;
  assign n25506 = n13437 ^ n11112 ^ n9767 ;
  assign n25507 = ( ~n24354 & n25505 ) | ( ~n24354 & n25506 ) | ( n25505 & n25506 ) ;
  assign n25508 = n19217 | n25507 ;
  assign n25509 = n25508 ^ n1168 ^ 1'b0 ;
  assign n25511 = n25510 ^ n25509 ^ n17154 ;
  assign n25512 = n5448 ^ n2783 ^ 1'b0 ;
  assign n25513 = n12152 & ~n25512 ;
  assign n25514 = n25511 & n25513 ;
  assign n25515 = n1875 & n15836 ;
  assign n25516 = n7969 | n10045 ;
  assign n25517 = n3068 | n25516 ;
  assign n25518 = ~n14576 & n25517 ;
  assign n25519 = n25515 & n25518 ;
  assign n25520 = n1868 & ~n19471 ;
  assign n25521 = n25519 & n25520 ;
  assign n25522 = n6889 ^ n758 ^ 1'b0 ;
  assign n25523 = n25522 ^ n3998 ^ 1'b0 ;
  assign n25524 = n4818 & n25523 ;
  assign n25525 = n9501 | n25524 ;
  assign n25526 = n3687 & n12598 ;
  assign n25527 = ~n271 & n25526 ;
  assign n25528 = n21002 & ~n25527 ;
  assign n25529 = ~n16326 & n25528 ;
  assign n25530 = ~n4495 & n16077 ;
  assign n25531 = ~n7798 & n25530 ;
  assign n25532 = ~n5100 & n25531 ;
  assign n25533 = n6366 & n9346 ;
  assign n25534 = n22299 ^ n16124 ^ 1'b0 ;
  assign n25535 = n14471 & ~n25534 ;
  assign n25536 = n6156 & ~n21165 ;
  assign n25537 = n25536 ^ n18336 ^ 1'b0 ;
  assign n25538 = n926 & n20732 ;
  assign n25539 = ~n25537 & n25538 ;
  assign n25540 = n11425 ^ n7844 ^ 1'b0 ;
  assign n25541 = n13626 & ~n25540 ;
  assign n25542 = n7066 & n25541 ;
  assign n25543 = n25542 ^ n6372 ^ 1'b0 ;
  assign n25544 = n8704 & n17540 ;
  assign n25545 = n13877 ^ n599 ^ 1'b0 ;
  assign n25546 = n25545 ^ n3798 ^ 1'b0 ;
  assign n25547 = n5155 | n25546 ;
  assign n25550 = n20732 ^ n5750 ^ 1'b0 ;
  assign n25551 = n23111 & n25550 ;
  assign n25552 = ~n1551 & n25551 ;
  assign n25548 = n11287 ^ n8846 ^ 1'b0 ;
  assign n25549 = n9465 | n25548 ;
  assign n25553 = n25552 ^ n25549 ^ 1'b0 ;
  assign n25554 = n22063 ^ n10441 ^ 1'b0 ;
  assign n25555 = n6602 | n14773 ;
  assign n25556 = n20369 | n25555 ;
  assign n25557 = n9472 ^ n729 ^ 1'b0 ;
  assign n25558 = n10776 & n11281 ;
  assign n25559 = x82 & ~n25558 ;
  assign n25562 = n933 & ~n8122 ;
  assign n25563 = n3185 | n18819 ;
  assign n25564 = ~n5805 & n25563 ;
  assign n25565 = n25562 & n25564 ;
  assign n25560 = n6683 & ~n13202 ;
  assign n25561 = n2896 | n25560 ;
  assign n25566 = n25565 ^ n25561 ^ 1'b0 ;
  assign n25567 = n19549 ^ n6943 ^ 1'b0 ;
  assign n25568 = n25567 ^ n11344 ^ 1'b0 ;
  assign n25569 = n2445 | n6636 ;
  assign n25570 = n25569 ^ n4160 ^ 1'b0 ;
  assign n25571 = n25570 ^ n3601 ^ 1'b0 ;
  assign n25572 = ~n8411 & n25571 ;
  assign n25573 = n25572 ^ n13000 ^ n9579 ;
  assign n25574 = n14122 & n14951 ;
  assign n25575 = n19196 | n24080 ;
  assign n25576 = n13266 ^ n6440 ^ 1'b0 ;
  assign n25577 = n5408 & n20616 ;
  assign n25578 = ~n25576 & n25577 ;
  assign n25579 = n25578 ^ n2988 ^ 1'b0 ;
  assign n25580 = n1922 & ~n4719 ;
  assign n25581 = n25580 ^ n557 ^ 1'b0 ;
  assign n25582 = n10050 ^ n550 ^ 1'b0 ;
  assign n25583 = n25581 & ~n25582 ;
  assign n25584 = n25583 ^ n18573 ^ n14397 ;
  assign n25585 = n25584 ^ n11711 ^ n10720 ;
  assign n25586 = n12990 ^ n11144 ^ 1'b0 ;
  assign n25587 = n9810 & n23485 ;
  assign n25591 = ~n1024 & n6762 ;
  assign n25588 = n2988 & ~n5025 ;
  assign n25589 = n25588 ^ n6001 ^ 1'b0 ;
  assign n25590 = n2462 | n25589 ;
  assign n25592 = n25591 ^ n25590 ^ n9956 ;
  assign n25593 = ( n981 & n13552 ) | ( n981 & ~n20170 ) | ( n13552 & ~n20170 ) ;
  assign n25594 = ( ~x100 & n18518 ) | ( ~x100 & n25593 ) | ( n18518 & n25593 ) ;
  assign n25595 = n9583 & n16712 ;
  assign n25596 = n15474 ^ n10319 ^ 1'b0 ;
  assign n25597 = n25595 & n25596 ;
  assign n25598 = n7569 | n9780 ;
  assign n25599 = n25598 ^ n10160 ^ 1'b0 ;
  assign n25600 = n22101 ^ n6561 ^ 1'b0 ;
  assign n25601 = n20987 ^ n17707 ^ n14756 ;
  assign n25602 = n25601 ^ n1247 ^ 1'b0 ;
  assign n25603 = n7047 ^ n829 ^ 1'b0 ;
  assign n25604 = ~n22133 & n25603 ;
  assign n25605 = ~n9842 & n25604 ;
  assign n25606 = n25605 ^ n6625 ^ 1'b0 ;
  assign n25607 = n11191 & n14266 ;
  assign n25608 = n25607 ^ n9813 ^ 1'b0 ;
  assign n25609 = n6628 ^ n6323 ^ n2325 ;
  assign n25610 = n25609 ^ n18057 ^ n9347 ;
  assign n25611 = n5575 & n17884 ;
  assign n25612 = n25611 ^ n4560 ^ 1'b0 ;
  assign n25613 = ~n12590 & n25612 ;
  assign n25614 = ~n2101 & n21695 ;
  assign n25615 = n15717 & n25614 ;
  assign n25616 = ~n5255 & n21910 ;
  assign n25617 = n12108 ^ n7393 ^ 1'b0 ;
  assign n25618 = n6075 | n25617 ;
  assign n25619 = n25618 ^ n12758 ^ n6368 ;
  assign n25620 = ~n9923 & n22906 ;
  assign n25621 = ~n25619 & n25620 ;
  assign n25622 = ( n25615 & n25616 ) | ( n25615 & n25621 ) | ( n25616 & n25621 ) ;
  assign n25624 = n14016 ^ n7973 ^ n2087 ;
  assign n25625 = n25624 ^ x45 ^ 1'b0 ;
  assign n25626 = n4510 & n25625 ;
  assign n25627 = n16634 & n25626 ;
  assign n25623 = n15262 | n20542 ;
  assign n25628 = n25627 ^ n25623 ^ 1'b0 ;
  assign n25629 = n25622 | n25628 ;
  assign n25630 = n20497 ^ n14504 ^ 1'b0 ;
  assign n25631 = n4191 & n25630 ;
  assign n25632 = n2483 ^ n686 ^ 1'b0 ;
  assign n25633 = n25632 ^ n7488 ^ 1'b0 ;
  assign n25634 = n25631 & n25633 ;
  assign n25635 = ~n4470 & n18922 ;
  assign n25636 = n25635 ^ n9891 ^ 1'b0 ;
  assign n25637 = ( n1474 & ~n10539 ) | ( n1474 & n25636 ) | ( ~n10539 & n25636 ) ;
  assign n25638 = n5895 ^ x108 ^ 1'b0 ;
  assign n25639 = ( n4296 & n25637 ) | ( n4296 & n25638 ) | ( n25637 & n25638 ) ;
  assign n25640 = n5932 & ~n25093 ;
  assign n25641 = n7270 & n25640 ;
  assign n25642 = ~n10969 & n25641 ;
  assign n25643 = n15741 | n25642 ;
  assign n25644 = n4413 ^ n2778 ^ 1'b0 ;
  assign n25645 = n20026 | n25644 ;
  assign n25646 = n3115 ^ n2217 ^ 1'b0 ;
  assign n25647 = ~n19778 & n25646 ;
  assign n25648 = n4832 | n13589 ;
  assign n25649 = n13487 ^ n5415 ^ 1'b0 ;
  assign n25650 = n25649 ^ n15001 ^ 1'b0 ;
  assign n25651 = n25650 ^ n9201 ^ n8276 ;
  assign n25652 = ( ~n10262 & n20749 ) | ( ~n10262 & n25651 ) | ( n20749 & n25651 ) ;
  assign n25653 = ~n4538 & n5993 ;
  assign n25654 = n16307 ^ n824 ^ 1'b0 ;
  assign n25655 = n5549 | n25654 ;
  assign n25656 = ~n4002 & n14316 ;
  assign n25657 = ~n25655 & n25656 ;
  assign n25658 = ~n9885 & n12201 ;
  assign n25659 = n5956 & n25658 ;
  assign n25660 = n13383 ^ n4828 ^ 1'b0 ;
  assign n25661 = ~n1653 & n25660 ;
  assign n25662 = ~n13966 & n25661 ;
  assign n25663 = n5997 & n25662 ;
  assign n25664 = n25663 ^ n15311 ^ 1'b0 ;
  assign n25665 = ~n25659 & n25664 ;
  assign n25666 = ~n7167 & n14903 ;
  assign n25667 = n7029 | n25666 ;
  assign n25668 = n16316 ^ n13533 ^ 1'b0 ;
  assign n25669 = n2026 | n25668 ;
  assign n25670 = n8529 ^ n5531 ^ 1'b0 ;
  assign n25671 = n4351 | n25670 ;
  assign n25672 = ( n2697 & n25669 ) | ( n2697 & n25671 ) | ( n25669 & n25671 ) ;
  assign n25673 = n2277 & ~n23452 ;
  assign n25674 = ~n13932 & n25673 ;
  assign n25675 = n19946 & n25674 ;
  assign n25676 = n5208 ^ n3183 ^ 1'b0 ;
  assign n25677 = n10267 & n25676 ;
  assign n25678 = n14119 ^ n6331 ^ 1'b0 ;
  assign n25679 = n5115 & ~n25678 ;
  assign n25680 = n25679 ^ n25659 ^ 1'b0 ;
  assign n25681 = n9365 ^ n1212 ^ 1'b0 ;
  assign n25682 = ~n7604 & n11610 ;
  assign n25683 = n25682 ^ x126 ^ 1'b0 ;
  assign n25684 = ~n2149 & n9394 ;
  assign n25685 = n22664 & n25684 ;
  assign n25686 = n17104 ^ n10543 ^ 1'b0 ;
  assign n25687 = n13988 | n25686 ;
  assign n25688 = n25687 ^ n20984 ^ 1'b0 ;
  assign n25689 = ( ~n4615 & n25685 ) | ( ~n4615 & n25688 ) | ( n25685 & n25688 ) ;
  assign n25690 = ~n693 & n2544 ;
  assign n25691 = n25690 ^ n9383 ^ 1'b0 ;
  assign n25693 = n531 ^ x7 ^ 1'b0 ;
  assign n25694 = ~n12701 & n25693 ;
  assign n25695 = n19664 & n25694 ;
  assign n25696 = n15756 ^ n8858 ^ 1'b0 ;
  assign n25697 = n25695 & ~n25696 ;
  assign n25692 = ~n1733 & n4029 ;
  assign n25698 = n25697 ^ n25692 ^ 1'b0 ;
  assign n25699 = n6294 & n17106 ;
  assign n25700 = n25699 ^ n9586 ^ 1'b0 ;
  assign n25701 = n15953 ^ n4302 ^ 1'b0 ;
  assign n25702 = ~n13388 & n25701 ;
  assign n25703 = n17250 & n20233 ;
  assign n25704 = ~n8807 & n20161 ;
  assign n25705 = n25704 ^ n17631 ^ 1'b0 ;
  assign n25706 = n2998 ^ n2278 ^ 1'b0 ;
  assign n25707 = n7204 & n10744 ;
  assign n25708 = ~n7204 & n25707 ;
  assign n25709 = ( n17681 & n19275 ) | ( n17681 & n25708 ) | ( n19275 & n25708 ) ;
  assign n25710 = n16129 | n25709 ;
  assign n25711 = n25710 ^ n1779 ^ 1'b0 ;
  assign n25712 = n14663 ^ n5986 ^ 1'b0 ;
  assign n25713 = n13644 & ~n25712 ;
  assign n25714 = n20386 ^ n5296 ^ 1'b0 ;
  assign n25715 = n25713 & n25714 ;
  assign n25716 = n25715 ^ n24723 ^ 1'b0 ;
  assign n25717 = n627 & n1009 ;
  assign n25718 = n25717 ^ n1773 ^ 1'b0 ;
  assign n25719 = n25718 ^ n14486 ^ n2953 ;
  assign n25720 = n17515 ^ n10296 ^ 1'b0 ;
  assign n25721 = n15484 & ~n25720 ;
  assign n25722 = n4773 ^ n2441 ^ 1'b0 ;
  assign n25723 = n25722 ^ n19958 ^ 1'b0 ;
  assign n25724 = n17855 & ~n25173 ;
  assign n25725 = n6101 & ~n21365 ;
  assign n25726 = n9406 ^ n5515 ^ 1'b0 ;
  assign n25727 = n11521 | n25726 ;
  assign n25728 = n12579 ^ n3051 ^ 1'b0 ;
  assign n25730 = n16402 ^ n9901 ^ 1'b0 ;
  assign n25729 = ~n1717 & n8276 ;
  assign n25731 = n25730 ^ n25729 ^ 1'b0 ;
  assign n25732 = ( n3271 & n5354 ) | ( n3271 & ~n12681 ) | ( n5354 & ~n12681 ) ;
  assign n25733 = ~n1036 & n4722 ;
  assign n25734 = ~n1010 & n25733 ;
  assign n25735 = n25732 & ~n25734 ;
  assign n25736 = n23062 ^ n8156 ^ 1'b0 ;
  assign n25737 = n5801 | n6329 ;
  assign n25738 = ~n7508 & n19070 ;
  assign n25739 = n25737 & n25738 ;
  assign n25740 = n25203 | n25739 ;
  assign n25741 = n25740 ^ n24291 ^ 1'b0 ;
  assign n25742 = n397 & ~n11645 ;
  assign n25743 = n8461 ^ n3847 ^ 1'b0 ;
  assign n25744 = n1001 & ~n25743 ;
  assign n25745 = n25744 ^ n19681 ^ 1'b0 ;
  assign n25746 = n12140 ^ x89 ^ 1'b0 ;
  assign n25747 = n25697 & n25746 ;
  assign n25748 = n4161 ^ n2266 ^ 1'b0 ;
  assign n25749 = n4870 & ~n20893 ;
  assign n25750 = ~n25748 & n25749 ;
  assign n25751 = n25750 ^ n12920 ^ 1'b0 ;
  assign n25752 = n25747 & ~n25751 ;
  assign n25753 = ~n1585 & n7245 ;
  assign n25754 = ~n5067 & n17181 ;
  assign n25755 = ~n19552 & n25754 ;
  assign n25756 = n19960 | n25755 ;
  assign n25757 = n25756 ^ n25475 ^ 1'b0 ;
  assign n25758 = ( n13446 & n18164 ) | ( n13446 & n24067 ) | ( n18164 & n24067 ) ;
  assign n25759 = n25758 ^ n6312 ^ 1'b0 ;
  assign n25760 = n24605 ^ n11178 ^ 1'b0 ;
  assign n25761 = n809 & n25760 ;
  assign n25762 = ( ~x123 & n3473 ) | ( ~x123 & n25761 ) | ( n3473 & n25761 ) ;
  assign n25763 = n2230 & n16574 ;
  assign n25764 = ( ~n8090 & n11647 ) | ( ~n8090 & n23600 ) | ( n11647 & n23600 ) ;
  assign n25765 = ~n1620 & n3475 ;
  assign n25766 = n25765 ^ n17668 ^ 1'b0 ;
  assign n25767 = n25764 & n25766 ;
  assign n25768 = ( ~n9423 & n25763 ) | ( ~n9423 & n25767 ) | ( n25763 & n25767 ) ;
  assign n25769 = n21218 ^ n12241 ^ n2130 ;
  assign n25775 = ~n12130 & n17953 ;
  assign n25776 = n25775 ^ n10796 ^ 1'b0 ;
  assign n25770 = ~n645 & n4593 ;
  assign n25771 = n2728 & n25770 ;
  assign n25772 = n25771 ^ n10070 ^ 1'b0 ;
  assign n25773 = n20403 | n25772 ;
  assign n25774 = n20384 | n25773 ;
  assign n25777 = n25776 ^ n25774 ^ 1'b0 ;
  assign n25778 = ~n10709 & n18729 ;
  assign n25779 = ( ~n473 & n17861 ) | ( ~n473 & n25778 ) | ( n17861 & n25778 ) ;
  assign n25782 = n1805 | n15453 ;
  assign n25783 = n25782 ^ n15539 ^ 1'b0 ;
  assign n25780 = n10886 ^ n5422 ^ n513 ;
  assign n25781 = n5592 & ~n25780 ;
  assign n25784 = n25783 ^ n25781 ^ n16650 ;
  assign n25785 = ( n5628 & n13117 ) | ( n5628 & ~n25784 ) | ( n13117 & ~n25784 ) ;
  assign n25786 = n12087 | n14940 ;
  assign n25787 = n1989 ^ x104 ^ 1'b0 ;
  assign n25788 = n20226 ^ n4425 ^ 1'b0 ;
  assign n25789 = n11175 | n25788 ;
  assign n25791 = n15246 ^ n13870 ^ 1'b0 ;
  assign n25790 = n16172 & ~n19963 ;
  assign n25792 = n25791 ^ n25790 ^ 1'b0 ;
  assign n25793 = n25792 ^ n11686 ^ 1'b0 ;
  assign n25794 = n19011 & ~n25793 ;
  assign n25795 = n25093 ^ n11203 ^ n7447 ;
  assign n25796 = n9838 ^ x176 ^ 1'b0 ;
  assign n25797 = n11420 ^ n8064 ^ 1'b0 ;
  assign n25798 = n1758 & ~n25797 ;
  assign n25799 = n3275 ^ n2685 ^ 1'b0 ;
  assign n25800 = n10867 & n25799 ;
  assign n25801 = n25798 & n25800 ;
  assign n25802 = n25801 ^ n7044 ^ 1'b0 ;
  assign n25803 = n25802 ^ n12212 ^ n12068 ;
  assign n25804 = ( ~n11351 & n18119 ) | ( ~n11351 & n25803 ) | ( n18119 & n25803 ) ;
  assign n25805 = n17740 ^ n2486 ^ 1'b0 ;
  assign n25806 = n13763 ^ n8352 ^ n5067 ;
  assign n25807 = n25806 ^ n17297 ^ 1'b0 ;
  assign n25808 = n25807 ^ n19047 ^ 1'b0 ;
  assign n25809 = ~n21396 & n25808 ;
  assign n25810 = n2831 | n11794 ;
  assign n25814 = n19301 ^ n17114 ^ n5046 ;
  assign n25811 = n4007 & ~n18744 ;
  assign n25812 = n25811 ^ n2670 ^ 1'b0 ;
  assign n25813 = n10617 & ~n25812 ;
  assign n25815 = n25814 ^ n25813 ^ n14566 ;
  assign n25816 = n3579 & n7477 ;
  assign n25817 = n5982 | n9981 ;
  assign n25818 = n25817 ^ n20957 ^ 1'b0 ;
  assign n25819 = n2359 & n3061 ;
  assign n25820 = n13883 ^ n2739 ^ n1762 ;
  assign n25821 = n25820 ^ n11024 ^ n3680 ;
  assign n25822 = n23393 ^ n18719 ^ 1'b0 ;
  assign n25823 = n16579 ^ n5752 ^ 1'b0 ;
  assign n25824 = n21151 | n25823 ;
  assign n25825 = n4881 & ~n9956 ;
  assign n25826 = n25825 ^ n3052 ^ 1'b0 ;
  assign n25827 = n24149 ^ n6995 ^ 1'b0 ;
  assign n25828 = n984 & n25827 ;
  assign n25829 = ~n1715 & n19532 ;
  assign n25830 = ~n25828 & n25829 ;
  assign n25831 = ( n721 & n3797 ) | ( n721 & n4729 ) | ( n3797 & n4729 ) ;
  assign n25833 = n2511 | n8893 ;
  assign n25832 = n256 & n17243 ;
  assign n25834 = n25833 ^ n25832 ^ 1'b0 ;
  assign n25835 = n3531 & ~n7861 ;
  assign n25836 = n4108 | n9708 ;
  assign n25837 = n25835 | n25836 ;
  assign n25838 = n16623 | n25837 ;
  assign n25839 = n8323 | n9968 ;
  assign n25840 = n3973 & ~n25839 ;
  assign n25841 = n25840 ^ n2067 ^ 1'b0 ;
  assign n25842 = n3310 & ~n18579 ;
  assign n25843 = n3438 ^ n2640 ^ x4 ;
  assign n25844 = n13741 & n25843 ;
  assign n25845 = ( ~n19957 & n25842 ) | ( ~n19957 & n25844 ) | ( n25842 & n25844 ) ;
  assign n25848 = n3985 & n11969 ;
  assign n25849 = n25848 ^ n2921 ^ 1'b0 ;
  assign n25850 = n25849 ^ n13035 ^ 1'b0 ;
  assign n25851 = n3126 & ~n25850 ;
  assign n25846 = n16344 ^ n11755 ^ 1'b0 ;
  assign n25847 = n5017 & ~n25846 ;
  assign n25852 = n25851 ^ n25847 ^ x115 ;
  assign n25853 = n19408 | n24329 ;
  assign n25854 = n25852 & ~n25853 ;
  assign n25855 = n1976 | n12660 ;
  assign n25856 = n1055 & ~n6363 ;
  assign n25857 = n10975 | n21452 ;
  assign n25858 = ~n3673 & n10434 ;
  assign n25859 = ~n2871 & n25858 ;
  assign n25860 = n25859 ^ n6141 ^ 1'b0 ;
  assign n25861 = ~n9369 & n19079 ;
  assign n25862 = n14513 ^ n2548 ^ n997 ;
  assign n25863 = ( ~n9074 & n22972 ) | ( ~n9074 & n24035 ) | ( n22972 & n24035 ) ;
  assign n25864 = n9126 ^ n8000 ^ 1'b0 ;
  assign n25867 = n1907 & n21740 ;
  assign n25865 = n18440 ^ n1636 ^ 1'b0 ;
  assign n25866 = n7121 | n25865 ;
  assign n25868 = n25867 ^ n25866 ^ 1'b0 ;
  assign n25869 = n17849 ^ n982 ^ 1'b0 ;
  assign n25870 = ~n476 & n1575 ;
  assign n25871 = ~n13859 & n24870 ;
  assign n25872 = n25871 ^ n5680 ^ 1'b0 ;
  assign n25873 = ~n2084 & n8310 ;
  assign n25874 = n25873 ^ n6232 ^ 1'b0 ;
  assign n25875 = n3988 & ~n25874 ;
  assign n25876 = n1033 | n14566 ;
  assign n25877 = n25876 ^ n6778 ^ 1'b0 ;
  assign n25878 = n25877 ^ n11103 ^ n2113 ;
  assign n25880 = n3718 & ~n5311 ;
  assign n25881 = n25880 ^ n14269 ^ n5503 ;
  assign n25879 = n8478 & ~n15560 ;
  assign n25882 = n25881 ^ n25879 ^ 1'b0 ;
  assign n25883 = n2650 | n9555 ;
  assign n25884 = n5314 & ~n25883 ;
  assign n25885 = n13469 ^ n11167 ^ 1'b0 ;
  assign n25886 = n15355 & ~n15822 ;
  assign n25887 = n8136 | n14561 ;
  assign n25888 = x187 & n25887 ;
  assign n25889 = n884 & ~n1368 ;
  assign n25890 = ~n1328 & n25889 ;
  assign n25891 = n25890 ^ n19675 ^ 1'b0 ;
  assign n25892 = n4535 & n25891 ;
  assign n25893 = ~n5820 & n22351 ;
  assign n25897 = ( ~n3473 & n3989 ) | ( ~n3473 & n12720 ) | ( n3989 & n12720 ) ;
  assign n25894 = n1886 | n9435 ;
  assign n25895 = n25894 ^ n12850 ^ n2765 ;
  assign n25896 = ~n9726 & n25895 ;
  assign n25898 = n25897 ^ n25896 ^ n11009 ;
  assign n25899 = n20840 ^ n9816 ^ 1'b0 ;
  assign n25900 = n463 & n25899 ;
  assign n25901 = n8780 ^ n541 ^ 1'b0 ;
  assign n25902 = ~n11561 & n22992 ;
  assign n25903 = n25902 ^ n20230 ^ 1'b0 ;
  assign n25904 = n12818 ^ n7636 ^ 1'b0 ;
  assign n25905 = n7214 ^ n2548 ^ 1'b0 ;
  assign n25906 = n25905 ^ n300 ^ 1'b0 ;
  assign n25907 = n25906 ^ n18465 ^ 1'b0 ;
  assign n25908 = n13220 & ~n25907 ;
  assign n25909 = n11167 | n17323 ;
  assign n25910 = n23954 ^ n585 ^ 1'b0 ;
  assign n25911 = ~n25909 & n25910 ;
  assign n25912 = n13571 ^ n10891 ^ 1'b0 ;
  assign n25914 = n1062 & ~n3734 ;
  assign n25913 = n10885 & n11077 ;
  assign n25915 = n25914 ^ n25913 ^ 1'b0 ;
  assign n25916 = ~n7924 & n25915 ;
  assign n25917 = n25916 ^ n13866 ^ 1'b0 ;
  assign n25918 = n7559 ^ n4984 ^ 1'b0 ;
  assign n25919 = n23101 ^ n19996 ^ 1'b0 ;
  assign n25920 = ~n25918 & n25919 ;
  assign n25921 = n25920 ^ n10661 ^ 1'b0 ;
  assign n25922 = ~n6080 & n14113 ;
  assign n25923 = n25922 ^ n18665 ^ 1'b0 ;
  assign n25924 = n25811 ^ n9420 ^ 1'b0 ;
  assign n25925 = n14679 ^ n12060 ^ 1'b0 ;
  assign n25926 = n19627 & ~n25925 ;
  assign n25927 = n11568 ^ n3198 ^ 1'b0 ;
  assign n25928 = ~n10913 & n25927 ;
  assign n25929 = ~n5065 & n25928 ;
  assign n25930 = n790 & ~n25929 ;
  assign n25931 = ~n5043 & n25930 ;
  assign n25932 = n25931 ^ n2990 ^ 1'b0 ;
  assign n25933 = n8471 & ~n25932 ;
  assign n25934 = n25933 ^ n13948 ^ 1'b0 ;
  assign n25935 = n22626 ^ n9913 ^ n349 ;
  assign n25936 = n25935 ^ n12275 ^ n6267 ;
  assign n25937 = n25936 ^ n6273 ^ 1'b0 ;
  assign n25938 = ( n835 & n5100 ) | ( n835 & n18935 ) | ( n5100 & n18935 ) ;
  assign n25939 = n11252 ^ n296 ^ 1'b0 ;
  assign n25940 = n18951 & n25939 ;
  assign n25951 = n24354 ^ n15002 ^ n8187 ;
  assign n25944 = n12902 & n14673 ;
  assign n25941 = n15002 & ~n20864 ;
  assign n25942 = n25941 ^ n3468 ^ 1'b0 ;
  assign n25943 = n3946 | n25942 ;
  assign n25945 = n25944 ^ n25943 ^ 1'b0 ;
  assign n25946 = ~n5535 & n16712 ;
  assign n25947 = n25946 ^ n2095 ^ 1'b0 ;
  assign n25948 = n25947 ^ x201 ^ 1'b0 ;
  assign n25949 = n13088 & n25948 ;
  assign n25950 = n25945 & n25949 ;
  assign n25952 = n25951 ^ n25950 ^ 1'b0 ;
  assign n25953 = n25952 ^ n8603 ^ 1'b0 ;
  assign n25954 = n24340 ^ n11852 ^ 1'b0 ;
  assign n25955 = ~n25953 & n25954 ;
  assign n25956 = n4328 & n21218 ;
  assign n25957 = n4976 & n25956 ;
  assign n25958 = ~n1350 & n12754 ;
  assign n25959 = n9170 ^ n1195 ^ 1'b0 ;
  assign n25960 = n10256 & n25959 ;
  assign n25961 = n25960 ^ n5598 ^ 1'b0 ;
  assign n25962 = n17104 & ~n25961 ;
  assign n25963 = n3081 | n20143 ;
  assign n25964 = n6515 & ~n20057 ;
  assign n25965 = n25964 ^ n2005 ^ 1'b0 ;
  assign n25966 = ( n3696 & n25963 ) | ( n3696 & n25965 ) | ( n25963 & n25965 ) ;
  assign n25971 = ( n1574 & n2291 ) | ( n1574 & ~n25187 ) | ( n2291 & ~n25187 ) ;
  assign n25967 = n2582 | n20706 ;
  assign n25968 = n25967 ^ n5550 ^ 1'b0 ;
  assign n25969 = n6866 & n25968 ;
  assign n25970 = n25969 ^ n329 ^ 1'b0 ;
  assign n25972 = n25971 ^ n25970 ^ 1'b0 ;
  assign n25975 = ~n1755 & n10085 ;
  assign n25973 = n6455 & n19889 ;
  assign n25974 = n17772 & n25973 ;
  assign n25976 = n25975 ^ n25974 ^ 1'b0 ;
  assign n25977 = n11328 ^ n11133 ^ 1'b0 ;
  assign n25978 = n15749 ^ n7523 ^ 1'b0 ;
  assign n25979 = n13303 ^ n6327 ^ n1969 ;
  assign n25980 = ( n4463 & ~n24829 ) | ( n4463 & n25979 ) | ( ~n24829 & n25979 ) ;
  assign n25981 = n18003 ^ n14035 ^ 1'b0 ;
  assign n25982 = n1925 & n4292 ;
  assign n25983 = n21616 | n25982 ;
  assign n25984 = n5013 & ~n25983 ;
  assign n25985 = n14092 ^ n3676 ^ 1'b0 ;
  assign n25986 = n3152 & ~n20561 ;
  assign n25987 = n25986 ^ n10472 ^ 1'b0 ;
  assign n25988 = n4031 & ~n14331 ;
  assign n25989 = n25988 ^ n6770 ^ 1'b0 ;
  assign n25990 = n25989 ^ n5986 ^ 1'b0 ;
  assign n25991 = n25990 ^ n5068 ^ 1'b0 ;
  assign n25992 = n24518 ^ n3848 ^ 1'b0 ;
  assign n25993 = n1365 ^ n1049 ^ 1'b0 ;
  assign n25994 = ( n2080 & n2749 ) | ( n2080 & n12765 ) | ( n2749 & n12765 ) ;
  assign n25995 = ~n527 & n25994 ;
  assign n25996 = n25995 ^ n14981 ^ 1'b0 ;
  assign n25997 = n5375 | n25996 ;
  assign n25998 = n25993 & ~n25997 ;
  assign n26001 = n871 & n10348 ;
  assign n25999 = n3352 | n6981 ;
  assign n26000 = n10541 & ~n25999 ;
  assign n26002 = n26001 ^ n26000 ^ 1'b0 ;
  assign n26008 = ~n1455 & n1597 ;
  assign n26009 = ~n1597 & n26008 ;
  assign n26010 = n4213 & ~n26009 ;
  assign n26011 = n26009 & n26010 ;
  assign n26005 = n8252 ^ n6802 ^ 1'b0 ;
  assign n26006 = ~n4990 & n26005 ;
  assign n26007 = ~n22795 & n26006 ;
  assign n26003 = n16305 & n22419 ;
  assign n26004 = ~n16305 & n26003 ;
  assign n26012 = n26011 ^ n26007 ^ n26004 ;
  assign n26013 = n13475 ^ n7377 ^ n6745 ;
  assign n26014 = ~n10606 & n15276 ;
  assign n26015 = n26014 ^ x108 ^ 1'b0 ;
  assign n26016 = n20448 ^ n12102 ^ 1'b0 ;
  assign n26017 = n9874 ^ n781 ^ 1'b0 ;
  assign n26018 = n4939 & n17049 ;
  assign n26019 = n4283 & n8551 ;
  assign n26020 = ~n4173 & n26019 ;
  assign n26021 = n7004 & n10411 ;
  assign n26022 = n26021 ^ n10818 ^ 1'b0 ;
  assign n26023 = ~n14969 & n15756 ;
  assign n26024 = n6690 & n11469 ;
  assign n26025 = ~n5994 & n26024 ;
  assign n26026 = n15502 ^ n3606 ^ 1'b0 ;
  assign n26027 = n16006 & ~n26026 ;
  assign n26028 = n21584 ^ n3775 ^ 1'b0 ;
  assign n26029 = n8374 & ~n18006 ;
  assign n26030 = n13380 ^ n7367 ^ 1'b0 ;
  assign n26031 = ~n26029 & n26030 ;
  assign n26032 = n26031 ^ n3465 ^ 1'b0 ;
  assign n26033 = ~n13616 & n26032 ;
  assign n26034 = n14547 & ~n21607 ;
  assign n26035 = ~n8515 & n23414 ;
  assign n26036 = n18980 & ~n26035 ;
  assign n26037 = n3100 | n24975 ;
  assign n26038 = n6724 ^ n802 ^ 1'b0 ;
  assign n26039 = n26037 & ~n26038 ;
  assign n26040 = n9380 ^ n6302 ^ 1'b0 ;
  assign n26041 = ( n11171 & ~n26039 ) | ( n11171 & n26040 ) | ( ~n26039 & n26040 ) ;
  assign n26042 = n634 & n24594 ;
  assign n26043 = ~n13069 & n26042 ;
  assign n26044 = n4772 ^ n407 ^ 1'b0 ;
  assign n26045 = n11591 & ~n26044 ;
  assign n26046 = n26045 ^ n9513 ^ 1'b0 ;
  assign n26047 = n26046 ^ n11355 ^ n3639 ;
  assign n26048 = n6542 & n26047 ;
  assign n26049 = n26048 ^ n22863 ^ 1'b0 ;
  assign n26050 = ( ~n1806 & n2846 ) | ( ~n1806 & n3839 ) | ( n2846 & n3839 ) ;
  assign n26051 = n7387 ^ n1577 ^ 1'b0 ;
  assign n26052 = n1814 & ~n12959 ;
  assign n26053 = ~n4915 & n26052 ;
  assign n26054 = n3361 & n5151 ;
  assign n26055 = n26054 ^ n1525 ^ 1'b0 ;
  assign n26056 = n1590 | n26055 ;
  assign n26059 = ~n7314 & n12903 ;
  assign n26060 = n3848 & n26059 ;
  assign n26057 = n11960 ^ n7264 ^ 1'b0 ;
  assign n26058 = ~n13017 & n26057 ;
  assign n26061 = n26060 ^ n26058 ^ n22816 ;
  assign n26062 = n10750 ^ n2567 ^ 1'b0 ;
  assign n26063 = n19581 & n26062 ;
  assign n26064 = n24116 ^ n16732 ^ 1'b0 ;
  assign n26065 = n20834 ^ n14862 ^ 1'b0 ;
  assign n26066 = n759 | n14070 ;
  assign n26067 = ( n14262 & n17028 ) | ( n14262 & ~n23990 ) | ( n17028 & ~n23990 ) ;
  assign n26068 = n7431 & n8933 ;
  assign n26069 = n26068 ^ n8539 ^ 1'b0 ;
  assign n26070 = ( ~n20969 & n21385 ) | ( ~n20969 & n26069 ) | ( n21385 & n26069 ) ;
  assign n26071 = n1155 & ~n16597 ;
  assign n26072 = n26071 ^ n752 ^ 1'b0 ;
  assign n26073 = n14551 | n19242 ;
  assign n26074 = n9138 ^ n6424 ^ 1'b0 ;
  assign n26075 = n16361 | n26074 ;
  assign n26076 = n26075 ^ n23812 ^ 1'b0 ;
  assign n26077 = n1526 & ~n3150 ;
  assign n26078 = ( n5453 & ~n9359 ) | ( n5453 & n26077 ) | ( ~n9359 & n26077 ) ;
  assign n26083 = n4442 ^ n2612 ^ n1085 ;
  assign n26079 = n21050 ^ n1006 ^ 1'b0 ;
  assign n26080 = n7604 ^ n7342 ^ 1'b0 ;
  assign n26081 = n11143 | n26080 ;
  assign n26082 = n26079 | n26081 ;
  assign n26084 = n26083 ^ n26082 ^ 1'b0 ;
  assign n26085 = n16639 ^ n16515 ^ 1'b0 ;
  assign n26086 = n26084 & ~n26085 ;
  assign n26087 = ( n3215 & n6729 ) | ( n3215 & ~n24688 ) | ( n6729 & ~n24688 ) ;
  assign n26088 = n443 & ~n10010 ;
  assign n26089 = ~n9375 & n26088 ;
  assign n26090 = ~n9795 & n26089 ;
  assign n26091 = n26087 & n26090 ;
  assign n26092 = n4738 & n23912 ;
  assign n26093 = n11083 & ~n26092 ;
  assign n26095 = n14178 ^ n6992 ^ n4819 ;
  assign n26096 = n7424 | n23547 ;
  assign n26097 = ( n6606 & n26095 ) | ( n6606 & ~n26096 ) | ( n26095 & ~n26096 ) ;
  assign n26094 = n1106 | n16606 ;
  assign n26098 = n26097 ^ n26094 ^ 1'b0 ;
  assign n26099 = n860 & ~n2774 ;
  assign n26100 = n22976 & ~n26099 ;
  assign n26101 = n18103 | n26100 ;
  assign n26102 = n1615 & ~n5090 ;
  assign n26103 = x181 & n11850 ;
  assign n26104 = n6709 & n26103 ;
  assign n26105 = n26104 ^ n18912 ^ 1'b0 ;
  assign n26106 = ~n599 & n5542 ;
  assign n26107 = n5742 | n8998 ;
  assign n26108 = n26107 ^ n19944 ^ 1'b0 ;
  assign n26109 = n1453 ^ n1370 ^ 1'b0 ;
  assign n26110 = n10206 & ~n11719 ;
  assign n26111 = ~n3706 & n26110 ;
  assign n26112 = ( n3617 & ~n4704 ) | ( n3617 & n4715 ) | ( ~n4704 & n4715 ) ;
  assign n26113 = ~n26111 & n26112 ;
  assign n26114 = n26113 ^ n5498 ^ 1'b0 ;
  assign n26115 = n2411 | n14610 ;
  assign n26116 = n8729 | n26115 ;
  assign n26117 = ( ~n1300 & n9148 ) | ( ~n1300 & n19704 ) | ( n9148 & n19704 ) ;
  assign n26118 = n843 & ~n14452 ;
  assign n26119 = n26118 ^ n14905 ^ 1'b0 ;
  assign n26120 = ( n15881 & ~n19669 ) | ( n15881 & n26119 ) | ( ~n19669 & n26119 ) ;
  assign n26121 = n12503 & n26120 ;
  assign n26122 = n6734 | n16550 ;
  assign n26123 = ( n7843 & n10090 ) | ( n7843 & ~n26122 ) | ( n10090 & ~n26122 ) ;
  assign n26124 = ( n1500 & n5187 ) | ( n1500 & ~n6349 ) | ( n5187 & ~n6349 ) ;
  assign n26125 = n26124 ^ n14092 ^ n498 ;
  assign n26126 = x114 & ~n26125 ;
  assign n26127 = n26126 ^ n9420 ^ n3732 ;
  assign n26128 = n10660 ^ n459 ^ 1'b0 ;
  assign n26129 = n8183 & ~n26128 ;
  assign n26130 = n26129 ^ n23542 ^ n7333 ;
  assign n26133 = n6851 & ~n14708 ;
  assign n26131 = n3652 & n5690 ;
  assign n26132 = n26131 ^ n8487 ^ 1'b0 ;
  assign n26134 = n26133 ^ n26132 ^ 1'b0 ;
  assign n26135 = n9964 & ~n15536 ;
  assign n26136 = ~n12006 & n26135 ;
  assign n26137 = ~n3015 & n12271 ;
  assign n26138 = n26137 ^ n12201 ^ 1'b0 ;
  assign n26139 = n19020 & ~n26138 ;
  assign n26140 = n23512 & n26139 ;
  assign n26141 = ( n3147 & ~n9572 ) | ( n3147 & n18595 ) | ( ~n9572 & n18595 ) ;
  assign n26142 = ( n3701 & n13399 ) | ( n3701 & ~n26141 ) | ( n13399 & ~n26141 ) ;
  assign n26146 = n5098 ^ n2830 ^ 1'b0 ;
  assign n26143 = n20378 ^ n6760 ^ 1'b0 ;
  assign n26144 = n15985 & ~n26143 ;
  assign n26145 = ~n20551 & n26144 ;
  assign n26147 = n26146 ^ n26145 ^ 1'b0 ;
  assign n26148 = n4412 | n25014 ;
  assign n26149 = n26148 ^ n14930 ^ 1'b0 ;
  assign n26150 = ( n3947 & n6310 ) | ( n3947 & ~n6804 ) | ( n6310 & ~n6804 ) ;
  assign n26151 = n26150 ^ n20061 ^ n11575 ;
  assign n26152 = ~n10012 & n15869 ;
  assign n26153 = n26152 ^ n16619 ^ n4161 ;
  assign n26155 = ( n3273 & n5573 ) | ( n3273 & ~n8545 ) | ( n5573 & ~n8545 ) ;
  assign n26156 = n26155 ^ n10349 ^ 1'b0 ;
  assign n26157 = n3321 & ~n17614 ;
  assign n26158 = n26156 & n26157 ;
  assign n26154 = n14280 & n25987 ;
  assign n26159 = n26158 ^ n26154 ^ 1'b0 ;
  assign n26160 = x250 & ~n1064 ;
  assign n26161 = n26160 ^ n8511 ^ 1'b0 ;
  assign n26162 = n26161 ^ n18793 ^ 1'b0 ;
  assign n26163 = n9072 & n26162 ;
  assign n26164 = ~n7068 & n26163 ;
  assign n26165 = n26164 ^ n8728 ^ 1'b0 ;
  assign n26166 = n5514 & ~n10839 ;
  assign n26167 = ~n7765 & n12121 ;
  assign n26168 = ~n10491 & n26167 ;
  assign n26169 = n7105 ^ n1119 ^ 1'b0 ;
  assign n26170 = n1145 & ~n26169 ;
  assign n26171 = n26170 ^ n12142 ^ 1'b0 ;
  assign n26172 = ~n19320 & n26171 ;
  assign n26173 = n26168 & n26172 ;
  assign n26174 = n3169 & n9213 ;
  assign n26175 = n14706 & n22491 ;
  assign n26176 = ~n26174 & n26175 ;
  assign n26181 = n7097 & ~n18025 ;
  assign n26177 = n22940 ^ n19668 ^ 1'b0 ;
  assign n26178 = n18771 ^ n9070 ^ n2577 ;
  assign n26179 = n26178 ^ n15450 ^ n304 ;
  assign n26180 = n26177 & n26179 ;
  assign n26182 = n26181 ^ n26180 ^ 1'b0 ;
  assign n26183 = n3307 | n9759 ;
  assign n26184 = n26183 ^ n2580 ^ 1'b0 ;
  assign n26185 = n4826 | n26184 ;
  assign n26186 = n7137 | n26185 ;
  assign n26187 = n6093 & ~n26186 ;
  assign n26188 = n26187 ^ n18483 ^ 1'b0 ;
  assign n26189 = ~n14564 & n17259 ;
  assign n26203 = n7672 ^ n2707 ^ 1'b0 ;
  assign n26204 = n9786 | n26203 ;
  assign n26200 = n21481 ^ n4464 ^ n2529 ;
  assign n26201 = ~n10225 & n26200 ;
  assign n26202 = ( n9281 & n10943 ) | ( n9281 & n26201 ) | ( n10943 & n26201 ) ;
  assign n26205 = n26204 ^ n26202 ^ 1'b0 ;
  assign n26190 = ~n2426 & n7790 ;
  assign n26191 = n26190 ^ n8474 ^ 1'b0 ;
  assign n26192 = n26191 ^ n8527 ^ n467 ;
  assign n26193 = n3933 & ~n12266 ;
  assign n26194 = n8851 | n26193 ;
  assign n26195 = n7988 | n26194 ;
  assign n26196 = n26195 ^ n20691 ^ 1'b0 ;
  assign n26197 = n4848 | n26196 ;
  assign n26198 = n26192 & ~n26197 ;
  assign n26199 = n26198 ^ n12363 ^ 1'b0 ;
  assign n26206 = n26205 ^ n26199 ^ n8345 ;
  assign n26207 = n1270 & n25218 ;
  assign n26208 = n26207 ^ n21784 ^ n19814 ;
  assign n26209 = n7221 & n14023 ;
  assign n26210 = ~n11422 & n26209 ;
  assign n26211 = n26210 ^ n4686 ^ 1'b0 ;
  assign n26212 = n15910 ^ n6383 ^ 1'b0 ;
  assign n26213 = ( n19326 & ~n19759 ) | ( n19326 & n22719 ) | ( ~n19759 & n22719 ) ;
  assign n26214 = n5244 & ~n26213 ;
  assign n26215 = n26214 ^ n15428 ^ 1'b0 ;
  assign n26216 = n3814 | n13732 ;
  assign n26217 = n1225 | n6602 ;
  assign n26218 = ~n1932 & n10085 ;
  assign n26219 = n25800 & ~n26218 ;
  assign n26220 = n26219 ^ n2467 ^ 1'b0 ;
  assign n26221 = ( n12228 & n26217 ) | ( n12228 & n26220 ) | ( n26217 & n26220 ) ;
  assign n26222 = n5924 | n24267 ;
  assign n26223 = n8415 ^ n8393 ^ 1'b0 ;
  assign n26224 = n1421 & ~n26223 ;
  assign n26225 = n26224 ^ n5203 ^ 1'b0 ;
  assign n26226 = n8407 ^ n6877 ^ 1'b0 ;
  assign n26227 = ~n15320 & n26226 ;
  assign n26228 = n26227 ^ n16307 ^ n7549 ;
  assign n26229 = n19854 ^ n11865 ^ 1'b0 ;
  assign n26230 = ~n20403 & n26229 ;
  assign n26231 = ~n16793 & n24706 ;
  assign n26232 = x114 & n25522 ;
  assign n26233 = n26232 ^ n24836 ^ 1'b0 ;
  assign n26234 = n407 & ~n4924 ;
  assign n26235 = n26234 ^ n9311 ^ 1'b0 ;
  assign n26236 = n19929 | n26235 ;
  assign n26237 = n12994 | n26236 ;
  assign n26238 = ~n7661 & n18611 ;
  assign n26239 = n5590 & ~n26238 ;
  assign n26240 = ~n16705 & n18639 ;
  assign n26241 = n4462 & n26240 ;
  assign n26242 = ~n21089 & n24052 ;
  assign n26243 = ( n4359 & n20845 ) | ( n4359 & n21190 ) | ( n20845 & n21190 ) ;
  assign n26244 = ( n1626 & n3972 ) | ( n1626 & n26243 ) | ( n3972 & n26243 ) ;
  assign n26245 = n11895 ^ n2766 ^ 1'b0 ;
  assign n26246 = ( ~n2531 & n17154 ) | ( ~n2531 & n26245 ) | ( n17154 & n26245 ) ;
  assign n26248 = n304 & n4385 ;
  assign n26249 = n26248 ^ n6593 ^ 1'b0 ;
  assign n26247 = ( n258 & n4058 ) | ( n258 & ~n9571 ) | ( n4058 & ~n9571 ) ;
  assign n26250 = n26249 ^ n26247 ^ 1'b0 ;
  assign n26251 = x111 | n23297 ;
  assign n26252 = n26251 ^ n25120 ^ n17038 ;
  assign n26253 = n12597 & ~n25052 ;
  assign n26254 = n15164 ^ n11849 ^ 1'b0 ;
  assign n26255 = n21761 | n26254 ;
  assign n26256 = n19247 & ~n26255 ;
  assign n26257 = n9605 & ~n14286 ;
  assign n26258 = n18937 ^ n9644 ^ n500 ;
  assign n26259 = n6906 | n26258 ;
  assign n26260 = n26259 ^ n23630 ^ 1'b0 ;
  assign n26261 = n4114 | n26260 ;
  assign n26262 = n8620 & ~n16311 ;
  assign n26263 = n6089 & n26262 ;
  assign n26266 = ( x182 & ~n1403 ) | ( x182 & n3425 ) | ( ~n1403 & n3425 ) ;
  assign n26264 = n7364 ^ n4045 ^ 1'b0 ;
  assign n26265 = n5649 & n26264 ;
  assign n26267 = n26266 ^ n26265 ^ n9161 ;
  assign n26268 = n3068 & n19389 ;
  assign n26269 = n26268 ^ n9489 ^ 1'b0 ;
  assign n26270 = n7972 & n14750 ;
  assign n26271 = n11339 ^ n6215 ^ 1'b0 ;
  assign n26272 = n4363 ^ n1970 ^ 1'b0 ;
  assign n26273 = ~n17400 & n26272 ;
  assign n26274 = n26273 ^ n10419 ^ n365 ;
  assign n26275 = n13421 ^ n6748 ^ 1'b0 ;
  assign n26276 = n26274 & ~n26275 ;
  assign n26277 = ( ~n6053 & n17911 ) | ( ~n6053 & n26276 ) | ( n17911 & n26276 ) ;
  assign n26278 = ~n12749 & n23592 ;
  assign n26279 = ~n12080 & n26278 ;
  assign n26280 = n26279 ^ n6614 ^ 1'b0 ;
  assign n26281 = n381 | n8088 ;
  assign n26282 = n21524 & ~n26281 ;
  assign n26283 = n10085 & n26282 ;
  assign n26284 = n23990 & n26283 ;
  assign n26285 = x125 & n8587 ;
  assign n26286 = ~n6394 & n26285 ;
  assign n26287 = n4608 | n16363 ;
  assign n26288 = n23450 | n26287 ;
  assign n26289 = ( n8622 & n10300 ) | ( n8622 & n11448 ) | ( n10300 & n11448 ) ;
  assign n26290 = n10262 ^ n6565 ^ 1'b0 ;
  assign n26291 = n26289 & ~n26290 ;
  assign n26292 = n26291 ^ n23152 ^ 1'b0 ;
  assign n26293 = n18938 & ~n22454 ;
  assign n26294 = n23532 ^ n11483 ^ n8229 ;
  assign n26295 = ( n10374 & ~n26261 ) | ( n10374 & n26294 ) | ( ~n26261 & n26294 ) ;
  assign n26297 = n17504 ^ n3926 ^ 1'b0 ;
  assign n26298 = ( n2540 & ~n5389 ) | ( n2540 & n8251 ) | ( ~n5389 & n8251 ) ;
  assign n26299 = ~n14563 & n17200 ;
  assign n26300 = ~n16100 & n26299 ;
  assign n26301 = ( n9178 & n26298 ) | ( n9178 & n26300 ) | ( n26298 & n26300 ) ;
  assign n26302 = n26297 & ~n26301 ;
  assign n26296 = n14310 ^ n14184 ^ n6642 ;
  assign n26303 = n26302 ^ n26296 ^ n18884 ;
  assign n26304 = n2124 | n2277 ;
  assign n26305 = n10516 & ~n26304 ;
  assign n26306 = ~n7679 & n8509 ;
  assign n26307 = n26305 & n26306 ;
  assign n26308 = n652 & n1565 ;
  assign n26309 = n18888 ^ n15986 ^ n15676 ;
  assign n26310 = n26308 & n26309 ;
  assign n26311 = ~n2558 & n22228 ;
  assign n26312 = n13436 & n15721 ;
  assign n26313 = n26312 ^ n3332 ^ 1'b0 ;
  assign n26314 = n11593 ^ n9259 ^ n8367 ;
  assign n26315 = n26314 ^ n17182 ^ 1'b0 ;
  assign n26316 = n4698 | n11863 ;
  assign n26317 = n3401 & ~n6614 ;
  assign n26318 = ~n12635 & n26317 ;
  assign n26319 = n26316 | n26318 ;
  assign n26320 = ~n4064 & n5757 ;
  assign n26321 = ~n5294 & n15739 ;
  assign n26322 = ~n26320 & n26321 ;
  assign n26323 = n11142 ^ n8794 ^ n1626 ;
  assign n26324 = n10558 | n22959 ;
  assign n26325 = n26324 ^ x160 ^ 1'b0 ;
  assign n26326 = n14325 ^ n13917 ^ n10029 ;
  assign n26327 = n26326 ^ n25849 ^ 1'b0 ;
  assign n26328 = n4828 & ~n5209 ;
  assign n26329 = n26328 ^ n16379 ^ n10130 ;
  assign n26330 = n9170 & n9585 ;
  assign n26331 = ( x178 & n17722 ) | ( x178 & n26330 ) | ( n17722 & n26330 ) ;
  assign n26332 = n13083 ^ n569 ^ 1'b0 ;
  assign n26336 = ( ~n6725 & n9672 ) | ( ~n6725 & n17303 ) | ( n9672 & n17303 ) ;
  assign n26333 = n1757 | n2061 ;
  assign n26334 = n26333 ^ n2436 ^ 1'b0 ;
  assign n26335 = n19737 & n26334 ;
  assign n26337 = n26336 ^ n26335 ^ 1'b0 ;
  assign n26338 = n1255 & n15550 ;
  assign n26339 = n12190 ^ n5179 ^ 1'b0 ;
  assign n26340 = n26339 ^ n6092 ^ 1'b0 ;
  assign n26341 = n10425 ^ n9844 ^ 1'b0 ;
  assign n26342 = ~n26340 & n26341 ;
  assign n26343 = n3405 & n19258 ;
  assign n26344 = n20362 ^ n14158 ^ n1023 ;
  assign n26345 = n9797 ^ n9361 ^ 1'b0 ;
  assign n26346 = n23786 & n26345 ;
  assign n26347 = n1304 ^ n1291 ^ 1'b0 ;
  assign n26348 = ~n1729 & n26347 ;
  assign n26349 = n26348 ^ n13494 ^ 1'b0 ;
  assign n26350 = n5167 & n6375 ;
  assign n26351 = n17985 ^ n10621 ^ n4777 ;
  assign n26352 = n26351 ^ n7360 ^ 1'b0 ;
  assign n26353 = n26350 & n26352 ;
  assign n26354 = ( n16103 & n17053 ) | ( n16103 & n26353 ) | ( n17053 & n26353 ) ;
  assign n26355 = n16131 & n26354 ;
  assign n26356 = ~n2858 & n3727 ;
  assign n26357 = n26356 ^ n5001 ^ 1'b0 ;
  assign n26358 = ~n15433 & n16278 ;
  assign n26359 = n5778 | n26358 ;
  assign n26360 = n9159 ^ n546 ^ 1'b0 ;
  assign n26361 = ~n2054 & n26360 ;
  assign n26362 = ~n5687 & n26361 ;
  assign n26363 = n26362 ^ n10553 ^ 1'b0 ;
  assign n26364 = n26359 & ~n26363 ;
  assign n26365 = n17836 ^ n11153 ^ n620 ;
  assign n26367 = ~n6051 & n13088 ;
  assign n26366 = ~n12341 & n16810 ;
  assign n26368 = n26367 ^ n26366 ^ 1'b0 ;
  assign n26369 = ( n7237 & n9282 ) | ( n7237 & n26368 ) | ( n9282 & n26368 ) ;
  assign n26370 = n1307 & ~n9183 ;
  assign n26372 = n2942 | n5295 ;
  assign n26373 = n26372 ^ n18577 ^ 1'b0 ;
  assign n26374 = n6161 ^ x220 ^ 1'b0 ;
  assign n26375 = n25123 & n26374 ;
  assign n26376 = n26375 ^ n26161 ^ 1'b0 ;
  assign n26377 = n26373 & ~n26376 ;
  assign n26371 = n13775 & n18953 ;
  assign n26378 = n26377 ^ n26371 ^ 1'b0 ;
  assign n26379 = n9556 ^ n2169 ^ 1'b0 ;
  assign n26380 = n1166 | n26379 ;
  assign n26381 = n12438 ^ n7767 ^ 1'b0 ;
  assign n26382 = n26381 ^ n14967 ^ 1'b0 ;
  assign n26383 = n5361 & ~n17377 ;
  assign n26384 = n26383 ^ n9603 ^ n397 ;
  assign n26385 = n549 | n6069 ;
  assign n26386 = n549 & ~n26385 ;
  assign n26387 = n1733 | n26386 ;
  assign n26388 = n13471 & ~n26387 ;
  assign n26389 = n26388 ^ n19102 ^ n2393 ;
  assign n26390 = n19706 ^ n3053 ^ 1'b0 ;
  assign n26391 = n1892 & ~n3293 ;
  assign n26392 = n26391 ^ n4649 ^ 1'b0 ;
  assign n26393 = ~n16732 & n26392 ;
  assign n26394 = n3475 & ~n12388 ;
  assign n26395 = n26394 ^ n718 ^ 1'b0 ;
  assign n26396 = n26395 ^ n20229 ^ 1'b0 ;
  assign n26397 = n14940 & ~n26396 ;
  assign n26398 = n16667 ^ n13697 ^ 1'b0 ;
  assign n26399 = n26398 ^ n8415 ^ 1'b0 ;
  assign n26400 = n14251 ^ n9757 ^ 1'b0 ;
  assign n26401 = n9371 | n26400 ;
  assign n26402 = n5334 ^ n3487 ^ n1069 ;
  assign n26403 = x87 & ~n26007 ;
  assign n26404 = ~n14606 & n26403 ;
  assign n26405 = n4298 | n5684 ;
  assign n26406 = n26405 ^ n25765 ^ 1'b0 ;
  assign n26407 = n26404 | n26406 ;
  assign n26408 = ( n18115 & n26402 ) | ( n18115 & ~n26407 ) | ( n26402 & ~n26407 ) ;
  assign n26409 = n3664 | n11310 ;
  assign n26410 = ( n5203 & ~n23788 ) | ( n5203 & n26409 ) | ( ~n23788 & n26409 ) ;
  assign n26411 = n9589 | n26410 ;
  assign n26412 = n26218 ^ n4557 ^ 1'b0 ;
  assign n26413 = ( n3311 & ~n7629 ) | ( n3311 & n7934 ) | ( ~n7629 & n7934 ) ;
  assign n26414 = n26413 ^ n8179 ^ 1'b0 ;
  assign n26415 = n1795 | n13744 ;
  assign n26416 = n26415 ^ n6831 ^ 1'b0 ;
  assign n26417 = n15271 & ~n26416 ;
  assign n26418 = ~n19566 & n26417 ;
  assign n26419 = ~n18784 & n22927 ;
  assign n26420 = n18718 ^ n5690 ^ 1'b0 ;
  assign n26421 = n26395 & ~n26420 ;
  assign n26422 = n3947 | n16702 ;
  assign n26423 = n26422 ^ n22854 ^ 1'b0 ;
  assign n26426 = ( ~n7649 & n11089 ) | ( ~n7649 & n14018 ) | ( n11089 & n14018 ) ;
  assign n26424 = n7701 ^ n4719 ^ 1'b0 ;
  assign n26425 = n6616 & n26424 ;
  assign n26427 = n26426 ^ n26425 ^ n3239 ;
  assign n26428 = n26427 ^ n14187 ^ 1'b0 ;
  assign n26429 = n15532 ^ n8637 ^ 1'b0 ;
  assign n26430 = n322 | n5890 ;
  assign n26431 = n25843 | n26430 ;
  assign n26432 = n4595 & n11550 ;
  assign n26433 = ( ~n1919 & n5257 ) | ( ~n1919 & n9987 ) | ( n5257 & n9987 ) ;
  assign n26434 = ( n323 & n7239 ) | ( n323 & n26433 ) | ( n7239 & n26433 ) ;
  assign n26435 = ~n395 & n5582 ;
  assign n26436 = ( n25428 & n25522 ) | ( n25428 & n26435 ) | ( n25522 & n26435 ) ;
  assign n26437 = n4418 | n12344 ;
  assign n26438 = n7121 & ~n14909 ;
  assign n26439 = n1596 & ~n24244 ;
  assign n26440 = n4520 & ~n16183 ;
  assign n26441 = n26440 ^ n11376 ^ 1'b0 ;
  assign n26442 = n26441 ^ n1690 ^ 1'b0 ;
  assign n26443 = n18114 & n26442 ;
  assign n26444 = n26443 ^ n16371 ^ 1'b0 ;
  assign n26446 = ~n4447 & n13456 ;
  assign n26447 = n13287 ^ n11593 ^ 1'b0 ;
  assign n26448 = n26447 ^ n3913 ^ 1'b0 ;
  assign n26449 = n26446 & n26448 ;
  assign n26445 = n13094 & n16373 ;
  assign n26450 = n26449 ^ n26445 ^ 1'b0 ;
  assign n26451 = n20866 | n26450 ;
  assign n26452 = n26451 ^ n1234 ^ 1'b0 ;
  assign n26453 = n25816 ^ n9944 ^ 1'b0 ;
  assign n26454 = n14842 | n26453 ;
  assign n26456 = n1197 & n4925 ;
  assign n26455 = n20943 ^ n14602 ^ n1861 ;
  assign n26457 = n26456 ^ n26455 ^ 1'b0 ;
  assign n26458 = ~n6207 & n26457 ;
  assign n26459 = n26458 ^ n939 ^ 1'b0 ;
  assign n26460 = ~n7632 & n8808 ;
  assign n26461 = n26460 ^ n8201 ^ 1'b0 ;
  assign n26462 = n24688 ^ n18498 ^ n8892 ;
  assign n26463 = n26461 | n26462 ;
  assign n26464 = n6453 & n26463 ;
  assign n26470 = n11386 & ~n15462 ;
  assign n26471 = ~n11386 & n26470 ;
  assign n26469 = n429 & n9342 ;
  assign n26465 = n3809 & ~n8528 ;
  assign n26466 = n8528 & n26465 ;
  assign n26467 = n21755 & ~n26466 ;
  assign n26468 = ~n21755 & n26467 ;
  assign n26472 = n26471 ^ n26469 ^ n26468 ;
  assign n26473 = n7581 & ~n13885 ;
  assign n26474 = n8305 & n26473 ;
  assign n26475 = n8677 & ~n17142 ;
  assign n26476 = n11474 ^ n743 ^ 1'b0 ;
  assign n26477 = n7029 ^ n5532 ^ 1'b0 ;
  assign n26478 = n26477 ^ n13739 ^ 1'b0 ;
  assign n26479 = n5420 & ~n26478 ;
  assign n26480 = ~n9606 & n24862 ;
  assign n26481 = n13523 & n26480 ;
  assign n26485 = n7721 ^ n6593 ^ 1'b0 ;
  assign n26482 = n16639 ^ n8457 ^ 1'b0 ;
  assign n26483 = n19629 & n26482 ;
  assign n26484 = n2228 & n26483 ;
  assign n26486 = n26485 ^ n26484 ^ 1'b0 ;
  assign n26487 = n1993 | n17400 ;
  assign n26488 = n26487 ^ n4034 ^ 1'b0 ;
  assign n26489 = n26488 ^ n6892 ^ n5159 ;
  assign n26490 = n2759 & n8531 ;
  assign n26491 = n26490 ^ n5751 ^ 1'b0 ;
  assign n26493 = n8519 ^ n4956 ^ x17 ;
  assign n26492 = n6438 | n9621 ;
  assign n26494 = n26493 ^ n26492 ^ n12612 ;
  assign n26495 = ~n26491 & n26494 ;
  assign n26496 = n26495 ^ n12464 ^ 1'b0 ;
  assign n26497 = ~n26489 & n26496 ;
  assign n26498 = n8667 ^ n6009 ^ 1'b0 ;
  assign n26499 = n7973 & n14128 ;
  assign n26500 = ~n489 & n25991 ;
  assign n26501 = n14331 ^ n8266 ^ n4514 ;
  assign n26502 = ~n24587 & n26501 ;
  assign n26505 = n13220 ^ n7437 ^ 1'b0 ;
  assign n26504 = n12379 ^ n10560 ^ 1'b0 ;
  assign n26503 = n5713 ^ n374 ^ 1'b0 ;
  assign n26506 = n26505 ^ n26504 ^ n26503 ;
  assign n26507 = n1585 & n3421 ;
  assign n26508 = n26507 ^ n1468 ^ 1'b0 ;
  assign n26509 = n26508 ^ n11385 ^ n4346 ;
  assign n26510 = n19901 & ~n26509 ;
  assign n26511 = n26510 ^ n19957 ^ 1'b0 ;
  assign n26512 = n4859 & ~n5246 ;
  assign n26513 = ~n5083 & n16920 ;
  assign n26514 = n1365 & ~n3147 ;
  assign n26515 = n6805 & n10372 ;
  assign n26516 = n16756 & n26515 ;
  assign n26517 = ~n11915 & n13923 ;
  assign n26518 = n5820 | n15194 ;
  assign n26519 = n9008 | n14259 ;
  assign n26520 = n26518 & n26519 ;
  assign n26521 = n26520 ^ n13411 ^ 1'b0 ;
  assign n26522 = n3770 ^ n1054 ^ 1'b0 ;
  assign n26523 = ~n2950 & n26522 ;
  assign n26524 = n26523 ^ n9747 ^ n7051 ;
  assign n26525 = n4982 ^ n2571 ^ n538 ;
  assign n26526 = n4242 & n26525 ;
  assign n26527 = n26526 ^ n5181 ^ 1'b0 ;
  assign n26528 = ( n22314 & ~n26524 ) | ( n22314 & n26527 ) | ( ~n26524 & n26527 ) ;
  assign n26529 = ~n11834 & n16624 ;
  assign n26530 = ( n8578 & ~n20912 ) | ( n8578 & n26529 ) | ( ~n20912 & n26529 ) ;
  assign n26531 = ( ~n5768 & n9260 ) | ( ~n5768 & n11537 ) | ( n9260 & n11537 ) ;
  assign n26532 = n26531 ^ n15622 ^ 1'b0 ;
  assign n26533 = n1831 & n3274 ;
  assign n26534 = n17519 & n26533 ;
  assign n26535 = n26534 ^ n12546 ^ n2217 ;
  assign n26536 = n26532 | n26535 ;
  assign n26537 = n3362 & ~n26536 ;
  assign n26539 = ( ~n2248 & n7565 ) | ( ~n2248 & n8755 ) | ( n7565 & n8755 ) ;
  assign n26538 = ~n6630 & n6956 ;
  assign n26540 = n26539 ^ n26538 ^ 1'b0 ;
  assign n26541 = ~n1041 & n2253 ;
  assign n26542 = n15190 & n26541 ;
  assign n26543 = n26540 & n26542 ;
  assign n26547 = n1768 & ~n2580 ;
  assign n26548 = ~n4723 & n26547 ;
  assign n26549 = n13316 | n26548 ;
  assign n26550 = n13048 & ~n26549 ;
  assign n26544 = n17259 ^ n5565 ^ n1726 ;
  assign n26545 = n14176 ^ n12848 ^ 1'b0 ;
  assign n26546 = n26544 & n26545 ;
  assign n26551 = n26550 ^ n26546 ^ 1'b0 ;
  assign n26552 = ( n3842 & n24457 ) | ( n3842 & n25476 ) | ( n24457 & n25476 ) ;
  assign n26553 = n21429 ^ n3901 ^ 1'b0 ;
  assign n26554 = n5624 | n26459 ;
  assign n26555 = n3618 & ~n26554 ;
  assign n26564 = n4062 & n15682 ;
  assign n26565 = n26564 ^ n9656 ^ 1'b0 ;
  assign n26566 = n19929 | n26565 ;
  assign n26567 = n19746 & ~n26566 ;
  assign n26568 = n26567 ^ n16341 ^ 1'b0 ;
  assign n26556 = n9490 ^ n4739 ^ 1'b0 ;
  assign n26557 = n21850 ^ n13324 ^ 1'b0 ;
  assign n26558 = n26556 & ~n26557 ;
  assign n26559 = n6025 ^ n3477 ^ 1'b0 ;
  assign n26560 = n2651 & ~n19990 ;
  assign n26561 = n26559 & ~n26560 ;
  assign n26562 = ~n26558 & n26561 ;
  assign n26563 = n22689 & ~n26562 ;
  assign n26569 = n26568 ^ n26563 ^ 1'b0 ;
  assign n26570 = n1106 | n4487 ;
  assign n26571 = n26570 ^ n19187 ^ 1'b0 ;
  assign n26572 = ~n854 & n26571 ;
  assign n26574 = ( x72 & ~x238 ) | ( x72 & n729 ) | ( ~x238 & n729 ) ;
  assign n26575 = n11765 ^ n6997 ^ 1'b0 ;
  assign n26576 = ~n10996 & n26575 ;
  assign n26577 = ~n9459 & n26576 ;
  assign n26578 = ~n26574 & n26577 ;
  assign n26573 = ~n789 & n15756 ;
  assign n26579 = n26578 ^ n26573 ^ n19300 ;
  assign n26580 = n12247 | n26579 ;
  assign n26581 = n26580 ^ n23178 ^ 1'b0 ;
  assign n26582 = ~n22433 & n26581 ;
  assign n26583 = ( n10934 & n12548 ) | ( n10934 & ~n14229 ) | ( n12548 & ~n14229 ) ;
  assign n26584 = n4762 ^ x57 ^ 1'b0 ;
  assign n26585 = n23632 | n26584 ;
  assign n26586 = n12918 ^ n1042 ^ 1'b0 ;
  assign n26587 = n19303 | n26586 ;
  assign n26588 = ( n1553 & ~n13946 ) | ( n1553 & n18667 ) | ( ~n13946 & n18667 ) ;
  assign n26589 = n9529 | n26588 ;
  assign n26595 = n5507 | n12372 ;
  assign n26596 = ( n2942 & ~n5154 ) | ( n2942 & n26595 ) | ( ~n5154 & n26595 ) ;
  assign n26592 = n10361 ^ n8087 ^ 1'b0 ;
  assign n26593 = n4275 | n26592 ;
  assign n26591 = n6950 & ~n7941 ;
  assign n26590 = n20397 ^ n11074 ^ 1'b0 ;
  assign n26594 = n26593 ^ n26591 ^ n26590 ;
  assign n26597 = n26596 ^ n26594 ^ n1121 ;
  assign n26598 = n3169 & n7322 ;
  assign n26599 = n7141 & n26598 ;
  assign n26600 = ( x118 & ~n3568 ) | ( x118 & n4322 ) | ( ~n3568 & n4322 ) ;
  assign n26601 = ( n2844 & n3099 ) | ( n2844 & ~n18005 ) | ( n3099 & ~n18005 ) ;
  assign n26602 = n15951 ^ n11810 ^ 1'b0 ;
  assign n26603 = ( n14505 & n26601 ) | ( n14505 & n26602 ) | ( n26601 & n26602 ) ;
  assign n26604 = n328 | n26603 ;
  assign n26605 = n26604 ^ n16789 ^ n9822 ;
  assign n26606 = n2883 & n26605 ;
  assign n26607 = ~n8862 & n26606 ;
  assign n26608 = ~n26600 & n26607 ;
  assign n26609 = n1268 & ~n5305 ;
  assign n26610 = n1261 ^ n455 ^ 1'b0 ;
  assign n26611 = n26609 & n26610 ;
  assign n26612 = ( ~n2497 & n5162 ) | ( ~n2497 & n22181 ) | ( n5162 & n22181 ) ;
  assign n26613 = n18398 ^ n8046 ^ 1'b0 ;
  assign n26614 = n1708 | n26613 ;
  assign n26615 = n907 & ~n26614 ;
  assign n26616 = n6801 & n26615 ;
  assign n26619 = n1328 & ~n2463 ;
  assign n26618 = n2932 | n6528 ;
  assign n26620 = n26619 ^ n26618 ^ 1'b0 ;
  assign n26621 = ( n5147 & n11863 ) | ( n5147 & n26620 ) | ( n11863 & n26620 ) ;
  assign n26617 = n6372 & ~n22651 ;
  assign n26622 = n26621 ^ n26617 ^ 1'b0 ;
  assign n26623 = n26616 | n26622 ;
  assign n26624 = ( ~n21320 & n26612 ) | ( ~n21320 & n26623 ) | ( n26612 & n26623 ) ;
  assign n26625 = n13256 ^ n6443 ^ n1791 ;
  assign n26626 = n3391 | n6772 ;
  assign n26627 = n26626 ^ n20098 ^ 1'b0 ;
  assign n26628 = ~n10633 & n12340 ;
  assign n26629 = n26628 ^ n3985 ^ 1'b0 ;
  assign n26630 = n26629 ^ n10566 ^ n2315 ;
  assign n26631 = n23620 ^ n5052 ^ 1'b0 ;
  assign n26632 = n7138 & ~n16133 ;
  assign n26633 = n26632 ^ n10198 ^ 1'b0 ;
  assign n26634 = n8393 ^ n7067 ^ 1'b0 ;
  assign n26635 = x67 & ~n2649 ;
  assign n26636 = n26635 ^ n19105 ^ 1'b0 ;
  assign n26637 = n12041 | n16752 ;
  assign n26638 = n26636 | n26637 ;
  assign n26639 = ( x141 & n5356 ) | ( x141 & ~n8683 ) | ( n5356 & ~n8683 ) ;
  assign n26643 = ( n8968 & ~n9453 ) | ( n8968 & n16087 ) | ( ~n9453 & n16087 ) ;
  assign n26641 = ~n8041 & n8282 ;
  assign n26642 = n26641 ^ n5247 ^ 1'b0 ;
  assign n26640 = n4319 ^ n3215 ^ 1'b0 ;
  assign n26644 = n26643 ^ n26642 ^ n26640 ;
  assign n26645 = ~n833 & n19552 ;
  assign n26646 = n26645 ^ n1022 ^ 1'b0 ;
  assign n26647 = n24866 ^ n2066 ^ 1'b0 ;
  assign n26648 = n26646 & n26647 ;
  assign n26649 = n7976 | n15992 ;
  assign n26650 = n26649 ^ n5824 ^ 1'b0 ;
  assign n26651 = n26650 ^ n13923 ^ 1'b0 ;
  assign n26652 = ~n1358 & n3947 ;
  assign n26653 = ~n3374 & n26652 ;
  assign n26654 = ~n2281 & n26653 ;
  assign n26655 = n19070 ^ n11956 ^ 1'b0 ;
  assign n26658 = n3239 ^ n1880 ^ 1'b0 ;
  assign n26659 = x57 & ~n26658 ;
  assign n26656 = n3307 ^ n1235 ^ n381 ;
  assign n26657 = n17356 | n26656 ;
  assign n26660 = n26659 ^ n26657 ^ 1'b0 ;
  assign n26661 = n16510 & n26660 ;
  assign n26662 = n16211 & n26661 ;
  assign n26663 = n10309 ^ n2422 ^ 1'b0 ;
  assign n26664 = n2351 & n26663 ;
  assign n26665 = ~n4170 & n26664 ;
  assign n26666 = n11681 & n26665 ;
  assign n26667 = n26666 ^ n15534 ^ n7133 ;
  assign n26668 = n13678 | n24811 ;
  assign n26669 = n26667 | n26668 ;
  assign n26670 = n11308 & ~n26669 ;
  assign n26671 = n7552 | n9132 ;
  assign n26672 = n5420 & n26671 ;
  assign n26673 = n5400 ^ n3208 ^ n610 ;
  assign n26674 = n1241 & ~n5560 ;
  assign n26675 = n20618 & n26674 ;
  assign n26676 = n9740 & ~n10241 ;
  assign n26677 = ~n7246 & n26676 ;
  assign n26678 = ~n8226 & n13853 ;
  assign n26679 = n26678 ^ n4831 ^ 1'b0 ;
  assign n26681 = n21999 ^ n14233 ^ 1'b0 ;
  assign n26680 = x174 & n16561 ;
  assign n26682 = n26681 ^ n26680 ^ 1'b0 ;
  assign n26683 = n604 & ~n12135 ;
  assign n26684 = n5412 & ~n7822 ;
  assign n26685 = n26684 ^ n10127 ^ 1'b0 ;
  assign n26686 = n26683 & n26685 ;
  assign n26687 = n16775 ^ n1907 ^ 1'b0 ;
  assign n26693 = ~n4035 & n5092 ;
  assign n26694 = n26693 ^ n13254 ^ 1'b0 ;
  assign n26691 = n5868 & ~n18387 ;
  assign n26689 = ~n4552 & n4829 ;
  assign n26690 = n474 & n26689 ;
  assign n26692 = n26691 ^ n26690 ^ 1'b0 ;
  assign n26688 = n11778 & n12480 ;
  assign n26695 = n26694 ^ n26692 ^ n26688 ;
  assign n26696 = n10956 ^ n6432 ^ 1'b0 ;
  assign n26697 = n26696 ^ n11903 ^ 1'b0 ;
  assign n26698 = ( n7760 & n19854 ) | ( n7760 & ~n22559 ) | ( n19854 & ~n22559 ) ;
  assign n26699 = n26698 ^ n2611 ^ n1495 ;
  assign n26700 = n10867 ^ n1271 ^ 1'b0 ;
  assign n26701 = n9981 | n26700 ;
  assign n26702 = n26701 ^ n14711 ^ n10643 ;
  assign n26703 = ( n1346 & ~n6147 ) | ( n1346 & n9274 ) | ( ~n6147 & n9274 ) ;
  assign n26704 = ( n4703 & n15649 ) | ( n4703 & ~n26703 ) | ( n15649 & ~n26703 ) ;
  assign n26705 = n26704 ^ n8678 ^ 1'b0 ;
  assign n26706 = n640 | n26705 ;
  assign n26707 = n22926 | n26706 ;
  assign n26708 = ( n1115 & ~n26702 ) | ( n1115 & n26707 ) | ( ~n26702 & n26707 ) ;
  assign n26709 = ( n5460 & n8678 ) | ( n5460 & n10868 ) | ( n8678 & n10868 ) ;
  assign n26710 = ( n3751 & ~n8734 ) | ( n3751 & n26709 ) | ( ~n8734 & n26709 ) ;
  assign n26711 = n11382 ^ n11072 ^ 1'b0 ;
  assign n26712 = ~n21015 & n26711 ;
  assign n26713 = n7378 & ~n23590 ;
  assign n26714 = n26713 ^ n4638 ^ 1'b0 ;
  assign n26715 = n530 & n15930 ;
  assign n26716 = n1339 | n24168 ;
  assign n26717 = n23741 & ~n26716 ;
  assign n26718 = n14841 ^ n5582 ^ 1'b0 ;
  assign n26719 = n5433 & ~n26718 ;
  assign n26720 = n9502 ^ n9496 ^ 1'b0 ;
  assign n26721 = n2968 & n26720 ;
  assign n26731 = ~n1934 & n3257 ;
  assign n26732 = ~n3257 & n26731 ;
  assign n26730 = n791 & ~n26652 ;
  assign n26733 = n26732 ^ n26730 ^ 1'b0 ;
  assign n26722 = n9764 ^ n1795 ^ 1'b0 ;
  assign n26723 = n24136 & n26722 ;
  assign n26724 = n1418 & ~n11875 ;
  assign n26725 = ( n11726 & n20522 ) | ( n11726 & ~n26724 ) | ( n20522 & ~n26724 ) ;
  assign n26726 = ~n13340 & n26725 ;
  assign n26727 = ~n26725 & n26726 ;
  assign n26728 = n26723 & ~n26727 ;
  assign n26729 = ~n26723 & n26728 ;
  assign n26734 = n26733 ^ n26729 ^ n9222 ;
  assign n26735 = n1130 & n6202 ;
  assign n26736 = ~n4173 & n15752 ;
  assign n26737 = ~n11223 & n22470 ;
  assign n26738 = ~n14078 & n26737 ;
  assign n26739 = n19029 | n26718 ;
  assign n26740 = n26739 ^ n23812 ^ 1'b0 ;
  assign n26741 = n13249 | n26740 ;
  assign n26742 = n5468 & n26741 ;
  assign n26743 = n5592 ^ n1645 ^ 1'b0 ;
  assign n26744 = n7026 & n14719 ;
  assign n26745 = ( n21740 & ~n26743 ) | ( n21740 & n26744 ) | ( ~n26743 & n26744 ) ;
  assign n26746 = n14620 ^ n5667 ^ n5592 ;
  assign n26747 = n26746 ^ n17700 ^ n9247 ;
  assign n26748 = ( n6961 & ~n25637 ) | ( n6961 & n26595 ) | ( ~n25637 & n26595 ) ;
  assign n26749 = n18933 ^ n17450 ^ 1'b0 ;
  assign n26750 = n5641 & n14068 ;
  assign n26751 = n26750 ^ n8674 ^ 1'b0 ;
  assign n26752 = n26751 ^ n20099 ^ 1'b0 ;
  assign n26753 = n26749 | n26752 ;
  assign n26754 = n5621 & n7621 ;
  assign n26755 = n26754 ^ n23741 ^ 1'b0 ;
  assign n26756 = n7544 ^ x37 ^ 1'b0 ;
  assign n26757 = n21835 ^ n16791 ^ 1'b0 ;
  assign n26758 = x171 & n26757 ;
  assign n26759 = n26758 ^ n12171 ^ n11848 ;
  assign n26760 = n22262 ^ n10271 ^ 1'b0 ;
  assign n26761 = n8889 | n26760 ;
  assign n26762 = n20035 | n20453 ;
  assign n26763 = n26762 ^ n10851 ^ 1'b0 ;
  assign n26764 = ( ~n4626 & n6001 ) | ( ~n4626 & n9621 ) | ( n6001 & n9621 ) ;
  assign n26765 = n13009 & n26764 ;
  assign n26766 = n8487 & n26765 ;
  assign n26768 = n6215 & n14804 ;
  assign n26767 = ~n21172 & n22571 ;
  assign n26769 = n26768 ^ n26767 ^ 1'b0 ;
  assign n26770 = n6101 | n26769 ;
  assign n26771 = n7244 ^ n1819 ^ 1'b0 ;
  assign n26772 = n19774 | n26771 ;
  assign n26774 = n1264 | n4787 ;
  assign n26773 = n633 & ~n10497 ;
  assign n26775 = n26774 ^ n26773 ^ 1'b0 ;
  assign n26776 = ~n3417 & n14787 ;
  assign n26781 = n2131 | n20584 ;
  assign n26782 = n26781 ^ n5376 ^ 1'b0 ;
  assign n26783 = n11689 & n26782 ;
  assign n26784 = ~n860 & n26783 ;
  assign n26777 = ( n13043 & n15937 ) | ( n13043 & n17339 ) | ( n15937 & n17339 ) ;
  assign n26778 = n5681 & ~n26777 ;
  assign n26779 = n26778 ^ n24824 ^ 1'b0 ;
  assign n26780 = n9998 | n26779 ;
  assign n26785 = n26784 ^ n26780 ^ 1'b0 ;
  assign n26786 = ~n19658 & n25698 ;
  assign n26787 = ( n4746 & ~n6698 ) | ( n4746 & n10521 ) | ( ~n6698 & n10521 ) ;
  assign n26788 = n2046 & ~n6899 ;
  assign n26789 = n26788 ^ n1189 ^ 1'b0 ;
  assign n26790 = n26789 ^ n22722 ^ n13156 ;
  assign n26791 = n3147 | n7341 ;
  assign n26792 = n26791 ^ n25914 ^ 1'b0 ;
  assign n26793 = n7490 & n26792 ;
  assign n26794 = ( n26787 & ~n26790 ) | ( n26787 & n26793 ) | ( ~n26790 & n26793 ) ;
  assign n26795 = n26636 | n26794 ;
  assign n26796 = n3472 & n9287 ;
  assign n26797 = n10267 | n24953 ;
  assign n26798 = n13817 & n23192 ;
  assign n26799 = n21681 ^ n18616 ^ 1'b0 ;
  assign n26800 = ~n22573 & n26799 ;
  assign n26801 = ~n26798 & n26800 ;
  assign n26802 = n26801 ^ n22504 ^ 1'b0 ;
  assign n26804 = n3756 | n14203 ;
  assign n26805 = n26804 ^ n20671 ^ 1'b0 ;
  assign n26803 = ~n3523 & n24169 ;
  assign n26806 = n26805 ^ n26803 ^ 1'b0 ;
  assign n26807 = n19991 | n26806 ;
  assign n26808 = n20662 ^ n13090 ^ 1'b0 ;
  assign n26810 = n7982 | n26805 ;
  assign n26809 = n19581 ^ n10753 ^ n539 ;
  assign n26811 = n26810 ^ n26809 ^ 1'b0 ;
  assign n26812 = n22338 | n26811 ;
  assign n26816 = n4462 ^ n3316 ^ 1'b0 ;
  assign n26814 = n3596 ^ n2346 ^ 1'b0 ;
  assign n26813 = n8107 | n14043 ;
  assign n26815 = n26814 ^ n26813 ^ 1'b0 ;
  assign n26817 = n26816 ^ n26815 ^ n13453 ;
  assign n26818 = n25374 | n26817 ;
  assign n26819 = n22351 & ~n26818 ;
  assign n26820 = n21526 ^ n2252 ^ 1'b0 ;
  assign n26821 = n26273 ^ n9950 ^ 1'b0 ;
  assign n26822 = n14259 ^ n3958 ^ 1'b0 ;
  assign n26823 = n7710 | n26822 ;
  assign n26824 = n26821 & ~n26823 ;
  assign n26825 = n1733 & ~n11152 ;
  assign n26826 = ( n2392 & n26581 ) | ( n2392 & n26825 ) | ( n26581 & n26825 ) ;
  assign n26827 = n24623 ^ n1846 ^ 1'b0 ;
  assign n26828 = n20455 & n26827 ;
  assign n26829 = n6081 | n11418 ;
  assign n26830 = n15062 ^ n10921 ^ 1'b0 ;
  assign n26831 = n26829 | n26830 ;
  assign n26832 = n1829 & ~n17542 ;
  assign n26833 = ( n2547 & n4002 ) | ( n2547 & n18906 ) | ( n4002 & n18906 ) ;
  assign n26834 = n11490 ^ n8029 ^ n6469 ;
  assign n26835 = n2475 & n26834 ;
  assign n26836 = n3106 & n20373 ;
  assign n26837 = n1582 & n26836 ;
  assign n26838 = ~n7980 & n26837 ;
  assign n26839 = n14605 & n18937 ;
  assign n26840 = n26838 & n26839 ;
  assign n26841 = n3141 & n6095 ;
  assign n26842 = n10275 ^ n5400 ^ 1'b0 ;
  assign n26843 = n6484 & n26842 ;
  assign n26844 = ~n22934 & n26843 ;
  assign n26845 = n26844 ^ n7749 ^ 1'b0 ;
  assign n26846 = n7877 ^ n3778 ^ n1102 ;
  assign n26847 = n26846 ^ n6600 ^ 1'b0 ;
  assign n26848 = n23459 ^ n8105 ^ 1'b0 ;
  assign n26849 = n26848 ^ n9553 ^ 1'b0 ;
  assign n26850 = n12348 & n16491 ;
  assign n26851 = n26850 ^ n25679 ^ 1'b0 ;
  assign n26852 = n8791 ^ n581 ^ 1'b0 ;
  assign n26853 = n26852 ^ n20662 ^ 1'b0 ;
  assign n26854 = n18950 | n26853 ;
  assign n26855 = n26854 ^ n2921 ^ 1'b0 ;
  assign n26856 = ( n18774 & ~n26851 ) | ( n18774 & n26855 ) | ( ~n26851 & n26855 ) ;
  assign n26857 = ~n11461 & n20283 ;
  assign n26858 = ~n12666 & n26155 ;
  assign n26859 = n5067 ^ n2875 ^ 1'b0 ;
  assign n26860 = ~n3536 & n26859 ;
  assign n26861 = n25202 ^ n16386 ^ n5491 ;
  assign n26862 = n19456 & n21133 ;
  assign n26863 = n3551 & n22022 ;
  assign n26864 = n26863 ^ n17003 ^ 1'b0 ;
  assign n26865 = ~n2384 & n18559 ;
  assign n26866 = n13356 ^ n7806 ^ n7603 ;
  assign n26867 = ( n9398 & n26126 ) | ( n9398 & ~n26866 ) | ( n26126 & ~n26866 ) ;
  assign n26868 = n26867 ^ n23406 ^ 1'b0 ;
  assign n26869 = n17226 | n26868 ;
  assign n26870 = ~n12603 & n21457 ;
  assign n26871 = n6177 & n26870 ;
  assign n26872 = n7719 & ~n26871 ;
  assign n26873 = n2807 & n26872 ;
  assign n26874 = n3213 ^ x75 ^ 1'b0 ;
  assign n26875 = ~n6672 & n26874 ;
  assign n26876 = n3207 | n20284 ;
  assign n26877 = ~n7795 & n26876 ;
  assign n26878 = ~n26875 & n26877 ;
  assign n26879 = n15694 ^ n2970 ^ n1314 ;
  assign n26880 = ~n17644 & n26879 ;
  assign n26881 = ( n26873 & n26878 ) | ( n26873 & n26880 ) | ( n26878 & n26880 ) ;
  assign n26882 = n3291 | n5122 ;
  assign n26883 = n19758 | n26882 ;
  assign n26884 = n26883 ^ n8477 ^ n8402 ;
  assign n26885 = n25632 ^ n13040 ^ 1'b0 ;
  assign n26886 = n26884 & n26885 ;
  assign n26887 = n21449 ^ n12189 ^ n5536 ;
  assign n26888 = n26887 ^ n14046 ^ 1'b0 ;
  assign n26889 = n18688 ^ x196 ^ 1'b0 ;
  assign n26890 = n11015 & n26889 ;
  assign n26891 = n26888 & n26890 ;
  assign n26897 = n6284 & n7727 ;
  assign n26898 = ~n4537 & n26897 ;
  assign n26899 = n26898 ^ n18396 ^ 1'b0 ;
  assign n26895 = n22281 ^ n700 ^ 1'b0 ;
  assign n26896 = n11951 | n26895 ;
  assign n26900 = n26899 ^ n26896 ^ 1'b0 ;
  assign n26892 = ~n15298 & n26704 ;
  assign n26893 = n908 & n26892 ;
  assign n26894 = n19166 & ~n26893 ;
  assign n26901 = n26900 ^ n26894 ^ 1'b0 ;
  assign n26902 = n9508 & n11140 ;
  assign n26903 = n6537 & ~n25766 ;
  assign n26904 = n26903 ^ n3019 ^ 1'b0 ;
  assign n26908 = n10506 | n17007 ;
  assign n26909 = n9744 | n26908 ;
  assign n26910 = ~n25029 & n26909 ;
  assign n26911 = n26910 ^ n20611 ^ 1'b0 ;
  assign n26905 = n23336 | n26805 ;
  assign n26906 = n26905 ^ n429 ^ 1'b0 ;
  assign n26907 = n26906 ^ n4975 ^ 1'b0 ;
  assign n26912 = n26911 ^ n26907 ^ n13738 ;
  assign n26913 = n25609 | n26912 ;
  assign n26914 = n23815 & ~n26913 ;
  assign n26915 = n14113 ^ n361 ^ 1'b0 ;
  assign n26916 = n4068 ^ n2149 ^ 1'b0 ;
  assign n26917 = ~n20061 & n26916 ;
  assign n26918 = n8509 & n20870 ;
  assign n26919 = ~n26917 & n26918 ;
  assign n26920 = n11743 ^ n7554 ^ 1'b0 ;
  assign n26921 = n1535 & ~n1711 ;
  assign n26922 = n26921 ^ n17609 ^ 1'b0 ;
  assign n26923 = n26922 ^ n387 ^ 1'b0 ;
  assign n26924 = n15980 ^ n4471 ^ 1'b0 ;
  assign n26925 = n8522 | n26924 ;
  assign n26926 = n1809 & n4335 ;
  assign n26927 = ~n25146 & n26926 ;
  assign n26928 = n15630 & ~n16040 ;
  assign n26929 = n26928 ^ n5898 ^ 1'b0 ;
  assign n26930 = n1748 & n15642 ;
  assign n26931 = ( n543 & n5923 ) | ( n543 & n26930 ) | ( n5923 & n26930 ) ;
  assign n26932 = n8964 ^ n854 ^ 1'b0 ;
  assign n26933 = n18150 & n26932 ;
  assign n26934 = n11915 & ~n26933 ;
  assign n26935 = n26934 ^ n15093 ^ 1'b0 ;
  assign n26936 = ~n7211 & n26935 ;
  assign n26937 = ( n10090 & n17642 ) | ( n10090 & n26523 ) | ( n17642 & n26523 ) ;
  assign n26938 = n26937 ^ n14123 ^ 1'b0 ;
  assign n26939 = n6323 & n15137 ;
  assign n26940 = n16026 ^ n3275 ^ 1'b0 ;
  assign n26941 = n26939 & ~n26940 ;
  assign n26942 = ~n7703 & n16770 ;
  assign n26943 = n1247 & n7329 ;
  assign n26944 = n19370 ^ n5607 ^ 1'b0 ;
  assign n26945 = n26187 ^ n16575 ^ 1'b0 ;
  assign n26946 = n10621 & n26945 ;
  assign n26947 = ~n26944 & n26946 ;
  assign n26948 = ~n11607 & n15413 ;
  assign n26949 = n26948 ^ n26642 ^ 1'b0 ;
  assign n26951 = n1166 | n11398 ;
  assign n26952 = n18270 | n26951 ;
  assign n26953 = n26952 ^ n7508 ^ 1'b0 ;
  assign n26950 = n12130 ^ n7041 ^ 1'b0 ;
  assign n26954 = n26953 ^ n26950 ^ n22883 ;
  assign n26955 = n5931 ^ n836 ^ 1'b0 ;
  assign n26956 = ~n5133 & n26955 ;
  assign n26957 = n14150 & n26956 ;
  assign n26959 = n7185 ^ n6153 ^ n4148 ;
  assign n26958 = ~n3354 & n5691 ;
  assign n26960 = n26959 ^ n26958 ^ 1'b0 ;
  assign n26961 = n2777 | n10109 ;
  assign n26962 = n11454 ^ n7986 ^ 1'b0 ;
  assign n26963 = n26962 ^ n1041 ^ 1'b0 ;
  assign n26964 = n26961 | n26963 ;
  assign n26965 = n26964 ^ n11066 ^ 1'b0 ;
  assign n26966 = n9375 & ~n18723 ;
  assign n26967 = ~n18425 & n26966 ;
  assign n26968 = ~n6459 & n13305 ;
  assign n26969 = n26968 ^ n2663 ^ 1'b0 ;
  assign n26970 = x42 & ~n26969 ;
  assign n26971 = n26970 ^ n19736 ^ 1'b0 ;
  assign n26972 = n1680 & ~n4027 ;
  assign n26973 = n5841 | n26972 ;
  assign n26974 = n14914 & ~n17504 ;
  assign n26975 = n2470 & n5363 ;
  assign n26976 = n26975 ^ n1152 ^ 1'b0 ;
  assign n26977 = n26976 ^ n10169 ^ 1'b0 ;
  assign n26978 = n543 & ~n26977 ;
  assign n26979 = n8711 | n26137 ;
  assign n26980 = n4941 & ~n7781 ;
  assign n26981 = ( n4537 & n6285 ) | ( n4537 & n26980 ) | ( n6285 & n26980 ) ;
  assign n26982 = x54 & ~n9316 ;
  assign n26983 = ~n8710 & n26982 ;
  assign n26984 = n2221 & ~n2436 ;
  assign n26985 = n25533 ^ n13829 ^ n5370 ;
  assign n26986 = ( n13452 & ~n21832 ) | ( n13452 & n26529 ) | ( ~n21832 & n26529 ) ;
  assign n26987 = n26202 ^ n24252 ^ n3032 ;
  assign n26988 = n26073 & ~n26987 ;
  assign n26989 = n26988 ^ n7520 ^ 1'b0 ;
  assign n26991 = n3398 ^ n301 ^ 1'b0 ;
  assign n26992 = ~n19169 & n26991 ;
  assign n26990 = n18014 & ~n24544 ;
  assign n26993 = n26992 ^ n26990 ^ 1'b0 ;
  assign n26994 = ( n7327 & n15265 ) | ( n7327 & ~n15475 ) | ( n15265 & ~n15475 ) ;
  assign n26995 = n25753 ^ n836 ^ 1'b0 ;
  assign n26996 = n24343 ^ n755 ^ 1'b0 ;
  assign n26999 = n3568 & ~n6066 ;
  assign n26998 = ~n8956 & n12753 ;
  assign n27000 = n26999 ^ n26998 ^ 1'b0 ;
  assign n27001 = n6294 | n27000 ;
  assign n27002 = n27001 ^ n24923 ^ 1'b0 ;
  assign n27003 = n18807 & n27002 ;
  assign n26997 = n11929 ^ n1671 ^ 1'b0 ;
  assign n27004 = n27003 ^ n26997 ^ 1'b0 ;
  assign n27005 = n983 & ~n1641 ;
  assign n27006 = ( n976 & n4917 ) | ( n976 & n7033 ) | ( n4917 & n7033 ) ;
  assign n27007 = n8231 & n17374 ;
  assign n27008 = n5057 & n27007 ;
  assign n27009 = ( n9166 & n23007 ) | ( n9166 & n27008 ) | ( n23007 & n27008 ) ;
  assign n27010 = n16914 ^ n13543 ^ 1'b0 ;
  assign n27011 = ~n26620 & n27010 ;
  assign n27012 = ~n1930 & n10245 ;
  assign n27013 = ~n27011 & n27012 ;
  assign n27014 = x117 & n14201 ;
  assign n27015 = ~n14201 & n27014 ;
  assign n27016 = n15034 | n27015 ;
  assign n27017 = n27013 & ~n27016 ;
  assign n27018 = n3079 & n18166 ;
  assign n27019 = x123 | n15063 ;
  assign n27020 = n14212 ^ n10241 ^ n8446 ;
  assign n27021 = ~n27019 & n27020 ;
  assign n27022 = ~n668 & n27021 ;
  assign n27023 = n4339 & ~n12720 ;
  assign n27024 = n13506 ^ n1388 ^ 1'b0 ;
  assign n27025 = n3850 | n27024 ;
  assign n27026 = n27025 ^ n24570 ^ n6447 ;
  assign n27027 = n17808 & n19254 ;
  assign n27028 = n18723 ^ n1848 ^ n1612 ;
  assign n27029 = n4168 | n9751 ;
  assign n27030 = n7890 & ~n15586 ;
  assign n27031 = n27029 & n27030 ;
  assign n27032 = n27031 ^ n8096 ^ 1'b0 ;
  assign n27033 = ~n3554 & n10122 ;
  assign n27034 = n3489 & ~n27033 ;
  assign n27035 = n27034 ^ n1231 ^ 1'b0 ;
  assign n27036 = n5647 ^ n3453 ^ n1190 ;
  assign n27037 = n338 & ~n27036 ;
  assign n27038 = ( n1119 & ~n1469 ) | ( n1119 & n3453 ) | ( ~n1469 & n3453 ) ;
  assign n27039 = n4196 & n27038 ;
  assign n27040 = n3545 ^ n2437 ^ 1'b0 ;
  assign n27041 = ( n3668 & n12708 ) | ( n3668 & ~n17128 ) | ( n12708 & ~n17128 ) ;
  assign n27042 = n9366 & n27041 ;
  assign n27043 = n27040 & n27042 ;
  assign n27044 = n24021 & ~n27043 ;
  assign n27045 = n11923 & n27044 ;
  assign n27046 = n14102 | n27045 ;
  assign n27047 = n27046 ^ n19076 ^ 1'b0 ;
  assign n27048 = n6672 ^ n5824 ^ n4587 ;
  assign n27049 = n27048 ^ n18561 ^ n7167 ;
  assign n27050 = n27049 ^ n7859 ^ 1'b0 ;
  assign n27051 = ( ~n1411 & n8446 ) | ( ~n1411 & n15646 ) | ( n8446 & n15646 ) ;
  assign n27052 = n27051 ^ n16465 ^ n2794 ;
  assign n27053 = n27052 ^ n1106 ^ 1'b0 ;
  assign n27054 = n27053 ^ n25187 ^ n5014 ;
  assign n27058 = ~n17038 & n25210 ;
  assign n27055 = n12644 ^ n1625 ^ 1'b0 ;
  assign n27056 = ( n574 & n4160 ) | ( n574 & n27055 ) | ( n4160 & n27055 ) ;
  assign n27057 = n12399 | n27056 ;
  assign n27059 = n27058 ^ n27057 ^ 1'b0 ;
  assign n27060 = ~n4618 & n16234 ;
  assign n27061 = n10363 ^ n8425 ^ 1'b0 ;
  assign n27062 = n4194 & ~n27061 ;
  assign n27063 = n27062 ^ x14 ^ 1'b0 ;
  assign n27064 = n3045 & n5841 ;
  assign n27065 = n20623 ^ n14135 ^ 1'b0 ;
  assign n27066 = ~n23623 & n27065 ;
  assign n27067 = x146 & n25612 ;
  assign n27068 = ( n1026 & n10950 ) | ( n1026 & n27067 ) | ( n10950 & n27067 ) ;
  assign n27069 = n9220 | n27068 ;
  assign n27070 = ~n1173 & n8255 ;
  assign n27071 = n27070 ^ n3472 ^ 1'b0 ;
  assign n27072 = n14187 & n27071 ;
  assign n27073 = n2914 & ~n27072 ;
  assign n27074 = ~n7500 & n8942 ;
  assign n27075 = n10736 & n27074 ;
  assign n27076 = n298 | n2231 ;
  assign n27077 = n27075 & ~n27076 ;
  assign n27078 = n2459 ^ n1768 ^ 1'b0 ;
  assign n27079 = ~n1019 & n27078 ;
  assign n27080 = n14528 ^ n8544 ^ 1'b0 ;
  assign n27081 = n5497 ^ n3152 ^ 1'b0 ;
  assign n27082 = n9813 & n27081 ;
  assign n27083 = n16012 ^ n13533 ^ 1'b0 ;
  assign n27084 = n6898 & n17598 ;
  assign n27085 = n27084 ^ n9622 ^ 1'b0 ;
  assign n27086 = ~n18881 & n27085 ;
  assign n27087 = ~n2971 & n27086 ;
  assign n27088 = ( n1413 & n27083 ) | ( n1413 & ~n27087 ) | ( n27083 & ~n27087 ) ;
  assign n27089 = ~n6341 & n25636 ;
  assign n27090 = n27089 ^ n16172 ^ 1'b0 ;
  assign n27091 = n27090 ^ n11993 ^ n2560 ;
  assign n27092 = x57 & ~n11019 ;
  assign n27093 = n4953 & n27092 ;
  assign n27094 = n4764 & n19759 ;
  assign n27095 = n27094 ^ n1771 ^ 1'b0 ;
  assign n27096 = n3601 ^ n2146 ^ n908 ;
  assign n27097 = n7377 & ~n27096 ;
  assign n27098 = n12171 & n27097 ;
  assign n27099 = n27098 ^ n10081 ^ n980 ;
  assign n27100 = ~n27095 & n27099 ;
  assign n27101 = n12648 & ~n24606 ;
  assign n27102 = n27100 & n27101 ;
  assign n27103 = n17200 & n23326 ;
  assign n27104 = n19304 & n20567 ;
  assign n27105 = ~n6774 & n27104 ;
  assign n27106 = ~x166 & n6156 ;
  assign n27107 = ( n5997 & ~n19127 ) | ( n5997 & n27106 ) | ( ~n19127 & n27106 ) ;
  assign n27108 = n17597 ^ n16668 ^ 1'b0 ;
  assign n27109 = n6651 & n27108 ;
  assign n27111 = n5278 | n11755 ;
  assign n27112 = n11713 ^ n10574 ^ 1'b0 ;
  assign n27113 = n27111 & ~n27112 ;
  assign n27110 = n13015 & ~n20841 ;
  assign n27114 = n27113 ^ n27110 ^ 1'b0 ;
  assign n27115 = n2009 & ~n27114 ;
  assign n27116 = n18638 & n22014 ;
  assign n27117 = ~n8982 & n27116 ;
  assign n27118 = n19156 | n27117 ;
  assign n27119 = n9551 & ~n14537 ;
  assign n27120 = n19523 & n27119 ;
  assign n27121 = n6522 & n27120 ;
  assign n27122 = n10820 & ~n27121 ;
  assign n27125 = n2761 | n8369 ;
  assign n27126 = n27125 ^ n2247 ^ 1'b0 ;
  assign n27124 = n3249 & ~n18835 ;
  assign n27127 = n27126 ^ n27124 ^ 1'b0 ;
  assign n27123 = n2806 | n24711 ;
  assign n27128 = n27127 ^ n27123 ^ 1'b0 ;
  assign n27129 = ( ~n2916 & n4563 ) | ( ~n2916 & n4654 ) | ( n4563 & n4654 ) ;
  assign n27130 = n4432 ^ n1605 ^ 1'b0 ;
  assign n27131 = ~n11705 & n27130 ;
  assign n27132 = n12510 | n27131 ;
  assign n27133 = n16189 ^ n11511 ^ n5096 ;
  assign n27134 = n7296 & ~n14949 ;
  assign n27135 = n1897 | n9324 ;
  assign n27136 = n27135 ^ n18720 ^ 1'b0 ;
  assign n27137 = n26619 & ~n27136 ;
  assign n27138 = ( n27133 & n27134 ) | ( n27133 & ~n27137 ) | ( n27134 & ~n27137 ) ;
  assign n27139 = n17892 ^ n8386 ^ n7687 ;
  assign n27141 = n6484 & ~n10516 ;
  assign n27142 = n27141 ^ n6887 ^ 1'b0 ;
  assign n27143 = n21173 ^ n3328 ^ 1'b0 ;
  assign n27144 = n12140 & ~n27143 ;
  assign n27145 = n27142 | n27144 ;
  assign n27140 = n7437 ^ n3829 ^ 1'b0 ;
  assign n27146 = n27145 ^ n27140 ^ 1'b0 ;
  assign n27147 = n20651 ^ n16185 ^ 1'b0 ;
  assign n27148 = n12755 & n15723 ;
  assign n27149 = n27147 & n27148 ;
  assign n27150 = n7312 & n26259 ;
  assign n27151 = n8959 | n17151 ;
  assign n27152 = n18390 | n27151 ;
  assign n27155 = n12074 | n18371 ;
  assign n27154 = n8709 & n17716 ;
  assign n27156 = n27155 ^ n27154 ^ 1'b0 ;
  assign n27153 = ~n12452 & n19419 ;
  assign n27157 = n27156 ^ n27153 ^ 1'b0 ;
  assign n27158 = n19278 ^ n18371 ^ 1'b0 ;
  assign n27159 = n8102 & ~n27158 ;
  assign n27160 = n18381 ^ n9831 ^ 1'b0 ;
  assign n27161 = n27159 & n27160 ;
  assign n27162 = n27161 ^ n13702 ^ n4303 ;
  assign n27163 = n17636 ^ n10093 ^ x191 ;
  assign n27164 = n27163 ^ n2460 ^ 1'b0 ;
  assign n27166 = ( n3453 & n5512 ) | ( n3453 & ~n22926 ) | ( n5512 & ~n22926 ) ;
  assign n27167 = n27166 ^ n21351 ^ 1'b0 ;
  assign n27165 = n20673 | n25868 ;
  assign n27168 = n27167 ^ n27165 ^ 1'b0 ;
  assign n27169 = n3367 & n8440 ;
  assign n27170 = n27169 ^ n3175 ^ 1'b0 ;
  assign n27171 = n14335 | n27170 ;
  assign n27172 = n23197 & ~n27171 ;
  assign n27173 = n17200 & ~n26851 ;
  assign n27174 = n27173 ^ n12394 ^ 1'b0 ;
  assign n27175 = n12190 ^ x109 ^ 1'b0 ;
  assign n27176 = n27175 ^ n8526 ^ 1'b0 ;
  assign n27177 = n6884 & n12974 ;
  assign n27178 = n27177 ^ n26888 ^ 1'b0 ;
  assign n27179 = n1025 & ~n2751 ;
  assign n27180 = n12580 | n16398 ;
  assign n27181 = n13679 & n15595 ;
  assign n27182 = x80 & ~n15994 ;
  assign n27183 = n27182 ^ n15034 ^ 1'b0 ;
  assign n27184 = n1374 & ~n27183 ;
  assign n27185 = n27184 ^ n463 ^ 1'b0 ;
  assign n27186 = n27181 | n27185 ;
  assign n27187 = n13036 | n16872 ;
  assign n27188 = n1142 & ~n27187 ;
  assign n27189 = n11361 ^ n8691 ^ 1'b0 ;
  assign n27190 = n8661 ^ n3793 ^ 1'b0 ;
  assign n27191 = n1046 & ~n27190 ;
  assign n27192 = n27191 ^ n11696 ^ 1'b0 ;
  assign n27193 = n1795 | n8929 ;
  assign n27194 = n8608 & ~n27193 ;
  assign n27195 = n7538 | n11405 ;
  assign n27196 = n26457 | n27195 ;
  assign n27197 = n27196 ^ n25694 ^ 1'b0 ;
  assign n27198 = ~n27194 & n27197 ;
  assign n27199 = n27198 ^ n4857 ^ 1'b0 ;
  assign n27200 = ( n18074 & n23168 ) | ( n18074 & ~n27199 ) | ( n23168 & ~n27199 ) ;
  assign n27201 = n8620 & ~n16014 ;
  assign n27202 = ~n1665 & n3108 ;
  assign n27203 = ~n4168 & n27202 ;
  assign n27204 = n3209 & ~n27203 ;
  assign n27205 = n6506 & n27204 ;
  assign n27206 = n2675 & ~n3299 ;
  assign n27207 = n27205 & n27206 ;
  assign n27208 = n27207 ^ n19470 ^ 1'b0 ;
  assign n27209 = n26551 & n27208 ;
  assign n27210 = n11300 & ~n18600 ;
  assign n27211 = n3588 & n27210 ;
  assign n27212 = n5132 & ~n27110 ;
  assign n27213 = n2134 | n8717 ;
  assign n27214 = n27213 ^ n8024 ^ 1'b0 ;
  assign n27215 = n27214 ^ x241 ^ 1'b0 ;
  assign n27216 = n27215 ^ n3386 ^ 1'b0 ;
  assign n27217 = n5038 | n27216 ;
  assign n27218 = n19070 ^ n15851 ^ 1'b0 ;
  assign n27219 = ( n2118 & n11459 ) | ( n2118 & ~n13895 ) | ( n11459 & ~n13895 ) ;
  assign n27220 = n13093 ^ n7464 ^ 1'b0 ;
  assign n27221 = n27219 & ~n27220 ;
  assign n27224 = ~n13774 & n18327 ;
  assign n27222 = n645 | n1425 ;
  assign n27223 = n1702 | n27222 ;
  assign n27225 = n27224 ^ n27223 ^ 1'b0 ;
  assign n27226 = ~n11457 & n14401 ;
  assign n27227 = ~n7044 & n27226 ;
  assign n27228 = n19742 ^ n16924 ^ n4859 ;
  assign n27229 = n1683 & n14146 ;
  assign n27230 = ~n10109 & n10151 ;
  assign n27231 = n27230 ^ n9591 ^ 1'b0 ;
  assign n27232 = n27231 ^ n5714 ^ 1'b0 ;
  assign n27233 = n4096 | n7233 ;
  assign n27234 = n27233 ^ n8207 ^ 1'b0 ;
  assign n27235 = n27234 ^ n380 ^ 1'b0 ;
  assign n27236 = n5678 & ~n27235 ;
  assign n27237 = n27236 ^ n8971 ^ 1'b0 ;
  assign n27238 = ( n2543 & ~n7686 ) | ( n2543 & n8250 ) | ( ~n7686 & n8250 ) ;
  assign n27239 = ~n10123 & n27238 ;
  assign n27240 = n19538 & n27239 ;
  assign n27241 = n17346 | n19540 ;
  assign n27242 = ( ~n8437 & n9121 ) | ( ~n8437 & n27241 ) | ( n9121 & n27241 ) ;
  assign n27246 = n547 & n21468 ;
  assign n27243 = n5482 ^ n4547 ^ n1034 ;
  assign n27244 = n23579 & n27243 ;
  assign n27245 = n27244 ^ n14796 ^ 1'b0 ;
  assign n27247 = n27246 ^ n27245 ^ 1'b0 ;
  assign n27248 = n6932 | n7348 ;
  assign n27249 = n27248 ^ n851 ^ 1'b0 ;
  assign n27250 = n19623 & ~n27249 ;
  assign n27251 = n7616 ^ n3074 ^ 1'b0 ;
  assign n27252 = n1182 & n20214 ;
  assign n27253 = n25593 & n27252 ;
  assign n27254 = n10315 & ~n27253 ;
  assign n27255 = n27254 ^ n13349 ^ 1'b0 ;
  assign n27256 = n12002 ^ n10391 ^ n9201 ;
  assign n27257 = n25502 ^ n22300 ^ 1'b0 ;
  assign n27258 = n3542 & ~n11223 ;
  assign n27259 = n4892 & ~n27258 ;
  assign n27260 = ~n2337 & n9726 ;
  assign n27261 = n19298 & ~n27260 ;
  assign n27262 = n27261 ^ n7339 ^ 1'b0 ;
  assign n27263 = n5200 & n5566 ;
  assign n27264 = n2313 & n16383 ;
  assign n27265 = n6098 & n27264 ;
  assign n27266 = n18274 ^ x177 ^ 1'b0 ;
  assign n27267 = ( n2667 & ~n9352 ) | ( n2667 & n27266 ) | ( ~n9352 & n27266 ) ;
  assign n27268 = n27267 ^ n21501 ^ 1'b0 ;
  assign n27269 = n27265 & n27268 ;
  assign n27270 = n9090 ^ x51 ^ 1'b0 ;
  assign n27271 = n5691 ^ n853 ^ 1'b0 ;
  assign n27272 = ( n6051 & n15915 ) | ( n6051 & ~n27271 ) | ( n15915 & ~n27271 ) ;
  assign n27273 = ~n27270 & n27272 ;
  assign n27278 = n10321 ^ n9298 ^ n6615 ;
  assign n27279 = n6234 & n27278 ;
  assign n27274 = n22048 ^ n5479 ^ 1'b0 ;
  assign n27275 = n8544 & ~n27274 ;
  assign n27276 = ~n7352 & n27275 ;
  assign n27277 = n23975 & ~n27276 ;
  assign n27280 = n27279 ^ n27277 ^ 1'b0 ;
  assign n27281 = n14768 ^ n4191 ^ 1'b0 ;
  assign n27282 = n1701 & n1999 ;
  assign n27283 = n27282 ^ n11764 ^ 1'b0 ;
  assign n27284 = n5646 | n7465 ;
  assign n27285 = n27283 & ~n27284 ;
  assign n27286 = n17806 ^ n15230 ^ 1'b0 ;
  assign n27287 = ~n21270 & n27286 ;
  assign n27288 = n704 & n27287 ;
  assign n27289 = x197 & ~n1546 ;
  assign n27290 = n27289 ^ n643 ^ 1'b0 ;
  assign n27291 = n12169 & ~n27290 ;
  assign n27292 = n27288 & n27291 ;
  assign n27293 = ( n12189 & n19617 ) | ( n12189 & n27292 ) | ( n19617 & n27292 ) ;
  assign n27294 = n18987 ^ n6882 ^ n5463 ;
  assign n27295 = n5684 & ~n7718 ;
  assign n27296 = ( n361 & ~n27294 ) | ( n361 & n27295 ) | ( ~n27294 & n27295 ) ;
  assign n27297 = n18622 & ~n27106 ;
  assign n27299 = n24833 ^ n9649 ^ 1'b0 ;
  assign n27300 = n2441 & ~n27299 ;
  assign n27298 = n1177 & ~n10657 ;
  assign n27301 = n27300 ^ n27298 ^ 1'b0 ;
  assign n27302 = n3947 | n6112 ;
  assign n27303 = n9645 | n19147 ;
  assign n27304 = n10333 ^ n5765 ^ 1'b0 ;
  assign n27305 = ( ~n3918 & n7598 ) | ( ~n3918 & n9393 ) | ( n7598 & n9393 ) ;
  assign n27306 = n2374 | n7118 ;
  assign n27307 = n27306 ^ n1737 ^ 1'b0 ;
  assign n27308 = ~n3422 & n27307 ;
  assign n27309 = n27308 ^ n1287 ^ 1'b0 ;
  assign n27310 = ( n429 & ~n7031 ) | ( n429 & n9615 ) | ( ~n7031 & n9615 ) ;
  assign n27311 = n8557 | n20899 ;
  assign n27312 = n27311 ^ n3218 ^ 1'b0 ;
  assign n27313 = n27310 | n27312 ;
  assign n27314 = n3297 & ~n27313 ;
  assign n27315 = n27314 ^ n3659 ^ 1'b0 ;
  assign n27316 = ( n23284 & n27309 ) | ( n23284 & n27315 ) | ( n27309 & n27315 ) ;
  assign n27317 = n16194 ^ n3182 ^ n1115 ;
  assign n27318 = n27317 ^ n6811 ^ 1'b0 ;
  assign n27319 = n27318 ^ n3682 ^ 1'b0 ;
  assign n27320 = ~n20868 & n27319 ;
  assign n27322 = ( ~n1232 & n3091 ) | ( ~n1232 & n12077 ) | ( n3091 & n12077 ) ;
  assign n27321 = n1911 | n16964 ;
  assign n27323 = n27322 ^ n27321 ^ 1'b0 ;
  assign n27324 = n657 & n4235 ;
  assign n27325 = ~n7190 & n17611 ;
  assign n27326 = n27325 ^ n20458 ^ 1'b0 ;
  assign n27327 = ( n7924 & n8270 ) | ( n7924 & ~n8859 ) | ( n8270 & ~n8859 ) ;
  assign n27335 = n5999 | n14580 ;
  assign n27330 = n2808 | n5672 ;
  assign n27331 = n27330 ^ n425 ^ 1'b0 ;
  assign n27328 = n5433 | n12317 ;
  assign n27329 = n27328 ^ x192 ^ 1'b0 ;
  assign n27332 = n27331 ^ n27329 ^ n486 ;
  assign n27333 = ~n5731 & n27332 ;
  assign n27334 = n27333 ^ n11548 ^ 1'b0 ;
  assign n27336 = n27335 ^ n27334 ^ 1'b0 ;
  assign n27337 = n19629 & ~n26825 ;
  assign n27338 = n10522 & ~n16874 ;
  assign n27339 = ~n3242 & n27338 ;
  assign n27340 = n1010 & ~n7613 ;
  assign n27341 = n27340 ^ n2829 ^ 1'b0 ;
  assign n27342 = ~n6191 & n18462 ;
  assign n27343 = n27342 ^ n8020 ^ 1'b0 ;
  assign n27344 = ~n3967 & n27343 ;
  assign n27346 = n15320 ^ n10736 ^ n1715 ;
  assign n27345 = ~n3189 & n9097 ;
  assign n27347 = n27346 ^ n27345 ^ n6901 ;
  assign n27348 = n27347 ^ n2781 ^ 1'b0 ;
  assign n27349 = n16848 ^ n2179 ^ n539 ;
  assign n27350 = n3638 & n20041 ;
  assign n27351 = n14362 | n27350 ;
  assign n27353 = n1129 & n3098 ;
  assign n27354 = n27353 ^ n4773 ^ 1'b0 ;
  assign n27352 = n4310 | n23548 ;
  assign n27355 = n27354 ^ n27352 ^ 1'b0 ;
  assign n27356 = n10444 ^ n3473 ^ n753 ;
  assign n27357 = n27356 ^ x98 ^ 1'b0 ;
  assign n27358 = n17632 ^ n4448 ^ 1'b0 ;
  assign n27359 = ~n27013 & n27358 ;
  assign n27360 = n27359 ^ n7544 ^ 1'b0 ;
  assign n27361 = ~x15 & n25667 ;
  assign n27362 = n27361 ^ n10214 ^ 1'b0 ;
  assign n27363 = n1892 & n2644 ;
  assign n27364 = n791 | n7580 ;
  assign n27365 = n27364 ^ n6558 ^ 1'b0 ;
  assign n27366 = n27365 ^ n18938 ^ n2699 ;
  assign n27367 = n11666 & n15881 ;
  assign n27368 = ( n674 & ~n1401 ) | ( n674 & n27367 ) | ( ~n1401 & n27367 ) ;
  assign n27369 = n21196 ^ n11920 ^ 1'b0 ;
  assign n27370 = n19633 ^ n15680 ^ 1'b0 ;
  assign n27371 = n9086 ^ x44 ^ 1'b0 ;
  assign n27372 = n27371 ^ n4089 ^ n314 ;
  assign n27373 = n24277 ^ n13268 ^ 1'b0 ;
  assign n27374 = n15115 ^ n8034 ^ 1'b0 ;
  assign n27375 = n2847 & n27374 ;
  assign n27376 = n27375 ^ n5093 ^ 1'b0 ;
  assign n27377 = n23898 & n27376 ;
  assign n27378 = n4080 ^ n2489 ^ 1'b0 ;
  assign n27379 = n19471 | n27378 ;
  assign n27380 = ~n8578 & n12595 ;
  assign n27381 = ~n6038 & n27380 ;
  assign n27382 = ( ~n2523 & n13093 ) | ( ~n2523 & n27381 ) | ( n13093 & n27381 ) ;
  assign n27385 = ~n9993 & n21787 ;
  assign n27386 = n11400 & n27385 ;
  assign n27383 = ~n11298 & n18355 ;
  assign n27384 = n21170 & n27383 ;
  assign n27387 = n27386 ^ n27384 ^ n25238 ;
  assign n27388 = n25102 ^ n9365 ^ 1'b0 ;
  assign n27389 = n13043 & ~n23736 ;
  assign n27390 = n17598 ^ n12184 ^ n10992 ;
  assign n27391 = n27389 & n27390 ;
  assign n27392 = n9496 ^ n1993 ^ 1'b0 ;
  assign n27393 = n12899 | n27392 ;
  assign n27394 = n14592 ^ n9537 ^ 1'b0 ;
  assign n27395 = ~n27393 & n27394 ;
  assign n27396 = n8346 & ~n19836 ;
  assign n27397 = ~n27395 & n27396 ;
  assign n27398 = n25221 ^ n3407 ^ 1'b0 ;
  assign n27399 = ~n19518 & n27398 ;
  assign n27400 = ~n2769 & n4606 ;
  assign n27401 = ~x47 & n27400 ;
  assign n27402 = n12693 | n27401 ;
  assign n27403 = n27402 ^ n10937 ^ n2736 ;
  assign n27404 = ( ~n4243 & n11771 ) | ( ~n4243 & n12690 ) | ( n11771 & n12690 ) ;
  assign n27405 = n7673 & n14095 ;
  assign n27406 = ~n1302 & n27405 ;
  assign n27407 = n2024 & n27406 ;
  assign n27409 = n4312 | n9606 ;
  assign n27408 = n7863 & n19627 ;
  assign n27410 = n27409 ^ n27408 ^ 1'b0 ;
  assign n27412 = n307 & ~n1293 ;
  assign n27413 = n27412 ^ n6692 ^ 1'b0 ;
  assign n27411 = ~n2425 & n10154 ;
  assign n27414 = n27413 ^ n27411 ^ 1'b0 ;
  assign n27415 = n27414 ^ n1323 ^ 1'b0 ;
  assign n27416 = n16651 & ~n27415 ;
  assign n27417 = n5296 ^ n2942 ^ 1'b0 ;
  assign n27418 = ( n5102 & ~n23336 ) | ( n5102 & n27417 ) | ( ~n23336 & n27417 ) ;
  assign n27419 = n27418 ^ n3824 ^ n338 ;
  assign n27420 = n12132 ^ n8033 ^ 1'b0 ;
  assign n27421 = n502 & ~n5194 ;
  assign n27422 = ~n286 & n27421 ;
  assign n27423 = n5642 & n27422 ;
  assign n27424 = n27423 ^ n13887 ^ n2637 ;
  assign n27425 = n27424 ^ n4503 ^ n347 ;
  assign n27426 = n27425 ^ n1442 ^ 1'b0 ;
  assign n27427 = n27426 ^ n4993 ^ 1'b0 ;
  assign n27428 = n3063 ^ n2421 ^ 1'b0 ;
  assign n27429 = n27428 ^ n12620 ^ 1'b0 ;
  assign n27430 = ~n2588 & n10490 ;
  assign n27431 = n8416 ^ n3985 ^ 1'b0 ;
  assign n27432 = n6715 & n20039 ;
  assign n27433 = n27432 ^ n22085 ^ 1'b0 ;
  assign n27434 = n27433 ^ n5145 ^ 1'b0 ;
  assign n27435 = ~n6292 & n18754 ;
  assign n27436 = ~n7208 & n27435 ;
  assign n27437 = n25376 ^ n23546 ^ 1'b0 ;
  assign n27438 = n4758 & n27437 ;
  assign n27439 = n27438 ^ n8261 ^ 1'b0 ;
  assign n27440 = ~n18098 & n27439 ;
  assign n27441 = n8965 ^ n6001 ^ 1'b0 ;
  assign n27442 = n1847 & ~n27441 ;
  assign n27445 = ( n8390 & ~n8899 ) | ( n8390 & n18351 ) | ( ~n8899 & n18351 ) ;
  assign n27446 = n27445 ^ n1425 ^ 1'b0 ;
  assign n27447 = n11878 | n27446 ;
  assign n27443 = n803 & ~n4413 ;
  assign n27444 = n10040 & n27443 ;
  assign n27448 = n27447 ^ n27444 ^ n23560 ;
  assign n27449 = n20031 ^ n19149 ^ n12590 ;
  assign n27450 = ( n8446 & n16732 ) | ( n8446 & n19783 ) | ( n16732 & n19783 ) ;
  assign n27451 = n15806 ^ x92 ^ 1'b0 ;
  assign n27452 = ( n11880 & n13122 ) | ( n11880 & n13590 ) | ( n13122 & n13590 ) ;
  assign n27453 = n10425 | n21779 ;
  assign n27454 = n15151 & ~n27453 ;
  assign n27455 = n3783 & ~n8374 ;
  assign n27456 = n27455 ^ n14843 ^ n2849 ;
  assign n27457 = n17424 & n27456 ;
  assign n27458 = n27457 ^ n1709 ^ 1'b0 ;
  assign n27459 = n1965 & n2676 ;
  assign n27460 = n27459 ^ x56 ^ 1'b0 ;
  assign n27461 = n27460 ^ n27332 ^ n3215 ;
  assign n27462 = n27461 ^ n6940 ^ 1'b0 ;
  assign n27463 = ~n27458 & n27462 ;
  assign n27464 = x197 & n23901 ;
  assign n27465 = n8931 & n20440 ;
  assign n27466 = n27464 & n27465 ;
  assign n27467 = n27466 ^ n14258 ^ n10922 ;
  assign n27468 = ( ~n2527 & n10781 ) | ( ~n2527 & n17163 ) | ( n10781 & n17163 ) ;
  assign n27469 = n2645 & ~n27468 ;
  assign n27470 = n21834 & n27469 ;
  assign n27471 = n19529 | n20734 ;
  assign n27472 = n20250 | n27471 ;
  assign n27473 = n15564 | n26330 ;
  assign n27474 = n12371 & ~n21071 ;
  assign n27475 = n27474 ^ n14551 ^ 1'b0 ;
  assign n27476 = n17758 ^ n4858 ^ 1'b0 ;
  assign n27477 = n14054 ^ n9286 ^ 1'b0 ;
  assign n27478 = ~n14971 & n27477 ;
  assign n27479 = n27478 ^ n1768 ^ 1'b0 ;
  assign n27480 = n6332 ^ n3386 ^ n686 ;
  assign n27481 = n23981 ^ n11969 ^ n1241 ;
  assign n27482 = ~n9398 & n27481 ;
  assign n27483 = n27480 & ~n27482 ;
  assign n27484 = n13966 ^ n11706 ^ 1'b0 ;
  assign n27485 = n10755 & ~n27484 ;
  assign n27486 = n6028 & n6904 ;
  assign n27487 = n27486 ^ n7745 ^ 1'b0 ;
  assign n27488 = ~n19368 & n27487 ;
  assign n27489 = n27485 | n27488 ;
  assign n27490 = n5594 ^ n3495 ^ 1'b0 ;
  assign n27491 = ~n9883 & n18276 ;
  assign n27492 = n27491 ^ n20269 ^ 1'b0 ;
  assign n27493 = ~n3901 & n17072 ;
  assign n27494 = n27493 ^ n20599 ^ 1'b0 ;
  assign n27495 = ( ~n13695 & n14102 ) | ( ~n13695 & n26124 ) | ( n14102 & n26124 ) ;
  assign n27496 = n19204 ^ n11052 ^ n5518 ;
  assign n27497 = n11628 & ~n27496 ;
  assign n27498 = n13154 & n27497 ;
  assign n27499 = n5419 & n12113 ;
  assign n27500 = n27499 ^ n14947 ^ 1'b0 ;
  assign n27501 = n20706 | n27500 ;
  assign n27502 = n572 & ~n11078 ;
  assign n27503 = n23468 ^ n6188 ^ 1'b0 ;
  assign n27504 = n18096 & n27503 ;
  assign n27505 = n17185 | n21326 ;
  assign n27506 = n11710 & ~n27505 ;
  assign n27507 = n7743 ^ n3526 ^ 1'b0 ;
  assign n27508 = n1013 & n27507 ;
  assign n27509 = n14586 | n27508 ;
  assign n27510 = n791 & n7363 ;
  assign n27511 = n27510 ^ n7458 ^ 1'b0 ;
  assign n27512 = n3831 & ~n17733 ;
  assign n27513 = n3154 & ~n8159 ;
  assign n27514 = n27513 ^ n16018 ^ n12853 ;
  assign n27515 = n4858 | n27514 ;
  assign n27516 = n8488 ^ n2020 ^ 1'b0 ;
  assign n27517 = n4954 | n13943 ;
  assign n27518 = n27517 ^ n13489 ^ 1'b0 ;
  assign n27519 = ( n2450 & n12931 ) | ( n2450 & ~n27518 ) | ( n12931 & ~n27518 ) ;
  assign n27520 = n5754 & n18069 ;
  assign n27521 = ~n27519 & n27520 ;
  assign n27522 = n9401 ^ n5641 ^ 1'b0 ;
  assign n27525 = n11037 & ~n23940 ;
  assign n27526 = n4599 & n27525 ;
  assign n27527 = n27526 ^ n6246 ^ 1'b0 ;
  assign n27523 = n12108 ^ n3010 ^ 1'b0 ;
  assign n27524 = n12462 | n27523 ;
  assign n27528 = n27527 ^ n27524 ^ n13746 ;
  assign n27529 = ( ~n4207 & n13566 ) | ( ~n4207 & n16610 ) | ( n13566 & n16610 ) ;
  assign n27530 = n27529 ^ n16187 ^ 1'b0 ;
  assign n27531 = n22605 ^ n1397 ^ 1'b0 ;
  assign n27532 = ~n10392 & n27531 ;
  assign n27533 = ~n13402 & n27532 ;
  assign n27534 = n27533 ^ n20119 ^ n13411 ;
  assign n27535 = x61 & n12155 ;
  assign n27536 = n15221 & ~n23401 ;
  assign n27537 = n2979 & ~n27536 ;
  assign n27538 = ~n14601 & n27537 ;
  assign n27539 = n23702 ^ n4850 ^ 1'b0 ;
  assign n27540 = n6810 & n22381 ;
  assign n27541 = ~n6810 & n27540 ;
  assign n27542 = n27541 ^ n21701 ^ 1'b0 ;
  assign n27543 = n11788 & ~n27542 ;
  assign n27544 = n5281 & n27543 ;
  assign n27545 = n12074 ^ n7007 ^ n4089 ;
  assign n27546 = n27545 ^ n5778 ^ 1'b0 ;
  assign n27547 = ~n19252 & n22261 ;
  assign n27548 = n27547 ^ n7854 ^ 1'b0 ;
  assign n27549 = n27548 ^ n5211 ^ 1'b0 ;
  assign n27550 = ~n27546 & n27549 ;
  assign n27551 = n8472 ^ n5232 ^ 1'b0 ;
  assign n27552 = n6041 & n23490 ;
  assign n27553 = n8520 & n24017 ;
  assign n27554 = n27553 ^ n19083 ^ 1'b0 ;
  assign n27555 = n21879 & ~n22822 ;
  assign n27556 = n27555 ^ n13004 ^ 1'b0 ;
  assign n27557 = n27556 ^ n26381 ^ n4915 ;
  assign n27558 = n7475 & n19732 ;
  assign n27559 = n27558 ^ n10745 ^ 1'b0 ;
  assign n27562 = n10175 ^ n6895 ^ 1'b0 ;
  assign n27563 = n17544 & ~n27562 ;
  assign n27564 = ~n737 & n27563 ;
  assign n27560 = n22461 ^ n11200 ^ 1'b0 ;
  assign n27561 = n12876 & n27560 ;
  assign n27565 = n27564 ^ n27561 ^ 1'b0 ;
  assign n27566 = n19759 ^ n4438 ^ 1'b0 ;
  assign n27567 = n2248 & ~n8102 ;
  assign n27568 = n23736 & n27567 ;
  assign n27569 = ~n7595 & n10274 ;
  assign n27570 = n16378 ^ n14644 ^ 1'b0 ;
  assign n27571 = n27570 ^ n18735 ^ 1'b0 ;
  assign n27572 = n27571 ^ n10497 ^ n6251 ;
  assign n27573 = ( n22444 & n27569 ) | ( n22444 & n27572 ) | ( n27569 & n27572 ) ;
  assign n27574 = n1558 | n4104 ;
  assign n27575 = n10099 & ~n27574 ;
  assign n27576 = n27575 ^ n26556 ^ n10983 ;
  assign n27577 = n8632 & ~n19641 ;
  assign n27578 = n27577 ^ n21173 ^ 1'b0 ;
  assign n27579 = n27578 ^ n9371 ^ 1'b0 ;
  assign n27580 = n24155 | n27579 ;
  assign n27581 = ~n2652 & n7988 ;
  assign n27582 = n16838 ^ n3388 ^ 1'b0 ;
  assign n27583 = ~n27581 & n27582 ;
  assign n27584 = n11157 ^ n10081 ^ 1'b0 ;
  assign n27585 = n11482 & n19052 ;
  assign n27586 = x76 & ~n19450 ;
  assign n27587 = n8098 | n16647 ;
  assign n27588 = n16827 ^ n1077 ^ 1'b0 ;
  assign n27589 = n12515 & ~n27588 ;
  assign n27590 = n22751 ^ n18645 ^ 1'b0 ;
  assign n27591 = n5464 & ~n27590 ;
  assign n27592 = ~n16697 & n27591 ;
  assign n27593 = ~n27589 & n27592 ;
  assign n27594 = n27593 ^ n13404 ^ 1'b0 ;
  assign n27595 = n24534 ^ n9039 ^ 1'b0 ;
  assign n27596 = n15542 & n27595 ;
  assign n27597 = n27594 & n27596 ;
  assign n27598 = n11573 | n14845 ;
  assign n27599 = ( n1122 & n19196 ) | ( n1122 & ~n27598 ) | ( n19196 & ~n27598 ) ;
  assign n27600 = n16732 ^ n13759 ^ 1'b0 ;
  assign n27601 = n3523 & ~n27031 ;
  assign n27602 = n27600 & ~n27601 ;
  assign n27603 = n3879 | n21630 ;
  assign n27604 = n27603 ^ n6089 ^ 1'b0 ;
  assign n27605 = n13695 & ~n27604 ;
  assign n27606 = n27605 ^ n5103 ^ 1'b0 ;
  assign n27607 = n23253 & n27606 ;
  assign n27608 = n5369 & ~n7109 ;
  assign n27609 = ~n22791 & n27608 ;
  assign n27610 = n19456 ^ n6915 ^ 1'b0 ;
  assign n27612 = n15522 ^ n6321 ^ 1'b0 ;
  assign n27613 = ~n2426 & n27612 ;
  assign n27614 = ~n11201 & n27613 ;
  assign n27611 = n1323 & ~n16408 ;
  assign n27615 = n27614 ^ n27611 ^ 1'b0 ;
  assign n27616 = n4446 & ~n25048 ;
  assign n27617 = n5264 ^ n4840 ^ 1'b0 ;
  assign n27618 = n21914 ^ n2336 ^ 1'b0 ;
  assign n27619 = n2258 | n21009 ;
  assign n27620 = n10973 & n13450 ;
  assign n27621 = n27620 ^ n11230 ^ 1'b0 ;
  assign n27622 = n3852 | n10099 ;
  assign n27623 = n27622 ^ n1941 ^ 1'b0 ;
  assign n27624 = n27623 ^ n12620 ^ 1'b0 ;
  assign n27625 = n14715 ^ n14154 ^ 1'b0 ;
  assign n27626 = n9463 & ~n27625 ;
  assign n27629 = n12007 ^ n2617 ^ x206 ;
  assign n27627 = n17387 ^ n10771 ^ 1'b0 ;
  assign n27628 = ~n16226 & n27627 ;
  assign n27630 = n27629 ^ n27628 ^ 1'b0 ;
  assign n27631 = ( n25193 & ~n27626 ) | ( n25193 & n27630 ) | ( ~n27626 & n27630 ) ;
  assign n27632 = n5153 & ~n9415 ;
  assign n27633 = n24858 ^ n12103 ^ 1'b0 ;
  assign n27634 = n6606 | n27633 ;
  assign n27635 = n24531 & ~n27634 ;
  assign n27636 = n14968 & n17699 ;
  assign n27637 = n27636 ^ n18280 ^ 1'b0 ;
  assign n27638 = n4078 | n14258 ;
  assign n27639 = n3547 | n27638 ;
  assign n27641 = n2578 & ~n5267 ;
  assign n27642 = x161 & n27641 ;
  assign n27640 = x195 & n23504 ;
  assign n27643 = n27642 ^ n27640 ^ 1'b0 ;
  assign n27644 = ( ~n23427 & n27639 ) | ( ~n23427 & n27643 ) | ( n27639 & n27643 ) ;
  assign n27645 = n4100 & ~n24726 ;
  assign n27646 = n26829 | n27238 ;
  assign n27647 = n27646 ^ n26906 ^ 1'b0 ;
  assign n27648 = ( n2730 & n19317 ) | ( n2730 & n27647 ) | ( n19317 & n27647 ) ;
  assign n27649 = ~n3141 & n23861 ;
  assign n27651 = ~n8427 & n8510 ;
  assign n27652 = n13657 & n27651 ;
  assign n27650 = n6696 & n11914 ;
  assign n27653 = n27652 ^ n27650 ^ 1'b0 ;
  assign n27654 = ~n7337 & n27653 ;
  assign n27655 = n27654 ^ n1228 ^ 1'b0 ;
  assign n27656 = n15277 | n22994 ;
  assign n27660 = n12221 ^ n11701 ^ n2548 ;
  assign n27661 = n3216 & ~n27660 ;
  assign n27662 = n27661 ^ n19746 ^ 1'b0 ;
  assign n27659 = ~n3195 & n9118 ;
  assign n27663 = n27662 ^ n27659 ^ 1'b0 ;
  assign n27657 = n10094 & ~n16127 ;
  assign n27658 = n5510 & ~n27657 ;
  assign n27664 = n27663 ^ n27658 ^ 1'b0 ;
  assign n27665 = n5968 & ~n25567 ;
  assign n27666 = n27665 ^ n16054 ^ 1'b0 ;
  assign n27667 = n13148 | n27666 ;
  assign n27668 = n20753 ^ n6998 ^ 1'b0 ;
  assign n27669 = ~n8636 & n9645 ;
  assign n27670 = n6721 & n27669 ;
  assign n27671 = n5386 ^ n4990 ^ n1369 ;
  assign n27672 = n27670 & n27671 ;
  assign n27673 = n12544 & ~n13592 ;
  assign n27674 = n4448 ^ n1858 ^ 1'b0 ;
  assign n27675 = n9421 | n25020 ;
  assign n27676 = n27675 ^ n4412 ^ 1'b0 ;
  assign n27679 = n4532 & n5590 ;
  assign n27680 = ~n6223 & n27679 ;
  assign n27677 = n7360 ^ n4900 ^ 1'b0 ;
  assign n27678 = n12937 | n27677 ;
  assign n27681 = n27680 ^ n27678 ^ n11140 ;
  assign n27682 = n3606 & n11610 ;
  assign n27683 = n27682 ^ n18238 ^ 1'b0 ;
  assign n27684 = n4595 & ~n24286 ;
  assign n27685 = x42 | n2350 ;
  assign n27686 = n27684 | n27685 ;
  assign n27687 = n5535 & n12150 ;
  assign n27688 = n27686 | n27687 ;
  assign n27689 = ~n3078 & n22006 ;
  assign n27690 = ~n3098 & n27689 ;
  assign n27691 = n11000 ^ n9045 ^ n2504 ;
  assign n27692 = ~n11184 & n27691 ;
  assign n27693 = n27692 ^ n20622 ^ 1'b0 ;
  assign n27694 = x73 & n14978 ;
  assign n27695 = n20020 ^ n4280 ^ 1'b0 ;
  assign n27696 = n18807 & ~n27695 ;
  assign n27697 = n1612 & ~n27696 ;
  assign n27698 = n22490 ^ n11376 ^ 1'b0 ;
  assign n27699 = x225 & ~n27698 ;
  assign n27700 = n27699 ^ n4175 ^ 1'b0 ;
  assign n27701 = n27697 | n27700 ;
  assign n27702 = n8509 ^ n7251 ^ 1'b0 ;
  assign n27703 = n14954 & ~n27702 ;
  assign n27704 = n13887 & n24985 ;
  assign n27705 = ~n27703 & n27704 ;
  assign n27706 = n4059 | n11219 ;
  assign n27707 = ~n1814 & n27706 ;
  assign n27708 = n5129 & ~n27707 ;
  assign n27709 = ( ~x81 & x159 ) | ( ~x81 & n12201 ) | ( x159 & n12201 ) ;
  assign n27710 = ~x100 & n22656 ;
  assign n27713 = n2556 & n18812 ;
  assign n27714 = ~n14995 & n27713 ;
  assign n27711 = n1209 & n2542 ;
  assign n27712 = n27711 ^ n20756 ^ 1'b0 ;
  assign n27715 = n27714 ^ n27712 ^ 1'b0 ;
  assign n27716 = n5772 | n27715 ;
  assign n27717 = n27716 ^ n1733 ^ 1'b0 ;
  assign n27718 = n11518 ^ n6995 ^ 1'b0 ;
  assign n27719 = n27718 ^ n16255 ^ 1'b0 ;
  assign n27720 = n8471 ^ n1297 ^ 1'b0 ;
  assign n27721 = n17713 ^ n3439 ^ 1'b0 ;
  assign n27722 = n1343 | n27721 ;
  assign n27723 = ( ~n13308 & n27720 ) | ( ~n13308 & n27722 ) | ( n27720 & n27722 ) ;
  assign n27724 = n10144 | n25228 ;
  assign n27725 = n15760 ^ n897 ^ 1'b0 ;
  assign n27726 = n4045 ^ n2053 ^ 1'b0 ;
  assign n27727 = n5194 ^ n1113 ^ 1'b0 ;
  assign n27728 = n15608 ^ n3320 ^ 1'b0 ;
  assign n27729 = ~n2412 & n27728 ;
  assign n27730 = ( n5490 & ~n11413 ) | ( n5490 & n27729 ) | ( ~n11413 & n27729 ) ;
  assign n27731 = n5155 ^ n4198 ^ 1'b0 ;
  assign n27732 = n1882 ^ n702 ^ 1'b0 ;
  assign n27733 = n18512 & n27732 ;
  assign n27734 = n27733 ^ n2640 ^ 1'b0 ;
  assign n27735 = n15637 & ~n17302 ;
  assign n27736 = n11416 & ~n27735 ;
  assign n27737 = n21789 ^ n17570 ^ n16245 ;
  assign n27738 = n13994 & ~n24595 ;
  assign n27739 = n25123 ^ n878 ^ 1'b0 ;
  assign n27740 = ~n16427 & n27739 ;
  assign n27741 = ~n20824 & n27740 ;
  assign n27742 = n27741 ^ n22856 ^ 1'b0 ;
  assign n27743 = n27341 ^ n26308 ^ 1'b0 ;
  assign n27744 = n13366 & ~n13500 ;
  assign n27745 = n27744 ^ n6591 ^ 1'b0 ;
  assign n27746 = n6653 & n27224 ;
  assign n27747 = n10059 & n27746 ;
  assign n27748 = ~n6636 & n8946 ;
  assign n27749 = n27748 ^ n14160 ^ 1'b0 ;
  assign n27750 = ~n27747 & n27749 ;
  assign n27751 = ~n11882 & n27750 ;
  assign n27752 = n6179 & n7164 ;
  assign n27753 = n27752 ^ n3923 ^ 1'b0 ;
  assign n27754 = ( ~n8115 & n8734 ) | ( ~n8115 & n27753 ) | ( n8734 & n27753 ) ;
  assign n27755 = n8354 & ~n27754 ;
  assign n27756 = n2227 ^ n490 ^ 1'b0 ;
  assign n27757 = ~n585 & n27756 ;
  assign n27758 = n27757 ^ n9632 ^ 1'b0 ;
  assign n27759 = n9731 & ~n27758 ;
  assign n27760 = n27759 ^ n26579 ^ 1'b0 ;
  assign n27761 = n5720 & ~n27760 ;
  assign n27762 = n26044 ^ n14572 ^ 1'b0 ;
  assign n27763 = n13517 | n27762 ;
  assign n27764 = n10859 | n11603 ;
  assign n27765 = n4259 & n19457 ;
  assign n27766 = n9901 | n9912 ;
  assign n27767 = n27766 ^ n19503 ^ 1'b0 ;
  assign n27768 = n6907 ^ n1540 ^ n300 ;
  assign n27769 = ( n4516 & ~n25601 ) | ( n4516 & n27768 ) | ( ~n25601 & n27768 ) ;
  assign n27770 = n7590 & ~n20844 ;
  assign n27771 = n27769 & n27770 ;
  assign n27772 = n8765 ^ n8587 ^ 1'b0 ;
  assign n27773 = n24610 & ~n27772 ;
  assign n27774 = n16488 & ~n20497 ;
  assign n27775 = n9881 & ~n12041 ;
  assign n27778 = n9178 ^ n2054 ^ 1'b0 ;
  assign n27779 = n7788 | n27778 ;
  assign n27780 = n27779 ^ n7636 ^ n4211 ;
  assign n27776 = n3773 ^ n2165 ^ 1'b0 ;
  assign n27777 = ~n15951 & n27776 ;
  assign n27781 = n27780 ^ n27777 ^ 1'b0 ;
  assign n27782 = n14775 ^ n10989 ^ 1'b0 ;
  assign n27783 = n5993 | n9897 ;
  assign n27784 = ~n17887 & n27783 ;
  assign n27785 = ~n19938 & n27784 ;
  assign n27786 = n27782 | n27785 ;
  assign n27787 = n3123 ^ n2600 ^ x148 ;
  assign n27788 = n3129 & n9374 ;
  assign n27789 = n6871 ^ n4038 ^ 1'b0 ;
  assign n27790 = n27788 & ~n27789 ;
  assign n27791 = n26505 ^ n23170 ^ 1'b0 ;
  assign n27792 = n3775 & n27791 ;
  assign n27795 = n13309 & ~n20790 ;
  assign n27793 = n3066 & n13041 ;
  assign n27794 = n16322 | n27793 ;
  assign n27796 = n27795 ^ n27794 ^ 1'b0 ;
  assign n27797 = ~n9498 & n17072 ;
  assign n27798 = n27797 ^ n6337 ^ 1'b0 ;
  assign n27799 = n27051 ^ n18073 ^ n301 ;
  assign n27800 = n27799 ^ n4208 ^ 1'b0 ;
  assign n27801 = n3459 ^ n2762 ^ 1'b0 ;
  assign n27802 = n15406 | n27801 ;
  assign n27803 = n6299 ^ n1306 ^ n580 ;
  assign n27804 = n27803 ^ n3955 ^ 1'b0 ;
  assign n27805 = n14835 ^ n14638 ^ 1'b0 ;
  assign n27806 = n5568 | n27805 ;
  assign n27807 = n17447 ^ n9982 ^ 1'b0 ;
  assign n27808 = ~n24595 & n27807 ;
  assign n27809 = n27406 & n27808 ;
  assign n27810 = ~n1648 & n14210 ;
  assign n27811 = n6470 & n27810 ;
  assign n27812 = n4100 ^ x8 ^ 1'b0 ;
  assign n27813 = n8194 & ~n27812 ;
  assign n27814 = ~n7296 & n27813 ;
  assign n27815 = ( n19596 & ~n22572 ) | ( n19596 & n27814 ) | ( ~n22572 & n27814 ) ;
  assign n27816 = n12625 ^ n1795 ^ 1'b0 ;
  assign n27817 = ~n10668 & n13284 ;
  assign n27818 = n27817 ^ n5813 ^ 1'b0 ;
  assign n27819 = n17285 | n20206 ;
  assign n27820 = n27818 & n27819 ;
  assign n27821 = n14344 ^ n10413 ^ 1'b0 ;
  assign n27822 = n4473 | n27821 ;
  assign n27823 = n16519 & ~n20540 ;
  assign n27824 = n27822 & n27823 ;
  assign n27825 = n17036 | n19105 ;
  assign n27826 = n2075 & ~n7665 ;
  assign n27827 = n14708 & n26178 ;
  assign n27828 = ( n10737 & n15483 ) | ( n10737 & ~n25914 ) | ( n15483 & ~n25914 ) ;
  assign n27829 = ~n4884 & n14145 ;
  assign n27830 = n27829 ^ n1054 ^ 1'b0 ;
  assign n27831 = n5939 & ~n24888 ;
  assign n27832 = n8405 | n18213 ;
  assign n27833 = x6 | n27832 ;
  assign n27834 = n5413 & n27833 ;
  assign n27835 = n27831 & n27834 ;
  assign n27836 = n9667 ^ n6493 ^ 1'b0 ;
  assign n27837 = n7857 ^ n3709 ^ n1431 ;
  assign n27838 = ( n19220 & n25931 ) | ( n19220 & ~n27837 ) | ( n25931 & ~n27837 ) ;
  assign n27839 = n9425 & n18282 ;
  assign n27840 = n4576 & n18390 ;
  assign n27841 = n27839 & n27840 ;
  assign n27842 = n4207 & ~n7378 ;
  assign n27843 = n27842 ^ n15797 ^ 1'b0 ;
  assign n27844 = n11163 | n23023 ;
  assign n27845 = n27844 ^ n2235 ^ 1'b0 ;
  assign n27846 = x150 & ~n26883 ;
  assign n27847 = ( ~n8222 & n10273 ) | ( ~n8222 & n24975 ) | ( n10273 & n24975 ) ;
  assign n27848 = n11530 & ~n18603 ;
  assign n27850 = n7052 & n24797 ;
  assign n27851 = n27850 ^ n2523 ^ 1'b0 ;
  assign n27849 = ~n766 & n6485 ;
  assign n27852 = n27851 ^ n27849 ^ 1'b0 ;
  assign n27853 = n27852 ^ n7619 ^ 1'b0 ;
  assign n27854 = n4534 | n16773 ;
  assign n27855 = n15081 & ~n27854 ;
  assign n27856 = n5512 ^ n4041 ^ n2846 ;
  assign n27857 = n16155 ^ n16060 ^ 1'b0 ;
  assign n27858 = x30 & ~n27857 ;
  assign n27859 = n14081 ^ n7693 ^ 1'b0 ;
  assign n27860 = n1801 | n5947 ;
  assign n27861 = n4768 ^ n607 ^ 1'b0 ;
  assign n27862 = n27860 & n27861 ;
  assign n27863 = n22779 ^ n19404 ^ 1'b0 ;
  assign n27864 = n3777 ^ n1795 ^ 1'b0 ;
  assign n27865 = n4602 | n27864 ;
  assign n27866 = ( n456 & ~n5996 ) | ( n456 & n12526 ) | ( ~n5996 & n12526 ) ;
  assign n27867 = n27865 & ~n27866 ;
  assign n27868 = n25575 ^ n12679 ^ 1'b0 ;
  assign n27869 = n27265 ^ n14422 ^ 1'b0 ;
  assign n27870 = n20755 & ~n27869 ;
  assign n27871 = n14102 ^ n5490 ^ 1'b0 ;
  assign n27872 = ~n7334 & n27871 ;
  assign n27873 = n27872 ^ n26545 ^ 1'b0 ;
  assign n27874 = n6998 & n27873 ;
  assign n27875 = n22206 ^ n918 ^ 1'b0 ;
  assign n27878 = n2996 & n4213 ;
  assign n27879 = n27878 ^ n19362 ^ 1'b0 ;
  assign n27880 = n27879 ^ n3627 ^ 1'b0 ;
  assign n27881 = ~n4146 & n27880 ;
  assign n27876 = ~n1483 & n18339 ;
  assign n27877 = n9750 & n27876 ;
  assign n27882 = n27881 ^ n27877 ^ 1'b0 ;
  assign n27883 = n13195 | n27882 ;
  assign n27884 = n22056 ^ n1192 ^ 1'b0 ;
  assign n27885 = n6085 & ~n10965 ;
  assign n27886 = n27885 ^ n20685 ^ 1'b0 ;
  assign n27887 = n27886 ^ n10879 ^ 1'b0 ;
  assign n27888 = n14533 ^ n739 ^ 1'b0 ;
  assign n27889 = n18997 | n27888 ;
  assign n27890 = n1980 & ~n27889 ;
  assign n27891 = ~n3884 & n27890 ;
  assign n27892 = n15202 & n20260 ;
  assign n27893 = n26601 ^ n18270 ^ 1'b0 ;
  assign n27894 = n9115 & ~n27893 ;
  assign n27895 = n15946 ^ n10050 ^ n9077 ;
  assign n27896 = n27895 ^ n3804 ^ 1'b0 ;
  assign n27897 = n8709 & ~n27896 ;
  assign n27898 = ~n4356 & n27897 ;
  assign n27899 = ( ~n3734 & n27894 ) | ( ~n3734 & n27898 ) | ( n27894 & n27898 ) ;
  assign n27900 = n21295 | n23019 ;
  assign n27901 = n1134 | n3625 ;
  assign n27902 = n3625 & ~n27901 ;
  assign n27903 = n27902 ^ n4719 ^ 1'b0 ;
  assign n27904 = ~n3651 & n27903 ;
  assign n27905 = n27904 ^ n13562 ^ 1'b0 ;
  assign n27908 = n11631 & n12802 ;
  assign n27909 = n27908 ^ n20657 ^ 1'b0 ;
  assign n27906 = n1342 | n8005 ;
  assign n27907 = n22604 & ~n27906 ;
  assign n27910 = n27909 ^ n27907 ^ n10183 ;
  assign n27911 = x58 & ~n27910 ;
  assign n27912 = ~n27905 & n27911 ;
  assign n27913 = n2816 | n25294 ;
  assign n27914 = ~n5244 & n20236 ;
  assign n27915 = ~n706 & n6323 ;
  assign n27916 = ~n27914 & n27915 ;
  assign n27917 = ( n6684 & n9339 ) | ( n6684 & n27916 ) | ( n9339 & n27916 ) ;
  assign n27918 = n9261 | n27917 ;
  assign n27919 = n27451 & ~n27918 ;
  assign n27920 = n17080 ^ n13844 ^ 1'b0 ;
  assign n27921 = n12417 & ~n27920 ;
  assign n27922 = n27921 ^ n1024 ^ 1'b0 ;
  assign n27923 = n27470 ^ n13293 ^ 1'b0 ;
  assign n27924 = n4489 & ~n27923 ;
  assign n27925 = n11086 & ~n12194 ;
  assign n27926 = ( n275 & n27049 ) | ( n275 & ~n27925 ) | ( n27049 & ~n27925 ) ;
  assign n27927 = n18332 ^ n1272 ^ 1'b0 ;
  assign n27928 = ~n5326 & n23780 ;
  assign n27929 = n21805 & n27928 ;
  assign n27930 = n27929 ^ n24862 ^ 1'b0 ;
  assign n27931 = n27930 ^ n11466 ^ 1'b0 ;
  assign n27932 = n22306 & n27931 ;
  assign n27933 = n8507 ^ n617 ^ 1'b0 ;
  assign n27934 = n27932 & n27933 ;
  assign n27935 = n12551 ^ x75 ^ 1'b0 ;
  assign n27936 = n24058 ^ n20764 ^ 1'b0 ;
  assign n27937 = n1667 ^ n1323 ^ 1'b0 ;
  assign n27938 = ~n27207 & n27937 ;
  assign n27940 = n9665 ^ x22 ^ 1'b0 ;
  assign n27939 = n5465 | n8372 ;
  assign n27941 = n27940 ^ n27939 ^ 1'b0 ;
  assign n27942 = n2930 & ~n8610 ;
  assign n27943 = ( ~n5384 & n13426 ) | ( ~n5384 & n27942 ) | ( n13426 & n27942 ) ;
  assign n27945 = n12832 ^ n1113 ^ 1'b0 ;
  assign n27946 = n18742 & n27945 ;
  assign n27944 = x8 & n4624 ;
  assign n27947 = n27946 ^ n27944 ^ 1'b0 ;
  assign n27948 = ( n2444 & n27943 ) | ( n2444 & n27947 ) | ( n27943 & n27947 ) ;
  assign n27949 = n25469 ^ n8775 ^ 1'b0 ;
  assign n27950 = n19217 ^ n9890 ^ n3657 ;
  assign n27951 = n27950 ^ x142 ^ 1'b0 ;
  assign n27952 = n27951 ^ n15649 ^ n14886 ;
  assign n27953 = n15165 ^ n14274 ^ 1'b0 ;
  assign n27954 = n27952 & ~n27953 ;
  assign n27955 = ~n1063 & n8295 ;
  assign n27956 = n8562 & n27955 ;
  assign n27957 = n15707 | n27956 ;
  assign n27958 = n24689 | n27957 ;
  assign n27959 = n1957 ^ n1865 ^ 1'b0 ;
  assign n27960 = ~n25855 & n27926 ;
  assign n27961 = n13146 ^ n7593 ^ 1'b0 ;
  assign n27962 = n15115 | n22924 ;
  assign n27964 = n18588 ^ n15926 ^ 1'b0 ;
  assign n27963 = n2029 & ~n6479 ;
  assign n27965 = n27964 ^ n27963 ^ n614 ;
  assign n27966 = ~n11534 & n21385 ;
  assign n27967 = n2180 & n27966 ;
  assign n27968 = ( n2002 & n12406 ) | ( n2002 & ~n27967 ) | ( n12406 & ~n27967 ) ;
  assign n27970 = ( ~n2132 & n4573 ) | ( ~n2132 & n4953 ) | ( n4573 & n4953 ) ;
  assign n27969 = n8002 & n15953 ;
  assign n27971 = n27970 ^ n27969 ^ 1'b0 ;
  assign n27973 = n2217 & n20440 ;
  assign n27974 = n27973 ^ n1735 ^ 1'b0 ;
  assign n27972 = n1730 & n24373 ;
  assign n27975 = n27974 ^ n27972 ^ 1'b0 ;
  assign n27978 = n1932 & ~n6459 ;
  assign n27979 = n27978 ^ n12301 ^ 1'b0 ;
  assign n27976 = n4648 & n5369 ;
  assign n27977 = n7151 & ~n27976 ;
  assign n27980 = n27979 ^ n27977 ^ n21828 ;
  assign n27981 = n27243 ^ n12741 ^ 1'b0 ;
  assign n27982 = n27981 ^ n14394 ^ 1'b0 ;
  assign n27983 = n15557 & ~n27982 ;
  assign n27984 = n4255 ^ n1401 ^ 1'b0 ;
  assign n27985 = n18454 & n27984 ;
  assign n27986 = n496 | n5008 ;
  assign n27987 = n10276 ^ n3608 ^ 1'b0 ;
  assign n27988 = n1376 & ~n27987 ;
  assign n27989 = ~n11242 & n27988 ;
  assign n27990 = n14490 | n25171 ;
  assign n27992 = n3126 & ~n10518 ;
  assign n27991 = n8996 ^ x11 ^ 1'b0 ;
  assign n27993 = n27992 ^ n27991 ^ 1'b0 ;
  assign n27994 = x0 | n27993 ;
  assign n27995 = n8735 & n20645 ;
  assign n27996 = n3920 & n6829 ;
  assign n27997 = n365 & n27996 ;
  assign n27998 = n2921 & ~n6370 ;
  assign n27999 = ~n1980 & n5576 ;
  assign n28000 = ~n2866 & n13944 ;
  assign n28001 = ~n27318 & n28000 ;
  assign n28002 = n9512 | n18506 ;
  assign n28006 = n4406 | n14208 ;
  assign n28003 = x247 & ~n16954 ;
  assign n28004 = n28003 ^ n11353 ^ 1'b0 ;
  assign n28005 = n2675 | n28004 ;
  assign n28007 = n28006 ^ n28005 ^ 1'b0 ;
  assign n28008 = ~n14945 & n19310 ;
  assign n28009 = ~n10572 & n28008 ;
  assign n28010 = ~n7021 & n28009 ;
  assign n28011 = n13632 ^ n3794 ^ n2797 ;
  assign n28012 = n4359 | n14102 ;
  assign n28013 = n18298 ^ n13169 ^ 1'b0 ;
  assign n28014 = n15695 ^ n11472 ^ 1'b0 ;
  assign n28015 = ( n11147 & n23698 ) | ( n11147 & n25464 ) | ( n23698 & n25464 ) ;
  assign n28016 = n2300 & n5313 ;
  assign n28017 = n24820 & n28016 ;
  assign n28018 = n4389 & n28017 ;
  assign n28019 = n19887 ^ n11961 ^ n3077 ;
  assign n28020 = n2766 & ~n28019 ;
  assign n28021 = n28020 ^ n11993 ^ 1'b0 ;
  assign n28022 = n4153 ^ n2844 ^ 1'b0 ;
  assign n28023 = n24995 & n28022 ;
  assign n28024 = n19946 ^ n2617 ^ 1'b0 ;
  assign n28025 = n11147 & ~n28024 ;
  assign n28026 = n28025 ^ n26534 ^ 1'b0 ;
  assign n28027 = n15418 ^ n14207 ^ 1'b0 ;
  assign n28028 = ~n4380 & n28027 ;
  assign n28029 = ~n7462 & n9502 ;
  assign n28030 = n10992 ^ n5850 ^ 1'b0 ;
  assign n28031 = n12029 & n19684 ;
  assign n28032 = n4371 & n28031 ;
  assign n28033 = n28030 & ~n28032 ;
  assign n28034 = ~n11878 & n28033 ;
  assign n28035 = n25299 & n28034 ;
  assign n28036 = n341 | n3324 ;
  assign n28037 = n28036 ^ n2243 ^ 1'b0 ;
  assign n28038 = n19649 & ~n26573 ;
  assign n28045 = n1415 | n10472 ;
  assign n28046 = n28045 ^ n15788 ^ 1'b0 ;
  assign n28040 = n2983 ^ n319 ^ 1'b0 ;
  assign n28041 = n13369 | n28040 ;
  assign n28042 = n24128 & ~n28041 ;
  assign n28043 = ~n5274 & n28042 ;
  assign n28044 = n14048 | n28043 ;
  assign n28047 = n28046 ^ n28044 ^ 1'b0 ;
  assign n28039 = ~n13000 & n16149 ;
  assign n28048 = n28047 ^ n28039 ^ 1'b0 ;
  assign n28049 = n14862 ^ n12620 ^ n3918 ;
  assign n28050 = n2194 & n12923 ;
  assign n28051 = n7004 | n13185 ;
  assign n28052 = n19852 & n28051 ;
  assign n28053 = n28052 ^ n5107 ^ 1'b0 ;
  assign n28054 = ~n7780 & n28053 ;
  assign n28055 = n13177 ^ n1180 ^ 1'b0 ;
  assign n28056 = n17009 & ~n28055 ;
  assign n28057 = n28056 ^ n17122 ^ n13302 ;
  assign n28058 = n12636 ^ n2743 ^ 1'b0 ;
  assign n28059 = n2057 & ~n9737 ;
  assign n28060 = ~n28058 & n28059 ;
  assign n28061 = n11351 & ~n20340 ;
  assign n28062 = n26137 & n28061 ;
  assign n28063 = ~n11124 & n23255 ;
  assign n28064 = ( n1113 & n12478 ) | ( n1113 & n28063 ) | ( n12478 & n28063 ) ;
  assign n28067 = n21484 ^ n5417 ^ 1'b0 ;
  assign n28065 = ~n458 & n16925 ;
  assign n28066 = ~n15126 & n28065 ;
  assign n28068 = n28067 ^ n28066 ^ n3104 ;
  assign n28071 = ~n15905 & n19473 ;
  assign n28072 = n28071 ^ n9343 ^ 1'b0 ;
  assign n28073 = n5811 | n28072 ;
  assign n28069 = n1553 & n10582 ;
  assign n28070 = n17114 & n28069 ;
  assign n28074 = n28073 ^ n28070 ^ 1'b0 ;
  assign n28077 = n3394 & ~n11428 ;
  assign n28075 = n15710 ^ n5841 ^ 1'b0 ;
  assign n28076 = n28075 ^ n2650 ^ 1'b0 ;
  assign n28078 = n28077 ^ n28076 ^ n8109 ;
  assign n28079 = n2530 | n3725 ;
  assign n28080 = n28079 ^ n3133 ^ 1'b0 ;
  assign n28081 = n26056 ^ n12656 ^ 1'b0 ;
  assign n28082 = n28080 | n28081 ;
  assign n28088 = n16019 ^ n5977 ^ n874 ;
  assign n28089 = n17985 ^ n1010 ^ 1'b0 ;
  assign n28090 = n14491 | n28089 ;
  assign n28091 = n28088 & ~n28090 ;
  assign n28092 = n28091 ^ n18773 ^ 1'b0 ;
  assign n28083 = n11878 ^ n7185 ^ 1'b0 ;
  assign n28084 = ~n27258 & n28083 ;
  assign n28085 = n28084 ^ n25618 ^ 1'b0 ;
  assign n28086 = n28085 ^ n17669 ^ 1'b0 ;
  assign n28087 = n8897 | n28086 ;
  assign n28093 = n28092 ^ n28087 ^ n20427 ;
  assign n28100 = x179 & n6479 ;
  assign n28101 = n28100 ^ n16148 ^ n7506 ;
  assign n28102 = n3233 | n7316 ;
  assign n28103 = ( n3869 & n14204 ) | ( n3869 & ~n28102 ) | ( n14204 & ~n28102 ) ;
  assign n28104 = ~n28101 & n28103 ;
  assign n28094 = n6484 ^ n1380 ^ 1'b0 ;
  assign n28095 = n4884 | n10348 ;
  assign n28096 = n28094 & ~n28095 ;
  assign n28097 = ~n3087 & n28096 ;
  assign n28098 = n9074 | n28097 ;
  assign n28099 = n26906 | n28098 ;
  assign n28105 = n28104 ^ n28099 ^ n759 ;
  assign n28106 = n6647 & n23035 ;
  assign n28107 = n28106 ^ n5037 ^ 1'b0 ;
  assign n28108 = n8229 & n13448 ;
  assign n28109 = n28108 ^ n10131 ^ 1'b0 ;
  assign n28110 = ( n25562 & ~n28107 ) | ( n25562 & n28109 ) | ( ~n28107 & n28109 ) ;
  assign n28111 = n28110 ^ n18943 ^ 1'b0 ;
  assign n28112 = n2959 ^ n1806 ^ 1'b0 ;
  assign n28113 = n14487 | n23905 ;
  assign n28114 = n28113 ^ n9755 ^ 1'b0 ;
  assign n28115 = n9693 & n28114 ;
  assign n28116 = ( ~n5850 & n13925 ) | ( ~n5850 & n23936 ) | ( n13925 & n23936 ) ;
  assign n28117 = n18330 | n26851 ;
  assign n28118 = ~n2226 & n6362 ;
  assign n28119 = ( n13556 & ~n28117 ) | ( n13556 & n28118 ) | ( ~n28117 & n28118 ) ;
  assign n28120 = n3215 ^ n1021 ^ n610 ;
  assign n28121 = n1919 & ~n28120 ;
  assign n28122 = n24845 ^ n24691 ^ 1'b0 ;
  assign n28123 = ~n7313 & n10944 ;
  assign n28124 = n28123 ^ n6756 ^ 1'b0 ;
  assign n28125 = n19169 | n28124 ;
  assign n28126 = n28125 ^ n1172 ^ 1'b0 ;
  assign n28127 = ~n6993 & n20161 ;
  assign n28128 = ~n6793 & n28127 ;
  assign n28129 = n6268 ^ n3714 ^ n607 ;
  assign n28130 = n28129 ^ n11161 ^ n1269 ;
  assign n28131 = n23492 ^ n15491 ^ 1'b0 ;
  assign n28132 = ~n1695 & n28131 ;
  assign n28133 = ~n28130 & n28132 ;
  assign n28134 = n28133 ^ n16438 ^ 1'b0 ;
  assign n28135 = n28134 ^ x7 ^ 1'b0 ;
  assign n28136 = ~n19636 & n28135 ;
  assign n28138 = n12165 ^ n3507 ^ 1'b0 ;
  assign n28137 = n13080 & n16659 ;
  assign n28139 = n28138 ^ n28137 ^ 1'b0 ;
  assign n28140 = n28046 ^ n10890 ^ n963 ;
  assign n28141 = ( n9362 & n27106 ) | ( n9362 & n28140 ) | ( n27106 & n28140 ) ;
  assign n28142 = n14510 ^ n13744 ^ 1'b0 ;
  assign n28143 = ~n9773 & n28142 ;
  assign n28144 = n28143 ^ n1592 ^ 1'b0 ;
  assign n28145 = ~n5133 & n14796 ;
  assign n28146 = x98 ^ x64 ^ 1'b0 ;
  assign n28147 = n28146 ^ n5130 ^ 1'b0 ;
  assign n28148 = n10624 | n28147 ;
  assign n28149 = ~n28145 & n28148 ;
  assign n28150 = n7399 ^ n5726 ^ 1'b0 ;
  assign n28151 = n23041 | n28150 ;
  assign n28152 = n28151 ^ n24997 ^ 1'b0 ;
  assign n28153 = n20688 & ~n27951 ;
  assign n28154 = n28153 ^ n16143 ^ 1'b0 ;
  assign n28155 = ~n9534 & n11531 ;
  assign n28156 = ~n2916 & n28155 ;
  assign n28157 = n28156 ^ n10782 ^ 1'b0 ;
  assign n28158 = n7675 ^ n4549 ^ 1'b0 ;
  assign n28159 = n6036 & n28158 ;
  assign n28160 = n28157 & n28159 ;
  assign n28161 = n28160 ^ n4618 ^ 1'b0 ;
  assign n28162 = n3973 ^ n940 ^ 1'b0 ;
  assign n28163 = n26539 & ~n28162 ;
  assign n28164 = n28163 ^ n12462 ^ 1'b0 ;
  assign n28165 = n7383 & n7476 ;
  assign n28166 = ( n593 & n22025 ) | ( n593 & n28165 ) | ( n22025 & n28165 ) ;
  assign n28167 = n24379 ^ n3972 ^ 1'b0 ;
  assign n28168 = n4696 ^ n4656 ^ 1'b0 ;
  assign n28169 = ~n27831 & n28168 ;
  assign n28170 = n10206 & n28169 ;
  assign n28171 = n28170 ^ n2739 ^ 1'b0 ;
  assign n28172 = ~n1147 & n24483 ;
  assign n28173 = n4170 | n13995 ;
  assign n28174 = n15874 & ~n22599 ;
  assign n28175 = n28174 ^ n13723 ^ 1'b0 ;
  assign n28176 = n21383 ^ n2922 ^ 1'b0 ;
  assign n28177 = n11837 ^ n4287 ^ n3716 ;
  assign n28178 = n24719 & ~n28177 ;
  assign n28179 = n28178 ^ x228 ^ 1'b0 ;
  assign n28180 = n1213 | n11457 ;
  assign n28181 = n27464 & ~n28180 ;
  assign n28182 = n28181 ^ n20146 ^ n4066 ;
  assign n28183 = n21515 ^ n8894 ^ 1'b0 ;
  assign n28184 = n6332 & ~n28183 ;
  assign n28186 = n3058 ^ x245 ^ 1'b0 ;
  assign n28185 = n6658 | n11349 ;
  assign n28187 = n28186 ^ n28185 ^ 1'b0 ;
  assign n28188 = n27246 ^ n7413 ^ 1'b0 ;
  assign n28189 = ~n18715 & n28188 ;
  assign n28190 = n11915 ^ n2197 ^ 1'b0 ;
  assign n28191 = n23547 & ~n28190 ;
  assign n28192 = ( n2351 & n15710 ) | ( n2351 & n21799 ) | ( n15710 & n21799 ) ;
  assign n28193 = x132 & n7544 ;
  assign n28194 = n14036 ^ x55 ^ 1'b0 ;
  assign n28195 = n17005 ^ n12712 ^ 1'b0 ;
  assign n28196 = n22114 & ~n28195 ;
  assign n28197 = n1613 | n2733 ;
  assign n28198 = n6398 | n28197 ;
  assign n28199 = n4913 & n28198 ;
  assign n28200 = n28199 ^ n16100 ^ 1'b0 ;
  assign n28201 = n2728 & ~n28200 ;
  assign n28202 = n28201 ^ n13913 ^ 1'b0 ;
  assign n28203 = n28202 ^ n9006 ^ 1'b0 ;
  assign n28204 = n8587 & ~n24407 ;
  assign n28205 = n25982 ^ n17813 ^ 1'b0 ;
  assign n28206 = x73 & n27860 ;
  assign n28208 = n23560 ^ n9663 ^ 1'b0 ;
  assign n28207 = n17492 & ~n18791 ;
  assign n28209 = n28208 ^ n28207 ^ 1'b0 ;
  assign n28210 = n28209 ^ n23427 ^ 1'b0 ;
  assign n28212 = n27731 ^ n7567 ^ n1559 ;
  assign n28211 = n11121 & n22096 ;
  assign n28213 = n28212 ^ n28211 ^ 1'b0 ;
  assign n28214 = n12074 & n16970 ;
  assign n28215 = ~n3881 & n12231 ;
  assign n28216 = n25975 ^ n7804 ^ 1'b0 ;
  assign n28217 = ( n14086 & ~n16466 ) | ( n14086 & n28216 ) | ( ~n16466 & n28216 ) ;
  assign n28218 = n28217 ^ n9327 ^ 1'b0 ;
  assign n28219 = ~n15115 & n28218 ;
  assign n28220 = n7695 & ~n26341 ;
  assign n28221 = n19535 ^ n12118 ^ n8899 ;
  assign n28222 = n4286 & ~n9131 ;
  assign n28223 = n28222 ^ n11251 ^ 1'b0 ;
  assign n28224 = n10097 & ~n16905 ;
  assign n28225 = n512 & ~n13196 ;
  assign n28226 = n20245 & n28225 ;
  assign n28227 = n854 & n1213 ;
  assign n28228 = ~n21370 & n28227 ;
  assign n28229 = n21040 ^ n1527 ^ 1'b0 ;
  assign n28230 = n5310 | n17769 ;
  assign n28231 = x188 | n12116 ;
  assign n28232 = n13471 & n28231 ;
  assign n28233 = ~n739 & n28232 ;
  assign n28234 = n28233 ^ n25186 ^ n9885 ;
  assign n28235 = n7643 & ~n9151 ;
  assign n28236 = n28235 ^ n21642 ^ 1'b0 ;
  assign n28237 = ~n1788 & n8683 ;
  assign n28238 = ~n7508 & n28237 ;
  assign n28239 = n14379 ^ n8927 ^ 1'b0 ;
  assign n28240 = ~n28238 & n28239 ;
  assign n28241 = n7673 & n10820 ;
  assign n28242 = n3175 & n28241 ;
  assign n28243 = n28051 ^ n1851 ^ 1'b0 ;
  assign n28244 = n8955 & ~n28243 ;
  assign n28245 = n673 & ~n8201 ;
  assign n28246 = ~n673 & n28245 ;
  assign n28247 = n2595 & ~n28246 ;
  assign n28248 = n1443 | n1761 ;
  assign n28249 = n28248 ^ n3910 ^ 1'b0 ;
  assign n28250 = n6314 | n15699 ;
  assign n28251 = n19916 & n20531 ;
  assign n28252 = ~n28250 & n28251 ;
  assign n28253 = n28249 | n28252 ;
  assign n28254 = n1453 & ~n28253 ;
  assign n28255 = n14917 & ~n16864 ;
  assign n28256 = n28255 ^ n20137 ^ 1'b0 ;
  assign n28257 = ~n19237 & n19695 ;
  assign n28258 = n1928 ^ n488 ^ 1'b0 ;
  assign n28259 = x121 & n28258 ;
  assign n28260 = n28257 | n28259 ;
  assign n28261 = n3316 & ~n28260 ;
  assign n28262 = n28261 ^ n9113 ^ 1'b0 ;
  assign n28263 = n10109 ^ n6625 ^ 1'b0 ;
  assign n28264 = ( n484 & n19511 ) | ( n484 & n28263 ) | ( n19511 & n28263 ) ;
  assign n28265 = n8527 & n9241 ;
  assign n28266 = n15680 & ~n28265 ;
  assign n28267 = n2416 & ~n28076 ;
  assign n28268 = n6501 ^ n4563 ^ 1'b0 ;
  assign n28269 = n15122 | n28268 ;
  assign n28275 = n5705 | n20010 ;
  assign n28276 = n28275 ^ n13781 ^ 1'b0 ;
  assign n28270 = n6225 ^ n2856 ^ n2712 ;
  assign n28271 = n12041 ^ n11163 ^ 1'b0 ;
  assign n28272 = n28270 & n28271 ;
  assign n28273 = n1435 & n28272 ;
  assign n28274 = n10771 & n28273 ;
  assign n28277 = n28276 ^ n28274 ^ n13473 ;
  assign n28278 = ~n3378 & n10605 ;
  assign n28279 = n28277 | n28278 ;
  assign n28280 = n8453 ^ n1703 ^ 1'b0 ;
  assign n28284 = n10922 ^ n1722 ^ x123 ;
  assign n28285 = n6648 ^ n994 ^ 1'b0 ;
  assign n28286 = n28284 & ~n28285 ;
  assign n28281 = n721 | n9956 ;
  assign n28282 = n28281 ^ n7306 ^ 1'b0 ;
  assign n28283 = n21835 & ~n28282 ;
  assign n28287 = n28286 ^ n28283 ^ 1'b0 ;
  assign n28288 = n28287 ^ n25649 ^ n10374 ;
  assign n28289 = n3077 ^ n1283 ^ 1'b0 ;
  assign n28290 = ~n5820 & n28289 ;
  assign n28291 = n28290 ^ n9816 ^ n4552 ;
  assign n28292 = n28291 ^ n24900 ^ n2586 ;
  assign n28293 = ~n8250 & n28292 ;
  assign n28298 = n7086 & ~n19757 ;
  assign n28299 = n28298 ^ n3338 ^ 1'b0 ;
  assign n28300 = n9398 | n28299 ;
  assign n28301 = n3317 | n28300 ;
  assign n28294 = n12215 ^ n3052 ^ n2993 ;
  assign n28295 = n4109 ^ n3814 ^ 1'b0 ;
  assign n28296 = n4626 | n28295 ;
  assign n28297 = n28294 & n28296 ;
  assign n28302 = n28301 ^ n28297 ^ n16952 ;
  assign n28303 = n4426 & n10963 ;
  assign n28304 = n28303 ^ n15303 ^ 1'b0 ;
  assign n28305 = n28302 & n28304 ;
  assign n28306 = ~n2460 & n13199 ;
  assign n28307 = n4967 & n28306 ;
  assign n28308 = n10979 & ~n28307 ;
  assign n28309 = ~n5677 & n8200 ;
  assign n28310 = ~n11519 & n28309 ;
  assign n28311 = ~n2214 & n28310 ;
  assign n28312 = ( n10669 & ~n13583 ) | ( n10669 & n25244 ) | ( ~n13583 & n25244 ) ;
  assign n28313 = n14730 & ~n28312 ;
  assign n28314 = n2962 & n5324 ;
  assign n28315 = ~n5324 & n28314 ;
  assign n28316 = n4331 & ~n28315 ;
  assign n28317 = n28315 & n28316 ;
  assign n28318 = ~n10265 & n20565 ;
  assign n28319 = n17458 | n18903 ;
  assign n28320 = ~n7185 & n10746 ;
  assign n28321 = n28320 ^ n24215 ^ 1'b0 ;
  assign n28322 = ~n28319 & n28321 ;
  assign n28323 = n23413 ^ n7584 ^ 1'b0 ;
  assign n28324 = n28323 ^ n5304 ^ 1'b0 ;
  assign n28325 = n28324 ^ n27196 ^ 1'b0 ;
  assign n28326 = n28325 ^ n8137 ^ n7170 ;
  assign n28327 = n25434 ^ n10298 ^ n1259 ;
  assign n28328 = ~n7799 & n22139 ;
  assign n28329 = n28328 ^ n23013 ^ 1'b0 ;
  assign n28330 = n10085 ^ n8320 ^ n5483 ;
  assign n28331 = ( ~n11170 & n14928 ) | ( ~n11170 & n28330 ) | ( n14928 & n28330 ) ;
  assign n28332 = ( ~n28327 & n28329 ) | ( ~n28327 & n28331 ) | ( n28329 & n28331 ) ;
  assign n28333 = n1304 & n4710 ;
  assign n28334 = ~n2727 & n2962 ;
  assign n28335 = n28334 ^ n8894 ^ 1'b0 ;
  assign n28336 = n11788 ^ n9457 ^ n985 ;
  assign n28337 = ( n4298 & ~n7477 ) | ( n4298 & n18149 ) | ( ~n7477 & n18149 ) ;
  assign n28339 = ~n1210 & n25018 ;
  assign n28340 = ~n13044 & n28339 ;
  assign n28341 = n28340 ^ n12058 ^ 1'b0 ;
  assign n28342 = ~n2425 & n28341 ;
  assign n28338 = n6102 & n15985 ;
  assign n28343 = n28342 ^ n28338 ^ 1'b0 ;
  assign n28344 = n14580 | n17507 ;
  assign n28345 = n13681 | n28344 ;
  assign n28346 = n22126 & n28345 ;
  assign n28347 = n28346 ^ n10027 ^ 1'b0 ;
  assign n28348 = ( n9569 & n21947 ) | ( n9569 & ~n28347 ) | ( n21947 & ~n28347 ) ;
  assign n28349 = n3138 & n9658 ;
  assign n28350 = n10901 & n28349 ;
  assign n28351 = ( n1409 & n7616 ) | ( n1409 & ~n28350 ) | ( n7616 & ~n28350 ) ;
  assign n28352 = n7223 & n13172 ;
  assign n28353 = n27212 ^ n27068 ^ 1'b0 ;
  assign n28354 = n22484 ^ n3804 ^ x70 ;
  assign n28355 = n18070 ^ n7074 ^ x8 ;
  assign n28356 = n8923 ^ n2621 ^ 1'b0 ;
  assign n28357 = n10116 | n15020 ;
  assign n28358 = n5085 ^ n3938 ^ n821 ;
  assign n28359 = n28358 ^ n23511 ^ 1'b0 ;
  assign n28360 = n2673 & n6677 ;
  assign n28361 = ~n17874 & n19581 ;
  assign n28362 = n28361 ^ n20676 ^ 1'b0 ;
  assign n28363 = n13805 & n24650 ;
  assign n28364 = n11821 ^ n3627 ^ 1'b0 ;
  assign n28365 = ~n559 & n28364 ;
  assign n28366 = ~n25638 & n28365 ;
  assign n28368 = n14366 ^ n9544 ^ 1'b0 ;
  assign n28367 = n286 | n1455 ;
  assign n28369 = n28368 ^ n28367 ^ n3283 ;
  assign n28370 = n27404 ^ n10919 ^ 1'b0 ;
  assign n28371 = n6216 & n28370 ;
  assign n28372 = ~n3296 & n20832 ;
  assign n28373 = n28372 ^ n12970 ^ 1'b0 ;
  assign n28374 = n3383 & n10724 ;
  assign n28376 = x229 & ~n15295 ;
  assign n28377 = n3261 & n28376 ;
  assign n28375 = n9871 & ~n20809 ;
  assign n28378 = n28377 ^ n28375 ^ 1'b0 ;
  assign n28379 = n16874 & ~n19587 ;
  assign n28380 = n8859 | n27705 ;
  assign n28381 = n28380 ^ n15284 ^ 1'b0 ;
  assign n28382 = n26049 ^ n2626 ^ 1'b0 ;
  assign n28383 = n1239 ^ x182 ^ 1'b0 ;
  assign n28384 = n10787 & n20243 ;
  assign n28385 = n9676 & n28384 ;
  assign n28386 = n17523 & ~n28385 ;
  assign n28387 = ~n28383 & n28386 ;
  assign n28388 = n5498 & n23151 ;
  assign n28389 = n3995 & n16285 ;
  assign n28390 = n28389 ^ n9072 ^ 1'b0 ;
  assign n28391 = n17677 ^ n17333 ^ 1'b0 ;
  assign n28392 = n4547 | n28391 ;
  assign n28393 = n7982 & n9540 ;
  assign n28397 = n5719 ^ n781 ^ 1'b0 ;
  assign n28394 = x125 & n16860 ;
  assign n28395 = n28394 ^ n1332 ^ 1'b0 ;
  assign n28396 = n28395 ^ n4271 ^ 1'b0 ;
  assign n28398 = n28397 ^ n28396 ^ 1'b0 ;
  assign n28399 = n9942 ^ n7828 ^ n4385 ;
  assign n28400 = n10900 & n28399 ;
  assign n28401 = n28400 ^ n3749 ^ 1'b0 ;
  assign n28402 = n1023 | n3454 ;
  assign n28403 = ~n14289 & n28402 ;
  assign n28404 = n2214 | n11191 ;
  assign n28405 = n28404 ^ n4480 ^ 1'b0 ;
  assign n28406 = n9949 & n23326 ;
  assign n28411 = n18454 ^ n688 ^ x251 ;
  assign n28409 = n2901 | n11169 ;
  assign n28410 = n28409 ^ n14017 ^ 1'b0 ;
  assign n28407 = n17081 | n17468 ;
  assign n28408 = n28407 ^ n12112 ^ 1'b0 ;
  assign n28412 = n28411 ^ n28410 ^ n28408 ;
  assign n28413 = n369 & ~n5178 ;
  assign n28414 = n28413 ^ n11124 ^ 1'b0 ;
  assign n28415 = n26244 ^ n18424 ^ 1'b0 ;
  assign n28416 = n8370 & n21419 ;
  assign n28417 = n13503 & n19575 ;
  assign n28418 = ~n10949 & n20603 ;
  assign n28419 = n28417 & n28418 ;
  assign n28420 = n5402 | n8912 ;
  assign n28421 = n28420 ^ n15572 ^ 1'b0 ;
  assign n28422 = n28419 & ~n28421 ;
  assign n28423 = ~n23783 & n28422 ;
  assign n28424 = ( n681 & n2038 ) | ( n681 & n9865 ) | ( n2038 & n9865 ) ;
  assign n28425 = n28296 ^ n9506 ^ 1'b0 ;
  assign n28426 = n13046 | n28425 ;
  assign n28427 = n28012 & ~n28426 ;
  assign n28428 = ~n2345 & n28427 ;
  assign n28429 = n1666 ^ n512 ^ 1'b0 ;
  assign n28430 = n13552 | n28429 ;
  assign n28431 = n7362 | n14876 ;
  assign n28432 = ~n6601 & n16534 ;
  assign n28433 = n23511 | n28432 ;
  assign n28434 = n27818 | n28433 ;
  assign n28435 = ( n366 & ~n453 ) | ( n366 & n10093 ) | ( ~n453 & n10093 ) ;
  assign n28436 = ( n4073 & n7915 ) | ( n4073 & n28435 ) | ( n7915 & n28435 ) ;
  assign n28437 = n16981 ^ n11183 ^ 1'b0 ;
  assign n28438 = ~n5677 & n28437 ;
  assign n28439 = ( ~n10512 & n28436 ) | ( ~n10512 & n28438 ) | ( n28436 & n28438 ) ;
  assign n28440 = n2206 & n6528 ;
  assign n28441 = n28440 ^ n26539 ^ 1'b0 ;
  assign n28443 = n5008 ^ n4312 ^ 1'b0 ;
  assign n28442 = n1491 & ~n15496 ;
  assign n28444 = n28443 ^ n28442 ^ 1'b0 ;
  assign n28445 = n7080 ^ n2402 ^ 1'b0 ;
  assign n28446 = n11966 ^ n11780 ^ 1'b0 ;
  assign n28447 = n9456 | n26422 ;
  assign n28448 = n28447 ^ n24775 ^ 1'b0 ;
  assign n28449 = n404 & n5752 ;
  assign n28450 = n28449 ^ n4171 ^ n4050 ;
  assign n28451 = ( n9844 & n13715 ) | ( n9844 & n19198 ) | ( n13715 & n19198 ) ;
  assign n28452 = n1768 & n8844 ;
  assign n28453 = n28452 ^ n25619 ^ n4094 ;
  assign n28454 = n28453 ^ n13543 ^ 1'b0 ;
  assign n28455 = n4242 ^ n3308 ^ 1'b0 ;
  assign n28456 = n18748 & n28455 ;
  assign n28457 = n673 | n6923 ;
  assign n28458 = n22289 & ~n28457 ;
  assign n28459 = ~n28456 & n28458 ;
  assign n28460 = n21057 ^ n13141 ^ 1'b0 ;
  assign n28463 = n14909 ^ n1415 ^ 1'b0 ;
  assign n28461 = n9545 ^ n9289 ^ 1'b0 ;
  assign n28462 = n4146 | n28461 ;
  assign n28464 = n28463 ^ n28462 ^ 1'b0 ;
  assign n28465 = n28460 & ~n28464 ;
  assign n28466 = n14994 ^ n3001 ^ 1'b0 ;
  assign n28467 = n6709 & n28466 ;
  assign n28468 = n25343 ^ x141 ^ 1'b0 ;
  assign n28469 = ( ~n353 & n5143 ) | ( ~n353 & n6447 ) | ( n5143 & n6447 ) ;
  assign n28470 = n10464 ^ n5077 ^ n1961 ;
  assign n28471 = n28470 ^ n20541 ^ n5303 ;
  assign n28472 = n1809 | n28471 ;
  assign n28473 = n8223 | n9178 ;
  assign n28474 = n28473 ^ n15450 ^ 1'b0 ;
  assign n28475 = n10424 | n28474 ;
  assign n28476 = n10366 ^ n9720 ^ 1'b0 ;
  assign n28477 = n28476 ^ n26740 ^ n8062 ;
  assign n28478 = n10203 ^ n9101 ^ 1'b0 ;
  assign n28479 = n432 | n7700 ;
  assign n28480 = n28479 ^ n3415 ^ 1'b0 ;
  assign n28481 = n28478 & n28480 ;
  assign n28482 = n10109 & n28481 ;
  assign n28483 = n28482 ^ n6305 ^ 1'b0 ;
  assign n28484 = n23560 ^ n12557 ^ 1'b0 ;
  assign n28485 = ~n12578 & n28438 ;
  assign n28486 = n23401 ^ n19753 ^ 1'b0 ;
  assign n28487 = n28485 & ~n28486 ;
  assign n28488 = ~n8793 & n25061 ;
  assign n28489 = n28488 ^ n4795 ^ 1'b0 ;
  assign n28490 = x253 & ~n28489 ;
  assign n28491 = n28490 ^ n18531 ^ 1'b0 ;
  assign n28492 = n16233 & n27494 ;
  assign n28493 = ~n12633 & n24043 ;
  assign n28494 = ~n8058 & n17708 ;
  assign n28495 = n28494 ^ n19467 ^ 1'b0 ;
  assign n28496 = n21856 | n28495 ;
  assign n28497 = n8271 | n28496 ;
  assign n28498 = ( x166 & n1279 ) | ( x166 & n3845 ) | ( n1279 & n3845 ) ;
  assign n28499 = ( n1079 & n17591 ) | ( n1079 & ~n25039 ) | ( n17591 & ~n25039 ) ;
  assign n28500 = ~n3481 & n4355 ;
  assign n28501 = n417 & n28500 ;
  assign n28502 = ~n19594 & n28501 ;
  assign n28503 = n23768 ^ n23494 ^ 1'b0 ;
  assign n28504 = n23901 | n28503 ;
  assign n28505 = ~n9392 & n13950 ;
  assign n28506 = n28505 ^ n5920 ^ 1'b0 ;
  assign n28507 = n7881 | n12238 ;
  assign n28508 = n12881 & ~n28507 ;
  assign n28509 = n24084 ^ n14454 ^ n5942 ;
  assign n28510 = ( n13366 & ~n28508 ) | ( n13366 & n28509 ) | ( ~n28508 & n28509 ) ;
  assign n28511 = n28510 ^ n25229 ^ 1'b0 ;
  assign n28512 = ~n28506 & n28511 ;
  assign n28513 = n16207 & ~n28512 ;
  assign n28514 = ( ~n1768 & n13313 ) | ( ~n1768 & n24228 ) | ( n13313 & n24228 ) ;
  assign n28515 = n24126 & ~n24407 ;
  assign n28516 = ~n648 & n10211 ;
  assign n28517 = n28516 ^ n4615 ^ 1'b0 ;
  assign n28518 = ~n10520 & n28517 ;
  assign n28519 = n15523 ^ n6313 ^ 1'b0 ;
  assign n28520 = n9813 & ~n28519 ;
  assign n28521 = n7476 & n28520 ;
  assign n28522 = n24252 & n28521 ;
  assign n28523 = n6548 | n13314 ;
  assign n28524 = ( ~n3777 & n4326 ) | ( ~n3777 & n22398 ) | ( n4326 & n22398 ) ;
  assign n28525 = n1208 | n1777 ;
  assign n28526 = n28525 ^ n3732 ^ 1'b0 ;
  assign n28527 = n28526 ^ n17350 ^ n1527 ;
  assign n28528 = x179 | n13580 ;
  assign n28529 = n28528 ^ n5988 ^ n1791 ;
  assign n28530 = ( n2224 & ~n5319 ) | ( n2224 & n14429 ) | ( ~n5319 & n14429 ) ;
  assign n28531 = n28530 ^ n11283 ^ 1'b0 ;
  assign n28532 = n23115 & n28531 ;
  assign n28533 = ~n28529 & n28532 ;
  assign n28534 = n9317 & ~n17527 ;
  assign n28535 = n28534 ^ n14986 ^ 1'b0 ;
  assign n28536 = n28535 ^ n28156 ^ 1'b0 ;
  assign n28537 = n28536 ^ n15585 ^ n11466 ;
  assign n28538 = n557 | n2462 ;
  assign n28539 = n2483 | n28538 ;
  assign n28540 = n4196 | n21274 ;
  assign n28541 = n9644 | n28540 ;
  assign n28542 = n13533 & ~n14972 ;
  assign n28543 = ~n28541 & n28542 ;
  assign n28544 = n10744 ^ n8246 ^ 1'b0 ;
  assign n28545 = n11467 & n28544 ;
  assign n28546 = n28545 ^ n18202 ^ 1'b0 ;
  assign n28547 = n18173 ^ n1024 ^ 1'b0 ;
  assign n28548 = n533 ^ x195 ^ 1'b0 ;
  assign n28549 = ~n6348 & n28548 ;
  assign n28550 = n5647 & ~n28549 ;
  assign n28551 = n25211 & n28550 ;
  assign n28553 = n10154 ^ n3016 ^ 1'b0 ;
  assign n28554 = n4119 & n20643 ;
  assign n28555 = n28553 & n28554 ;
  assign n28552 = n10053 ^ n9437 ^ 1'b0 ;
  assign n28556 = n28555 ^ n28552 ^ 1'b0 ;
  assign n28557 = n7235 & ~n8897 ;
  assign n28558 = n15018 & n28557 ;
  assign n28559 = n28558 ^ n20263 ^ n2816 ;
  assign n28561 = ~n798 & n8176 ;
  assign n28562 = n2120 & n28561 ;
  assign n28560 = n8151 | n17287 ;
  assign n28563 = n28562 ^ n28560 ^ n6668 ;
  assign n28564 = n12012 ^ n7008 ^ 1'b0 ;
  assign n28565 = n28564 ^ n28443 ^ n12261 ;
  assign n28566 = n12808 ^ n9282 ^ 1'b0 ;
  assign n28567 = n19633 | n28566 ;
  assign n28568 = n2656 | n20261 ;
  assign n28569 = n18045 & ~n28568 ;
  assign n28570 = n6953 & n22064 ;
  assign n28571 = n5537 & n28570 ;
  assign n28572 = n22413 & ~n24781 ;
  assign n28573 = ~n21434 & n28572 ;
  assign n28574 = n17524 & n20580 ;
  assign n28575 = n8539 | n21028 ;
  assign n28576 = ~n15240 & n28575 ;
  assign n28577 = n25480 ^ n20187 ^ 1'b0 ;
  assign n28578 = ~n28576 & n28577 ;
  assign n28579 = n18101 ^ n6303 ^ 1'b0 ;
  assign n28580 = n28579 ^ n4289 ^ 1'b0 ;
  assign n28581 = n3769 & n18376 ;
  assign n28582 = n19695 & n28581 ;
  assign n28583 = n21692 ^ n8205 ^ 1'b0 ;
  assign n28585 = n25109 ^ n18735 ^ 1'b0 ;
  assign n28584 = n5840 | n20362 ;
  assign n28586 = n28585 ^ n28584 ^ 1'b0 ;
  assign n28587 = n4242 ^ n1571 ^ 1'b0 ;
  assign n28588 = ~n22056 & n28587 ;
  assign n28589 = n28588 ^ n22392 ^ n10429 ;
  assign n28590 = n2918 & n28589 ;
  assign n28591 = n3241 & ~n9084 ;
  assign n28592 = n18589 & ~n28591 ;
  assign n28593 = n28592 ^ n7966 ^ 1'b0 ;
  assign n28594 = n7080 ^ n6684 ^ 1'b0 ;
  assign n28595 = n7260 & ~n28594 ;
  assign n28596 = ~n3008 & n25390 ;
  assign n28597 = n28596 ^ n17106 ^ 1'b0 ;
  assign n28598 = ~n7083 & n12393 ;
  assign n28599 = n28598 ^ n9575 ^ 1'b0 ;
  assign n28600 = n14798 ^ n2706 ^ 1'b0 ;
  assign n28601 = ~n9646 & n14677 ;
  assign n28602 = n4060 & n28601 ;
  assign n28603 = n12341 | n14122 ;
  assign n28604 = n28603 ^ n5590 ^ 1'b0 ;
  assign n28605 = ~n10553 & n18757 ;
  assign n28606 = n28605 ^ n3301 ^ 1'b0 ;
  assign n28607 = n11913 & ~n28606 ;
  assign n28608 = n28607 ^ n19422 ^ 1'b0 ;
  assign n28609 = n28604 & n28608 ;
  assign n28610 = n4541 & n15869 ;
  assign n28611 = n24066 ^ n21367 ^ 1'b0 ;
  assign n28612 = n14719 & n28611 ;
  assign n28613 = n28612 ^ n14262 ^ 1'b0 ;
  assign n28614 = n1524 & n28613 ;
  assign n28615 = n26111 ^ n1777 ^ 1'b0 ;
  assign n28616 = n14835 ^ n3951 ^ n1526 ;
  assign n28617 = x158 & ~n8055 ;
  assign n28618 = n28617 ^ n877 ^ 1'b0 ;
  assign n28619 = n16262 ^ n1271 ^ 1'b0 ;
  assign n28620 = n28618 & n28619 ;
  assign n28621 = n28616 & n28620 ;
  assign n28622 = n28621 ^ n10214 ^ 1'b0 ;
  assign n28623 = n13487 ^ n6683 ^ n1865 ;
  assign n28624 = ( ~n15924 & n25607 ) | ( ~n15924 & n27917 ) | ( n25607 & n27917 ) ;
  assign n28625 = n1192 | n12749 ;
  assign n28626 = n2555 & n3292 ;
  assign n28627 = ( n2735 & ~n15893 ) | ( n2735 & n28626 ) | ( ~n15893 & n28626 ) ;
  assign n28628 = n28627 ^ n15629 ^ 1'b0 ;
  assign n28629 = n26140 ^ n6713 ^ 1'b0 ;
  assign n28630 = ~n17595 & n18996 ;
  assign n28633 = n12744 ^ n11864 ^ 1'b0 ;
  assign n28631 = n11415 ^ n6614 ^ 1'b0 ;
  assign n28632 = n20243 & ~n28631 ;
  assign n28634 = n28633 ^ n28632 ^ n6526 ;
  assign n28635 = n12885 ^ n8201 ^ n5934 ;
  assign n28636 = ~n5257 & n15659 ;
  assign n28637 = n28636 ^ n5461 ^ 1'b0 ;
  assign n28638 = ~n18924 & n28637 ;
  assign n28639 = n28638 ^ n5038 ^ 1'b0 ;
  assign n28640 = n7277 & ~n11371 ;
  assign n28641 = n10839 & ~n27581 ;
  assign n28642 = ~n28640 & n28641 ;
  assign n28643 = n28642 ^ n11657 ^ 1'b0 ;
  assign n28644 = n26244 ^ n5369 ^ 1'b0 ;
  assign n28645 = n28643 & n28644 ;
  assign n28646 = n3543 & ~n6831 ;
  assign n28647 = n16604 | n28646 ;
  assign n28648 = n28647 ^ n5016 ^ 1'b0 ;
  assign n28649 = n1145 & n18942 ;
  assign n28650 = n1285 & n28649 ;
  assign n28651 = ( n28001 & ~n28648 ) | ( n28001 & n28650 ) | ( ~n28648 & n28650 ) ;
  assign n28652 = n24502 ^ n20119 ^ n8830 ;
  assign n28653 = n17666 | n25456 ;
  assign n28654 = ~n9666 & n28653 ;
  assign n28655 = ~n2047 & n28654 ;
  assign n28656 = n12627 ^ n7734 ^ 1'b0 ;
  assign n28657 = n28656 ^ n11446 ^ 1'b0 ;
  assign n28658 = n18296 & ~n28657 ;
  assign n28659 = n11133 & ~n26318 ;
  assign n28660 = n18473 & n28659 ;
  assign n28661 = n15668 | n16367 ;
  assign n28662 = n28660 & ~n28661 ;
  assign n28663 = n18618 & ~n24504 ;
  assign n28664 = ~n19285 & n28663 ;
  assign n28665 = n10411 & n28664 ;
  assign n28666 = n20768 ^ n8503 ^ n4529 ;
  assign n28667 = n2687 | n28666 ;
  assign n28668 = n28470 ^ n5057 ^ n3451 ;
  assign n28669 = n989 | n8955 ;
  assign n28670 = n21681 & ~n28669 ;
  assign n28672 = n9874 & ~n26574 ;
  assign n28673 = n2653 & n28672 ;
  assign n28671 = n2853 & n3700 ;
  assign n28674 = n28673 ^ n28671 ^ 1'b0 ;
  assign n28675 = n7336 ^ n2209 ^ 1'b0 ;
  assign n28676 = n28674 & n28675 ;
  assign n28677 = n2962 & ~n28676 ;
  assign n28678 = ( n516 & n1739 ) | ( n516 & n28677 ) | ( n1739 & n28677 ) ;
  assign n28679 = n28670 | n28678 ;
  assign n28680 = n26548 ^ n12576 ^ 1'b0 ;
  assign n28681 = ( ~n5356 & n9015 ) | ( ~n5356 & n16002 ) | ( n9015 & n16002 ) ;
  assign n28682 = n28680 & n28681 ;
  assign n28683 = ~n3586 & n14095 ;
  assign n28684 = x221 & n28683 ;
  assign n28685 = n28682 & n28684 ;
  assign n28686 = n9255 | n28685 ;
  assign n28687 = ~n8775 & n11857 ;
  assign n28688 = n2810 | n28687 ;
  assign n28689 = n28688 ^ n6119 ^ 1'b0 ;
  assign n28690 = n28689 ^ n21153 ^ 1'b0 ;
  assign n28691 = n21069 | n28690 ;
  assign n28692 = n13679 ^ n3095 ^ 1'b0 ;
  assign n28693 = n28692 ^ n1249 ^ 1'b0 ;
  assign n28697 = n5546 | n25765 ;
  assign n28696 = ( n12977 & ~n15939 ) | ( n12977 & n20771 ) | ( ~n15939 & n20771 ) ;
  assign n28698 = n28697 ^ n28696 ^ n12934 ;
  assign n28694 = n6060 | n9398 ;
  assign n28695 = n22285 | n28694 ;
  assign n28699 = n28698 ^ n28695 ^ 1'b0 ;
  assign n28700 = ~n4607 & n10882 ;
  assign n28701 = n28700 ^ n17499 ^ 1'b0 ;
  assign n28702 = ~n4826 & n6537 ;
  assign n28703 = n28702 ^ n2210 ^ 1'b0 ;
  assign n28704 = n8179 & n28703 ;
  assign n28705 = n10371 ^ n1464 ^ 1'b0 ;
  assign n28706 = n4491 & ~n28705 ;
  assign n28707 = ( n14286 & n28704 ) | ( n14286 & n28706 ) | ( n28704 & n28706 ) ;
  assign n28708 = n19791 ^ n8283 ^ 1'b0 ;
  assign n28709 = n8370 & n28708 ;
  assign n28710 = n17958 & ~n21109 ;
  assign n28711 = n28710 ^ n7067 ^ 1'b0 ;
  assign n28712 = n28711 ^ n10097 ^ 1'b0 ;
  assign n28713 = n5720 | n28712 ;
  assign n28714 = n17398 & ~n28713 ;
  assign n28715 = n28714 ^ n1192 ^ 1'b0 ;
  assign n28716 = n18591 & n18660 ;
  assign n28717 = n14408 & n28716 ;
  assign n28718 = n12937 & ~n17969 ;
  assign n28719 = n9616 & n27378 ;
  assign n28720 = n28719 ^ n358 ^ 1'b0 ;
  assign n28721 = n580 & n28720 ;
  assign n28722 = n7887 ^ n5703 ^ 1'b0 ;
  assign n28723 = n17395 & ~n28722 ;
  assign n28724 = n570 & n20514 ;
  assign n28725 = n18047 ^ n14887 ^ 1'b0 ;
  assign n28726 = n28725 ^ n15161 ^ 1'b0 ;
  assign n28727 = n6884 & ~n14122 ;
  assign n28728 = n28727 ^ n18593 ^ 1'b0 ;
  assign n28729 = ~n9514 & n10374 ;
  assign n28730 = n22885 ^ n5304 ^ 1'b0 ;
  assign n28731 = ~n7783 & n28730 ;
  assign n28732 = n25533 & n28731 ;
  assign n28733 = n28729 & n28732 ;
  assign n28734 = n4547 ^ n3933 ^ n3195 ;
  assign n28735 = n15175 & n19891 ;
  assign n28736 = n28734 & n28735 ;
  assign n28737 = n11529 ^ n1521 ^ 1'b0 ;
  assign n28738 = ~n6856 & n28737 ;
  assign n28739 = n12815 & n20847 ;
  assign n28740 = ~n3954 & n28739 ;
  assign n28741 = ~n1177 & n28740 ;
  assign n28742 = n6047 & ~n8900 ;
  assign n28743 = n19841 ^ n10763 ^ 1'b0 ;
  assign n28744 = n5135 & ~n12183 ;
  assign n28745 = ( n7298 & ~n8813 ) | ( n7298 & n28744 ) | ( ~n8813 & n28744 ) ;
  assign n28746 = n8295 ^ n4007 ^ 1'b0 ;
  assign n28747 = ~n28745 & n28746 ;
  assign n28748 = n28747 ^ n27796 ^ 1'b0 ;
  assign n28749 = n27680 | n28748 ;
  assign n28750 = ( n3384 & n6884 ) | ( n3384 & n9286 ) | ( n6884 & n9286 ) ;
  assign n28751 = n1967 | n23452 ;
  assign n28752 = n28751 ^ n1442 ^ 1'b0 ;
  assign n28753 = n7420 | n12429 ;
  assign n28754 = n7097 & n7448 ;
  assign n28755 = n28754 ^ n1879 ^ 1'b0 ;
  assign n28756 = n21838 ^ n15719 ^ 1'b0 ;
  assign n28757 = ~n28755 & n28756 ;
  assign n28758 = n2355 & ~n9530 ;
  assign n28759 = ~n28757 & n28758 ;
  assign n28760 = n666 & ~n26871 ;
  assign n28761 = n19876 & n28760 ;
  assign n28762 = ( n10166 & n24147 ) | ( n10166 & ~n26525 ) | ( n24147 & ~n26525 ) ;
  assign n28763 = ~x119 & n19721 ;
  assign n28764 = ~n6962 & n18518 ;
  assign n28765 = n28764 ^ n23087 ^ 1'b0 ;
  assign n28766 = ( n1242 & n4986 ) | ( n1242 & n22242 ) | ( n4986 & n22242 ) ;
  assign n28767 = ~n12538 & n27411 ;
  assign n28768 = ~x165 & n28767 ;
  assign n28769 = n22338 ^ n7088 ^ 1'b0 ;
  assign n28770 = n1228 | n12006 ;
  assign n28771 = n15550 ^ n12882 ^ n1370 ;
  assign n28772 = ( n6636 & n24177 ) | ( n6636 & ~n25631 ) | ( n24177 & ~n25631 ) ;
  assign n28773 = n20035 ^ n14002 ^ 1'b0 ;
  assign n28774 = n8813 & ~n28773 ;
  assign n28775 = n21851 | n26756 ;
  assign n28776 = n6892 | n28775 ;
  assign n28777 = n19688 ^ n18270 ^ 1'b0 ;
  assign n28778 = ~n6602 & n28777 ;
  assign n28779 = n697 & n12525 ;
  assign n28780 = ( n1665 & n28501 ) | ( n1665 & ~n28779 ) | ( n28501 & ~n28779 ) ;
  assign n28781 = n13725 ^ n1214 ^ 1'b0 ;
  assign n28782 = n28780 | n28781 ;
  assign n28784 = ( ~n18874 & n20635 ) | ( ~n18874 & n23936 ) | ( n20635 & n23936 ) ;
  assign n28785 = n26789 & ~n28784 ;
  assign n28786 = n28785 ^ n9640 ^ 1'b0 ;
  assign n28783 = n11281 | n24876 ;
  assign n28787 = n28786 ^ n28783 ^ 1'b0 ;
  assign n28788 = ( ~n2489 & n9073 ) | ( ~n2489 & n13649 ) | ( n9073 & n13649 ) ;
  assign n28789 = n28788 ^ n22346 ^ 1'b0 ;
  assign n28790 = n28789 ^ n20957 ^ n15793 ;
  assign n28791 = n998 & n1358 ;
  assign n28792 = ( n11755 & n24451 ) | ( n11755 & ~n28791 ) | ( n24451 & ~n28791 ) ;
  assign n28794 = n8119 ^ n6246 ^ 1'b0 ;
  assign n28793 = ~n1856 & n2829 ;
  assign n28795 = n28794 ^ n28793 ^ 1'b0 ;
  assign n28796 = n1991 & n7668 ;
  assign n28797 = n28796 ^ n19602 ^ 1'b0 ;
  assign n28798 = n3617 ^ x187 ^ 1'b0 ;
  assign n28799 = ~n760 & n28480 ;
  assign n28800 = n28799 ^ n11686 ^ 1'b0 ;
  assign n28801 = n28798 & ~n28800 ;
  assign n28802 = n28801 ^ n1741 ^ 1'b0 ;
  assign n28803 = n16494 ^ n5769 ^ n4473 ;
  assign n28804 = n1697 | n5085 ;
  assign n28805 = n28804 ^ n5952 ^ 1'b0 ;
  assign n28806 = ~n12317 & n28805 ;
  assign n28807 = ( ~n1180 & n28803 ) | ( ~n1180 & n28806 ) | ( n28803 & n28806 ) ;
  assign n28808 = ( n10512 & ~n13448 ) | ( n10512 & n15548 ) | ( ~n13448 & n15548 ) ;
  assign n28809 = n28808 ^ n15369 ^ 1'b0 ;
  assign n28810 = n15920 ^ n1709 ^ 1'b0 ;
  assign n28811 = ~n26633 & n28810 ;
  assign n28812 = n643 | n11910 ;
  assign n28813 = n28812 ^ n23265 ^ n16683 ;
  assign n28814 = ~n7469 & n28813 ;
  assign n28815 = n28814 ^ n19055 ^ 1'b0 ;
  assign n28816 = n20098 ^ n11153 ^ n4182 ;
  assign n28817 = n8256 | n22191 ;
  assign n28818 = n27404 ^ n7367 ^ n7007 ;
  assign n28819 = n2226 | n5067 ;
  assign n28820 = n17416 ^ n3403 ^ 1'b0 ;
  assign n28821 = ~n28819 & n28820 ;
  assign n28822 = n28588 ^ n6361 ^ 1'b0 ;
  assign n28823 = n7523 & n28822 ;
  assign n28824 = n22912 & n28823 ;
  assign n28825 = n28824 ^ n10701 ^ 1'b0 ;
  assign n28826 = n18109 | n24252 ;
  assign n28827 = n25355 | n28826 ;
  assign n28828 = n28827 ^ n13542 ^ 1'b0 ;
  assign n28829 = n11442 ^ n4073 ^ 1'b0 ;
  assign n28830 = n28828 | n28829 ;
  assign n28831 = n22348 ^ n401 ^ 1'b0 ;
  assign n28832 = n21928 ^ n20165 ^ n7587 ;
  assign n28833 = ~n2172 & n25940 ;
  assign n28834 = n20738 & n28833 ;
  assign n28835 = n28832 | n28834 ;
  assign n28836 = n28831 & ~n28835 ;
  assign n28837 = ~n4034 & n7214 ;
  assign n28838 = n6745 & n28837 ;
  assign n28839 = n5366 & ~n28838 ;
  assign n28840 = n8912 ^ n4804 ^ 1'b0 ;
  assign n28841 = n5298 & ~n6770 ;
  assign n28842 = n28841 ^ n21495 ^ 1'b0 ;
  assign n28843 = n18886 & n23714 ;
  assign n28844 = ~n27315 & n28843 ;
  assign n28845 = n23377 ^ n1347 ^ 1'b0 ;
  assign n28846 = n22146 ^ n11133 ^ 1'b0 ;
  assign n28847 = n28845 & ~n28846 ;
  assign n28848 = n25773 ^ n14639 ^ 1'b0 ;
  assign n28849 = n28847 | n28848 ;
  assign n28850 = n6088 | n7383 ;
  assign n28851 = n28850 ^ n21326 ^ 1'b0 ;
  assign n28852 = n1038 | n13128 ;
  assign n28853 = n1776 & ~n1920 ;
  assign n28854 = n19631 ^ n19601 ^ n8367 ;
  assign n28855 = ( n17761 & n19909 ) | ( n17761 & ~n28854 ) | ( n19909 & ~n28854 ) ;
  assign n28856 = n19855 ^ n1024 ^ 1'b0 ;
  assign n28857 = n14493 ^ n9266 ^ 1'b0 ;
  assign n28858 = n28856 & ~n28857 ;
  assign n28859 = n28858 ^ n6896 ^ 1'b0 ;
  assign n28860 = n28859 ^ n16621 ^ 1'b0 ;
  assign n28861 = ~n2484 & n6389 ;
  assign n28862 = ~n9581 & n28861 ;
  assign n28863 = n28862 ^ n8200 ^ n7155 ;
  assign n28864 = n11383 & ~n16877 ;
  assign n28865 = ~n28863 & n28864 ;
  assign n28866 = n10759 & n28865 ;
  assign n28867 = n8121 | n28866 ;
  assign n28868 = n24247 | n28867 ;
  assign n28869 = n23869 ^ n20964 ^ 1'b0 ;
  assign n28870 = n17072 & n28869 ;
  assign n28871 = n28870 ^ n1277 ^ x244 ;
  assign n28878 = n4829 ^ n2967 ^ 1'b0 ;
  assign n28872 = n23869 ^ n11786 ^ n6705 ;
  assign n28873 = n28872 ^ n20645 ^ n11505 ;
  assign n28874 = n23962 | n28873 ;
  assign n28875 = n28874 ^ n3097 ^ 1'b0 ;
  assign n28876 = ~n4405 & n8194 ;
  assign n28877 = ~n28875 & n28876 ;
  assign n28879 = n28878 ^ n28877 ^ 1'b0 ;
  assign n28880 = n1423 | n18413 ;
  assign n28881 = n24831 | n28880 ;
  assign n28882 = n28881 ^ n25263 ^ n5341 ;
  assign n28883 = n18418 ^ n4808 ^ 1'b0 ;
  assign n28884 = ( n2548 & ~n7653 ) | ( n2548 & n23418 ) | ( ~n7653 & n23418 ) ;
  assign n28885 = n16769 | n28884 ;
  assign n28886 = n28885 ^ n27499 ^ n4582 ;
  assign n28887 = n28886 ^ n23954 ^ 1'b0 ;
  assign n28889 = ~x73 & n6892 ;
  assign n28890 = n21757 & n28889 ;
  assign n28888 = n11006 | n15722 ;
  assign n28891 = n28890 ^ n28888 ^ 1'b0 ;
  assign n28892 = n963 | n11147 ;
  assign n28893 = n15031 | n28892 ;
  assign n28894 = n28893 ^ n8009 ^ 1'b0 ;
  assign n28895 = n28891 | n28894 ;
  assign n28896 = n15713 ^ n9260 ^ 1'b0 ;
  assign n28897 = n8161 | n28896 ;
  assign n28898 = n11950 ^ n3293 ^ 1'b0 ;
  assign n28899 = n1619 & n28898 ;
  assign n28900 = n21949 & n28899 ;
  assign n28901 = n13441 ^ n1722 ^ 1'b0 ;
  assign n28902 = ~n19531 & n28901 ;
  assign n28903 = n21898 ^ n9552 ^ n8394 ;
  assign n28904 = n28903 ^ n3683 ^ 1'b0 ;
  assign n28905 = ~n28299 & n28904 ;
  assign n28906 = n6193 | n15128 ;
  assign n28907 = n2203 & ~n11722 ;
  assign n28908 = ( n7198 & n28906 ) | ( n7198 & ~n28907 ) | ( n28906 & ~n28907 ) ;
  assign n28909 = n8688 ^ n8100 ^ 1'b0 ;
  assign n28910 = n6596 & n28909 ;
  assign n28911 = n10661 ^ x42 ^ 1'b0 ;
  assign n28912 = n28910 & ~n28911 ;
  assign n28913 = n28912 ^ n19232 ^ n6697 ;
  assign n28914 = n27558 ^ n3782 ^ 1'b0 ;
  assign n28915 = n24870 & n28914 ;
  assign n28916 = n23456 & n28915 ;
  assign n28917 = n4723 | n13527 ;
  assign n28918 = n27144 & n28917 ;
  assign n28919 = n3903 & n28918 ;
  assign n28920 = n9241 | n28919 ;
  assign n28921 = n9666 ^ n886 ^ 1'b0 ;
  assign n28922 = n13556 ^ n7127 ^ 1'b0 ;
  assign n28923 = n11407 & ~n28922 ;
  assign n28924 = ~n872 & n16646 ;
  assign n28925 = x75 & n28924 ;
  assign n28926 = n8666 & n28925 ;
  assign n28927 = ~n9776 & n25758 ;
  assign n28928 = n18260 | n28927 ;
  assign n28929 = n28928 ^ n21638 ^ 1'b0 ;
  assign n28930 = n28875 ^ n21788 ^ n6969 ;
  assign n28931 = n10212 ^ n6709 ^ 1'b0 ;
  assign n28932 = n17769 ^ n5154 ^ 1'b0 ;
  assign n28933 = ~n11590 & n28932 ;
  assign n28934 = n28933 ^ n27788 ^ 1'b0 ;
  assign n28935 = n2390 & ~n6307 ;
  assign n28936 = n14510 | n28935 ;
  assign n28937 = n28936 ^ n6264 ^ 1'b0 ;
  assign n28938 = n28934 & n28937 ;
  assign n28939 = ~n3391 & n8083 ;
  assign n28940 = n28939 ^ n12630 ^ 1'b0 ;
  assign n28941 = n2449 & ~n7821 ;
  assign n28942 = ~n25619 & n28941 ;
  assign n28943 = n16542 | n28942 ;
  assign n28944 = n28943 ^ n22696 ^ 1'b0 ;
  assign n28945 = n17469 & ~n20392 ;
  assign n28946 = ~n12338 & n28945 ;
  assign n28947 = n28944 | n28946 ;
  assign n28948 = n6075 ^ n686 ^ 1'b0 ;
  assign n28949 = n13860 & ~n28948 ;
  assign n28950 = ~n16398 & n28949 ;
  assign n28951 = ( n1142 & n1155 ) | ( n1142 & ~n16557 ) | ( n1155 & ~n16557 ) ;
  assign n28952 = n11935 | n28951 ;
  assign n28953 = n23687 & ~n28952 ;
  assign n28954 = n17446 ^ n7573 ^ n463 ;
  assign n28955 = n1372 & ~n28954 ;
  assign n28956 = n17687 ^ n13802 ^ 1'b0 ;
  assign n28957 = n8948 & ~n10525 ;
  assign n28958 = ~x160 & n28957 ;
  assign n28959 = ( n1073 & n4450 ) | ( n1073 & ~n4879 ) | ( n4450 & ~n4879 ) ;
  assign n28960 = n1339 | n28959 ;
  assign n28961 = ~n2914 & n3024 ;
  assign n28962 = n2914 & n28961 ;
  assign n28964 = n5640 | n8148 ;
  assign n28965 = n8148 & ~n28964 ;
  assign n28963 = n15574 & n18724 ;
  assign n28966 = n28965 ^ n28963 ^ 1'b0 ;
  assign n28967 = ~n28962 & n28966 ;
  assign n28968 = ~n984 & n20868 ;
  assign n28969 = ~n2054 & n28968 ;
  assign n28970 = n28969 ^ n5129 ^ n2524 ;
  assign n28971 = n1930 | n10314 ;
  assign n28972 = n28971 ^ n4335 ^ 1'b0 ;
  assign n28973 = n28972 ^ n4499 ^ n3625 ;
  assign n28974 = ~n9751 & n26884 ;
  assign n28975 = ~n28973 & n28974 ;
  assign n28976 = n4066 | n8280 ;
  assign n28977 = n10016 & ~n28976 ;
  assign n28978 = n28975 & n28977 ;
  assign n28979 = ~n13195 & n26005 ;
  assign n28980 = n17122 & n28979 ;
  assign n28981 = n5341 | n6480 ;
  assign n28982 = n28981 ^ n19733 ^ 1'b0 ;
  assign n28983 = n28982 ^ n19087 ^ 1'b0 ;
  assign n28984 = n14891 ^ n679 ^ 1'b0 ;
  assign n28985 = n19510 ^ n5849 ^ 1'b0 ;
  assign n28986 = n7946 | n28985 ;
  assign n28987 = ( n2218 & ~n3905 ) | ( n2218 & n5418 ) | ( ~n3905 & n5418 ) ;
  assign n28988 = n7912 | n28987 ;
  assign n28989 = ~n7512 & n8386 ;
  assign n28990 = ~n4363 & n28989 ;
  assign n28991 = n19736 | n28990 ;
  assign n28992 = n14947 | n28991 ;
  assign n28993 = ~n6440 & n28992 ;
  assign n28994 = n20440 ^ n12635 ^ n12118 ;
  assign n28995 = n13036 ^ n5269 ^ 1'b0 ;
  assign n28996 = n12853 ^ n9475 ^ 1'b0 ;
  assign n28997 = ( n21419 & n28995 ) | ( n21419 & n28996 ) | ( n28995 & n28996 ) ;
  assign n28998 = n10653 ^ n2922 ^ 1'b0 ;
  assign n28999 = n28997 & n28998 ;
  assign n29000 = ( n963 & n20774 ) | ( n963 & ~n21787 ) | ( n20774 & ~n21787 ) ;
  assign n29001 = ( n11781 & n14697 ) | ( n11781 & ~n23168 ) | ( n14697 & ~n23168 ) ;
  assign n29002 = n5778 ^ n1741 ^ 1'b0 ;
  assign n29003 = ~n9942 & n29002 ;
  assign n29004 = n10590 & n28770 ;
  assign n29005 = n11509 & n29004 ;
  assign n29006 = x11 & ~n1995 ;
  assign n29007 = n29006 ^ n13220 ^ 1'b0 ;
  assign n29008 = n3926 | n29007 ;
  assign n29009 = ~n1880 & n4375 ;
  assign n29010 = n29009 ^ n14227 ^ 1'b0 ;
  assign n29011 = ~n3233 & n29010 ;
  assign n29012 = ~n2963 & n29011 ;
  assign n29013 = n29012 ^ n18718 ^ 1'b0 ;
  assign n29014 = ~n2234 & n29013 ;
  assign n29015 = ( n16803 & ~n29008 ) | ( n16803 & n29014 ) | ( ~n29008 & n29014 ) ;
  assign n29016 = n28203 ^ n11365 ^ n4553 ;
  assign n29018 = n1589 | n7934 ;
  assign n29019 = n29018 ^ n5577 ^ 1'b0 ;
  assign n29017 = n737 & n22665 ;
  assign n29020 = n29019 ^ n29017 ^ 1'b0 ;
  assign n29021 = n698 | n29020 ;
  assign n29022 = n3270 & n14589 ;
  assign n29023 = n6606 & n29022 ;
  assign n29024 = n16392 & ~n17178 ;
  assign n29026 = n18757 ^ n15955 ^ 1'b0 ;
  assign n29027 = n12685 | n29026 ;
  assign n29028 = n20952 & ~n29027 ;
  assign n29025 = n7356 & n12346 ;
  assign n29029 = n29028 ^ n29025 ^ n5083 ;
  assign n29030 = n19993 ^ n15311 ^ n7708 ;
  assign n29031 = n29030 ^ n21526 ^ n17230 ;
  assign n29032 = n25291 & n29031 ;
  assign n29033 = n18061 ^ n9502 ^ 1'b0 ;
  assign n29034 = n17775 ^ n16494 ^ n14006 ;
  assign n29035 = ~n29033 & n29034 ;
  assign n29036 = n6473 & ~n13363 ;
  assign n29037 = ~n22406 & n29036 ;
  assign n29038 = n5730 ^ n5242 ^ 1'b0 ;
  assign n29039 = n563 | n29038 ;
  assign n29040 = ~n12526 & n18427 ;
  assign n29041 = ~n16325 & n29040 ;
  assign n29042 = ( n9326 & ~n17313 ) | ( n9326 & n29041 ) | ( ~n17313 & n29041 ) ;
  assign n29043 = n9059 & n10963 ;
  assign n29044 = n29042 & n29043 ;
  assign n29046 = n2282 & n2791 ;
  assign n29045 = n6966 & n25537 ;
  assign n29047 = n29046 ^ n29045 ^ 1'b0 ;
  assign n29048 = ~n4096 & n18940 ;
  assign n29049 = n29048 ^ n4282 ^ 1'b0 ;
  assign n29050 = n27487 ^ n6831 ^ 1'b0 ;
  assign n29051 = n29050 ^ n12069 ^ 1'b0 ;
  assign n29052 = n5477 ^ n2194 ^ 1'b0 ;
  assign n29053 = n29052 ^ n24415 ^ 1'b0 ;
  assign n29055 = n14743 ^ n6739 ^ 1'b0 ;
  assign n29056 = n1158 & ~n29055 ;
  assign n29054 = n21000 ^ n7924 ^ n6614 ;
  assign n29057 = n29056 ^ n29054 ^ n26334 ;
  assign n29058 = n11640 | n19714 ;
  assign n29059 = n8643 & ~n26681 ;
  assign n29060 = n14338 ^ n11823 ^ 1'b0 ;
  assign n29061 = n17563 | n29060 ;
  assign n29062 = n13807 & n25570 ;
  assign n29063 = n29062 ^ n17873 ^ 1'b0 ;
  assign n29064 = ~n1858 & n18924 ;
  assign n29065 = ( n1218 & ~n2548 ) | ( n1218 & n4743 ) | ( ~n2548 & n4743 ) ;
  assign n29066 = n29065 ^ n15421 ^ 1'b0 ;
  assign n29067 = n3312 | n29066 ;
  assign n29068 = n24145 | n29067 ;
  assign n29069 = n27977 ^ n24955 ^ n23533 ;
  assign n29070 = n8530 | n10324 ;
  assign n29071 = n4643 | n29070 ;
  assign n29072 = ~n18385 & n29071 ;
  assign n29073 = n8497 & n9264 ;
  assign n29074 = ~x58 & n29073 ;
  assign n29075 = n29074 ^ n8044 ^ 1'b0 ;
  assign n29076 = n3804 | n29075 ;
  assign n29077 = n1181 & ~n3160 ;
  assign n29078 = n29076 & n29077 ;
  assign n29079 = n1479 & n8622 ;
  assign n29080 = n6385 ^ n1829 ^ 1'b0 ;
  assign n29081 = n27782 | n29080 ;
  assign n29082 = n29079 & ~n29081 ;
  assign n29083 = n29082 ^ n27907 ^ 1'b0 ;
  assign n29084 = ~n2476 & n7963 ;
  assign n29085 = n10657 & n29084 ;
  assign n29086 = n18805 ^ n16851 ^ 1'b0 ;
  assign n29087 = n15484 & ~n29086 ;
  assign n29088 = n28117 ^ n18808 ^ 1'b0 ;
  assign n29089 = n11686 & n29088 ;
  assign n29090 = ~n727 & n4120 ;
  assign n29091 = ~n4120 & n29090 ;
  assign n29092 = n16715 & n29091 ;
  assign n29097 = ~n824 & n5083 ;
  assign n29098 = n4369 & n29097 ;
  assign n29099 = n29098 ^ n11840 ^ 1'b0 ;
  assign n29093 = n11772 ^ n9330 ^ n4719 ;
  assign n29094 = n16416 ^ n10917 ^ 1'b0 ;
  assign n29095 = ~n29093 & n29094 ;
  assign n29096 = ~n7932 & n29095 ;
  assign n29100 = n29099 ^ n29096 ^ 1'b0 ;
  assign n29101 = n29092 | n29100 ;
  assign n29102 = n1601 | n29101 ;
  assign n29103 = n4858 ^ n3791 ^ 1'b0 ;
  assign n29104 = n5373 & n29103 ;
  assign n29105 = n18723 & ~n29104 ;
  assign n29109 = ~n3506 & n9953 ;
  assign n29106 = n18082 ^ n10385 ^ 1'b0 ;
  assign n29107 = n29106 ^ n10997 ^ n2394 ;
  assign n29108 = ~n24316 & n29107 ;
  assign n29110 = n29109 ^ n29108 ^ 1'b0 ;
  assign n29111 = n1590 & ~n11672 ;
  assign n29112 = n4371 | n9833 ;
  assign n29113 = n29112 ^ n3985 ^ 1'b0 ;
  assign n29114 = n23269 & ~n29113 ;
  assign n29115 = ( n17297 & n22809 ) | ( n17297 & n23751 ) | ( n22809 & n23751 ) ;
  assign n29116 = n29115 ^ n17506 ^ 1'b0 ;
  assign n29117 = ~n19287 & n29116 ;
  assign n29118 = n4614 ^ n4274 ^ 1'b0 ;
  assign n29123 = n18283 ^ n4775 ^ 1'b0 ;
  assign n29119 = n7013 & n22314 ;
  assign n29120 = n6778 & n29119 ;
  assign n29121 = n11536 | n29120 ;
  assign n29122 = n14324 | n29121 ;
  assign n29124 = n29123 ^ n29122 ^ n14079 ;
  assign n29125 = n10781 ^ n3518 ^ 1'b0 ;
  assign n29126 = n543 & ~n29125 ;
  assign n29127 = n2440 | n29126 ;
  assign n29128 = n10310 & n17243 ;
  assign n29129 = n29128 ^ n979 ^ 1'b0 ;
  assign n29130 = n372 & n20216 ;
  assign n29131 = n12279 | n29130 ;
  assign n29132 = n28680 ^ n7426 ^ n5538 ;
  assign n29133 = n15049 | n29132 ;
  assign n29134 = n2107 | n17516 ;
  assign n29135 = n29134 ^ n7334 ^ n4030 ;
  assign n29136 = ( n3859 & n24095 ) | ( n3859 & ~n24797 ) | ( n24095 & ~n24797 ) ;
  assign n29137 = n29136 ^ n14472 ^ 1'b0 ;
  assign n29138 = n7769 | n29137 ;
  assign n29139 = ( n4774 & n6555 ) | ( n4774 & ~n29138 ) | ( n6555 & ~n29138 ) ;
  assign n29140 = n9105 ^ n1285 ^ 1'b0 ;
  assign n29141 = n17034 ^ n4255 ^ n624 ;
  assign n29142 = n29141 ^ n21225 ^ 1'b0 ;
  assign n29143 = ~n29140 & n29142 ;
  assign n29144 = n29143 ^ n19508 ^ 1'b0 ;
  assign n29145 = n21343 ^ n16087 ^ 1'b0 ;
  assign n29146 = n29145 ^ n10488 ^ 1'b0 ;
  assign n29147 = n27759 & n29146 ;
  assign n29148 = n5514 | n27458 ;
  assign n29149 = n29147 | n29148 ;
  assign n29150 = n1421 & n13274 ;
  assign n29151 = n29150 ^ n8480 ^ 1'b0 ;
  assign n29152 = n29151 ^ n27614 ^ 1'b0 ;
  assign n29153 = n14439 | n24096 ;
  assign n29155 = n8815 ^ n2532 ^ 1'b0 ;
  assign n29156 = n29155 ^ n10484 ^ 1'b0 ;
  assign n29157 = ~n5730 & n29156 ;
  assign n29154 = ~n4931 & n8719 ;
  assign n29158 = n29157 ^ n29154 ^ 1'b0 ;
  assign n29159 = n29158 ^ n13475 ^ 1'b0 ;
  assign n29160 = n12600 & ~n12631 ;
  assign n29161 = n10237 | n27356 ;
  assign n29162 = n29161 ^ n2038 ^ 1'b0 ;
  assign n29163 = ( n5840 & ~n29160 ) | ( n5840 & n29162 ) | ( ~n29160 & n29162 ) ;
  assign n29164 = n29163 ^ n6381 ^ 1'b0 ;
  assign n29165 = n3670 & ~n19852 ;
  assign n29166 = n29165 ^ n26020 ^ 1'b0 ;
  assign n29167 = n28935 | n29166 ;
  assign n29168 = x174 & n7356 ;
  assign n29169 = n29168 ^ n5836 ^ 1'b0 ;
  assign n29170 = n17304 ^ n7685 ^ 1'b0 ;
  assign n29171 = ( n2483 & n21681 ) | ( n2483 & ~n29170 ) | ( n21681 & ~n29170 ) ;
  assign n29172 = n29169 & ~n29171 ;
  assign n29173 = n2821 | n19210 ;
  assign n29174 = n3193 | n29173 ;
  assign n29175 = ( n5246 & n15697 ) | ( n5246 & n29174 ) | ( n15697 & n29174 ) ;
  assign n29176 = ~n4531 & n29175 ;
  assign n29177 = ~n6309 & n17230 ;
  assign n29178 = n29177 ^ n10913 ^ 1'b0 ;
  assign n29179 = ( n9867 & n10305 ) | ( n9867 & ~n11357 ) | ( n10305 & ~n11357 ) ;
  assign n29180 = ~n5355 & n29179 ;
  assign n29181 = n14158 & n21295 ;
  assign n29182 = n28976 & n29181 ;
  assign n29183 = n7603 & ~n8695 ;
  assign n29184 = n29183 ^ n9551 ^ 1'b0 ;
  assign n29185 = ~n26508 & n29184 ;
  assign n29186 = n4707 ^ n2223 ^ 1'b0 ;
  assign n29187 = n731 | n29186 ;
  assign n29188 = ~n9500 & n29187 ;
  assign n29189 = n29188 ^ n10662 ^ n2276 ;
  assign n29190 = ( x247 & n4171 ) | ( x247 & ~n26247 ) | ( n4171 & ~n26247 ) ;
  assign n29191 = n4839 ^ n4548 ^ n3733 ;
  assign n29192 = n29191 ^ n24799 ^ 1'b0 ;
  assign n29193 = n5765 & n21089 ;
  assign n29194 = ( n4460 & n13009 ) | ( n4460 & ~n17591 ) | ( n13009 & ~n17591 ) ;
  assign n29195 = n4750 ^ n4521 ^ 1'b0 ;
  assign n29196 = n8187 & ~n29195 ;
  assign n29197 = n11929 ^ n1697 ^ 1'b0 ;
  assign n29198 = n13223 | n29197 ;
  assign n29199 = n15280 | n29198 ;
  assign n29200 = n29199 ^ n2184 ^ 1'b0 ;
  assign n29201 = n29200 ^ n3294 ^ 1'b0 ;
  assign n29202 = n14095 ^ n13162 ^ n4696 ;
  assign n29203 = n29202 ^ n19451 ^ 1'b0 ;
  assign n29204 = n7693 | n23044 ;
  assign n29205 = n29204 ^ n10378 ^ 1'b0 ;
  assign n29206 = n5981 | n19876 ;
  assign n29207 = n29206 ^ x106 ^ 1'b0 ;
  assign n29209 = n13309 ^ n2819 ^ x103 ;
  assign n29210 = n29209 ^ n1779 ^ 1'b0 ;
  assign n29208 = n8495 & ~n16454 ;
  assign n29211 = n29210 ^ n29208 ^ 1'b0 ;
  assign n29212 = n29211 ^ n1435 ^ 1'b0 ;
  assign n29213 = n29207 & n29212 ;
  assign n29214 = ~n6481 & n29213 ;
  assign n29215 = n1984 & n27709 ;
  assign n29216 = n29215 ^ n7861 ^ 1'b0 ;
  assign n29217 = n23845 ^ n1325 ^ 1'b0 ;
  assign n29218 = ( n10424 & ~n13231 ) | ( n10424 & n29217 ) | ( ~n13231 & n29217 ) ;
  assign n29219 = n1669 & n22452 ;
  assign n29220 = n29219 ^ n5694 ^ 1'b0 ;
  assign n29221 = n19944 & n29220 ;
  assign n29222 = n20036 & n29221 ;
  assign n29223 = n29222 ^ n692 ^ 1'b0 ;
  assign n29224 = n5666 & n29223 ;
  assign n29225 = n22983 ^ n5744 ^ 1'b0 ;
  assign n29226 = ~n12182 & n29225 ;
  assign n29227 = n6438 & ~n20958 ;
  assign n29228 = n29227 ^ n11284 ^ 1'b0 ;
  assign n29229 = n5710 | n6704 ;
  assign n29230 = n29229 ^ n17352 ^ 1'b0 ;
  assign n29231 = n2462 | n3907 ;
  assign n29232 = ( ~n5067 & n8691 ) | ( ~n5067 & n29231 ) | ( n8691 & n29231 ) ;
  assign n29233 = n23144 & n23628 ;
  assign n29234 = ~n28051 & n29233 ;
  assign n29235 = ~n1259 & n6544 ;
  assign n29236 = n14456 ^ n2739 ^ 1'b0 ;
  assign n29237 = ~n4887 & n8496 ;
  assign n29238 = n21369 & n29237 ;
  assign n29239 = n29238 ^ n12753 ^ 1'b0 ;
  assign n29240 = n4954 & n8999 ;
  assign n29241 = n24206 ^ n6253 ^ 1'b0 ;
  assign n29242 = n29240 & ~n29241 ;
  assign n29243 = n29242 ^ n8725 ^ n2420 ;
  assign n29244 = ~n9014 & n25889 ;
  assign n29245 = n17985 & n29244 ;
  assign n29247 = n2969 & ~n28711 ;
  assign n29246 = n1528 & ~n10685 ;
  assign n29248 = n29247 ^ n29246 ^ n20912 ;
  assign n29249 = n29248 ^ n16807 ^ n9028 ;
  assign n29250 = ~n5410 & n20603 ;
  assign n29251 = ~n2091 & n29250 ;
  assign n29252 = n11767 ^ n9067 ^ 1'b0 ;
  assign n29253 = ~n29251 & n29252 ;
  assign n29254 = ~n29249 & n29253 ;
  assign n29255 = n10262 | n21757 ;
  assign n29256 = n29255 ^ n6338 ^ 1'b0 ;
  assign n29257 = n20088 ^ x182 ^ 1'b0 ;
  assign n29258 = n29256 & n29257 ;
  assign n29259 = ~n9236 & n24818 ;
  assign n29260 = n25537 ^ n23546 ^ n5491 ;
  assign n29261 = ( n9900 & n10267 ) | ( n9900 & n12697 ) | ( n10267 & n12697 ) ;
  assign n29262 = ( ~n5755 & n19202 ) | ( ~n5755 & n29261 ) | ( n19202 & n29261 ) ;
  assign n29263 = n5381 ^ n2248 ^ 1'b0 ;
  assign n29264 = n29263 ^ n3061 ^ 1'b0 ;
  assign n29265 = n26486 ^ n8998 ^ 1'b0 ;
  assign n29266 = n26869 | n29265 ;
  assign n29267 = n4729 & n13778 ;
  assign n29268 = n27428 & n29267 ;
  assign n29269 = n27722 ^ n5452 ^ n1900 ;
  assign n29270 = n16489 & ~n29269 ;
  assign n29271 = n5646 & n17907 ;
  assign n29272 = n18258 & n29271 ;
  assign n29273 = ~n16408 & n16971 ;
  assign n29274 = n29273 ^ n26001 ^ 1'b0 ;
  assign n29276 = n5594 ^ n2824 ^ 1'b0 ;
  assign n29277 = n6281 & ~n29276 ;
  assign n29275 = n10405 ^ n10066 ^ 1'b0 ;
  assign n29278 = n29277 ^ n29275 ^ 1'b0 ;
  assign n29280 = n22206 ^ n8317 ^ n5125 ;
  assign n29279 = n20565 & n28072 ;
  assign n29281 = n29280 ^ n29279 ^ n3961 ;
  assign n29282 = n20392 ^ n4527 ^ 1'b0 ;
  assign n29283 = n6051 & n29282 ;
  assign n29284 = n29283 ^ n19276 ^ 1'b0 ;
  assign n29285 = n3231 & ~n9227 ;
  assign n29286 = n2806 | n5471 ;
  assign n29287 = n29286 ^ n5762 ^ 1'b0 ;
  assign n29288 = n29287 ^ n5830 ^ 1'b0 ;
  assign n29289 = ~n7394 & n29288 ;
  assign n29290 = n13883 ^ n4867 ^ 1'b0 ;
  assign n29291 = n29289 & n29290 ;
  assign n29292 = n29285 & n29291 ;
  assign n29293 = n7696 & n14584 ;
  assign n29294 = n15119 ^ n5006 ^ 1'b0 ;
  assign n29295 = n6970 & ~n29294 ;
  assign n29296 = n22869 & ~n23470 ;
  assign n29297 = ~n1475 & n26308 ;
  assign n29298 = n1475 & n29297 ;
  assign n29299 = n668 & n2194 ;
  assign n29300 = ~n668 & n29299 ;
  assign n29301 = n29300 ^ n8376 ^ 1'b0 ;
  assign n29302 = n29298 | n29301 ;
  assign n29303 = n29298 & ~n29302 ;
  assign n29304 = n1236 & n1587 ;
  assign n29305 = ~n1587 & n29304 ;
  assign n29306 = ~n1277 & n1677 ;
  assign n29307 = n1277 & n29306 ;
  assign n29308 = n1349 & ~n1974 ;
  assign n29309 = n29307 & n29308 ;
  assign n29310 = n1266 & n29309 ;
  assign n29311 = ~n29305 & n29310 ;
  assign n29312 = n21921 & n29311 ;
  assign n29313 = n29303 | n29312 ;
  assign n29314 = n15648 & ~n29313 ;
  assign n29315 = n7477 & n20918 ;
  assign n29316 = n13552 ^ n1194 ^ 1'b0 ;
  assign n29317 = n7428 & n20737 ;
  assign n29318 = n18718 ^ n12176 ^ 1'b0 ;
  assign n29319 = n27948 & n29318 ;
  assign n29320 = n3721 ^ n3326 ^ 1'b0 ;
  assign n29321 = n12604 ^ n2735 ^ 1'b0 ;
  assign n29322 = n11594 | n24269 ;
  assign n29323 = n11630 & ~n29322 ;
  assign n29324 = n16199 ^ n2047 ^ 1'b0 ;
  assign n29325 = ~n2838 & n29324 ;
  assign n29326 = n29325 ^ n9773 ^ 1'b0 ;
  assign n29327 = n1557 & n29326 ;
  assign n29328 = n29327 ^ n13725 ^ 1'b0 ;
  assign n29329 = n28347 ^ n11488 ^ 1'b0 ;
  assign n29330 = ~n7788 & n10911 ;
  assign n29331 = n2311 & ~n25986 ;
  assign n29332 = n8665 & n29331 ;
  assign n29333 = n29332 ^ n2371 ^ 1'b0 ;
  assign n29334 = n7962 | n10960 ;
  assign n29335 = n712 & ~n29334 ;
  assign n29336 = n29335 ^ n3702 ^ 1'b0 ;
  assign n29337 = n3782 & n29336 ;
  assign n29338 = ~n10958 & n19847 ;
  assign n29339 = n5798 & n29338 ;
  assign n29340 = n1651 & ~n5788 ;
  assign n29341 = n17560 & n29340 ;
  assign n29342 = n14414 & n16953 ;
  assign n29343 = ~n1036 & n8309 ;
  assign n29344 = n21494 ^ n3374 ^ 1'b0 ;
  assign n29345 = ~n21461 & n29344 ;
  assign n29346 = ~n29343 & n29345 ;
  assign n29347 = n29346 ^ n9141 ^ 1'b0 ;
  assign n29348 = n1073 & n5154 ;
  assign n29349 = n29347 & ~n29348 ;
  assign n29350 = n16868 ^ n407 ^ 1'b0 ;
  assign n29351 = n2286 & ~n29350 ;
  assign n29352 = n29351 ^ n8425 ^ 1'b0 ;
  assign n29353 = n7369 & ~n29352 ;
  assign n29354 = ~n347 & n24174 ;
  assign n29355 = n29354 ^ n14689 ^ 1'b0 ;
  assign n29356 = n8215 & n10132 ;
  assign n29357 = n29356 ^ n22380 ^ 1'b0 ;
  assign n29358 = n24272 ^ n21000 ^ n15054 ;
  assign n29359 = n14509 ^ n12974 ^ n5196 ;
  assign n29360 = n9526 | n25193 ;
  assign n29361 = n1166 | n2178 ;
  assign n29362 = n29361 ^ n2340 ^ 1'b0 ;
  assign n29363 = n29362 ^ n28119 ^ 1'b0 ;
  assign n29364 = n26867 ^ n20995 ^ 1'b0 ;
  assign n29365 = n20060 & ~n26866 ;
  assign n29366 = ~n16354 & n29365 ;
  assign n29367 = n4271 & n21280 ;
  assign n29369 = n3750 ^ n1473 ^ 1'b0 ;
  assign n29370 = n3918 & n29369 ;
  assign n29371 = n9548 | n29370 ;
  assign n29368 = ~n17272 & n26994 ;
  assign n29372 = n29371 ^ n29368 ^ 1'b0 ;
  assign n29373 = n1597 | n2967 ;
  assign n29374 = ~n18190 & n29373 ;
  assign n29375 = ~n1200 & n16732 ;
  assign n29376 = n29375 ^ n849 ^ 1'b0 ;
  assign n29377 = ( ~n14549 & n29374 ) | ( ~n14549 & n29376 ) | ( n29374 & n29376 ) ;
  assign n29378 = n7556 ^ n508 ^ 1'b0 ;
  assign n29379 = ~n10411 & n29378 ;
  assign n29380 = n19409 ^ n6019 ^ 1'b0 ;
  assign n29386 = x102 & ~n6213 ;
  assign n29387 = ~n12489 & n29386 ;
  assign n29388 = ~n5072 & n29387 ;
  assign n29382 = n1569 & n22079 ;
  assign n29383 = n20203 & n29382 ;
  assign n29384 = n29383 ^ n15276 ^ n5596 ;
  assign n29381 = n24909 ^ n9401 ^ n5584 ;
  assign n29385 = n29384 ^ n29381 ^ 1'b0 ;
  assign n29389 = n29388 ^ n29385 ^ 1'b0 ;
  assign n29390 = n9188 & n21271 ;
  assign n29391 = n29390 ^ x221 ^ 1'b0 ;
  assign n29392 = n3618 | n18096 ;
  assign n29393 = ( ~n5720 & n29391 ) | ( ~n5720 & n29392 ) | ( n29391 & n29392 ) ;
  assign n29395 = n8592 | n19326 ;
  assign n29394 = n15721 & ~n21908 ;
  assign n29396 = n29395 ^ n29394 ^ 1'b0 ;
  assign n29397 = n8556 & n10702 ;
  assign n29398 = ~n2248 & n29397 ;
  assign n29399 = n27350 & ~n28549 ;
  assign n29400 = n29398 & n29399 ;
  assign n29401 = n27481 ^ n2322 ^ 1'b0 ;
  assign n29402 = ~n1698 & n29401 ;
  assign n29403 = ~n28476 & n29402 ;
  assign n29404 = n29403 ^ n19131 ^ 1'b0 ;
  assign n29405 = ~n4714 & n6318 ;
  assign n29406 = ~n6810 & n29405 ;
  assign n29407 = n4951 ^ x18 ^ 1'b0 ;
  assign n29408 = n5113 | n29407 ;
  assign n29409 = n29408 ^ n12835 ^ n985 ;
  assign n29410 = n18228 ^ n15363 ^ 1'b0 ;
  assign n29411 = n8674 & n29410 ;
  assign n29412 = n16362 ^ n8078 ^ 1'b0 ;
  assign n29413 = ~n982 & n5678 ;
  assign n29414 = n6622 & n29413 ;
  assign n29415 = ~n5962 & n21182 ;
  assign n29416 = n29415 ^ x227 ^ 1'b0 ;
  assign n29417 = n22191 ^ n17855 ^ 1'b0 ;
  assign n29418 = n6462 & n19107 ;
  assign n29419 = n18378 ^ n10941 ^ 1'b0 ;
  assign n29420 = n7603 & ~n29419 ;
  assign n29421 = ~n24343 & n29420 ;
  assign n29422 = x48 | n1585 ;
  assign n29423 = n15442 ^ n2539 ^ 1'b0 ;
  assign n29424 = ~n26652 & n29423 ;
  assign n29425 = n3727 | n5173 ;
  assign n29426 = ( n29422 & ~n29424 ) | ( n29422 & n29425 ) | ( ~n29424 & n29425 ) ;
  assign n29427 = n28177 ^ n5678 ^ 1'b0 ;
  assign n29428 = n13340 | n29427 ;
  assign n29429 = n29428 ^ n11379 ^ n11198 ;
  assign n29430 = n13792 ^ n6327 ^ 1'b0 ;
  assign n29431 = n6131 | n19418 ;
  assign n29432 = n18449 | n29431 ;
  assign n29433 = n14996 & ~n29432 ;
  assign n29434 = n2014 & n18594 ;
  assign n29435 = ~n27739 & n29434 ;
  assign n29436 = n11941 | n12160 ;
  assign n29437 = n29436 ^ n22955 ^ 1'b0 ;
  assign n29441 = n8554 ^ n304 ^ 1'b0 ;
  assign n29442 = n15963 & ~n29441 ;
  assign n29438 = n12012 & n14396 ;
  assign n29439 = n29438 ^ n13040 ^ 1'b0 ;
  assign n29440 = n11833 & n29439 ;
  assign n29443 = n29442 ^ n29440 ^ x187 ;
  assign n29444 = ~n3504 & n8572 ;
  assign n29445 = ~n18648 & n29444 ;
  assign n29446 = n1344 & n6982 ;
  assign n29447 = n978 & n29446 ;
  assign n29448 = n29445 | n29447 ;
  assign n29449 = n5433 & ~n29448 ;
  assign n29450 = ~x178 & n2560 ;
  assign n29451 = n29450 ^ n23027 ^ 1'b0 ;
  assign n29452 = n9546 & ~n29451 ;
  assign n29453 = ~n731 & n23392 ;
  assign n29454 = n9087 & n20101 ;
  assign n29455 = n10512 & n29454 ;
  assign n29456 = n29455 ^ n25734 ^ n15784 ;
  assign n29458 = ~n7532 & n17668 ;
  assign n29457 = n2573 & ~n4095 ;
  assign n29459 = n29458 ^ n29457 ^ 1'b0 ;
  assign n29460 = n29459 ^ n23571 ^ n9667 ;
  assign n29461 = n26081 ^ n2068 ^ 1'b0 ;
  assign n29462 = n9280 | n29461 ;
  assign n29464 = n4251 | n6375 ;
  assign n29465 = ( ~n8603 & n19230 ) | ( ~n8603 & n29464 ) | ( n19230 & n29464 ) ;
  assign n29463 = n28744 ^ n9606 ^ 1'b0 ;
  assign n29466 = n29465 ^ n29463 ^ n8791 ;
  assign n29467 = ~n22394 & n29466 ;
  assign n29468 = n17980 & n29467 ;
  assign n29469 = n4286 | n4521 ;
  assign n29470 = n431 | n9015 ;
  assign n29471 = n29469 & ~n29470 ;
  assign n29472 = ~n1304 & n29471 ;
  assign n29473 = n19601 & ~n23286 ;
  assign n29474 = n29473 ^ n10617 ^ 1'b0 ;
  assign n29475 = n6884 & n10717 ;
  assign n29476 = ~n1911 & n8997 ;
  assign n29477 = n29476 ^ n4826 ^ 1'b0 ;
  assign n29478 = n29477 ^ n20987 ^ 1'b0 ;
  assign n29480 = n559 ^ n429 ^ 1'b0 ;
  assign n29481 = n5027 | n29480 ;
  assign n29482 = ( n2970 & n6257 ) | ( n2970 & ~n29481 ) | ( n6257 & ~n29481 ) ;
  assign n29483 = ( ~n3517 & n13992 ) | ( ~n3517 & n29482 ) | ( n13992 & n29482 ) ;
  assign n29479 = n1024 & n2486 ;
  assign n29484 = n29483 ^ n29479 ^ 1'b0 ;
  assign n29485 = n14123 & n25384 ;
  assign n29486 = n29485 ^ n1427 ^ 1'b0 ;
  assign n29487 = n29486 ^ n5816 ^ 1'b0 ;
  assign n29488 = n21021 ^ n15988 ^ 1'b0 ;
  assign n29493 = n2144 ^ n2061 ^ 1'b0 ;
  assign n29494 = n29493 ^ n5643 ^ 1'b0 ;
  assign n29495 = n474 & ~n29494 ;
  assign n29491 = ~n9482 & n13309 ;
  assign n29492 = n29491 ^ n7073 ^ 1'b0 ;
  assign n29489 = n12008 ^ n3174 ^ 1'b0 ;
  assign n29490 = n13679 & ~n29489 ;
  assign n29496 = n29495 ^ n29492 ^ n29490 ;
  assign n29498 = n18194 ^ n16761 ^ 1'b0 ;
  assign n29499 = n25358 & n29498 ;
  assign n29497 = ( n2355 & n5949 ) | ( n2355 & ~n14411 ) | ( n5949 & ~n14411 ) ;
  assign n29500 = n29499 ^ n29497 ^ n25539 ;
  assign n29501 = ( n12077 & n17548 ) | ( n12077 & n21702 ) | ( n17548 & n21702 ) ;
  assign n29502 = ( n15812 & n19554 ) | ( n15812 & ~n29501 ) | ( n19554 & ~n29501 ) ;
  assign n29503 = n10092 & n11713 ;
  assign n29504 = n29503 ^ n9339 ^ 1'b0 ;
  assign n29510 = ( n1780 & ~n8044 ) | ( n1780 & n11885 ) | ( ~n8044 & n11885 ) ;
  assign n29505 = n15727 & ~n18306 ;
  assign n29506 = x35 & ~n18030 ;
  assign n29507 = n29505 & n29506 ;
  assign n29508 = ( n14646 & ~n20369 ) | ( n14646 & n29507 ) | ( ~n20369 & n29507 ) ;
  assign n29509 = n26560 | n29508 ;
  assign n29511 = n29510 ^ n29509 ^ 1'b0 ;
  assign n29512 = n15705 | n15909 ;
  assign n29513 = n29512 ^ n2008 ^ 1'b0 ;
  assign n29514 = n8555 & n29513 ;
  assign n29515 = n16332 ^ n15956 ^ 1'b0 ;
  assign n29516 = n2106 & n16485 ;
  assign n29517 = ( n2525 & n29515 ) | ( n2525 & n29516 ) | ( n29515 & n29516 ) ;
  assign n29518 = n7578 & ~n22959 ;
  assign n29519 = n3841 & ~n12867 ;
  assign n29520 = n29519 ^ n3056 ^ 1'b0 ;
  assign n29521 = n13777 & ~n16998 ;
  assign n29522 = n5762 & n29521 ;
  assign n29523 = n19480 & ~n22619 ;
  assign n29524 = n27780 & n29523 ;
  assign n29525 = n26577 ^ n18418 ^ 1'b0 ;
  assign n29526 = ( n13668 & n14042 ) | ( n13668 & ~n29525 ) | ( n14042 & ~n29525 ) ;
  assign n29527 = ( n7431 & n11056 ) | ( n7431 & ~n27536 ) | ( n11056 & ~n27536 ) ;
  assign n29528 = n23865 ^ n7523 ^ 1'b0 ;
  assign n29529 = n2558 | n13920 ;
  assign n29530 = n4727 ^ n3615 ^ 1'b0 ;
  assign n29531 = n18951 & ~n29530 ;
  assign n29532 = n29531 ^ n15676 ^ 1'b0 ;
  assign n29533 = n23814 ^ n3293 ^ 1'b0 ;
  assign n29534 = n14477 & n29533 ;
  assign n29535 = n12106 & n29534 ;
  assign n29536 = n29535 ^ n2855 ^ 1'b0 ;
  assign n29538 = n11397 ^ n308 ^ 1'b0 ;
  assign n29537 = ~n3785 & n4236 ;
  assign n29539 = n29538 ^ n29537 ^ 1'b0 ;
  assign n29540 = n3058 | n13846 ;
  assign n29541 = ~x67 & n29540 ;
  assign n29542 = n29541 ^ n17228 ^ n10310 ;
  assign n29543 = n22446 ^ n8386 ^ 1'b0 ;
  assign n29544 = x55 & n29543 ;
  assign n29545 = ( n574 & ~n29542 ) | ( n574 & n29544 ) | ( ~n29542 & n29544 ) ;
  assign n29546 = n18638 ^ n12494 ^ 1'b0 ;
  assign n29547 = n29546 ^ n25093 ^ n10543 ;
  assign n29548 = n2362 | n26961 ;
  assign n29549 = n29548 ^ n16001 ^ 1'b0 ;
  assign n29550 = n8645 ^ n516 ^ 1'b0 ;
  assign n29553 = n7695 ^ n7617 ^ 1'b0 ;
  assign n29551 = n8630 ^ n1590 ^ 1'b0 ;
  assign n29552 = ( n1362 & n15252 ) | ( n1362 & n29551 ) | ( n15252 & n29551 ) ;
  assign n29554 = n29553 ^ n29552 ^ n8026 ;
  assign n29555 = ~n4594 & n12415 ;
  assign n29556 = n29555 ^ n7369 ^ 1'b0 ;
  assign n29557 = ~n6207 & n29556 ;
  assign n29558 = n1348 & n20695 ;
  assign n29559 = n11810 & n29558 ;
  assign n29560 = ~n29557 & n29559 ;
  assign n29561 = n10103 & n19112 ;
  assign n29562 = n29117 ^ n9455 ^ 1'b0 ;
  assign n29563 = n29561 & ~n29562 ;
  assign n29564 = ( n1151 & ~n2169 ) | ( n1151 & n10014 ) | ( ~n2169 & n10014 ) ;
  assign n29565 = ( ~n6207 & n14498 ) | ( ~n6207 & n29564 ) | ( n14498 & n29564 ) ;
  assign n29566 = n3043 & n6372 ;
  assign n29567 = n661 | n10097 ;
  assign n29568 = ( n18457 & n29566 ) | ( n18457 & n29567 ) | ( n29566 & n29567 ) ;
  assign n29569 = ~n5598 & n9226 ;
  assign n29570 = ~n18975 & n29569 ;
  assign n29571 = ~n21079 & n29570 ;
  assign n29575 = n14728 ^ n9956 ^ 1'b0 ;
  assign n29576 = n29575 ^ n15140 ^ 1'b0 ;
  assign n29577 = n2054 & ~n29576 ;
  assign n29573 = ~n2257 & n6082 ;
  assign n29572 = n7353 | n12568 ;
  assign n29574 = n29573 ^ n29572 ^ 1'b0 ;
  assign n29578 = n29577 ^ n29574 ^ 1'b0 ;
  assign n29579 = n19200 ^ n9222 ^ 1'b0 ;
  assign n29580 = ( x184 & ~n9302 ) | ( x184 & n29579 ) | ( ~n9302 & n29579 ) ;
  assign n29581 = n7946 & ~n11746 ;
  assign n29582 = ( n453 & n7145 ) | ( n453 & ~n8564 ) | ( n7145 & ~n8564 ) ;
  assign n29583 = n15998 & ~n29582 ;
  assign n29584 = n29583 ^ n9307 ^ 1'b0 ;
  assign n29585 = n3508 & n9743 ;
  assign n29586 = n5037 ^ n4331 ^ n745 ;
  assign n29587 = n24450 ^ n1992 ^ 1'b0 ;
  assign n29588 = n29587 ^ n4001 ^ 1'b0 ;
  assign n29589 = n29586 & n29588 ;
  assign n29590 = ~n9939 & n19232 ;
  assign n29591 = n29590 ^ n5927 ^ 1'b0 ;
  assign n29592 = n29591 ^ n15520 ^ 1'b0 ;
  assign n29593 = ~n2292 & n29592 ;
  assign n29594 = n29593 ^ n7055 ^ 1'b0 ;
  assign n29595 = ~n22040 & n29594 ;
  assign n29596 = n8651 ^ n7484 ^ 1'b0 ;
  assign n29597 = ~n9102 & n29596 ;
  assign n29598 = n4198 & ~n29597 ;
  assign n29599 = n17216 ^ n8025 ^ 1'b0 ;
  assign n29600 = n29598 | n29599 ;
  assign n29601 = n8161 ^ n6616 ^ 1'b0 ;
  assign n29602 = n13161 & ~n17733 ;
  assign n29603 = ~n29601 & n29602 ;
  assign n29604 = n17028 & n17240 ;
  assign n29605 = n29604 ^ n8720 ^ n8345 ;
  assign n29608 = n24882 ^ n12538 ^ 1'b0 ;
  assign n29606 = n2850 & ~n20692 ;
  assign n29607 = n29606 ^ n16483 ^ 1'b0 ;
  assign n29609 = n29608 ^ n29607 ^ n15618 ;
  assign n29610 = n2353 | n9435 ;
  assign n29611 = n14604 & n29610 ;
  assign n29612 = ~n21411 & n29611 ;
  assign n29613 = n29612 ^ n9545 ^ 1'b0 ;
  assign n29614 = n15520 | n29613 ;
  assign n29615 = n6618 & n16077 ;
  assign n29616 = n29615 ^ n8722 ^ 1'b0 ;
  assign n29617 = n29616 ^ n11524 ^ 1'b0 ;
  assign n29618 = n9938 | n29617 ;
  assign n29619 = n29618 ^ n4207 ^ 1'b0 ;
  assign n29620 = ~n18616 & n27629 ;
  assign n29621 = ~n28861 & n29620 ;
  assign n29622 = n11328 & n15803 ;
  assign n29623 = n7571 & n29622 ;
  assign n29624 = n17339 ^ n10126 ^ n2581 ;
  assign n29625 = n26378 ^ n21953 ^ n5091 ;
  assign n29626 = n4693 & n13637 ;
  assign n29627 = n16662 & n29626 ;
  assign n29628 = ~n1935 & n29124 ;
  assign n29629 = n29627 & n29628 ;
  assign n29631 = n14873 ^ n13603 ^ 1'b0 ;
  assign n29630 = n5740 & n10421 ;
  assign n29632 = n29631 ^ n29630 ^ 1'b0 ;
  assign n29633 = n14976 ^ n6683 ^ n2688 ;
  assign n29634 = n12155 | n29633 ;
  assign n29635 = n1802 | n29634 ;
  assign n29636 = ~n2518 & n21658 ;
  assign n29640 = n5541 | n7064 ;
  assign n29641 = n29640 ^ n8659 ^ 1'b0 ;
  assign n29639 = ~x66 & n2981 ;
  assign n29642 = n29641 ^ n29639 ^ n939 ;
  assign n29637 = ~n23297 & n24874 ;
  assign n29638 = ~n5210 & n29637 ;
  assign n29643 = n29642 ^ n29638 ^ n25698 ;
  assign n29644 = ~n10962 & n16512 ;
  assign n29645 = n29644 ^ n7781 ^ 1'b0 ;
  assign n29646 = n29645 ^ n7348 ^ 1'b0 ;
  assign n29647 = ( n3998 & ~n20935 ) | ( n3998 & n29646 ) | ( ~n20935 & n29646 ) ;
  assign n29648 = n20899 | n22741 ;
  assign n29649 = n29648 ^ n13799 ^ 1'b0 ;
  assign n29650 = n4840 & ~n29385 ;
  assign n29651 = n16812 & n23912 ;
  assign n29652 = n17802 & ~n29651 ;
  assign n29653 = n29652 ^ n1865 ^ 1'b0 ;
  assign n29655 = ~n6901 & n17666 ;
  assign n29656 = n29655 ^ n10227 ^ 1'b0 ;
  assign n29654 = n1475 | n3761 ;
  assign n29657 = n29656 ^ n29654 ^ 1'b0 ;
  assign n29658 = n9692 & n12717 ;
  assign n29659 = n29658 ^ n10093 ^ 1'b0 ;
  assign n29660 = n28550 ^ n315 ^ 1'b0 ;
  assign n29661 = n5719 & ~n29660 ;
  assign n29662 = n1665 | n24882 ;
  assign n29663 = n24046 ^ n8165 ^ n4388 ;
  assign n29664 = n11357 ^ n11147 ^ 1'b0 ;
  assign n29665 = ~n23477 & n29664 ;
  assign n29666 = n29665 ^ n28972 ^ 1'b0 ;
  assign n29667 = n26744 ^ n20590 ^ 1'b0 ;
  assign n29668 = n20941 | n29667 ;
  assign n29669 = n21695 ^ n3134 ^ 1'b0 ;
  assign n29670 = ~n29668 & n29669 ;
  assign n29671 = n13793 ^ n7106 ^ 1'b0 ;
  assign n29672 = n19946 | n29671 ;
  assign n29673 = n29672 ^ n10637 ^ 1'b0 ;
  assign n29674 = n14905 ^ n7734 ^ 1'b0 ;
  assign n29675 = x1 & ~n29674 ;
  assign n29676 = ( n1097 & n8366 ) | ( n1097 & n27749 ) | ( n8366 & n27749 ) ;
  assign n29677 = n26469 ^ n25473 ^ 1'b0 ;
  assign n29678 = n2765 | n29677 ;
  assign n29679 = n26461 & ~n29678 ;
  assign n29680 = n29679 ^ n21121 ^ 1'b0 ;
  assign n29681 = n6401 ^ n4907 ^ 1'b0 ;
  assign n29682 = n4480 | n29681 ;
  assign n29683 = n17450 & n26095 ;
  assign n29684 = n15812 & n29683 ;
  assign n29685 = n29684 ^ n6290 ^ 1'b0 ;
  assign n29687 = ~n3449 & n4913 ;
  assign n29688 = ~n2907 & n12213 ;
  assign n29689 = ~n29687 & n29688 ;
  assign n29686 = n22367 ^ n10563 ^ n4047 ;
  assign n29690 = n29689 ^ n29686 ^ n14687 ;
  assign n29691 = n8152 & ~n27877 ;
  assign n29692 = n15198 & n29691 ;
  assign n29693 = ~n10517 & n29692 ;
  assign n29694 = n13217 & ~n19741 ;
  assign n29695 = n29693 & n29694 ;
  assign n29696 = ~n526 & n7359 ;
  assign n29697 = ~n3808 & n29651 ;
  assign n29698 = n11571 ^ n11391 ^ 1'b0 ;
  assign n29699 = n29698 ^ n9163 ^ 1'b0 ;
  assign n29701 = n3641 & n14187 ;
  assign n29700 = n1029 & ~n5310 ;
  assign n29702 = n29701 ^ n29700 ^ 1'b0 ;
  assign n29703 = ~n14756 & n17847 ;
  assign n29704 = n3888 & n29703 ;
  assign n29705 = n15504 ^ n14405 ^ n3147 ;
  assign n29706 = n4701 | n29705 ;
  assign n29707 = ~n7718 & n23024 ;
  assign n29708 = n29707 ^ n23688 ^ 1'b0 ;
  assign n29709 = n5927 | n13235 ;
  assign n29710 = n29709 ^ n19992 ^ 1'b0 ;
  assign n29711 = n27732 ^ n26326 ^ 1'b0 ;
  assign n29712 = n22307 & ~n29711 ;
  assign n29713 = ~n7170 & n29712 ;
  assign n29714 = x129 | n24343 ;
  assign n29715 = n14981 & ~n29714 ;
  assign n29716 = n19906 ^ n16654 ^ 1'b0 ;
  assign n29717 = n11713 & n21374 ;
  assign n29718 = n29717 ^ n6867 ^ 1'b0 ;
  assign n29719 = ( n17333 & n25203 ) | ( n17333 & n26186 ) | ( n25203 & n26186 ) ;
  assign n29720 = ( n704 & ~n5184 ) | ( n704 & n10576 ) | ( ~n5184 & n10576 ) ;
  assign n29721 = n7937 | n18480 ;
  assign n29722 = ( n6352 & n29720 ) | ( n6352 & ~n29721 ) | ( n29720 & ~n29721 ) ;
  assign n29723 = n8053 | n16440 ;
  assign n29724 = n29723 ^ n6500 ^ 1'b0 ;
  assign n29725 = ~n3944 & n8800 ;
  assign n29726 = ~n26578 & n29725 ;
  assign n29727 = ( n3832 & n21085 ) | ( n3832 & ~n29726 ) | ( n21085 & ~n29726 ) ;
  assign n29728 = n29724 | n29727 ;
  assign n29729 = n20658 & ~n29728 ;
  assign n29730 = n27946 ^ n4382 ^ 1'b0 ;
  assign n29731 = n5292 | n29730 ;
  assign n29732 = n4549 & ~n29731 ;
  assign n29733 = n14481 ^ n1166 ^ n500 ;
  assign n29734 = n24825 & n29733 ;
  assign n29735 = n11396 ^ n926 ^ 1'b0 ;
  assign n29736 = n3704 & ~n29735 ;
  assign n29737 = n1671 & ~n12663 ;
  assign n29738 = ~n11222 & n29737 ;
  assign n29739 = n29510 ^ n18752 ^ 1'b0 ;
  assign n29740 = n3903 ^ n3662 ^ 1'b0 ;
  assign n29741 = ( ~n18786 & n22564 ) | ( ~n18786 & n29740 ) | ( n22564 & n29740 ) ;
  assign n29742 = n23147 & ~n29741 ;
  assign n29743 = n29742 ^ n26244 ^ 1'b0 ;
  assign n29744 = n10023 | n25391 ;
  assign n29745 = n29744 ^ n14449 ^ 1'b0 ;
  assign n29746 = n24268 ^ n20705 ^ 1'b0 ;
  assign n29747 = n13035 ^ n7732 ^ 1'b0 ;
  assign n29748 = n29747 ^ n12739 ^ n6322 ;
  assign n29749 = n3273 ^ n2781 ^ 1'b0 ;
  assign n29750 = n12277 | n29749 ;
  assign n29751 = n4917 ^ n1932 ^ 1'b0 ;
  assign n29752 = n19622 & ~n29751 ;
  assign n29753 = ~n15749 & n29752 ;
  assign n29754 = ~n23704 & n26815 ;
  assign n29755 = n4759 | n29754 ;
  assign n29756 = n29755 ^ n405 ^ 1'b0 ;
  assign n29757 = n20987 ^ n9104 ^ 1'b0 ;
  assign n29758 = n29601 & ~n29757 ;
  assign n29759 = n18156 ^ n2008 ^ 1'b0 ;
  assign n29760 = n2098 | n28942 ;
  assign n29761 = n17136 | n26968 ;
  assign n29762 = n26127 ^ n14247 ^ 1'b0 ;
  assign n29763 = ~n4179 & n29762 ;
  assign n29764 = n790 & ~n5523 ;
  assign n29765 = ~n24084 & n29764 ;
  assign n29766 = n29188 ^ n4800 ^ 1'b0 ;
  assign n29767 = n11719 | n29766 ;
  assign n29768 = x162 & n4950 ;
  assign n29769 = n29768 ^ n8055 ^ 1'b0 ;
  assign n29770 = ~n13008 & n27111 ;
  assign n29771 = n8825 | n22759 ;
  assign n29772 = n19409 | n29771 ;
  assign n29773 = n2431 | n29580 ;
  assign n29774 = n24546 ^ n4918 ^ 1'b0 ;
  assign n29775 = n2829 & ~n29774 ;
  assign n29776 = n16269 ^ n5421 ^ 1'b0 ;
  assign n29777 = n4971 | n29776 ;
  assign n29778 = n12355 & n29777 ;
  assign n29779 = n19798 ^ n6066 ^ 1'b0 ;
  assign n29780 = ~n5469 & n29779 ;
  assign n29781 = n8165 & ~n19142 ;
  assign n29782 = n29781 ^ n7433 ^ 1'b0 ;
  assign n29783 = ( n29778 & n29780 ) | ( n29778 & n29782 ) | ( n29780 & n29782 ) ;
  assign n29784 = ~n6122 & n16252 ;
  assign n29785 = n28475 ^ n21750 ^ 1'b0 ;
  assign n29786 = n18963 | n29785 ;
  assign n29787 = n9960 | n15795 ;
  assign n29789 = n22374 ^ n12376 ^ n10331 ;
  assign n29788 = n3104 | n21770 ;
  assign n29790 = n29789 ^ n29788 ^ 1'b0 ;
  assign n29791 = n8808 ^ n6371 ^ 1'b0 ;
  assign n29792 = n10368 & ~n29791 ;
  assign n29794 = n733 | n785 ;
  assign n29795 = n29794 ^ x123 ^ 1'b0 ;
  assign n29796 = n29795 ^ n19310 ^ 1'b0 ;
  assign n29793 = n9517 & n10671 ;
  assign n29797 = n29796 ^ n29793 ^ 1'b0 ;
  assign n29798 = n29797 ^ n15726 ^ 1'b0 ;
  assign n29799 = n29792 & n29798 ;
  assign n29800 = n3295 & ~n25277 ;
  assign n29801 = n8726 ^ n5896 ^ 1'b0 ;
  assign n29802 = ~n15618 & n29801 ;
  assign n29804 = ~n6314 & n24134 ;
  assign n29803 = ( n4200 & n16667 ) | ( n4200 & n27384 ) | ( n16667 & n27384 ) ;
  assign n29805 = n29804 ^ n29803 ^ n13692 ;
  assign n29806 = n3831 & ~n22092 ;
  assign n29807 = n19861 & n29806 ;
  assign n29808 = n5502 ^ n607 ^ 1'b0 ;
  assign n29809 = n2765 & ~n29808 ;
  assign n29810 = n29809 ^ n7402 ^ 1'b0 ;
  assign n29811 = n13982 ^ n7658 ^ 1'b0 ;
  assign n29812 = ~n918 & n2241 ;
  assign n29813 = n29812 ^ n5011 ^ 1'b0 ;
  assign n29814 = n29811 & ~n29813 ;
  assign n29815 = n10592 & n14625 ;
  assign n29816 = n29815 ^ n5205 ^ 1'b0 ;
  assign n29817 = n17887 ^ n10313 ^ 1'b0 ;
  assign n29819 = ( n2176 & ~n3798 ) | ( n2176 & n5443 ) | ( ~n3798 & n5443 ) ;
  assign n29818 = x146 & ~n15455 ;
  assign n29820 = n29819 ^ n29818 ^ 1'b0 ;
  assign n29821 = n8512 ^ n4876 ^ 1'b0 ;
  assign n29822 = n23696 & n29821 ;
  assign n29823 = ~n2380 & n8966 ;
  assign n29824 = n29823 ^ n26067 ^ 1'b0 ;
  assign n29825 = n2252 & n26204 ;
  assign n29826 = n18536 & n29414 ;
  assign n29827 = n1902 | n8312 ;
  assign n29828 = n3786 | n8457 ;
  assign n29829 = n3501 | n29828 ;
  assign n29830 = n29829 ^ x179 ^ 1'b0 ;
  assign n29831 = n3128 & n29830 ;
  assign n29832 = n29831 ^ n4168 ^ 1'b0 ;
  assign n29834 = n18935 ^ n5920 ^ 1'b0 ;
  assign n29833 = n12697 ^ n4768 ^ 1'b0 ;
  assign n29835 = n29834 ^ n29833 ^ n18604 ;
  assign n29836 = n3464 & n3817 ;
  assign n29841 = n10699 | n25890 ;
  assign n29842 = n24272 & ~n29841 ;
  assign n29837 = ~n18935 & n23081 ;
  assign n29838 = n7645 ^ n2575 ^ 1'b0 ;
  assign n29839 = n29838 ^ n14518 ^ n274 ;
  assign n29840 = n29837 & n29839 ;
  assign n29843 = n29842 ^ n29840 ^ 1'b0 ;
  assign n29844 = n13860 ^ n4264 ^ 1'b0 ;
  assign n29845 = n21675 & n29844 ;
  assign n29846 = n12363 & n27910 ;
  assign n29847 = n2956 & ~n4800 ;
  assign n29848 = n29847 ^ x168 ^ 1'b0 ;
  assign n29849 = ~n18079 & n29848 ;
  assign n29850 = n5962 | n20325 ;
  assign n29851 = n4328 | n29850 ;
  assign n29852 = ~n2733 & n15047 ;
  assign n29853 = n29852 ^ n6611 ^ 1'b0 ;
  assign n29854 = ( n22018 & n29851 ) | ( n22018 & n29853 ) | ( n29851 & n29853 ) ;
  assign n29855 = n7310 | n29854 ;
  assign n29856 = n29849 | n29855 ;
  assign n29857 = ~n5577 & n7128 ;
  assign n29858 = n29857 ^ n4165 ^ 1'b0 ;
  assign n29859 = n9661 & ~n29858 ;
  assign n29860 = n997 | n23292 ;
  assign n29861 = n4557 & ~n5094 ;
  assign n29862 = n29861 ^ n3743 ^ 1'b0 ;
  assign n29863 = n29862 ^ n23459 ^ 1'b0 ;
  assign n29864 = n13134 | n29863 ;
  assign n29865 = n4194 & ~n8519 ;
  assign n29866 = n7172 ^ n3743 ^ 1'b0 ;
  assign n29867 = ~n904 & n29866 ;
  assign n29868 = n3954 & n29867 ;
  assign n29869 = n7782 | n12679 ;
  assign n29870 = n12948 & ~n29869 ;
  assign n29871 = n6205 ^ n6176 ^ 1'b0 ;
  assign n29872 = ( n6760 & n25964 ) | ( n6760 & ~n29871 ) | ( n25964 & ~n29871 ) ;
  assign n29873 = n29872 ^ n6555 ^ 1'b0 ;
  assign n29874 = ~n3342 & n29873 ;
  assign n29875 = n1182 & n20563 ;
  assign n29876 = n20945 & n29875 ;
  assign n29877 = n11053 ^ n473 ^ 1'b0 ;
  assign n29878 = ~n29876 & n29877 ;
  assign n29879 = ~n3470 & n9224 ;
  assign n29880 = n29879 ^ n17426 ^ 1'b0 ;
  assign n29881 = n16521 & ~n18338 ;
  assign n29882 = n29881 ^ n8830 ^ 1'b0 ;
  assign n29883 = ~n4498 & n28280 ;
  assign n29884 = n29883 ^ n12929 ^ 1'b0 ;
  assign n29888 = n7088 ^ n1113 ^ 1'b0 ;
  assign n29885 = n4456 ^ n3794 ^ 1'b0 ;
  assign n29886 = n3520 & n29885 ;
  assign n29887 = ~n11176 & n29886 ;
  assign n29889 = n29888 ^ n29887 ^ 1'b0 ;
  assign n29890 = n2829 | n21409 ;
  assign n29891 = ~n10621 & n23330 ;
  assign n29892 = n1692 & ~n6870 ;
  assign n29893 = n6981 & n29892 ;
  assign n29894 = n1909 | n9583 ;
  assign n29895 = n27642 ^ n9984 ^ n3551 ;
  assign n29896 = n14350 & n29895 ;
  assign n29897 = n29896 ^ n11593 ^ 1'b0 ;
  assign n29898 = ( ~n2465 & n8594 ) | ( ~n2465 & n24148 ) | ( n8594 & n24148 ) ;
  assign n29904 = n17032 ^ n5896 ^ 1'b0 ;
  assign n29900 = n15649 ^ n8337 ^ 1'b0 ;
  assign n29901 = ~n8363 & n29900 ;
  assign n29902 = n4622 | n29901 ;
  assign n29903 = n29902 ^ n6034 ^ 1'b0 ;
  assign n29899 = n26043 ^ n14814 ^ 1'b0 ;
  assign n29905 = n29904 ^ n29903 ^ n29899 ;
  assign n29906 = n16083 & n28757 ;
  assign n29907 = ( n978 & ~n4650 ) | ( n978 & n7429 ) | ( ~n4650 & n7429 ) ;
  assign n29908 = ( ~n3685 & n9948 ) | ( ~n3685 & n29907 ) | ( n9948 & n29907 ) ;
  assign n29909 = n29908 ^ n8567 ^ 1'b0 ;
  assign n29910 = n21286 & ~n29909 ;
  assign n29911 = n29910 ^ n22015 ^ 1'b0 ;
  assign n29912 = n1136 | n29911 ;
  assign n29913 = n16908 ^ n3389 ^ 1'b0 ;
  assign n29915 = n3691 & n20595 ;
  assign n29914 = n1130 & n10766 ;
  assign n29916 = n29915 ^ n29914 ^ n2749 ;
  assign n29919 = n6170 | n16923 ;
  assign n29917 = n1882 | n5884 ;
  assign n29918 = n24669 | n29917 ;
  assign n29920 = n29919 ^ n29918 ^ 1'b0 ;
  assign n29921 = ( ~n7027 & n15690 ) | ( ~n7027 & n16205 ) | ( n15690 & n16205 ) ;
  assign n29922 = n980 ^ n428 ^ 1'b0 ;
  assign n29923 = n14304 | n29922 ;
  assign n29924 = n16093 | n16105 ;
  assign n29925 = n7320 ^ n980 ^ 1'b0 ;
  assign n29926 = n451 & ~n29925 ;
  assign n29927 = n11641 ^ n8601 ^ 1'b0 ;
  assign n29928 = n29926 & ~n29927 ;
  assign n29929 = n1553 & n29928 ;
  assign n29930 = n29929 ^ n8585 ^ 1'b0 ;
  assign n29932 = n2956 ^ x22 ^ 1'b0 ;
  assign n29931 = n24017 & ~n24258 ;
  assign n29933 = n29932 ^ n29931 ^ n24006 ;
  assign n29934 = n23332 ^ n1325 ^ 1'b0 ;
  assign n29937 = n9636 ^ n5538 ^ n376 ;
  assign n29938 = ~n4150 & n29937 ;
  assign n29935 = n26976 ^ n10128 ^ 1'b0 ;
  assign n29936 = ~n10019 & n29935 ;
  assign n29939 = n29938 ^ n29936 ^ 1'b0 ;
  assign n29940 = n22070 ^ n7756 ^ 1'b0 ;
  assign n29941 = n7492 ^ n1150 ^ 1'b0 ;
  assign n29942 = n25540 ^ n3760 ^ 1'b0 ;
  assign n29943 = n672 & n12572 ;
  assign n29944 = n14555 ^ n3237 ^ 1'b0 ;
  assign n29945 = n983 | n2547 ;
  assign n29946 = n29945 ^ n2959 ^ 1'b0 ;
  assign n29947 = ~n11772 & n29946 ;
  assign n29948 = n14780 ^ n706 ^ 1'b0 ;
  assign n29949 = n29947 | n29948 ;
  assign n29950 = n3413 & ~n20130 ;
  assign n29951 = n15577 ^ n7974 ^ 1'b0 ;
  assign n29952 = ~n2422 & n29951 ;
  assign n29953 = n6445 ^ n610 ^ 1'b0 ;
  assign n29954 = n27478 ^ n24208 ^ 1'b0 ;
  assign n29955 = n6279 | n29954 ;
  assign n29956 = n29955 ^ n20407 ^ n9542 ;
  assign n29957 = ( n2213 & n9744 ) | ( n2213 & ~n23430 ) | ( n9744 & ~n23430 ) ;
  assign n29958 = ~n6494 & n12815 ;
  assign n29959 = n9804 & ~n29958 ;
  assign n29960 = n19512 ^ n17626 ^ 1'b0 ;
  assign n29961 = ( n4313 & n29959 ) | ( n4313 & n29960 ) | ( n29959 & n29960 ) ;
  assign n29962 = n26293 & ~n29032 ;
  assign n29963 = n4243 & n29962 ;
  assign n29964 = n15020 & n16415 ;
  assign n29965 = ~n22659 & n29964 ;
  assign n29966 = n29965 ^ n21877 ^ 1'b0 ;
  assign n29967 = ~n3551 & n14224 ;
  assign n29971 = n668 & ~n25849 ;
  assign n29968 = ~n5432 & n18158 ;
  assign n29969 = n29968 ^ n15747 ^ 1'b0 ;
  assign n29970 = n29969 ^ n6842 ^ n2578 ;
  assign n29972 = n29971 ^ n29970 ^ 1'b0 ;
  assign n29973 = ~n9099 & n29972 ;
  assign n29974 = ~n2910 & n3764 ;
  assign n29975 = ~n8813 & n29188 ;
  assign n29976 = n16106 ^ n3973 ^ 1'b0 ;
  assign n29977 = n7007 & ~n29976 ;
  assign n29978 = ~n10055 & n21374 ;
  assign n29979 = n29978 ^ n21515 ^ 1'b0 ;
  assign n29980 = ( n20570 & ~n29126 ) | ( n20570 & n29979 ) | ( ~n29126 & n29979 ) ;
  assign n29981 = n2885 & ~n15893 ;
  assign n29982 = n29981 ^ n6382 ^ 1'b0 ;
  assign n29983 = n14175 & ~n29982 ;
  assign n29984 = n29983 ^ n8035 ^ n2796 ;
  assign n29985 = ~n7254 & n10973 ;
  assign n29986 = n5253 | n22735 ;
  assign n29987 = n29986 ^ n10348 ^ 1'b0 ;
  assign n29988 = ~n1515 & n14330 ;
  assign n29989 = ~n19668 & n29988 ;
  assign n29990 = n5984 & n29989 ;
  assign n29991 = ~n14746 & n17598 ;
  assign n29992 = n29991 ^ n26624 ^ 1'b0 ;
  assign n29993 = n13007 & ~n24618 ;
  assign n29994 = ~n28535 & n29993 ;
  assign n29995 = n26656 ^ n14486 ^ 1'b0 ;
  assign n29996 = ( n4705 & n27694 ) | ( n4705 & ~n29995 ) | ( n27694 & ~n29995 ) ;
  assign n29997 = n9883 ^ n4108 ^ 1'b0 ;
  assign n29998 = n5221 & ~n29997 ;
  assign n30000 = ~n7569 & n12373 ;
  assign n30001 = n30000 ^ n7253 ^ n1377 ;
  assign n30002 = n30001 ^ n8848 ^ 1'b0 ;
  assign n29999 = ~n14620 & n23212 ;
  assign n30003 = n30002 ^ n29999 ^ 1'b0 ;
  assign n30004 = n5522 & n8468 ;
  assign n30005 = n26353 ^ n19696 ^ 1'b0 ;
  assign n30006 = n10378 | n12881 ;
  assign n30007 = ~n9504 & n30006 ;
  assign n30008 = n13543 & n30007 ;
  assign n30009 = x21 & ~n15053 ;
  assign n30010 = ~x21 & n30009 ;
  assign n30011 = n10078 & n30010 ;
  assign n30012 = n3567 | n15316 ;
  assign n30013 = n30012 ^ n5637 ^ 1'b0 ;
  assign n30014 = n16331 & n26515 ;
  assign n30015 = n24056 ^ n16343 ^ 1'b0 ;
  assign n30016 = n30015 ^ n27916 ^ 1'b0 ;
  assign n30017 = n3905 | n30016 ;
  assign n30018 = n13948 & n21965 ;
  assign n30019 = n30018 ^ n2357 ^ 1'b0 ;
  assign n30020 = ~n2318 & n17055 ;
  assign n30021 = n30019 & ~n30020 ;
  assign n30022 = ~n16276 & n23869 ;
  assign n30023 = n4279 & ~n24046 ;
  assign n30024 = n13752 & n22526 ;
  assign n30025 = ~n17932 & n30024 ;
  assign n30026 = n18058 | n19836 ;
  assign n30027 = n30025 & n30026 ;
  assign n30028 = n30027 ^ n4364 ^ 1'b0 ;
  assign n30029 = n23879 & ~n30028 ;
  assign n30030 = n28652 ^ n2791 ^ 1'b0 ;
  assign n30031 = n3302 & ~n19810 ;
  assign n30032 = n15833 & n30031 ;
  assign n30033 = n30032 ^ n19287 ^ 1'b0 ;
  assign n30038 = ( n1514 & n7811 ) | ( n1514 & n9960 ) | ( n7811 & n9960 ) ;
  assign n30036 = ~n12790 & n15159 ;
  assign n30037 = n11569 & n30036 ;
  assign n30039 = n30038 ^ n30037 ^ 1'b0 ;
  assign n30034 = n5117 & ~n14231 ;
  assign n30035 = ~n27480 & n30034 ;
  assign n30040 = n30039 ^ n30035 ^ 1'b0 ;
  assign n30041 = n15341 & n21003 ;
  assign n30042 = n9028 & n30041 ;
  assign n30043 = n29466 ^ n8438 ^ 1'b0 ;
  assign n30044 = n30043 ^ n5724 ^ 1'b0 ;
  assign n30045 = n4284 & ~n30044 ;
  assign n30049 = ~n10265 & n14884 ;
  assign n30046 = n1124 | n18274 ;
  assign n30047 = n4802 & ~n30046 ;
  assign n30048 = n9822 & ~n30047 ;
  assign n30050 = n30049 ^ n30048 ^ 1'b0 ;
  assign n30051 = n19901 & n24327 ;
  assign n30052 = n30051 ^ n9579 ^ 1'b0 ;
  assign n30059 = n23432 ^ n15190 ^ 1'b0 ;
  assign n30060 = ~n14441 & n30059 ;
  assign n30061 = n30060 ^ n8791 ^ 1'b0 ;
  assign n30054 = n8966 ^ n4789 ^ 1'b0 ;
  assign n30055 = n3526 & ~n30054 ;
  assign n30053 = n3642 | n18667 ;
  assign n30056 = n30055 ^ n30053 ^ 1'b0 ;
  assign n30057 = n7630 & n30056 ;
  assign n30058 = n4425 & n30057 ;
  assign n30062 = n30061 ^ n30058 ^ n1830 ;
  assign n30063 = n4398 | n17485 ;
  assign n30064 = ~n14346 & n30063 ;
  assign n30065 = n26642 & n30064 ;
  assign n30066 = n8305 | n15516 ;
  assign n30067 = n30066 ^ n9513 ^ 1'b0 ;
  assign n30068 = n30067 ^ n11066 ^ 1'b0 ;
  assign n30069 = n5487 & n19668 ;
  assign n30070 = n21223 ^ n12193 ^ 1'b0 ;
  assign n30071 = n20119 ^ n4699 ^ 1'b0 ;
  assign n30075 = n3263 ^ n758 ^ 1'b0 ;
  assign n30072 = n319 & ~n10968 ;
  assign n30073 = n3178 & n28677 ;
  assign n30074 = n30072 & n30073 ;
  assign n30076 = n30075 ^ n30074 ^ 1'b0 ;
  assign n30077 = n4058 & n12472 ;
  assign n30078 = x26 & ~n1788 ;
  assign n30079 = ~n28272 & n30078 ;
  assign n30080 = n770 & ~n30079 ;
  assign n30081 = n28280 ^ n9500 ^ n1228 ;
  assign n30082 = n28069 & ~n30081 ;
  assign n30083 = n1168 & ~n8430 ;
  assign n30084 = n30083 ^ n16612 ^ n6233 ;
  assign n30085 = n4072 | n12601 ;
  assign n30086 = n16186 | n30085 ;
  assign n30087 = n808 & ~n3051 ;
  assign n30088 = ~n18158 & n30087 ;
  assign n30089 = n30088 ^ n1572 ^ 1'b0 ;
  assign n30090 = n30089 ^ n14677 ^ n12004 ;
  assign n30091 = n28468 ^ n17808 ^ 1'b0 ;
  assign n30092 = n13989 ^ n4945 ^ 1'b0 ;
  assign n30094 = n4466 | n12718 ;
  assign n30095 = n30094 ^ n8608 ^ 1'b0 ;
  assign n30093 = n18853 | n29145 ;
  assign n30096 = n30095 ^ n30093 ^ 1'b0 ;
  assign n30097 = n22096 ^ n2384 ^ 1'b0 ;
  assign n30098 = ~n6868 & n30097 ;
  assign n30101 = n6729 & ~n13641 ;
  assign n30099 = n2012 & ~n5029 ;
  assign n30100 = n30099 ^ n25673 ^ n23311 ;
  assign n30102 = n30101 ^ n30100 ^ n8667 ;
  assign n30103 = n7146 ^ n5857 ^ n2652 ;
  assign n30104 = n30103 ^ n16536 ^ 1'b0 ;
  assign n30105 = ~n5027 & n16060 ;
  assign n30106 = n5693 & n30105 ;
  assign n30107 = n17744 | n24413 ;
  assign n30108 = n30107 ^ n13590 ^ 1'b0 ;
  assign n30109 = n6813 | n14895 ;
  assign n30110 = n30109 ^ n9540 ^ 1'b0 ;
  assign n30111 = n30110 ^ n24461 ^ 1'b0 ;
  assign n30112 = x65 & n3166 ;
  assign n30113 = ~n2962 & n30112 ;
  assign n30114 = ( n16324 & ~n18559 ) | ( n16324 & n30113 ) | ( ~n18559 & n30113 ) ;
  assign n30115 = n11529 ^ n1596 ^ 1'b0 ;
  assign n30116 = n4194 & ~n5463 ;
  assign n30117 = n30116 ^ n24030 ^ 1'b0 ;
  assign n30118 = n13243 ^ n4213 ^ 1'b0 ;
  assign n30119 = ( n10753 & n10888 ) | ( n10753 & ~n20922 ) | ( n10888 & ~n20922 ) ;
  assign n30120 = n11503 & n30119 ;
  assign n30121 = n2151 & n26519 ;
  assign n30122 = n9701 & ~n12419 ;
  assign n30123 = n30122 ^ n28067 ^ n14891 ;
  assign n30124 = x220 | n1880 ;
  assign n30125 = n30124 ^ n4931 ^ 1'b0 ;
  assign n30126 = ~n2614 & n14424 ;
  assign n30127 = ~n17233 & n30126 ;
  assign n30128 = n15808 | n30127 ;
  assign n30129 = n2226 & ~n30128 ;
  assign n30130 = n17030 ^ n9334 ^ 1'b0 ;
  assign n30131 = n27426 & ~n30130 ;
  assign n30132 = n30131 ^ n5800 ^ 1'b0 ;
  assign n30133 = n26491 ^ n20977 ^ 1'b0 ;
  assign n30134 = n22035 | n30133 ;
  assign n30135 = n2305 & ~n11872 ;
  assign n30136 = n30135 ^ n28257 ^ n18280 ;
  assign n30137 = n14967 ^ n5242 ^ 1'b0 ;
  assign n30138 = n1122 & ~n30137 ;
  assign n30139 = n21217 | n24568 ;
  assign n30140 = ~n15695 & n23659 ;
  assign n30141 = n1515 | n4029 ;
  assign n30142 = n30141 ^ n25048 ^ 1'b0 ;
  assign n30143 = n9201 ^ n2483 ^ 1'b0 ;
  assign n30144 = n2235 & n6594 ;
  assign n30145 = n30144 ^ n10530 ^ 1'b0 ;
  assign n30146 = n9338 ^ n7685 ^ 1'b0 ;
  assign n30147 = n30146 ^ n20314 ^ n9217 ;
  assign n30148 = n9480 & ~n30147 ;
  assign n30149 = n30148 ^ n14254 ^ 1'b0 ;
  assign n30150 = ~n4378 & n17645 ;
  assign n30151 = n6265 & n30150 ;
  assign n30152 = n9591 ^ n1902 ^ 1'b0 ;
  assign n30153 = ~n9247 & n30152 ;
  assign n30154 = n10665 ^ n1869 ^ 1'b0 ;
  assign n30155 = ~n15610 & n30154 ;
  assign n30156 = n28614 ^ n17230 ^ 1'b0 ;
  assign n30157 = ( n2582 & n15846 ) | ( n2582 & n22127 ) | ( n15846 & n22127 ) ;
  assign n30161 = n10383 | n26031 ;
  assign n30158 = n3702 & n4004 ;
  assign n30159 = n30158 ^ n527 ^ 1'b0 ;
  assign n30160 = n11836 & ~n30159 ;
  assign n30162 = n30161 ^ n30160 ^ n23151 ;
  assign n30163 = n14224 & n29721 ;
  assign n30164 = n30163 ^ n8114 ^ 1'b0 ;
  assign n30165 = n9708 & ~n30164 ;
  assign n30166 = n451 & ~n1941 ;
  assign n30167 = ~n20763 & n30166 ;
  assign n30170 = n20345 ^ n18294 ^ n5916 ;
  assign n30171 = n18289 & ~n30170 ;
  assign n30172 = n30171 ^ n17601 ^ 1'b0 ;
  assign n30168 = x40 & x225 ;
  assign n30169 = n30168 ^ n2728 ^ 1'b0 ;
  assign n30173 = n30172 ^ n30169 ^ 1'b0 ;
  assign n30174 = n9356 ^ n5722 ^ 1'b0 ;
  assign n30175 = n15932 ^ n6621 ^ n2644 ;
  assign n30176 = n30175 ^ n17755 ^ 1'b0 ;
  assign n30177 = n30174 & n30176 ;
  assign n30178 = ( ~x22 & n2534 ) | ( ~x22 & n24116 ) | ( n2534 & n24116 ) ;
  assign n30179 = n30178 ^ n19083 ^ 1'b0 ;
  assign n30180 = n7381 & n30179 ;
  assign n30181 = n30180 ^ n9622 ^ 1'b0 ;
  assign n30182 = ~n2332 & n26943 ;
  assign n30183 = n20828 & n30182 ;
  assign n30185 = n7573 & ~n17071 ;
  assign n30186 = n19722 & n30185 ;
  assign n30184 = ~n22951 & n25905 ;
  assign n30187 = n30186 ^ n30184 ^ n20809 ;
  assign n30188 = ~n6176 & n25914 ;
  assign n30189 = n2722 & ~n3875 ;
  assign n30190 = n30189 ^ n12680 ^ n9222 ;
  assign n30191 = ( n6584 & n30188 ) | ( n6584 & n30190 ) | ( n30188 & n30190 ) ;
  assign n30192 = ~x116 & n6938 ;
  assign n30193 = ( ~n20823 & n30161 ) | ( ~n20823 & n30192 ) | ( n30161 & n30192 ) ;
  assign n30194 = n1259 | n4306 ;
  assign n30195 = n30194 ^ n2818 ^ 1'b0 ;
  assign n30196 = ~n26298 & n30195 ;
  assign n30197 = n14969 & ~n22367 ;
  assign n30198 = n30197 ^ n24904 ^ n1448 ;
  assign n30199 = n30196 & n30198 ;
  assign n30200 = n19180 & n30199 ;
  assign n30201 = n9780 & ~n29582 ;
  assign n30202 = n14877 & n30201 ;
  assign n30203 = n30202 ^ n3506 ^ 1'b0 ;
  assign n30204 = n7199 & n10144 ;
  assign n30205 = n30204 ^ n9475 ^ 1'b0 ;
  assign n30206 = n648 & n30205 ;
  assign n30207 = n12291 ^ n277 ^ 1'b0 ;
  assign n30208 = ~n28443 & n30207 ;
  assign n30209 = ( n13996 & ~n28959 ) | ( n13996 & n30208 ) | ( ~n28959 & n30208 ) ;
  assign n30210 = n30209 ^ n7972 ^ 1'b0 ;
  assign n30211 = n16974 ^ n6189 ^ 1'b0 ;
  assign n30212 = n2315 & n30211 ;
  assign n30215 = n12373 ^ n9364 ^ 1'b0 ;
  assign n30216 = n5314 | n30215 ;
  assign n30213 = n26498 ^ n2441 ^ 1'b0 ;
  assign n30214 = n6693 & n30213 ;
  assign n30217 = n30216 ^ n30214 ^ n20452 ;
  assign n30218 = ( n8497 & ~n18498 ) | ( n8497 & n30217 ) | ( ~n18498 & n30217 ) ;
  assign n30219 = n28280 ^ n21275 ^ 1'b0 ;
  assign n30220 = ~n12377 & n30219 ;
  assign n30221 = n9885 ^ n6628 ^ 1'b0 ;
  assign n30222 = n30221 ^ n28541 ^ 1'b0 ;
  assign n30223 = n915 & ~n25394 ;
  assign n30224 = n16845 ^ n7191 ^ 1'b0 ;
  assign n30225 = n14631 & ~n30224 ;
  assign n30226 = n11072 ^ n9805 ^ 1'b0 ;
  assign n30227 = n14216 | n30226 ;
  assign n30228 = ( n5198 & n18373 ) | ( n5198 & ~n30227 ) | ( n18373 & ~n30227 ) ;
  assign n30229 = n30228 ^ n8833 ^ 1'b0 ;
  assign n30230 = n30225 & n30229 ;
  assign n30231 = n29684 ^ n8423 ^ 1'b0 ;
  assign n30232 = n23213 ^ n10192 ^ 1'b0 ;
  assign n30233 = n13189 & n30232 ;
  assign n30234 = ~n25824 & n30233 ;
  assign n30235 = n19308 & n30234 ;
  assign n30236 = n6602 | n14567 ;
  assign n30237 = n30236 ^ n9099 ^ 1'b0 ;
  assign n30238 = ~n17270 & n22992 ;
  assign n30239 = n3624 & n30238 ;
  assign n30240 = n20737 ^ n13832 ^ 1'b0 ;
  assign n30241 = n5387 & ~n5461 ;
  assign n30242 = ~n28683 & n30241 ;
  assign n30243 = n15671 & ~n17038 ;
  assign n30244 = n17209 ^ n4995 ^ 1'b0 ;
  assign n30245 = n12194 | n30244 ;
  assign n30246 = n30243 | n30245 ;
  assign n30247 = n30246 ^ n6203 ^ 1'b0 ;
  assign n30248 = n7815 ^ n5879 ^ 1'b0 ;
  assign n30249 = n1993 | n5243 ;
  assign n30250 = n30249 ^ n4148 ^ 1'b0 ;
  assign n30251 = ~n803 & n30250 ;
  assign n30252 = n2372 & n30251 ;
  assign n30253 = n20591 ^ n933 ^ 1'b0 ;
  assign n30254 = n30253 ^ n28914 ^ 1'b0 ;
  assign n30255 = ( n5507 & ~n21069 ) | ( n5507 & n28598 ) | ( ~n21069 & n28598 ) ;
  assign n30256 = n30255 ^ n3185 ^ 1'b0 ;
  assign n30257 = n12282 | n18189 ;
  assign n30258 = n30257 ^ n29046 ^ 1'b0 ;
  assign n30259 = n30258 ^ n9331 ^ 1'b0 ;
  assign n30260 = n19820 & ~n24465 ;
  assign n30261 = n28394 ^ n26599 ^ 1'b0 ;
  assign n30262 = n30260 & ~n30261 ;
  assign n30263 = ~n11351 & n12715 ;
  assign n30264 = n14957 & ~n30263 ;
  assign n30265 = n7200 ^ n3170 ^ 1'b0 ;
  assign n30266 = n6058 ^ n305 ^ 1'b0 ;
  assign n30267 = n30265 | n30266 ;
  assign n30268 = n10091 & ~n29263 ;
  assign n30269 = n10312 & n30268 ;
  assign n30270 = n29569 ^ n6624 ^ 1'b0 ;
  assign n30271 = ~n5103 & n30270 ;
  assign n30272 = n26567 ^ n8898 ^ n8897 ;
  assign n30273 = x167 & ~n4278 ;
  assign n30274 = ~n7219 & n30273 ;
  assign n30275 = n30274 ^ n10288 ^ n7172 ;
  assign n30276 = n26656 ^ n23199 ^ n14481 ;
  assign n30277 = ~n10978 & n12798 ;
  assign n30278 = n14269 ^ n9175 ^ 1'b0 ;
  assign n30279 = ~n1970 & n30278 ;
  assign n30280 = n8062 ^ n560 ^ 1'b0 ;
  assign n30281 = ( n2289 & ~n9695 ) | ( n2289 & n30280 ) | ( ~n9695 & n30280 ) ;
  assign n30282 = n21185 ^ n9576 ^ 1'b0 ;
  assign n30283 = n11236 & ~n30282 ;
  assign n30284 = n25368 ^ n11830 ^ 1'b0 ;
  assign n30285 = n19264 | n30284 ;
  assign n30286 = n6801 & n10786 ;
  assign n30287 = n29754 ^ n3710 ^ 1'b0 ;
  assign n30288 = ( n9946 & ~n12293 ) | ( n9946 & n13297 ) | ( ~n12293 & n13297 ) ;
  assign n30289 = n28550 ^ n2210 ^ 1'b0 ;
  assign n30290 = ~n1514 & n20320 ;
  assign n30291 = n30290 ^ n5675 ^ 1'b0 ;
  assign n30292 = n10867 ^ n5980 ^ 1'b0 ;
  assign n30293 = n19855 & n30292 ;
  assign n30294 = n2118 & n14469 ;
  assign n30295 = n13662 ^ n1762 ^ 1'b0 ;
  assign n30296 = n13768 & n30295 ;
  assign n30297 = n30296 ^ n10781 ^ 1'b0 ;
  assign n30298 = n15990 ^ n4326 ^ 1'b0 ;
  assign n30299 = n5025 ^ n3554 ^ 1'b0 ;
  assign n30300 = n22503 ^ n20866 ^ 1'b0 ;
  assign n30301 = x37 & ~n4594 ;
  assign n30302 = n30301 ^ n15593 ^ 1'b0 ;
  assign n30303 = n27558 ^ n14218 ^ 1'b0 ;
  assign n30304 = n16791 & ~n30303 ;
  assign n30305 = n13292 & n16474 ;
  assign n30306 = n25224 ^ n6558 ^ n2441 ;
  assign n30307 = ( n7802 & n11134 ) | ( n7802 & ~n24119 ) | ( n11134 & ~n24119 ) ;
  assign n30308 = ~x170 & n25949 ;
  assign n30309 = n19046 ^ n766 ^ 1'b0 ;
  assign n30310 = n30308 & ~n30309 ;
  assign n30311 = ~n12914 & n13649 ;
  assign n30312 = ~n30310 & n30311 ;
  assign n30313 = n13758 & n16612 ;
  assign n30314 = ~n5010 & n30313 ;
  assign n30315 = n7208 & ~n30314 ;
  assign n30316 = n30315 ^ n1972 ^ 1'b0 ;
  assign n30317 = n7843 & n23049 ;
  assign n30318 = n30317 ^ n14113 ^ 1'b0 ;
  assign n30319 = n8819 & ~n24117 ;
  assign n30321 = n6865 & n10964 ;
  assign n30320 = n18270 ^ n17642 ^ 1'b0 ;
  assign n30322 = n30321 ^ n30320 ^ 1'b0 ;
  assign n30323 = ~n21922 & n23186 ;
  assign n30324 = n16254 ^ n2673 ^ x59 ;
  assign n30325 = n18691 ^ n12977 ^ 1'b0 ;
  assign n30326 = n3993 ^ x203 ^ 1'b0 ;
  assign n30327 = ~n23343 & n29787 ;
  assign n30328 = n3664 & ~n10915 ;
  assign n30329 = n755 & n15307 ;
  assign n30330 = n10405 & n26648 ;
  assign n30331 = n1900 ^ n1215 ^ 1'b0 ;
  assign n30332 = n4407 & ~n16229 ;
  assign n30333 = n30332 ^ n23151 ^ 1'b0 ;
  assign n30334 = n10970 & ~n16631 ;
  assign n30335 = ( n1213 & ~n8229 ) | ( n1213 & n9263 ) | ( ~n8229 & n9263 ) ;
  assign n30336 = n17437 & ~n30335 ;
  assign n30337 = ~n3504 & n5775 ;
  assign n30338 = ~n24156 & n30337 ;
  assign n30339 = n10699 ^ n2680 ^ 1'b0 ;
  assign n30340 = ~n30338 & n30339 ;
  assign n30341 = n25819 ^ n10976 ^ 1'b0 ;
  assign n30342 = n3066 & ~n18716 ;
  assign n30343 = n18945 ^ n17483 ^ 1'b0 ;
  assign n30344 = n30343 ^ n11043 ^ n6808 ;
  assign n30345 = ~n20425 & n30344 ;
  assign n30346 = n25393 ^ n24089 ^ 1'b0 ;
  assign n30347 = n12473 ^ n3283 ^ 1'b0 ;
  assign n30348 = ~n9916 & n14354 ;
  assign n30349 = ( n6851 & n23660 ) | ( n6851 & ~n30348 ) | ( n23660 & ~n30348 ) ;
  assign n30350 = n1821 & n20879 ;
  assign n30351 = n30350 ^ n15320 ^ 1'b0 ;
  assign n30352 = n30349 & n30351 ;
  assign n30353 = n23242 ^ n5209 ^ 1'b0 ;
  assign n30356 = x80 & ~n3608 ;
  assign n30357 = ~n1701 & n30356 ;
  assign n30354 = n2712 | n19641 ;
  assign n30355 = n12642 & ~n30354 ;
  assign n30358 = n30357 ^ n30355 ^ n1489 ;
  assign n30359 = n27653 ^ n1070 ^ 1'b0 ;
  assign n30360 = n18156 & ~n30359 ;
  assign n30361 = n3554 & ~n20804 ;
  assign n30362 = n30361 ^ n29155 ^ n10336 ;
  assign n30363 = ~n7856 & n24512 ;
  assign n30364 = n30363 ^ n21229 ^ 1'b0 ;
  assign n30365 = ~n4342 & n26350 ;
  assign n30366 = n30365 ^ n3797 ^ 1'b0 ;
  assign n30367 = n13763 | n22549 ;
  assign n30368 = n30366 & n30367 ;
  assign n30369 = ~n8613 & n8850 ;
  assign n30370 = n29351 ^ n9120 ^ n6750 ;
  assign n30371 = ~n8086 & n30370 ;
  assign n30372 = n8833 ^ n5525 ^ 1'b0 ;
  assign n30373 = n1270 & n13950 ;
  assign n30374 = n30373 ^ n6643 ^ 1'b0 ;
  assign n30375 = n30374 ^ n14079 ^ 1'b0 ;
  assign n30376 = n14518 ^ n13664 ^ 1'b0 ;
  assign n30377 = n8342 | n30376 ;
  assign n30378 = ( ~n27594 & n30375 ) | ( ~n27594 & n30377 ) | ( n30375 & n30377 ) ;
  assign n30379 = n6558 | n22859 ;
  assign n30380 = n21073 ^ x36 ^ 1'b0 ;
  assign n30381 = n11174 & n17447 ;
  assign n30382 = n4973 & n30381 ;
  assign n30384 = n6814 ^ n6683 ^ 1'b0 ;
  assign n30385 = n16460 | n30384 ;
  assign n30383 = n29645 ^ n19278 ^ n7006 ;
  assign n30386 = n30385 ^ n30383 ^ 1'b0 ;
  assign n30387 = ~n3847 & n30386 ;
  assign n30388 = n15714 ^ n3485 ^ 1'b0 ;
  assign n30389 = n22375 ^ n8584 ^ 1'b0 ;
  assign n30390 = n30388 | n30389 ;
  assign n30391 = n19117 & ~n30390 ;
  assign n30392 = ~n30387 & n30391 ;
  assign n30393 = n12773 & ~n27510 ;
  assign n30394 = n30393 ^ n16855 ^ 1'b0 ;
  assign n30395 = ~n17518 & n30394 ;
  assign n30397 = n4284 ^ n1625 ^ n296 ;
  assign n30396 = ~n16189 & n27194 ;
  assign n30398 = n30397 ^ n30396 ^ 1'b0 ;
  assign n30399 = ~n17941 & n30398 ;
  assign n30400 = n10551 ^ n1509 ^ 1'b0 ;
  assign n30401 = ( n2600 & ~n30399 ) | ( n2600 & n30400 ) | ( ~n30399 & n30400 ) ;
  assign n30402 = n30401 ^ n14591 ^ n11188 ;
  assign n30403 = n25638 | n30402 ;
  assign n30404 = ~n6196 & n7371 ;
  assign n30405 = n30404 ^ n21122 ^ n16348 ;
  assign n30406 = n3570 ^ n3077 ^ 1'b0 ;
  assign n30407 = ( n2357 & n13316 ) | ( n2357 & n30406 ) | ( n13316 & n30406 ) ;
  assign n30408 = n4542 & ~n30407 ;
  assign n30409 = ~n9835 & n15941 ;
  assign n30410 = ~n9088 & n30409 ;
  assign n30411 = ~n14869 & n30410 ;
  assign n30412 = ( n13066 & n20604 ) | ( n13066 & ~n24672 ) | ( n20604 & ~n24672 ) ;
  assign n30413 = n21770 | n25446 ;
  assign n30414 = n20788 & ~n23004 ;
  assign n30415 = n20206 ^ n8474 ^ 1'b0 ;
  assign n30416 = n15768 ^ n13464 ^ 1'b0 ;
  assign n30417 = n8395 & n11509 ;
  assign n30418 = ( n8415 & n23941 ) | ( n8415 & n30417 ) | ( n23941 & n30417 ) ;
  assign n30419 = ~n6034 & n18937 ;
  assign n30420 = n6665 | n21161 ;
  assign n30421 = ( n6501 & n30419 ) | ( n6501 & ~n30420 ) | ( n30419 & ~n30420 ) ;
  assign n30422 = n8264 | n13705 ;
  assign n30423 = n20011 ^ n10432 ^ 1'b0 ;
  assign n30424 = n4283 & ~n30423 ;
  assign n30425 = n30422 & n30424 ;
  assign n30426 = n11136 & n12231 ;
  assign n30427 = ~n4376 & n10391 ;
  assign n30428 = n15107 & n20950 ;
  assign n30429 = n30427 & n30428 ;
  assign n30430 = n6232 & n10783 ;
  assign n30431 = n30430 ^ n26562 ^ 1'b0 ;
  assign n30432 = n5223 & ~n8266 ;
  assign n30433 = ~n30431 & n30432 ;
  assign n30434 = n16070 & ~n16187 ;
  assign n30435 = ~n5644 & n30434 ;
  assign n30436 = n27779 & n30435 ;
  assign n30437 = ( n2344 & ~n3261 ) | ( n2344 & n15150 ) | ( ~n3261 & n15150 ) ;
  assign n30438 = n25221 ^ n21783 ^ 1'b0 ;
  assign n30439 = n18518 & ~n30438 ;
  assign n30440 = ( n1663 & ~n4753 ) | ( n1663 & n12289 ) | ( ~n4753 & n12289 ) ;
  assign n30442 = n11786 ^ n6233 ^ 1'b0 ;
  assign n30443 = n16962 | n30442 ;
  assign n30441 = n8774 ^ n1234 ^ 1'b0 ;
  assign n30444 = n30443 ^ n30441 ^ n11728 ;
  assign n30445 = n18964 ^ n1291 ^ 1'b0 ;
  assign n30446 = n6727 | n30445 ;
  assign n30447 = n6704 | n28597 ;
  assign n30448 = n30447 ^ n17967 ^ 1'b0 ;
  assign n30449 = n15005 ^ n2737 ^ 1'b0 ;
  assign n30450 = ~n10657 & n30449 ;
  assign n30451 = ~n6780 & n14531 ;
  assign n30452 = ~n474 & n30451 ;
  assign n30453 = n21817 & ~n26683 ;
  assign n30454 = n21458 ^ n12867 ^ 1'b0 ;
  assign n30455 = n8565 & n17281 ;
  assign n30456 = ~n10947 & n30455 ;
  assign n30457 = n1769 | n5054 ;
  assign n30458 = n30456 & ~n30457 ;
  assign n30459 = n867 & n17558 ;
  assign n30460 = ~n10293 & n30459 ;
  assign n30464 = n16168 ^ n10830 ^ 1'b0 ;
  assign n30465 = ( ~n10264 & n12966 ) | ( ~n10264 & n30464 ) | ( n12966 & n30464 ) ;
  assign n30461 = ~n833 & n11353 ;
  assign n30462 = ~n2031 & n30461 ;
  assign n30463 = n30462 ^ n13895 ^ n5637 ;
  assign n30466 = n30465 ^ n30463 ^ 1'b0 ;
  assign n30467 = n30466 ^ n19586 ^ n5765 ;
  assign n30468 = ~n4776 & n7918 ;
  assign n30469 = n21229 & n30468 ;
  assign n30470 = n30469 ^ n23533 ^ 1'b0 ;
  assign n30471 = ( n998 & ~n11963 ) | ( n998 & n26636 ) | ( ~n11963 & n26636 ) ;
  assign n30472 = n19481 ^ n16943 ^ 1'b0 ;
  assign n30473 = n2652 ^ n1869 ^ 1'b0 ;
  assign n30474 = n13533 & ~n30473 ;
  assign n30475 = ~n14412 & n30474 ;
  assign n30476 = n25543 ^ n21768 ^ 1'b0 ;
  assign n30477 = ~n2365 & n6292 ;
  assign n30478 = ( n10944 & n15390 ) | ( n10944 & n29657 ) | ( n15390 & n29657 ) ;
  assign n30483 = n12361 ^ n2930 ^ 1'b0 ;
  assign n30479 = n8844 ^ n6194 ^ 1'b0 ;
  assign n30480 = n14856 & ~n30479 ;
  assign n30481 = ( ~n23111 & n25275 ) | ( ~n23111 & n30480 ) | ( n25275 & n30480 ) ;
  assign n30482 = ( n7206 & ~n10915 ) | ( n7206 & n30481 ) | ( ~n10915 & n30481 ) ;
  assign n30484 = n30483 ^ n30482 ^ 1'b0 ;
  assign n30485 = n18267 & n27527 ;
  assign n30486 = n25269 & n30485 ;
  assign n30487 = ( n9642 & ~n17869 ) | ( n9642 & n30486 ) | ( ~n17869 & n30486 ) ;
  assign n30488 = n1442 & ~n19890 ;
  assign n30489 = ~n25475 & n30488 ;
  assign n30490 = n402 | n20847 ;
  assign n30491 = ( n20988 & ~n23688 ) | ( n20988 & n30490 ) | ( ~n23688 & n30490 ) ;
  assign n30492 = n29100 & ~n30491 ;
  assign n30493 = ( n13230 & n23101 ) | ( n13230 & ~n25694 ) | ( n23101 & ~n25694 ) ;
  assign n30494 = n6068 | n7110 ;
  assign n30495 = n2518 | n16838 ;
  assign n30496 = n13366 & n21828 ;
  assign n30497 = ~n2275 & n24684 ;
  assign n30498 = n30497 ^ n15142 ^ 1'b0 ;
  assign n30501 = n11282 | n18767 ;
  assign n30499 = n606 & n10408 ;
  assign n30500 = n30499 ^ n28506 ^ 1'b0 ;
  assign n30502 = n30501 ^ n30500 ^ 1'b0 ;
  assign n30503 = ( ~n3150 & n16282 ) | ( ~n3150 & n18918 ) | ( n16282 & n18918 ) ;
  assign n30504 = n11954 ^ n9236 ^ n7752 ;
  assign n30505 = n27242 | n30504 ;
  assign n30506 = n11332 ^ n3374 ^ 1'b0 ;
  assign n30507 = n30505 & ~n30506 ;
  assign n30508 = ~n15887 & n26298 ;
  assign n30509 = n30508 ^ n13280 ^ 1'b0 ;
  assign n30510 = n12083 ^ n6103 ^ 1'b0 ;
  assign n30511 = n24062 & ~n30510 ;
  assign n30512 = ( ~n7719 & n13651 ) | ( ~n7719 & n20161 ) | ( n13651 & n20161 ) ;
  assign n30513 = n1705 & ~n30512 ;
  assign n30514 = n30513 ^ n17588 ^ n8356 ;
  assign n30515 = n14558 ^ n11069 ^ 1'b0 ;
  assign n30516 = n8919 | n30515 ;
  assign n30517 = n3954 | n30516 ;
  assign n30518 = n20362 ^ n18610 ^ n9139 ;
  assign n30519 = n1752 & ~n11918 ;
  assign n30520 = ~n30518 & n30519 ;
  assign n30521 = ( n1801 & ~n30517 ) | ( n1801 & n30520 ) | ( ~n30517 & n30520 ) ;
  assign n30522 = n1544 & n8850 ;
  assign n30523 = n1486 & ~n30522 ;
  assign n30524 = n14638 ^ n3869 ^ n3618 ;
  assign n30525 = n12415 ^ n6853 ^ 1'b0 ;
  assign n30526 = n30524 & ~n30525 ;
  assign n30527 = ~n536 & n20770 ;
  assign n30528 = n4772 | n22484 ;
  assign n30529 = n20651 ^ n10810 ^ n462 ;
  assign n30530 = ~n531 & n20559 ;
  assign n30531 = n30529 & n30530 ;
  assign n30532 = n30531 ^ n8128 ^ n2055 ;
  assign n30533 = n2536 & ~n30532 ;
  assign n30534 = n30533 ^ n5232 ^ 1'b0 ;
  assign n30535 = n401 & ~n20285 ;
  assign n30536 = n12396 & ~n30535 ;
  assign n30537 = n30536 ^ n2939 ^ 1'b0 ;
  assign n30538 = n6352 & ~n9930 ;
  assign n30539 = n20837 ^ x165 ^ 1'b0 ;
  assign n30540 = n30539 ^ n12047 ^ 1'b0 ;
  assign n30541 = ~n19091 & n30540 ;
  assign n30542 = ~n30538 & n30541 ;
  assign n30543 = n22469 ^ n14429 ^ n2232 ;
  assign n30544 = ~n16827 & n20795 ;
  assign n30545 = n3714 & n30544 ;
  assign n30546 = ~n30543 & n30545 ;
  assign n30547 = x1 & n1484 ;
  assign n30548 = ~n732 & n30547 ;
  assign n30549 = n16134 ^ n6186 ^ 1'b0 ;
  assign n30550 = ~n30548 & n30549 ;
  assign n30551 = ( x217 & ~n4658 ) | ( x217 & n12047 ) | ( ~n4658 & n12047 ) ;
  assign n30552 = n15001 & n21912 ;
  assign n30553 = n15370 ^ n10300 ^ 1'b0 ;
  assign n30554 = ~n6591 & n10315 ;
  assign n30563 = n10525 ^ n8032 ^ 1'b0 ;
  assign n30564 = n10636 ^ n4641 ^ 1'b0 ;
  assign n30565 = n30563 & ~n30564 ;
  assign n30555 = ~n5835 & n22490 ;
  assign n30556 = n1677 & n30555 ;
  assign n30557 = n30556 ^ n11824 ^ 1'b0 ;
  assign n30558 = ~n8760 & n30557 ;
  assign n30559 = ~n15307 & n30558 ;
  assign n30560 = n880 | n30559 ;
  assign n30561 = n22031 | n30560 ;
  assign n30562 = n30561 ^ n19180 ^ n12140 ;
  assign n30566 = n30565 ^ n30562 ^ 1'b0 ;
  assign n30567 = n30554 | n30566 ;
  assign n30568 = n30567 ^ n3958 ^ 1'b0 ;
  assign n30569 = ~n24889 & n30568 ;
  assign n30570 = n4797 ^ n2004 ^ 1'b0 ;
  assign n30571 = ~n21481 & n30570 ;
  assign n30572 = n21630 ^ n519 ^ 1'b0 ;
  assign n30573 = n16140 | n23155 ;
  assign n30574 = ~n30572 & n30573 ;
  assign n30575 = n3246 & n30574 ;
  assign n30576 = ~n7269 & n9047 ;
  assign n30577 = n30576 ^ n968 ^ 1'b0 ;
  assign n30578 = n16839 ^ n1230 ^ 1'b0 ;
  assign n30579 = ~n30577 & n30578 ;
  assign n30580 = n10515 ^ n10438 ^ 1'b0 ;
  assign n30581 = n4562 & ~n17782 ;
  assign n30582 = n16811 & n25973 ;
  assign n30583 = n3600 & n15360 ;
  assign n30584 = n30583 ^ n5231 ^ 1'b0 ;
  assign n30585 = n3244 | n26305 ;
  assign n30587 = n6242 & n13583 ;
  assign n30586 = n12408 & ~n19677 ;
  assign n30588 = n30587 ^ n30586 ^ 1'b0 ;
  assign n30589 = ( n15317 & ~n18831 ) | ( n15317 & n21717 ) | ( ~n18831 & n21717 ) ;
  assign n30590 = n22215 ^ n1208 ^ 1'b0 ;
  assign n30591 = ~n20328 & n30590 ;
  assign n30592 = ~n23057 & n27111 ;
  assign n30593 = n30592 ^ n18043 ^ 1'b0 ;
  assign n30594 = n1703 & ~n19616 ;
  assign n30595 = n19863 | n30594 ;
  assign n30596 = n24835 & ~n30595 ;
  assign n30597 = n3995 & ~n20328 ;
  assign n30598 = n6314 & n30597 ;
  assign n30599 = n2281 | n30598 ;
  assign n30600 = n22408 & ~n30599 ;
  assign n30601 = n926 & n12319 ;
  assign n30602 = n30601 ^ n19281 ^ n2592 ;
  assign n30603 = n30600 | n30602 ;
  assign n30604 = n10198 ^ n9585 ^ 1'b0 ;
  assign n30605 = ~n12335 & n25091 ;
  assign n30606 = n8340 ^ x58 ^ 1'b0 ;
  assign n30607 = ~n23428 & n30606 ;
  assign n30608 = ~n30605 & n30607 ;
  assign n30609 = n30608 ^ n23567 ^ 1'b0 ;
  assign n30610 = n27468 | n29384 ;
  assign n30611 = n17589 ^ n2272 ^ 1'b0 ;
  assign n30612 = n9139 & n13685 ;
  assign n30613 = n30612 ^ n6756 ^ 1'b0 ;
  assign n30614 = n429 & n30613 ;
  assign n30615 = n24757 ^ n15055 ^ 1'b0 ;
  assign n30616 = n9072 & ~n30615 ;
  assign n30617 = ~n1750 & n5341 ;
  assign n30618 = ( n7799 & n26047 ) | ( n7799 & ~n30617 ) | ( n26047 & ~n30617 ) ;
  assign n30619 = n9099 | n19308 ;
  assign n30620 = ( n4001 & n6550 ) | ( n4001 & ~n30619 ) | ( n6550 & ~n30619 ) ;
  assign n30621 = n12725 | n14751 ;
  assign n30622 = n5535 & ~n30621 ;
  assign n30623 = ~n5661 & n14502 ;
  assign n30624 = n30623 ^ n5658 ^ 1'b0 ;
  assign n30625 = n24743 ^ n6421 ^ 1'b0 ;
  assign n30626 = n26224 & n30625 ;
  assign n30627 = x39 & n16534 ;
  assign n30628 = n6558 & n30627 ;
  assign n30629 = n30628 ^ n25269 ^ 1'b0 ;
  assign n30630 = ( n2264 & n14139 ) | ( n2264 & ~n23826 ) | ( n14139 & ~n23826 ) ;
  assign n30631 = n22099 ^ n15998 ^ n7367 ;
  assign n30632 = n2870 | n19244 ;
  assign n30633 = n30632 ^ n17755 ^ 1'b0 ;
  assign n30634 = n18459 | n20409 ;
  assign n30635 = n8377 & ~n30634 ;
  assign n30636 = ~n9032 & n21493 ;
  assign n30637 = n7352 & ~n8389 ;
  assign n30638 = n1483 & n30637 ;
  assign n30639 = ~n5656 & n17172 ;
  assign n30640 = n5285 & ~n25403 ;
  assign n30641 = n20458 & n23512 ;
  assign n30642 = n25186 ^ n5634 ^ 1'b0 ;
  assign n30643 = n13442 & n30642 ;
  assign n30644 = n8339 & n14294 ;
  assign n30645 = n30644 ^ n14299 ^ 1'b0 ;
  assign n30646 = ~n11838 & n20820 ;
  assign n30647 = x157 & n3460 ;
  assign n30648 = ~x157 & n30647 ;
  assign n30649 = ~n2361 & n30648 ;
  assign n30650 = ( ~n1235 & n12219 ) | ( ~n1235 & n30649 ) | ( n12219 & n30649 ) ;
  assign n30651 = n24465 ^ n12743 ^ 1'b0 ;
  assign n30652 = ~n30650 & n30651 ;
  assign n30653 = n22006 & n30652 ;
  assign n30654 = ~n30652 & n30653 ;
  assign n30655 = n12219 & n22139 ;
  assign n30656 = n30655 ^ n14040 ^ 1'b0 ;
  assign n30657 = n30656 ^ n5085 ^ 1'b0 ;
  assign n30658 = n12987 | n20883 ;
  assign n30659 = n30657 | n30658 ;
  assign n30660 = n3767 & ~n19828 ;
  assign n30661 = ( ~n3540 & n19526 ) | ( ~n3540 & n28110 ) | ( n19526 & n28110 ) ;
  assign n30662 = n4323 & n9404 ;
  assign n30663 = n30662 ^ n867 ^ 1'b0 ;
  assign n30664 = ( n4698 & n26031 ) | ( n4698 & ~n30663 ) | ( n26031 & ~n30663 ) ;
  assign n30665 = ( ~n7028 & n17062 ) | ( ~n7028 & n30664 ) | ( n17062 & n30664 ) ;
  assign n30666 = n12612 ^ n12176 ^ 1'b0 ;
  assign n30667 = n10245 & ~n30666 ;
  assign n30668 = n30667 ^ n15676 ^ 1'b0 ;
  assign n30669 = n6501 & ~n8395 ;
  assign n30670 = n24416 & n30669 ;
  assign n30671 = n1181 & n13048 ;
  assign n30672 = n4947 & n30671 ;
  assign n30673 = n9489 ^ n2748 ^ 1'b0 ;
  assign n30674 = ~n729 & n30673 ;
  assign n30675 = n10137 & ~n22483 ;
  assign n30676 = n30675 ^ n4276 ^ 1'b0 ;
  assign n30678 = ~n2484 & n22114 ;
  assign n30679 = n30678 ^ n9971 ^ 1'b0 ;
  assign n30677 = n6613 ^ x12 ^ 1'b0 ;
  assign n30680 = n30679 ^ n30677 ^ n1330 ;
  assign n30681 = n13635 ^ n5509 ^ 1'b0 ;
  assign n30682 = n7830 & ~n30681 ;
  assign n30683 = ( n11575 & ~n30680 ) | ( n11575 & n30682 ) | ( ~n30680 & n30682 ) ;
  assign n30684 = n2480 & ~n14435 ;
  assign n30685 = n1758 & ~n10520 ;
  assign n30686 = n10265 & n30685 ;
  assign n30687 = n14587 & ~n15564 ;
  assign n30689 = n4824 | n6192 ;
  assign n30688 = n7338 & ~n11529 ;
  assign n30690 = n30689 ^ n30688 ^ 1'b0 ;
  assign n30691 = ( n21652 & n23622 ) | ( n21652 & ~n30690 ) | ( n23622 & ~n30690 ) ;
  assign n30692 = n2558 & n21578 ;
  assign n30693 = ( n12671 & n23901 ) | ( n12671 & ~n30692 ) | ( n23901 & ~n30692 ) ;
  assign n30694 = n19751 ^ n15915 ^ 1'b0 ;
  assign n30695 = ~n7668 & n17316 ;
  assign n30696 = n15793 ^ n6947 ^ 1'b0 ;
  assign n30697 = n30695 & ~n30696 ;
  assign n30698 = n30697 ^ n16870 ^ 1'b0 ;
  assign n30699 = n24689 ^ n24593 ^ n8378 ;
  assign n30700 = n30699 ^ n5648 ^ 1'b0 ;
  assign n30701 = n308 | n30700 ;
  assign n30702 = n28209 ^ n9802 ^ 1'b0 ;
  assign n30703 = n21559 ^ n15366 ^ n681 ;
  assign n30705 = n2425 | n18253 ;
  assign n30706 = n30705 ^ n6756 ^ 1'b0 ;
  assign n30704 = n19209 & ~n23050 ;
  assign n30707 = n30706 ^ n30704 ^ 1'b0 ;
  assign n30708 = n30707 ^ n17091 ^ 1'b0 ;
  assign n30709 = n20259 ^ n4542 ^ 1'b0 ;
  assign n30710 = n23390 ^ n1453 ^ 1'b0 ;
  assign n30711 = ~n349 & n2501 ;
  assign n30712 = n30711 ^ n9692 ^ 1'b0 ;
  assign n30713 = n20382 ^ n19992 ^ 1'b0 ;
  assign n30714 = n15009 | n30713 ;
  assign n30715 = n10002 ^ n2019 ^ 1'b0 ;
  assign n30716 = n30715 ^ n18114 ^ n2085 ;
  assign n30717 = n8282 & ~n13114 ;
  assign n30718 = n9553 & n30717 ;
  assign n30719 = n30718 ^ n9009 ^ 1'b0 ;
  assign n30720 = n1996 & n25911 ;
  assign n30721 = n29082 ^ n6240 ^ n5497 ;
  assign n30722 = n7954 ^ n3812 ^ n3603 ;
  assign n30723 = n5562 & n30722 ;
  assign n30724 = ~n12078 & n19151 ;
  assign n30725 = ~n5641 & n30724 ;
  assign n30726 = n10276 ^ n2002 ^ 1'b0 ;
  assign n30727 = n4261 & ~n30726 ;
  assign n30728 = ~n23592 & n30727 ;
  assign n30729 = n30725 & n30728 ;
  assign n30730 = n2468 | n17200 ;
  assign n30731 = n19134 & n30571 ;
  assign n30732 = n30730 & n30731 ;
  assign n30733 = n16642 ^ n6242 ^ 1'b0 ;
  assign n30734 = n472 & ~n21873 ;
  assign n30735 = ~n660 & n30734 ;
  assign n30736 = n18385 ^ n10490 ^ 1'b0 ;
  assign n30737 = n12617 & n17028 ;
  assign n30738 = n30737 ^ n3997 ^ 1'b0 ;
  assign n30739 = ~n1038 & n30738 ;
  assign n30740 = n3801 & ~n30739 ;
  assign n30741 = ~n17350 & n30740 ;
  assign n30742 = n3552 | n12372 ;
  assign n30743 = n30742 ^ n7191 ^ 1'b0 ;
  assign n30744 = n10755 & n18218 ;
  assign n30745 = ( n2332 & ~n30743 ) | ( n2332 & n30744 ) | ( ~n30743 & n30744 ) ;
  assign n30746 = ~n5970 & n23971 ;
  assign n30747 = n14476 & n24817 ;
  assign n30748 = ~n1826 & n11764 ;
  assign n30749 = n30748 ^ n10066 ^ 1'b0 ;
  assign n30750 = n6257 | n30749 ;
  assign n30753 = x45 & ~n2853 ;
  assign n30754 = n17485 ^ n7766 ^ 1'b0 ;
  assign n30755 = ( n23546 & n30753 ) | ( n23546 & ~n30754 ) | ( n30753 & ~n30754 ) ;
  assign n30751 = ~n3420 & n3611 ;
  assign n30752 = n30751 ^ n9052 ^ 1'b0 ;
  assign n30756 = n30755 ^ n30752 ^ 1'b0 ;
  assign n30757 = n1233 & ~n6417 ;
  assign n30758 = n30757 ^ n5892 ^ 1'b0 ;
  assign n30759 = ~n675 & n9722 ;
  assign n30760 = n30759 ^ n2214 ^ 1'b0 ;
  assign n30761 = ( n16883 & n30410 ) | ( n16883 & n30760 ) | ( n30410 & n30760 ) ;
  assign n30762 = ( x63 & n30758 ) | ( x63 & n30761 ) | ( n30758 & n30761 ) ;
  assign n30763 = x67 & ~n8001 ;
  assign n30764 = n2120 & n30763 ;
  assign n30765 = n1760 & ~n30764 ;
  assign n30766 = n9891 ^ n6756 ^ 1'b0 ;
  assign n30767 = n7056 & ~n30766 ;
  assign n30768 = n7568 ^ n5008 ^ 1'b0 ;
  assign n30769 = ( n12069 & n30767 ) | ( n12069 & n30768 ) | ( n30767 & n30768 ) ;
  assign n30770 = n27212 ^ n9567 ^ 1'b0 ;
  assign n30771 = ~n30146 & n30770 ;
  assign n30773 = n29530 ^ n14035 ^ 1'b0 ;
  assign n30774 = n10886 & ~n30773 ;
  assign n30772 = n5532 ^ n2272 ^ 1'b0 ;
  assign n30775 = n30774 ^ n30772 ^ 1'b0 ;
  assign n30776 = n11667 & n30775 ;
  assign n30777 = ~n5535 & n27318 ;
  assign n30778 = n30777 ^ n27267 ^ 1'b0 ;
  assign n30779 = ( n3818 & ~n21481 ) | ( n3818 & n23755 ) | ( ~n21481 & n23755 ) ;
  assign n30780 = n12510 & n15981 ;
  assign n30781 = n30780 ^ n7943 ^ n6455 ;
  assign n30782 = n17230 & ~n30781 ;
  assign n30783 = n9039 ^ n1040 ^ 1'b0 ;
  assign n30784 = ~n18620 & n30783 ;
  assign n30785 = ~n18442 & n30784 ;
  assign n30786 = ~n28881 & n30785 ;
  assign n30787 = n6394 ^ n2138 ^ 1'b0 ;
  assign n30788 = n10248 & ~n12980 ;
  assign n30789 = ( n8603 & ~n16286 ) | ( n8603 & n30788 ) | ( ~n16286 & n30788 ) ;
  assign n30790 = ( n8437 & n11134 ) | ( n8437 & n30789 ) | ( n11134 & n30789 ) ;
  assign n30791 = ( n6808 & n7070 ) | ( n6808 & ~n27170 ) | ( n7070 & ~n27170 ) ;
  assign n30792 = n1356 | n4813 ;
  assign n30793 = n30792 ^ n11396 ^ 1'b0 ;
  assign n30794 = n11365 & ~n30793 ;
  assign n30795 = n15571 & n30794 ;
  assign n30796 = n1228 & n14802 ;
  assign n30797 = n30796 ^ n1683 ^ 1'b0 ;
  assign n30798 = n21400 & ~n30797 ;
  assign n30799 = n24984 | n25750 ;
  assign n30802 = n1683 & n4513 ;
  assign n30803 = n30802 ^ n6174 ^ 1'b0 ;
  assign n30800 = n2726 ^ n2019 ^ 1'b0 ;
  assign n30801 = ~n1302 & n30800 ;
  assign n30804 = n30803 ^ n30801 ^ n5846 ;
  assign n30805 = n14481 | n15955 ;
  assign n30806 = ~n4827 & n18296 ;
  assign n30807 = n1404 & n30806 ;
  assign n30808 = n9544 ^ n6375 ^ 1'b0 ;
  assign n30809 = ~n9247 & n30808 ;
  assign n30810 = n30809 ^ n1551 ^ 1'b0 ;
  assign n30811 = n30810 ^ n10497 ^ 1'b0 ;
  assign n30812 = ~n30807 & n30811 ;
  assign n30814 = ( n2712 & n3764 ) | ( n2712 & n5060 ) | ( n3764 & n5060 ) ;
  assign n30813 = n14631 | n25343 ;
  assign n30815 = n30814 ^ n30813 ^ n17060 ;
  assign n30816 = ( ~n3606 & n7584 ) | ( ~n3606 & n20641 ) | ( n7584 & n20641 ) ;
  assign n30817 = n1733 | n10354 ;
  assign n30818 = n30026 | n30817 ;
  assign n30819 = n5859 & n22999 ;
  assign n30820 = n14723 & n23106 ;
  assign n30821 = n10816 | n22221 ;
  assign n30822 = n19533 & n30821 ;
  assign n30823 = n18191 & n25803 ;
  assign n30824 = ( n4769 & n7523 ) | ( n4769 & n10404 ) | ( n7523 & n10404 ) ;
  assign n30825 = x247 & n13165 ;
  assign n30826 = n30824 & n30825 ;
  assign n30828 = n17458 | n23595 ;
  assign n30827 = n4450 & n12760 ;
  assign n30829 = n30828 ^ n30827 ^ 1'b0 ;
  assign n30830 = n22109 ^ n10125 ^ 1'b0 ;
  assign n30831 = n1209 & ~n10718 ;
  assign n30832 = n30831 ^ n11337 ^ 1'b0 ;
  assign n30833 = n4286 & n23865 ;
  assign n30834 = n12803 & n30833 ;
  assign n30835 = n27048 ^ n2371 ^ 1'b0 ;
  assign n30836 = ~n11742 & n30835 ;
  assign n30837 = n7636 & n30836 ;
  assign n30838 = ~n2264 & n30837 ;
  assign n30839 = n28026 | n30838 ;
  assign n30840 = n30839 ^ n1731 ^ 1'b0 ;
  assign n30844 = ~n2332 & n3920 ;
  assign n30845 = ~n8815 & n30844 ;
  assign n30846 = n30845 ^ n21828 ^ n5645 ;
  assign n30841 = n7946 | n9622 ;
  assign n30842 = n30841 ^ n4383 ^ 1'b0 ;
  assign n30843 = n7429 & ~n30842 ;
  assign n30847 = n30846 ^ n30843 ^ 1'b0 ;
  assign n30848 = ( n2797 & n5217 ) | ( n2797 & n16552 ) | ( n5217 & n16552 ) ;
  assign n30849 = n30848 ^ n25966 ^ 1'b0 ;
  assign n30850 = n19440 & n30849 ;
  assign n30851 = n1442 & n13488 ;
  assign n30852 = ( n16651 & n19549 ) | ( n16651 & ~n30851 ) | ( n19549 & ~n30851 ) ;
  assign n30853 = n8516 ^ n6990 ^ n6401 ;
  assign n30854 = n18610 & n30853 ;
  assign n30855 = n3917 & ~n10460 ;
  assign n30856 = n30855 ^ n8477 ^ 1'b0 ;
  assign n30857 = n3695 & n20908 ;
  assign n30858 = n7127 | n30857 ;
  assign n30859 = n4335 | n30858 ;
  assign n30860 = ~n28443 & n30859 ;
  assign n30861 = n14006 & n30860 ;
  assign n30862 = n8701 | n10574 ;
  assign n30863 = n30862 ^ n5176 ^ 1'b0 ;
  assign n30864 = ~n15669 & n22228 ;
  assign n30865 = n30864 ^ n2531 ^ 1'b0 ;
  assign n30866 = ~n30863 & n30865 ;
  assign n30867 = n13319 | n30866 ;
  assign n30868 = n30861 & ~n30867 ;
  assign n30869 = n19629 ^ n1125 ^ 1'b0 ;
  assign n30870 = n11342 & n21915 ;
  assign n30871 = ~n3899 & n15780 ;
  assign n30872 = ( n12142 & n30870 ) | ( n12142 & n30871 ) | ( n30870 & n30871 ) ;
  assign n30873 = n9895 & ~n30872 ;
  assign n30874 = n30869 & n30873 ;
  assign n30875 = ~n6336 & n10262 ;
  assign n30876 = ~n12283 & n30875 ;
  assign n30877 = n22514 ^ n22385 ^ 1'b0 ;
  assign n30878 = ~n30876 & n30877 ;
  assign n30879 = n1311 | n15111 ;
  assign n30880 = n30879 ^ n29754 ^ n14399 ;
  assign n30881 = ~n626 & n19583 ;
  assign n30882 = n30881 ^ n20774 ^ 1'b0 ;
  assign n30883 = n9733 | n20022 ;
  assign n30884 = n5724 & ~n30883 ;
  assign n30885 = n19226 | n30884 ;
  assign n30886 = ( ~n2224 & n30882 ) | ( ~n2224 & n30885 ) | ( n30882 & n30885 ) ;
  assign n30887 = n17400 ^ n12061 ^ n11141 ;
  assign n30888 = ( ~n6212 & n19195 ) | ( ~n6212 & n30887 ) | ( n19195 & n30887 ) ;
  assign n30889 = n8505 & ~n21138 ;
  assign n30890 = n5302 ^ n4876 ^ 1'b0 ;
  assign n30891 = n5230 | n8009 ;
  assign n30892 = n30891 ^ n29210 ^ 1'b0 ;
  assign n30893 = n8550 | n21822 ;
  assign n30894 = n30893 ^ n15701 ^ 1'b0 ;
  assign n30895 = n25456 ^ n21922 ^ 1'b0 ;
  assign n30896 = n16169 & ~n30895 ;
  assign n30897 = n11111 & n30896 ;
  assign n30898 = n21229 & ~n27818 ;
  assign n30899 = n11878 | n11976 ;
  assign n30900 = n30898 & ~n30899 ;
  assign n30901 = ( n12185 & n13083 ) | ( n12185 & n23211 ) | ( n13083 & n23211 ) ;
  assign n30902 = n15874 & n30901 ;
  assign n30903 = n30902 ^ n18638 ^ 1'b0 ;
  assign n30904 = n15756 | n16870 ;
  assign n30905 = n10003 & ~n30904 ;
  assign n30906 = n14300 ^ n4899 ^ 1'b0 ;
  assign n30907 = ~n11380 & n30906 ;
  assign n30908 = ( n21941 & n24500 ) | ( n21941 & n25438 ) | ( n24500 & n25438 ) ;
  assign n30909 = n15785 & ~n19912 ;
  assign n30910 = n2971 | n20288 ;
  assign n30911 = n329 | n20019 ;
  assign n30912 = n8584 | n30911 ;
  assign n30913 = n30912 ^ n2272 ^ 1'b0 ;
  assign n30914 = n14240 ^ n11719 ^ n7308 ;
  assign n30915 = n17665 & ~n18424 ;
  assign n30916 = n3760 & ~n5042 ;
  assign n30917 = n6734 | n22317 ;
  assign n30918 = n4024 & ~n30917 ;
  assign n30919 = n13216 ^ n6966 ^ 1'b0 ;
  assign n30920 = ( n30916 & ~n30918 ) | ( n30916 & n30919 ) | ( ~n30918 & n30919 ) ;
  assign n30921 = n25046 ^ n5850 ^ n462 ;
  assign n30922 = ~n1170 & n27131 ;
  assign n30923 = n18591 & n30922 ;
  assign n30928 = ~n5264 & n12606 ;
  assign n30929 = ( n3773 & n10400 ) | ( n3773 & n30928 ) | ( n10400 & n30928 ) ;
  assign n30925 = n26340 ^ n5888 ^ 1'b0 ;
  assign n30924 = n22538 ^ n20010 ^ 1'b0 ;
  assign n30926 = n30925 ^ n30924 ^ 1'b0 ;
  assign n30927 = n725 & n30926 ;
  assign n30930 = n30929 ^ n30927 ^ 1'b0 ;
  assign n30931 = n29586 & ~n30930 ;
  assign n30932 = n18805 & n22833 ;
  assign n30933 = ~n713 & n10083 ;
  assign n30934 = ~n14583 & n30933 ;
  assign n30936 = n5227 | n8340 ;
  assign n30937 = ~n3808 & n30936 ;
  assign n30938 = n5300 & n30937 ;
  assign n30935 = n14828 ^ n8011 ^ 1'b0 ;
  assign n30939 = n30938 ^ n30935 ^ 1'b0 ;
  assign n30940 = ~n1996 & n11989 ;
  assign n30941 = n30940 ^ n18626 ^ n10234 ;
  assign n30942 = n11767 ^ n2667 ^ 1'b0 ;
  assign n30943 = n30942 ^ n30067 ^ n5172 ;
  assign n30944 = ~n3554 & n30253 ;
  assign n30945 = n10755 ^ n7820 ^ 1'b0 ;
  assign n30946 = ~n5001 & n30945 ;
  assign n30947 = n30944 & n30946 ;
  assign n30948 = n5832 ^ n5125 ^ n304 ;
  assign n30949 = n5714 | n30948 ;
  assign n30950 = n24865 ^ n20710 ^ 1'b0 ;
  assign n30951 = n11843 & n30950 ;
  assign n30952 = n358 & n3923 ;
  assign n30953 = ~n3923 & n30952 ;
  assign n30954 = n5343 & n21504 ;
  assign n30955 = n30953 & n30954 ;
  assign n30956 = n5469 | n30955 ;
  assign n30957 = n5469 & ~n30956 ;
  assign n30958 = n4654 | n30957 ;
  assign n30959 = n30957 & ~n30958 ;
  assign n30960 = n3772 & n13240 ;
  assign n30961 = ~n13240 & n30960 ;
  assign n30962 = ~n30959 & n30961 ;
  assign n30964 = n1941 | n6349 ;
  assign n30965 = n1941 & ~n30964 ;
  assign n30966 = ~n2002 & n13377 ;
  assign n30967 = n2002 & n30966 ;
  assign n30968 = n30965 | n30967 ;
  assign n30969 = n30965 & ~n30968 ;
  assign n30963 = n7756 | n13159 ;
  assign n30970 = n30969 ^ n30963 ^ 1'b0 ;
  assign n30971 = n13350 ^ n5408 ^ 1'b0 ;
  assign n30972 = ~n3954 & n26334 ;
  assign n30973 = n3954 & n30972 ;
  assign n30974 = n30971 & ~n30973 ;
  assign n30975 = ~n30971 & n30974 ;
  assign n30978 = n13563 ^ n1571 ^ 1'b0 ;
  assign n30979 = n5396 & ~n30978 ;
  assign n30980 = n30978 & n30979 ;
  assign n30981 = n12609 | n30980 ;
  assign n30982 = n12609 & ~n30981 ;
  assign n30976 = n7190 ^ n4651 ^ 1'b0 ;
  assign n30977 = n795 | n30976 ;
  assign n30983 = n30982 ^ n30977 ^ 1'b0 ;
  assign n30984 = ~n30975 & n30983 ;
  assign n30985 = ( n30962 & n30970 ) | ( n30962 & n30984 ) | ( n30970 & n30984 ) ;
  assign n30986 = n7508 & n28823 ;
  assign n30987 = n25540 ^ n6966 ^ 1'b0 ;
  assign n30988 = ~n4034 & n21081 ;
  assign n30989 = ~n22951 & n30988 ;
  assign n30990 = n4521 | n12934 ;
  assign n30991 = ~n7333 & n26265 ;
  assign n30992 = ~n11689 & n30991 ;
  assign n30993 = n18167 ^ n16567 ^ 1'b0 ;
  assign n30994 = n30992 & ~n30993 ;
  assign n30995 = ( n11268 & n17687 ) | ( n11268 & ~n18605 ) | ( n17687 & ~n18605 ) ;
  assign n30996 = ~n2080 & n30995 ;
  assign n30997 = n16586 & n30996 ;
  assign n30998 = n8963 | n20141 ;
  assign n30999 = n15756 & ~n30998 ;
  assign n31000 = n5766 | n10012 ;
  assign n31001 = n31000 ^ n25655 ^ n24079 ;
  assign n31002 = n26319 ^ n11219 ^ n4668 ;
  assign n31003 = n19137 ^ n7334 ^ 1'b0 ;
  assign n31004 = n31003 ^ n19376 ^ n14326 ;
  assign n31005 = n31004 ^ n13263 ^ 1'b0 ;
  assign n31006 = n3439 & ~n7185 ;
  assign n31007 = n4086 ^ n385 ^ 1'b0 ;
  assign n31008 = n432 & ~n31007 ;
  assign n31009 = n31008 ^ n15649 ^ 1'b0 ;
  assign n31010 = n31006 & n31009 ;
  assign n31011 = n23202 ^ n6972 ^ 1'b0 ;
  assign n31012 = n15440 | n31011 ;
  assign n31013 = n15333 | n31012 ;
  assign n31014 = n31013 ^ n29230 ^ 1'b0 ;
  assign n31015 = n7509 ^ n4060 ^ 1'b0 ;
  assign n31016 = n19135 ^ n8416 ^ 1'b0 ;
  assign n31017 = ( n13162 & n16781 ) | ( n13162 & n31016 ) | ( n16781 & n31016 ) ;
  assign n31018 = n4607 & n31017 ;
  assign n31020 = n7645 ^ n1997 ^ 1'b0 ;
  assign n31021 = n12952 | n31020 ;
  assign n31019 = n13277 ^ n3587 ^ 1'b0 ;
  assign n31022 = n31021 ^ n31019 ^ 1'b0 ;
  assign n31023 = n29149 ^ n9177 ^ 1'b0 ;
  assign n31024 = n5170 | n31023 ;
  assign n31025 = n31024 ^ n27346 ^ 1'b0 ;
  assign n31026 = n24198 ^ n4500 ^ n3081 ;
  assign n31028 = n27127 ^ n9396 ^ n3175 ;
  assign n31027 = n1509 & n23131 ;
  assign n31029 = n31028 ^ n31027 ^ x98 ;
  assign n31030 = n27083 & ~n31029 ;
  assign n31031 = n20057 ^ n1565 ^ 1'b0 ;
  assign n31032 = ~n15552 & n17716 ;
  assign n31033 = n31032 ^ n21419 ^ 1'b0 ;
  assign n31034 = n16540 ^ n8789 ^ 1'b0 ;
  assign n31035 = n11721 ^ n5699 ^ n3769 ;
  assign n31036 = n1354 | n13611 ;
  assign n31037 = n20397 | n31036 ;
  assign n31038 = n2082 & n15984 ;
  assign n31039 = n31038 ^ n1090 ^ 1'b0 ;
  assign n31040 = n6967 | n13499 ;
  assign n31041 = n31040 ^ n25488 ^ 1'b0 ;
  assign n31042 = ( ~n2149 & n8348 ) | ( ~n2149 & n11956 ) | ( n8348 & n11956 ) ;
  assign n31043 = n31042 ^ n13894 ^ 1'b0 ;
  assign n31044 = x168 & n981 ;
  assign n31045 = ~n981 & n31044 ;
  assign n31046 = n1053 & ~n12215 ;
  assign n31047 = n31045 & n31046 ;
  assign n31048 = n1348 & n31047 ;
  assign n31049 = ~n7473 & n31048 ;
  assign n31050 = n1837 | n31049 ;
  assign n31051 = n31050 ^ n7293 ^ 1'b0 ;
  assign n31052 = ( ~n7151 & n9275 ) | ( ~n7151 & n31051 ) | ( n9275 & n31051 ) ;
  assign n31053 = n31052 ^ n19722 ^ n9469 ;
  assign n31054 = ~n22330 & n25828 ;
  assign n31055 = n31054 ^ n4862 ^ 1'b0 ;
  assign n31056 = n31055 ^ n27077 ^ 1'b0 ;
  assign n31057 = ~n31053 & n31056 ;
  assign n31058 = n1323 & n4469 ;
  assign n31059 = n28749 | n31058 ;
  assign n31060 = n26878 & ~n31059 ;
  assign n31061 = n17069 ^ n5228 ^ 1'b0 ;
  assign n31062 = n17026 & n31061 ;
  assign n31063 = n5176 & ~n8201 ;
  assign n31064 = n30557 & n31063 ;
  assign n31065 = ~n31062 & n31064 ;
  assign n31066 = n31065 ^ n4242 ^ 1'b0 ;
  assign n31067 = n20188 ^ n12165 ^ 1'b0 ;
  assign n31068 = ~n9977 & n31067 ;
  assign n31072 = n6442 & n17500 ;
  assign n31073 = ~n14693 & n31072 ;
  assign n31069 = n2969 & n30689 ;
  assign n31070 = ( ~n5805 & n17204 ) | ( ~n5805 & n31069 ) | ( n17204 & n31069 ) ;
  assign n31071 = ( n11915 & n19135 ) | ( n11915 & ~n31070 ) | ( n19135 & ~n31070 ) ;
  assign n31074 = n31073 ^ n31071 ^ 1'b0 ;
  assign n31075 = n3099 & n3182 ;
  assign n31076 = n14743 ^ n10250 ^ 1'b0 ;
  assign n31077 = n17129 ^ n890 ^ 1'b0 ;
  assign n31078 = n11452 ^ n11175 ^ 1'b0 ;
  assign n31079 = n6365 & ~n31078 ;
  assign n31080 = n18003 ^ n16148 ^ n4739 ;
  assign n31081 = ( n1650 & ~n7310 ) | ( n1650 & n24332 ) | ( ~n7310 & n24332 ) ;
  assign n31082 = ~n26493 & n31081 ;
  assign n31083 = n15837 ^ n5151 ^ 1'b0 ;
  assign n31084 = n7754 | n31083 ;
  assign n31085 = n15919 | n31084 ;
  assign n31086 = n31082 & ~n31085 ;
  assign n31087 = n12705 ^ n10132 ^ 1'b0 ;
  assign n31088 = ~n27137 & n31087 ;
  assign n31089 = n18134 ^ n4473 ^ 1'b0 ;
  assign n31090 = n15744 & ~n20429 ;
  assign n31091 = n18879 & n31090 ;
  assign n31092 = n24843 ^ n9087 ^ n1627 ;
  assign n31093 = n5272 & ~n31092 ;
  assign n31094 = n10223 ^ n1266 ^ 1'b0 ;
  assign n31095 = n1724 & n2851 ;
  assign n31096 = n31095 ^ n18805 ^ 1'b0 ;
  assign n31097 = ~n4378 & n31096 ;
  assign n31098 = n31097 ^ n29019 ^ 1'b0 ;
  assign n31099 = n22984 ^ n12503 ^ 1'b0 ;
  assign n31100 = n17243 & ~n31099 ;
  assign n31101 = n8120 ^ n2680 ^ 1'b0 ;
  assign n31102 = n1000 & n31101 ;
  assign n31103 = n28663 ^ n27944 ^ 1'b0 ;
  assign n31104 = n10859 | n28677 ;
  assign n31105 = n29124 ^ n18357 ^ 1'b0 ;
  assign n31106 = n9047 & n31105 ;
  assign n31107 = n2651 & ~n17351 ;
  assign n31108 = n31107 ^ n7603 ^ 1'b0 ;
  assign n31109 = n31108 ^ n20202 ^ n15398 ;
  assign n31110 = n4132 | n13272 ;
  assign n31111 = n31110 ^ n31092 ^ n1210 ;
  assign n31112 = n560 & ~n10940 ;
  assign n31113 = n9130 & n31112 ;
  assign n31114 = n8069 | n15281 ;
  assign n31115 = n31114 ^ n18968 ^ 1'b0 ;
  assign n31116 = n13784 & ~n31115 ;
  assign n31117 = n9033 & n11252 ;
  assign n31118 = ~n6012 & n31117 ;
  assign n31119 = n1067 | n18119 ;
  assign n31120 = n5735 & n11426 ;
  assign n31121 = n21153 ^ n5178 ^ 1'b0 ;
  assign n31122 = n16581 & n18723 ;
  assign n31123 = n6589 & ~n30757 ;
  assign n31124 = n18468 & n31123 ;
  assign n31125 = n19654 & n31124 ;
  assign n31126 = n17232 | n31125 ;
  assign n31127 = n15300 & ~n31126 ;
  assign n31128 = n18479 ^ n14303 ^ n8886 ;
  assign n31129 = n31128 ^ n5701 ^ 1'b0 ;
  assign n31130 = ~n6255 & n31129 ;
  assign n31131 = n12680 | n21682 ;
  assign n31138 = n5641 & n13467 ;
  assign n31139 = ~n13467 & n31138 ;
  assign n31132 = n4366 | n18003 ;
  assign n31133 = ~n6314 & n31132 ;
  assign n31134 = ~n31132 & n31133 ;
  assign n31135 = n2492 | n18642 ;
  assign n31136 = n269 | n31135 ;
  assign n31137 = ~n31134 & n31136 ;
  assign n31140 = n31139 ^ n31137 ^ 1'b0 ;
  assign n31141 = n1843 & n5014 ;
  assign n31142 = ~n5014 & n31141 ;
  assign n31143 = n2513 & ~n31142 ;
  assign n31144 = n31142 & n31143 ;
  assign n31145 = n31144 ^ n13443 ^ 1'b0 ;
  assign n31146 = n31140 & n31145 ;
  assign n31147 = n2754 & n31146 ;
  assign n31148 = ~n31146 & n31147 ;
  assign n31149 = n30474 ^ n2339 ^ n296 ;
  assign n31150 = x13 & ~n2131 ;
  assign n31151 = ~n31149 & n31150 ;
  assign n31152 = ~n9068 & n12018 ;
  assign n31154 = n3804 | n26829 ;
  assign n31155 = n31154 ^ n16107 ^ 1'b0 ;
  assign n31153 = n13390 ^ n7876 ^ 1'b0 ;
  assign n31156 = n31155 ^ n31153 ^ 1'b0 ;
  assign n31157 = n26049 & ~n31156 ;
  assign n31158 = ~n2618 & n16933 ;
  assign n31159 = n10149 & n23391 ;
  assign n31160 = n15988 & n31159 ;
  assign n31161 = n20442 ^ n19512 ^ 1'b0 ;
  assign n31162 = ~n5793 & n5872 ;
  assign n31163 = n31162 ^ n16741 ^ 1'b0 ;
  assign n31164 = n14142 ^ n5661 ^ 1'b0 ;
  assign n31165 = n16980 | n31164 ;
  assign n31166 = ( ~n3212 & n3352 ) | ( ~n3212 & n31165 ) | ( n3352 & n31165 ) ;
  assign n31167 = ~n1023 & n6988 ;
  assign n31168 = n13510 & n31167 ;
  assign n31169 = n12699 & n31168 ;
  assign n31170 = n17473 ^ n1453 ^ 1'b0 ;
  assign n31171 = n13995 & ~n28689 ;
  assign n31172 = ~n4731 & n31171 ;
  assign n31173 = ~n25011 & n31172 ;
  assign n31174 = n4211 | n22497 ;
  assign n31175 = n24198 ^ n1777 ^ n531 ;
  assign n31176 = ~n14992 & n31175 ;
  assign n31177 = ( n11066 & ~n31174 ) | ( n11066 & n31176 ) | ( ~n31174 & n31176 ) ;
  assign n31178 = n19659 ^ n6080 ^ n1928 ;
  assign n31179 = n31178 ^ n26301 ^ n1926 ;
  assign n31180 = n7694 & n10757 ;
  assign n31181 = ~n7046 & n31180 ;
  assign n31182 = n31181 ^ n13990 ^ 1'b0 ;
  assign n31183 = n25140 ^ n19561 ^ 1'b0 ;
  assign n31184 = n17209 | n31183 ;
  assign n31185 = n22870 | n25542 ;
  assign n31186 = n14207 & n31185 ;
  assign n31187 = n20443 ^ n3073 ^ 1'b0 ;
  assign n31188 = ( n858 & n7767 ) | ( n858 & ~n31187 ) | ( n7767 & ~n31187 ) ;
  assign n31189 = n31188 ^ n16438 ^ 1'b0 ;
  assign n31190 = n31189 ^ n26334 ^ n18112 ;
  assign n31191 = n28588 ^ n12640 ^ 1'b0 ;
  assign n31192 = n25205 ^ n20889 ^ 1'b0 ;
  assign n31193 = n16460 & ~n22566 ;
  assign n31194 = ~n4259 & n31193 ;
  assign n31195 = n17146 | n31194 ;
  assign n31196 = n26177 ^ n25715 ^ 1'b0 ;
  assign n31197 = n20890 & ~n31196 ;
  assign n31198 = n3714 | n28552 ;
  assign n31199 = n31198 ^ n21170 ^ 1'b0 ;
  assign n31200 = n3041 & ~n28959 ;
  assign n31201 = n31200 ^ n23571 ^ 1'b0 ;
  assign n31202 = n29862 ^ n14922 ^ 1'b0 ;
  assign n31203 = ~n21846 & n31202 ;
  assign n31204 = ~n17414 & n31203 ;
  assign n31205 = n31201 & n31204 ;
  assign n31206 = n31205 ^ n25410 ^ 1'b0 ;
  assign n31207 = ~n11163 & n27926 ;
  assign n31208 = n31207 ^ n10576 ^ 1'b0 ;
  assign n31209 = n25798 ^ n8940 ^ 1'b0 ;
  assign n31210 = ( ~n4398 & n17264 ) | ( ~n4398 & n31209 ) | ( n17264 & n31209 ) ;
  assign n31211 = n2246 & ~n11066 ;
  assign n31212 = n13446 & n18779 ;
  assign n31213 = n7101 & n31212 ;
  assign n31214 = n19511 ^ n12145 ^ n4550 ;
  assign n31216 = n12248 ^ x229 ^ 1'b0 ;
  assign n31217 = n2512 | n31216 ;
  assign n31215 = n4127 & ~n11415 ;
  assign n31218 = n31217 ^ n31215 ^ n18203 ;
  assign n31219 = n15703 & n19105 ;
  assign n31220 = n3850 | n11070 ;
  assign n31221 = n14587 | n31220 ;
  assign n31222 = n31221 ^ n12874 ^ 1'b0 ;
  assign n31223 = n31219 & n31222 ;
  assign n31224 = n14286 ^ n2100 ^ 1'b0 ;
  assign n31226 = ~x161 & n15747 ;
  assign n31225 = ~n15699 & n16026 ;
  assign n31227 = n31226 ^ n31225 ^ n26848 ;
  assign n31228 = n21268 | n26560 ;
  assign n31229 = n17268 | n31228 ;
  assign n31230 = ~n17878 & n24669 ;
  assign n31231 = n20160 & ~n31230 ;
  assign n31232 = ~n23207 & n31231 ;
  assign n31233 = ~n4540 & n29754 ;
  assign n31234 = n12707 ^ n8381 ^ 1'b0 ;
  assign n31235 = n6364 | n31234 ;
  assign n31236 = ( n5326 & n6147 ) | ( n5326 & ~n30169 ) | ( n6147 & ~n30169 ) ;
  assign n31237 = n31236 ^ n4743 ^ 1'b0 ;
  assign n31238 = n3469 & n16761 ;
  assign n31239 = n10832 & ~n31238 ;
  assign n31240 = n10183 ^ n10051 ^ n3405 ;
  assign n31241 = n25944 & n31240 ;
  assign n31242 = n10284 & n21015 ;
  assign n31243 = ~n24183 & n31242 ;
  assign n31244 = n5944 ^ n5373 ^ 1'b0 ;
  assign n31245 = n31243 | n31244 ;
  assign n31246 = n29796 ^ n7091 ^ 1'b0 ;
  assign n31247 = n27940 & n31246 ;
  assign n31248 = ~n1719 & n29361 ;
  assign n31249 = n18014 & n31248 ;
  assign n31250 = n19860 ^ n6184 ^ 1'b0 ;
  assign n31251 = n31249 & n31250 ;
  assign n31252 = n31251 ^ n14250 ^ 1'b0 ;
  assign n31253 = n9329 | n31252 ;
  assign n31254 = n19078 ^ n5685 ^ 1'b0 ;
  assign n31259 = n14965 & n16199 ;
  assign n31255 = n20464 ^ n11160 ^ 1'b0 ;
  assign n31256 = n842 & n31255 ;
  assign n31257 = ~n10471 & n31256 ;
  assign n31258 = n31257 ^ n3316 ^ 1'b0 ;
  assign n31260 = n31259 ^ n31258 ^ 1'b0 ;
  assign n31261 = n12985 ^ n4276 ^ 1'b0 ;
  assign n31262 = n25450 ^ n4646 ^ 1'b0 ;
  assign n31263 = n31261 & ~n31262 ;
  assign n31264 = ( ~n13201 & n14212 ) | ( ~n13201 & n31263 ) | ( n14212 & n31263 ) ;
  assign n31265 = n1782 | n2732 ;
  assign n31266 = n18169 & ~n22328 ;
  assign n31268 = n9479 ^ n5832 ^ 1'b0 ;
  assign n31269 = n7068 & ~n31268 ;
  assign n31267 = ~n7776 & n10028 ;
  assign n31270 = n31269 ^ n31267 ^ 1'b0 ;
  assign n31271 = ~n26636 & n30856 ;
  assign n31272 = n31271 ^ n3300 ^ 1'b0 ;
  assign n31273 = ~n6082 & n29849 ;
  assign n31275 = ~n7245 & n17754 ;
  assign n31276 = ~n23592 & n31275 ;
  assign n31274 = n3038 | n10502 ;
  assign n31277 = n31276 ^ n31274 ^ 1'b0 ;
  assign n31278 = n14569 & n29174 ;
  assign n31279 = n22822 & n31278 ;
  assign n31280 = n31279 ^ n7393 ^ n1319 ;
  assign n31282 = n23732 ^ n16075 ^ n9296 ;
  assign n31281 = n8616 | n14178 ;
  assign n31283 = n31282 ^ n31281 ^ n17668 ;
  assign n31284 = n19389 & n31283 ;
  assign n31285 = n8517 | n13254 ;
  assign n31286 = n31285 ^ n11458 ^ 1'b0 ;
  assign n31287 = n4293 & n20448 ;
  assign n31288 = n6889 & n14254 ;
  assign n31289 = n533 & n31288 ;
  assign n31290 = ( n4153 & n4620 ) | ( n4153 & ~n31289 ) | ( n4620 & ~n31289 ) ;
  assign n31291 = ~n5354 & n31290 ;
  assign n31292 = n10917 ^ n9214 ^ x70 ;
  assign n31293 = ~n1615 & n14474 ;
  assign n31294 = n4903 & n31293 ;
  assign n31295 = n31294 ^ n21021 ^ 1'b0 ;
  assign n31296 = n21572 & ~n31295 ;
  assign n31297 = n2806 | n19654 ;
  assign n31298 = n31297 ^ n7021 ^ 1'b0 ;
  assign n31299 = n5115 | n12446 ;
  assign n31300 = ( n31296 & n31298 ) | ( n31296 & n31299 ) | ( n31298 & n31299 ) ;
  assign n31301 = n354 & n9331 ;
  assign n31302 = n27781 | n31301 ;
  assign n31303 = n31302 ^ n26601 ^ 1'b0 ;
  assign n31304 = n6438 | n14421 ;
  assign n31305 = n13184 & ~n31304 ;
  assign n31306 = n2726 | n31305 ;
  assign n31307 = n14078 ^ n7619 ^ n6102 ;
  assign n31308 = n3797 | n31307 ;
  assign n31312 = ~n20310 & n29593 ;
  assign n31309 = n11547 ^ n8805 ^ 1'b0 ;
  assign n31310 = n8893 & n31309 ;
  assign n31311 = n5317 & n31310 ;
  assign n31313 = n31312 ^ n31311 ^ 1'b0 ;
  assign n31314 = n16644 & ~n21964 ;
  assign n31315 = n5887 | n15634 ;
  assign n31316 = n31314 | n31315 ;
  assign n31317 = n7370 & n12368 ;
  assign n31318 = n31317 ^ n14848 ^ 1'b0 ;
  assign n31319 = n17689 & n30517 ;
  assign n31320 = n31319 ^ n19516 ^ n16464 ;
  assign n31321 = ~n16093 & n26675 ;
  assign n31322 = n12692 ^ n8487 ^ n7223 ;
  assign n31323 = n5890 ^ n3504 ^ 1'b0 ;
  assign n31324 = n31323 ^ n5072 ^ 1'b0 ;
  assign n31325 = ~n31322 & n31324 ;
  assign n31326 = n31325 ^ n970 ^ 1'b0 ;
  assign n31327 = n17692 & n31326 ;
  assign n31328 = n2815 | n3844 ;
  assign n31329 = n31328 ^ n1108 ^ 1'b0 ;
  assign n31330 = ~n6406 & n31329 ;
  assign n31331 = n4926 ^ n714 ^ 1'b0 ;
  assign n31332 = n2228 & n13408 ;
  assign n31333 = n17973 ^ n8961 ^ 1'b0 ;
  assign n31334 = n1532 | n31333 ;
  assign n31335 = n31334 ^ n2824 ^ 1'b0 ;
  assign n31336 = ~n31332 & n31335 ;
  assign n31337 = n5865 ^ n1027 ^ 1'b0 ;
  assign n31338 = n4373 | n26252 ;
  assign n31339 = n31337 | n31338 ;
  assign n31340 = n31339 ^ n13063 ^ 1'b0 ;
  assign n31341 = n5420 | n10392 ;
  assign n31342 = ~n5703 & n31341 ;
  assign n31343 = n18454 & ~n21980 ;
  assign n31344 = ~n31342 & n31343 ;
  assign n31345 = ( n1268 & n3523 ) | ( n1268 & ~n6468 ) | ( n3523 & ~n6468 ) ;
  assign n31346 = x36 & ~n604 ;
  assign n31347 = n18302 & n31346 ;
  assign n31348 = n31347 ^ n18465 ^ 1'b0 ;
  assign n31354 = n13835 ^ n4263 ^ 1'b0 ;
  assign n31352 = n15955 | n16161 ;
  assign n31353 = n31352 ^ n25897 ^ 1'b0 ;
  assign n31349 = n6604 ^ n1330 ^ 1'b0 ;
  assign n31350 = n22914 ^ n21548 ^ 1'b0 ;
  assign n31351 = n31349 | n31350 ;
  assign n31355 = n31354 ^ n31353 ^ n31351 ;
  assign n31356 = n5219 ^ x41 ^ 1'b0 ;
  assign n31357 = n10891 & n31356 ;
  assign n31358 = ( n6010 & n6627 ) | ( n6010 & ~n17704 ) | ( n6627 & ~n17704 ) ;
  assign n31359 = n31358 ^ n19393 ^ n3098 ;
  assign n31360 = n8667 | n15607 ;
  assign n31361 = n31360 ^ n5194 ^ 1'b0 ;
  assign n31362 = n19260 & n31361 ;
  assign n31363 = n269 & n3091 ;
  assign n31364 = n31363 ^ n9353 ^ 1'b0 ;
  assign n31365 = n18516 ^ n6403 ^ 1'b0 ;
  assign n31366 = n18665 | n31365 ;
  assign n31367 = n31364 | n31366 ;
  assign n31368 = n25189 ^ n5947 ^ 1'b0 ;
  assign n31369 = ( ~n4900 & n23693 ) | ( ~n4900 & n25661 ) | ( n23693 & n25661 ) ;
  assign n31370 = ~n3675 & n7083 ;
  assign n31371 = n13697 & n31370 ;
  assign n31372 = ~n2787 & n7318 ;
  assign n31373 = n22661 ^ n18643 ^ 1'b0 ;
  assign n31374 = n5599 & n31097 ;
  assign n31375 = n31374 ^ n19217 ^ 1'b0 ;
  assign n31376 = n1546 | n17364 ;
  assign n31377 = n31376 ^ n8303 ^ 1'b0 ;
  assign n31378 = n18047 | n21058 ;
  assign n31379 = n20633 ^ n14935 ^ 1'b0 ;
  assign n31380 = x174 & ~n2361 ;
  assign n31381 = n18163 & n31380 ;
  assign n31382 = n2958 & ~n31381 ;
  assign n31383 = n31382 ^ n23752 ^ 1'b0 ;
  assign n31384 = n17150 & ~n31383 ;
  assign n31385 = n23546 & n31384 ;
  assign n31386 = n22414 & ~n27819 ;
  assign n31389 = n22293 ^ n21835 ^ n17872 ;
  assign n31387 = n2850 ^ n2130 ^ 1'b0 ;
  assign n31388 = n24168 | n31387 ;
  assign n31390 = n31389 ^ n31388 ^ 1'b0 ;
  assign n31391 = n21528 ^ n2921 ^ 1'b0 ;
  assign n31392 = n5997 | n31391 ;
  assign n31393 = n17300 & n21836 ;
  assign n31394 = ~n10186 & n31393 ;
  assign n31395 = ~n5720 & n25830 ;
  assign n31396 = n8830 & n15930 ;
  assign n31397 = n31396 ^ n11577 ^ 1'b0 ;
  assign n31398 = n31397 ^ n9177 ^ n3115 ;
  assign n31399 = ( n913 & n9529 ) | ( n913 & ~n31398 ) | ( n9529 & ~n31398 ) ;
  assign n31400 = x7 & n16623 ;
  assign n31401 = n1665 & n31400 ;
  assign n31402 = n3058 & n3495 ;
  assign n31403 = n14675 ^ n10571 ^ n3453 ;
  assign n31404 = n4059 & n10455 ;
  assign n31405 = x45 & n31404 ;
  assign n31406 = ~n31403 & n31405 ;
  assign n31407 = ( n1521 & ~n5927 ) | ( n1521 & n10122 ) | ( ~n5927 & n10122 ) ;
  assign n31408 = n6798 & n31407 ;
  assign n31409 = n21017 & n31408 ;
  assign n31410 = n6869 & ~n8921 ;
  assign n31411 = n10321 & ~n20855 ;
  assign n31412 = n14476 & n31411 ;
  assign n31413 = n31412 ^ n3681 ^ 1'b0 ;
  assign n31417 = n7643 ^ n3550 ^ n1258 ;
  assign n31418 = n4207 & ~n5140 ;
  assign n31419 = ~n31417 & n31418 ;
  assign n31416 = n1033 | n5725 ;
  assign n31420 = n31419 ^ n31416 ^ 1'b0 ;
  assign n31414 = ( x155 & n606 ) | ( x155 & ~n7672 ) | ( n606 & ~n7672 ) ;
  assign n31415 = n14036 & n31414 ;
  assign n31421 = n31420 ^ n31415 ^ 1'b0 ;
  assign n31422 = n12601 & n31421 ;
  assign n31423 = ~n17296 & n31422 ;
  assign n31424 = ( n3477 & n5515 ) | ( n3477 & ~n27253 ) | ( n5515 & ~n27253 ) ;
  assign n31425 = n27783 ^ n12201 ^ 1'b0 ;
  assign n31426 = ~n8828 & n31425 ;
  assign n31427 = ( ~n385 & n5762 ) | ( ~n385 & n26166 ) | ( n5762 & n26166 ) ;
  assign n31428 = n5143 | n31427 ;
  assign n31429 = ~n17213 & n25263 ;
  assign n31430 = ~n26973 & n31429 ;
  assign n31432 = n10990 ^ n1548 ^ 1'b0 ;
  assign n31431 = n13757 & n22150 ;
  assign n31433 = n31432 ^ n31431 ^ 1'b0 ;
  assign n31434 = ~n11666 & n31433 ;
  assign n31435 = n19863 & ~n30147 ;
  assign n31436 = n3171 & ~n27634 ;
  assign n31437 = n17626 ^ n11719 ^ 1'b0 ;
  assign n31438 = n18425 ^ n9425 ^ 1'b0 ;
  assign n31439 = n451 & ~n813 ;
  assign n31440 = n31439 ^ n2595 ^ 1'b0 ;
  assign n31441 = n31440 ^ n25306 ^ n6731 ;
  assign n31444 = n22863 ^ n369 ^ 1'b0 ;
  assign n31442 = n4765 ^ n1987 ^ 1'b0 ;
  assign n31443 = ~n1339 & n31442 ;
  assign n31445 = n31444 ^ n31443 ^ n29631 ;
  assign n31446 = n21638 ^ n10122 ^ 1'b0 ;
  assign n31447 = ~n791 & n28250 ;
  assign n31448 = ~n13801 & n31447 ;
  assign n31449 = n31448 ^ n16352 ^ 1'b0 ;
  assign n31450 = n11553 & n18095 ;
  assign n31451 = ( n8998 & n13635 ) | ( n8998 & n17364 ) | ( n13635 & n17364 ) ;
  assign n31452 = n1630 & ~n31451 ;
  assign n31453 = ( n1233 & ~n1631 ) | ( n1233 & n13785 ) | ( ~n1631 & n13785 ) ;
  assign n31454 = n12051 | n31453 ;
  assign n31455 = n31454 ^ n11281 ^ 1'b0 ;
  assign n31456 = n16390 ^ n11974 ^ 1'b0 ;
  assign n31457 = n27788 & n31456 ;
  assign n31458 = n547 & n24836 ;
  assign n31459 = n14697 & n31458 ;
  assign n31460 = n15155 & n19298 ;
  assign n31461 = n2521 & n25009 ;
  assign n31462 = ~n29915 & n31461 ;
  assign n31463 = n5531 ^ x118 ^ 1'b0 ;
  assign n31464 = n31463 ^ n13758 ^ 1'b0 ;
  assign n31465 = n30501 & n31464 ;
  assign n31467 = ~n4742 & n13383 ;
  assign n31468 = ~n4862 & n31467 ;
  assign n31466 = n2223 & n7774 ;
  assign n31469 = n31468 ^ n31466 ^ 1'b0 ;
  assign n31470 = n31469 ^ n21733 ^ 1'b0 ;
  assign n31471 = ( n4636 & n8213 ) | ( n4636 & ~n23311 ) | ( n8213 & ~n23311 ) ;
  assign n31472 = n9853 ^ n9672 ^ 1'b0 ;
  assign n31473 = ( n21482 & ~n31471 ) | ( n21482 & n31472 ) | ( ~n31471 & n31472 ) ;
  assign n31474 = n16491 ^ n4815 ^ 1'b0 ;
  assign n31475 = n15614 | n31474 ;
  assign n31476 = n31475 ^ n963 ^ 1'b0 ;
  assign n31477 = n31476 ^ n2900 ^ 1'b0 ;
  assign n31478 = n13685 ^ n8906 ^ 1'b0 ;
  assign n31479 = n31478 ^ n30689 ^ 1'b0 ;
  assign n31480 = n2259 | n31479 ;
  assign n31481 = n10444 & n31480 ;
  assign n31482 = n31481 ^ x66 ^ 1'b0 ;
  assign n31483 = n21443 & n24882 ;
  assign n31484 = n31483 ^ n20920 ^ 1'b0 ;
  assign n31485 = n10947 & n16722 ;
  assign n31486 = n3246 | n12048 ;
  assign n31487 = n31485 | n31486 ;
  assign n31488 = n29464 ^ n12265 ^ 1'b0 ;
  assign n31489 = n31487 & ~n31488 ;
  assign n31490 = ~n3141 & n9457 ;
  assign n31491 = n995 & ~n31490 ;
  assign n31492 = n725 & ~n12611 ;
  assign n31493 = n31492 ^ n24136 ^ 1'b0 ;
  assign n31494 = n31493 ^ n9198 ^ 1'b0 ;
  assign n31495 = n5289 & ~n22429 ;
  assign n31496 = n14304 ^ n10218 ^ 1'b0 ;
  assign n31497 = n3638 & n31496 ;
  assign n31498 = ~n4889 & n31497 ;
  assign n31499 = ~n301 & n23687 ;
  assign n31500 = n27401 ^ n15105 ^ 1'b0 ;
  assign n31501 = ~n2239 & n4980 ;
  assign n31502 = n2239 & n31501 ;
  assign n31503 = ~n3778 & n31502 ;
  assign n31504 = ~n2195 & n3270 ;
  assign n31505 = ~n3270 & n31504 ;
  assign n31506 = n9483 | n31505 ;
  assign n31507 = n9316 | n31506 ;
  assign n31508 = n31507 ^ n733 ^ 1'b0 ;
  assign n31509 = n31503 | n31508 ;
  assign n31510 = n31503 & ~n31509 ;
  assign n31511 = n31510 ^ n16343 ^ n5855 ;
  assign n31512 = n892 | n30916 ;
  assign n31513 = n31512 ^ n18805 ^ 1'b0 ;
  assign n31514 = x172 & ~n14117 ;
  assign n31515 = n31514 ^ n23656 ^ 1'b0 ;
  assign n31516 = ~n3469 & n25888 ;
  assign n31518 = n6060 ^ n2219 ^ n1906 ;
  assign n31517 = n10639 ^ n5895 ^ x229 ;
  assign n31519 = n31518 ^ n31517 ^ 1'b0 ;
  assign n31520 = n31519 ^ n6241 ^ n5825 ;
  assign n31521 = n646 & n29187 ;
  assign n31522 = n29985 ^ n20124 ^ 1'b0 ;
  assign n31523 = n3598 & n31522 ;
  assign n31525 = n9686 & n17428 ;
  assign n31526 = ( n8965 & ~n13837 ) | ( n8965 & n31525 ) | ( ~n13837 & n31525 ) ;
  assign n31524 = n18290 & ~n19773 ;
  assign n31527 = n31526 ^ n31524 ^ 1'b0 ;
  assign n31528 = n10702 ^ n2077 ^ 1'b0 ;
  assign n31529 = n31528 ^ n31030 ^ 1'b0 ;
  assign n31530 = n26675 ^ n12956 ^ 1'b0 ;
  assign n31531 = n29413 & ~n31530 ;
  assign n31532 = n1103 | n4470 ;
  assign n31533 = x7 | n31532 ;
  assign n31534 = n903 & ~n7255 ;
  assign n31535 = ~n31533 & n31534 ;
  assign n31536 = ( ~n4456 & n5683 ) | ( ~n4456 & n31535 ) | ( n5683 & n31535 ) ;
  assign n31539 = n10182 | n20883 ;
  assign n31540 = n31539 ^ n7067 ^ 1'b0 ;
  assign n31537 = n19686 ^ n6705 ^ 1'b0 ;
  assign n31538 = n18528 & n31537 ;
  assign n31541 = n31540 ^ n31538 ^ 1'b0 ;
  assign n31542 = ~n20133 & n30130 ;
  assign n31543 = n4480 | n31542 ;
  assign n31544 = ( n8957 & n19776 ) | ( n8957 & ~n27814 ) | ( n19776 & ~n27814 ) ;
  assign n31545 = n10612 ^ n2095 ^ 1'b0 ;
  assign n31546 = n31544 | n31545 ;
  assign n31547 = ~n13846 & n24153 ;
  assign n31548 = n5968 ^ n915 ^ 1'b0 ;
  assign n31549 = n17929 ^ n4758 ^ 1'b0 ;
  assign n31550 = n31548 & ~n31549 ;
  assign n31551 = ( ~n5952 & n14396 ) | ( ~n5952 & n24129 ) | ( n14396 & n24129 ) ;
  assign n31552 = n16540 | n31551 ;
  assign n31553 = n3680 ^ x7 ^ 1'b0 ;
  assign n31554 = n4386 | n31553 ;
  assign n31555 = n3732 & ~n10422 ;
  assign n31557 = ( n9771 & n18805 ) | ( n9771 & ~n20030 ) | ( n18805 & ~n20030 ) ;
  assign n31558 = n22476 | n31557 ;
  assign n31559 = n18459 | n31558 ;
  assign n31560 = n31559 ^ n18683 ^ n2437 ;
  assign n31556 = n3817 & n13372 ;
  assign n31561 = n31560 ^ n31556 ^ 1'b0 ;
  assign n31562 = n10501 | n18600 ;
  assign n31563 = n13362 & n18164 ;
  assign n31564 = n9884 | n27215 ;
  assign n31565 = n27265 ^ n342 ^ 1'b0 ;
  assign n31566 = n6922 | n31565 ;
  assign n31567 = n7450 ^ n2368 ^ 1'b0 ;
  assign n31568 = n25558 & ~n29084 ;
  assign n31569 = ~n428 & n981 ;
  assign n31570 = n14229 ^ n13004 ^ 1'b0 ;
  assign n31571 = n20465 | n31570 ;
  assign n31572 = n3911 & ~n9520 ;
  assign n31573 = ~x138 & n1129 ;
  assign n31574 = ~n9895 & n31573 ;
  assign n31575 = n31574 ^ n13757 ^ n6856 ;
  assign n31576 = ~n6330 & n18452 ;
  assign n31577 = n8069 & n31576 ;
  assign n31578 = ~n9241 & n31577 ;
  assign n31579 = n6668 & n7271 ;
  assign n31580 = n31579 ^ n17967 ^ 1'b0 ;
  assign n31581 = n8235 & n9390 ;
  assign n31582 = n15555 ^ n14253 ^ 1'b0 ;
  assign n31583 = n31581 | n31582 ;
  assign n31584 = ~n423 & n28051 ;
  assign n31585 = n13501 ^ n5916 ^ n3620 ;
  assign n31586 = n31585 ^ n12393 ^ 1'b0 ;
  assign n31587 = ~n6126 & n25568 ;
  assign n31588 = n20591 & ~n23297 ;
  assign n31589 = n4375 | n31588 ;
  assign n31590 = n21116 ^ n19235 ^ 1'b0 ;
  assign n31591 = n19633 ^ n7411 ^ 1'b0 ;
  assign n31592 = n31591 ^ n2486 ^ x132 ;
  assign n31593 = n6153 | n25269 ;
  assign n31594 = ( n14300 & n27348 ) | ( n14300 & ~n31593 ) | ( n27348 & ~n31593 ) ;
  assign n31595 = ~n2935 & n3878 ;
  assign n31596 = n31595 ^ n23066 ^ 1'b0 ;
  assign n31597 = n26853 ^ n12614 ^ 1'b0 ;
  assign n31598 = n10293 & n14171 ;
  assign n31599 = ( n5835 & n9269 ) | ( n5835 & n22160 ) | ( n9269 & n22160 ) ;
  assign n31600 = n31599 ^ n24436 ^ n7264 ;
  assign n31601 = n3528 & ~n31600 ;
  assign n31602 = n16843 ^ n11376 ^ 1'b0 ;
  assign n31603 = ~n12406 & n13623 ;
  assign n31604 = n8929 | n31603 ;
  assign n31605 = n1886 | n31604 ;
  assign n31606 = n31605 ^ n5408 ^ 1'b0 ;
  assign n31607 = ~n7174 & n11699 ;
  assign n31608 = n31607 ^ n20443 ^ 1'b0 ;
  assign n31609 = ~n21515 & n31608 ;
  assign n31610 = n4312 | n6502 ;
  assign n31611 = n4326 | n31610 ;
  assign n31612 = ~n18973 & n31611 ;
  assign n31613 = n31612 ^ n26829 ^ 1'b0 ;
  assign n31614 = n12692 & ~n31613 ;
  assign n31615 = n11920 & ~n19748 ;
  assign n31616 = ~n10138 & n16501 ;
  assign n31617 = n16627 ^ n7954 ^ 1'b0 ;
  assign n31618 = ( ~n17748 & n23387 ) | ( ~n17748 & n31617 ) | ( n23387 & n31617 ) ;
  assign n31619 = n28589 ^ n6921 ^ 1'b0 ;
  assign n31620 = n20388 & n31619 ;
  assign n31621 = n22947 & ~n31511 ;
  assign n31628 = n22335 ^ n6730 ^ 1'b0 ;
  assign n31629 = n21869 & n31628 ;
  assign n31630 = n31629 ^ n19066 ^ 1'b0 ;
  assign n31622 = x71 & ~n5888 ;
  assign n31623 = n25990 ^ n6808 ^ 1'b0 ;
  assign n31624 = n10742 & n31623 ;
  assign n31625 = n31622 & n31624 ;
  assign n31626 = n31625 ^ n3126 ^ 1'b0 ;
  assign n31627 = n518 & ~n31626 ;
  assign n31631 = n31630 ^ n31627 ^ 1'b0 ;
  assign n31632 = n26099 ^ n19863 ^ n6341 ;
  assign n31633 = n25811 ^ n16087 ^ 1'b0 ;
  assign n31634 = n445 & n1880 ;
  assign n31635 = x136 & n31634 ;
  assign n31636 = n31635 ^ n3195 ^ 1'b0 ;
  assign n31637 = ( n24342 & n31633 ) | ( n24342 & ~n31636 ) | ( n31633 & ~n31636 ) ;
  assign n31638 = n13955 ^ n11694 ^ 1'b0 ;
  assign n31639 = n31638 ^ n24035 ^ 1'b0 ;
  assign n31640 = n4097 & n31639 ;
  assign n31641 = ~n1613 & n31640 ;
  assign n31642 = n6932 & n31641 ;
  assign n31643 = n16500 ^ n2264 ^ 1'b0 ;
  assign n31644 = n7831 | n31643 ;
  assign n31646 = ( n6784 & n15164 ) | ( n6784 & ~n29419 ) | ( n15164 & ~n29419 ) ;
  assign n31645 = n1246 & n8293 ;
  assign n31647 = n31646 ^ n31645 ^ n23349 ;
  assign n31648 = n6589 & ~n11219 ;
  assign n31649 = n31648 ^ n12319 ^ 1'b0 ;
  assign n31650 = n21953 & n31649 ;
  assign n31651 = ( ~x76 & n22273 ) | ( ~x76 & n31650 ) | ( n22273 & n31650 ) ;
  assign n31652 = n2302 ^ n1339 ^ 1'b0 ;
  assign n31653 = ~n8635 & n25730 ;
  assign n31654 = n13416 ^ n7708 ^ 1'b0 ;
  assign n31655 = n19863 & ~n31654 ;
  assign n31656 = n31655 ^ n29466 ^ n8001 ;
  assign n31657 = n31653 & n31656 ;
  assign n31658 = ~n3943 & n31657 ;
  assign n31659 = n15627 & n21750 ;
  assign n31660 = ~n9249 & n24320 ;
  assign n31661 = ~n2757 & n31660 ;
  assign n31662 = n1031 & n9330 ;
  assign n31663 = n31662 ^ n19131 ^ 1'b0 ;
  assign n31664 = ( n3716 & n11974 ) | ( n3716 & n14971 ) | ( n11974 & n14971 ) ;
  assign n31665 = ~n27071 & n30097 ;
  assign n31666 = n12749 & n14777 ;
  assign n31667 = n6798 & ~n11874 ;
  assign n31668 = n31667 ^ n8461 ^ 1'b0 ;
  assign n31669 = n31668 ^ n12368 ^ 1'b0 ;
  assign n31670 = n31669 ^ n4907 ^ 1'b0 ;
  assign n31671 = n1590 ^ n847 ^ 1'b0 ;
  assign n31672 = ( x254 & ~n11383 ) | ( x254 & n31671 ) | ( ~n11383 & n31671 ) ;
  assign n31673 = n27498 ^ n2519 ^ 1'b0 ;
  assign n31674 = n8888 & n11131 ;
  assign n31676 = n6889 | n27393 ;
  assign n31675 = n2190 | n7767 ;
  assign n31677 = n31676 ^ n31675 ^ 1'b0 ;
  assign n31678 = ~n612 & n18087 ;
  assign n31679 = n11384 | n27217 ;
  assign n31680 = n31679 ^ n20511 ^ 1'b0 ;
  assign n31681 = n24219 ^ n13245 ^ 1'b0 ;
  assign n31682 = n14775 & ~n19716 ;
  assign n31683 = ~n1506 & n31682 ;
  assign n31684 = ( n31676 & ~n31681 ) | ( n31676 & n31683 ) | ( ~n31681 & n31683 ) ;
  assign n31685 = n24899 & ~n26667 ;
  assign n31686 = x36 & n11072 ;
  assign n31687 = n7260 ^ n7106 ^ 1'b0 ;
  assign n31688 = n31686 & ~n31687 ;
  assign n31689 = n3254 ^ n3003 ^ 1'b0 ;
  assign n31690 = n31688 & ~n31689 ;
  assign n31691 = n3415 | n3424 ;
  assign n31694 = n11810 | n12943 ;
  assign n31692 = n3449 | n19325 ;
  assign n31693 = ~n14991 & n31692 ;
  assign n31695 = n31694 ^ n31693 ^ 1'b0 ;
  assign n31696 = n24447 ^ n15312 ^ 1'b0 ;
  assign n31697 = n1880 | n31696 ;
  assign n31698 = n1403 & n20509 ;
  assign n31699 = ~n9890 & n31698 ;
  assign n31700 = n8739 & ~n22832 ;
  assign n31701 = ( x138 & n31699 ) | ( x138 & ~n31700 ) | ( n31699 & ~n31700 ) ;
  assign n31702 = n2312 | n18252 ;
  assign n31703 = n31702 ^ n15045 ^ 1'b0 ;
  assign n31704 = n20407 ^ x146 ^ 1'b0 ;
  assign n31705 = n9844 ^ n1017 ^ 1'b0 ;
  assign n31706 = ( ~n6526 & n10522 ) | ( ~n6526 & n31705 ) | ( n10522 & n31705 ) ;
  assign n31707 = x81 | n20943 ;
  assign n31708 = n8485 | n28528 ;
  assign n31709 = n5573 | n25722 ;
  assign n31710 = n3316 & ~n31709 ;
  assign n31711 = n23401 & n31710 ;
  assign n31712 = n17333 & ~n31711 ;
  assign n31713 = n21702 ^ n6440 ^ n5799 ;
  assign n31714 = n31713 ^ n24836 ^ 1'b0 ;
  assign n31715 = ( n1062 & n22103 ) | ( n1062 & ~n28323 ) | ( n22103 & ~n28323 ) ;
  assign n31716 = n6720 & ~n22832 ;
  assign n31717 = n31716 ^ n24708 ^ 1'b0 ;
  assign n31718 = n17903 ^ n10532 ^ 1'b0 ;
  assign n31719 = n25989 & ~n31718 ;
  assign n31720 = n20056 ^ n15449 ^ 1'b0 ;
  assign n31721 = n6852 & n16239 ;
  assign n31722 = n6795 & n31721 ;
  assign n31723 = ( n28453 & ~n31720 ) | ( n28453 & n31722 ) | ( ~n31720 & n31722 ) ;
  assign n31724 = n8083 ^ n1289 ^ 1'b0 ;
  assign n31725 = n31724 ^ n11165 ^ 1'b0 ;
  assign n31726 = n5465 ^ n3465 ^ 1'b0 ;
  assign n31727 = n3013 | n31726 ;
  assign n31728 = n3666 | n4677 ;
  assign n31729 = n984 & ~n7888 ;
  assign n31730 = ( n6898 & n31728 ) | ( n6898 & ~n31729 ) | ( n31728 & ~n31729 ) ;
  assign n31731 = n30793 ^ n12015 ^ n11621 ;
  assign n31732 = n16507 | n17875 ;
  assign n31733 = n12087 ^ n7087 ^ 1'b0 ;
  assign n31734 = n4892 | n18945 ;
  assign n31735 = n26258 ^ n22434 ^ n6152 ;
  assign n31736 = n15653 ^ n6164 ^ 1'b0 ;
  assign n31742 = n29630 ^ n10168 ^ 1'b0 ;
  assign n31737 = ~n1418 & n25877 ;
  assign n31738 = n7879 | n31737 ;
  assign n31739 = n30809 | n31738 ;
  assign n31740 = n23900 & n31739 ;
  assign n31741 = ~n1587 & n31740 ;
  assign n31743 = n31742 ^ n31741 ^ 1'b0 ;
  assign n31744 = n16070 ^ x83 ^ 1'b0 ;
  assign n31745 = n31093 ^ n917 ^ 1'b0 ;
  assign n31746 = n24847 ^ n1685 ^ 1'b0 ;
  assign n31747 = n7578 | n12542 ;
  assign n31748 = ( n15990 & n20912 ) | ( n15990 & ~n31747 ) | ( n20912 & ~n31747 ) ;
  assign n31749 = n9456 & ~n27819 ;
  assign n31750 = n19521 & n26573 ;
  assign n31751 = n31750 ^ n31082 ^ 1'b0 ;
  assign n31752 = ( n3967 & n15028 ) | ( n3967 & ~n31751 ) | ( n15028 & ~n31751 ) ;
  assign n31753 = ( n1622 & ~n15193 ) | ( n1622 & n31752 ) | ( ~n15193 & n31752 ) ;
  assign n31754 = n31753 ^ n8214 ^ 1'b0 ;
  assign n31755 = n11808 | n31754 ;
  assign n31756 = n520 & n25425 ;
  assign n31757 = n28598 & n31756 ;
  assign n31758 = n7675 & n31757 ;
  assign n31759 = n14758 | n15957 ;
  assign n31760 = ~n3647 & n31759 ;
  assign n31761 = n10621 & n30189 ;
  assign n31762 = n21364 ^ n1250 ^ 1'b0 ;
  assign n31763 = n23532 ^ n10130 ^ 1'b0 ;
  assign n31764 = n15714 & ~n27647 ;
  assign n31765 = ~n11863 & n31764 ;
  assign n31769 = n3728 ^ n2556 ^ n1418 ;
  assign n31770 = n31769 ^ n2667 ^ 1'b0 ;
  assign n31771 = n5864 & ~n31770 ;
  assign n31766 = n9506 & ~n19135 ;
  assign n31767 = n31766 ^ n19030 ^ 1'b0 ;
  assign n31768 = n4418 & ~n31767 ;
  assign n31772 = n31771 ^ n31768 ^ 1'b0 ;
  assign n31775 = n3383 ^ n2678 ^ n749 ;
  assign n31773 = n6403 & n8780 ;
  assign n31774 = n4666 & ~n31773 ;
  assign n31776 = n31775 ^ n31774 ^ 1'b0 ;
  assign n31777 = n12562 ^ n4435 ^ 1'b0 ;
  assign n31778 = n15703 & ~n21017 ;
  assign n31779 = n31778 ^ n28959 ^ 1'b0 ;
  assign n31780 = ( n2517 & n8345 ) | ( n2517 & n15946 ) | ( n8345 & n15946 ) ;
  assign n31781 = n25105 ^ n18604 ^ n13203 ;
  assign n31782 = ( n1380 & n13511 ) | ( n1380 & ~n27533 ) | ( n13511 & ~n27533 ) ;
  assign n31783 = n31782 ^ n1168 ^ 1'b0 ;
  assign n31784 = n21071 ^ n2214 ^ 1'b0 ;
  assign n31785 = ~n31783 & n31784 ;
  assign n31786 = n11956 | n14891 ;
  assign n31787 = n28960 ^ n27665 ^ 1'b0 ;
  assign n31788 = n13945 & ~n18953 ;
  assign n31789 = n27833 ^ n9287 ^ n1486 ;
  assign n31790 = n31789 ^ n24645 ^ 1'b0 ;
  assign n31791 = n11945 | n15756 ;
  assign n31792 = n22658 & ~n31791 ;
  assign n31793 = n31792 ^ n14473 ^ 1'b0 ;
  assign n31794 = n5231 & ~n25403 ;
  assign n31795 = n19645 & n31794 ;
  assign n31796 = ~n15751 & n25233 ;
  assign n31797 = n31796 ^ n15030 ^ 1'b0 ;
  assign n31798 = ~n2431 & n7360 ;
  assign n31799 = ~n4038 & n31798 ;
  assign n31800 = ~n1093 & n10688 ;
  assign n31801 = n31800 ^ n2120 ^ 1'b0 ;
  assign n31802 = n5833 | n13656 ;
  assign n31803 = n5680 | n31802 ;
  assign n31804 = n3967 ^ n2259 ^ 1'b0 ;
  assign n31805 = ( n326 & ~n20957 ) | ( n326 & n27421 ) | ( ~n20957 & n27421 ) ;
  assign n31806 = n8602 | n15153 ;
  assign n31807 = n23474 | n31806 ;
  assign n31808 = ~n10513 & n19429 ;
  assign n31809 = n31808 ^ n6432 ^ 1'b0 ;
  assign n31810 = n15338 & ~n31809 ;
  assign n31811 = n17903 & n31810 ;
  assign n31812 = n13373 & ~n15550 ;
  assign n31813 = n31812 ^ n7584 ^ 1'b0 ;
  assign n31814 = ~n19444 & n31813 ;
  assign n31820 = n1553 & ~n18404 ;
  assign n31821 = n31820 ^ n2534 ^ 1'b0 ;
  assign n31822 = n31821 ^ n2257 ^ 1'b0 ;
  assign n31823 = ~n2483 & n31822 ;
  assign n31824 = n31823 ^ n17348 ^ 1'b0 ;
  assign n31825 = ~n14057 & n31824 ;
  assign n31815 = n16307 | n18156 ;
  assign n31816 = n6516 & ~n21867 ;
  assign n31817 = ~n16105 & n31816 ;
  assign n31818 = n6869 & ~n31817 ;
  assign n31819 = ~n31815 & n31818 ;
  assign n31826 = n31825 ^ n31819 ^ n9201 ;
  assign n31827 = n19940 ^ n12522 ^ 1'b0 ;
  assign n31828 = n1974 & ~n15561 ;
  assign n31829 = n17670 ^ n10850 ^ 1'b0 ;
  assign n31830 = n3845 & ~n28012 ;
  assign n31834 = ~n1323 & n4124 ;
  assign n31833 = n4722 & ~n13683 ;
  assign n31831 = n2131 | n10529 ;
  assign n31832 = n31831 ^ n10050 ^ 1'b0 ;
  assign n31835 = n31834 ^ n31833 ^ n31832 ;
  assign n31839 = n27052 ^ n5528 ^ 1'b0 ;
  assign n31840 = ~n8760 & n31839 ;
  assign n31836 = n3344 & ~n16004 ;
  assign n31837 = ~n3189 & n31836 ;
  assign n31838 = n31837 ^ n20325 ^ 1'b0 ;
  assign n31841 = n31840 ^ n31838 ^ n8039 ;
  assign n31842 = n8037 | n25140 ;
  assign n31843 = n11745 | n31842 ;
  assign n31844 = n21109 ^ n9811 ^ 1'b0 ;
  assign n31845 = n12460 & ~n15572 ;
  assign n31846 = n31845 ^ n29350 ^ n28663 ;
  assign n31847 = n29466 & ~n31846 ;
  assign n31848 = n31847 ^ n22785 ^ 1'b0 ;
  assign n31849 = ~n15418 & n21755 ;
  assign n31851 = n6193 ^ n835 ^ 1'b0 ;
  assign n31850 = ( ~n3362 & n8755 ) | ( ~n3362 & n29212 ) | ( n8755 & n29212 ) ;
  assign n31852 = n31851 ^ n31850 ^ 1'b0 ;
  assign n31853 = n9178 & n29052 ;
  assign n31854 = n31853 ^ n994 ^ 1'b0 ;
  assign n31855 = n31854 ^ n10824 ^ 1'b0 ;
  assign n31856 = n31476 & n31855 ;
  assign n31857 = n3431 | n20983 ;
  assign n31858 = n19432 & ~n31857 ;
  assign n31859 = n19457 & n31858 ;
  assign n31860 = ~n4767 & n14498 ;
  assign n31861 = ~n20019 & n31860 ;
  assign n31862 = n31861 ^ n10921 ^ 1'b0 ;
  assign n31863 = n26540 | n31862 ;
  assign n31864 = n1377 & ~n3343 ;
  assign n31865 = ~n1377 & n31864 ;
  assign n31866 = n8933 & ~n31865 ;
  assign n31867 = ~n2605 & n31866 ;
  assign n31868 = n18008 ^ n8993 ^ 1'b0 ;
  assign n31869 = n15919 ^ n2544 ^ 1'b0 ;
  assign n31870 = ~n8860 & n10855 ;
  assign n31871 = n31870 ^ n25099 ^ 1'b0 ;
  assign n31872 = n31869 & ~n31871 ;
  assign n31873 = n31872 ^ n1970 ^ 1'b0 ;
  assign n31874 = n11163 & ~n30918 ;
  assign n31875 = n31874 ^ n15790 ^ 1'b0 ;
  assign n31876 = n12899 ^ n7033 ^ 1'b0 ;
  assign n31877 = ~n18380 & n31876 ;
  assign n31878 = n16299 | n31877 ;
  assign n31879 = n16267 ^ n16087 ^ n7503 ;
  assign n31882 = n16305 ^ n6126 ^ n5376 ;
  assign n31880 = n5445 | n7869 ;
  assign n31881 = n31880 ^ n9026 ^ 1'b0 ;
  assign n31883 = n31882 ^ n31881 ^ 1'b0 ;
  assign n31884 = ~n18161 & n27324 ;
  assign n31885 = n6682 & n18699 ;
  assign n31886 = n31885 ^ n5050 ^ 1'b0 ;
  assign n31887 = n20960 & n26297 ;
  assign n31888 = n14976 & n31887 ;
  assign n31889 = ~n399 & n23043 ;
  assign n31890 = n10961 ^ n6400 ^ n2340 ;
  assign n31891 = ~n2827 & n31890 ;
  assign n31892 = n5162 ^ n3415 ^ n3103 ;
  assign n31893 = n31892 ^ n4773 ^ 1'b0 ;
  assign n31894 = n6914 & ~n25989 ;
  assign n31895 = n4222 & ~n22367 ;
  assign n31896 = n31895 ^ n15668 ^ 1'b0 ;
  assign n31897 = n17776 & n24526 ;
  assign n31898 = n3937 ^ n2504 ^ 1'b0 ;
  assign n31899 = n10737 & ~n31898 ;
  assign n31900 = n21015 & n31899 ;
  assign n31901 = n10143 ^ n4948 ^ n481 ;
  assign n31902 = n30225 ^ n2547 ^ 1'b0 ;
  assign n31903 = n9999 | n16704 ;
  assign n31904 = n16754 | n31903 ;
  assign n31905 = n31904 ^ n8086 ^ 1'b0 ;
  assign n31906 = n4821 | n26652 ;
  assign n31907 = n29651 & ~n31906 ;
  assign n31908 = n8999 & n14350 ;
  assign n31909 = n31908 ^ n5415 ^ 1'b0 ;
  assign n31910 = ~n7324 & n27807 ;
  assign n31911 = ~n10068 & n18058 ;
  assign n31912 = n31911 ^ n3624 ^ 1'b0 ;
  assign n31913 = n31910 | n31912 ;
  assign n31914 = n31913 ^ n9121 ^ 1'b0 ;
  assign n31915 = n14222 & ~n14790 ;
  assign n31916 = n31915 ^ n6236 ^ 1'b0 ;
  assign n31917 = n31914 & ~n31916 ;
  assign n31918 = n8627 | n13641 ;
  assign n31919 = n14587 & ~n31918 ;
  assign n31920 = ~n8381 & n31919 ;
  assign n31921 = n19742 | n20688 ;
  assign n31922 = n1164 & n31921 ;
  assign n31923 = n9167 ^ n1380 ^ n1003 ;
  assign n31924 = ~n31559 & n31923 ;
  assign n31926 = n21071 ^ x243 ^ 1'b0 ;
  assign n31925 = ~n16103 & n17497 ;
  assign n31927 = n31926 ^ n31925 ^ 1'b0 ;
  assign n31928 = n16291 & ~n31927 ;
  assign n31929 = n31928 ^ n9093 ^ 1'b0 ;
  assign n31930 = n7644 ^ n5499 ^ 1'b0 ;
  assign n31931 = ~n24341 & n31930 ;
  assign n31932 = ( ~n7910 & n30542 ) | ( ~n7910 & n31931 ) | ( n30542 & n31931 ) ;
  assign n31933 = n6970 & n24601 ;
  assign n31934 = n31933 ^ n13605 ^ 1'b0 ;
  assign n31935 = n10164 ^ n8187 ^ 1'b0 ;
  assign n31936 = ( ~n5019 & n8170 ) | ( ~n5019 & n13823 ) | ( n8170 & n13823 ) ;
  assign n31937 = n31936 ^ n3903 ^ 1'b0 ;
  assign n31938 = n31935 & n31937 ;
  assign n31939 = ~n7658 & n31938 ;
  assign n31940 = n31934 & ~n31939 ;
  assign n31941 = n31940 ^ n23240 ^ 1'b0 ;
  assign n31943 = ~n10192 & n21739 ;
  assign n31944 = n31943 ^ n27196 ^ 1'b0 ;
  assign n31942 = n16839 & ~n22237 ;
  assign n31945 = n31944 ^ n31942 ^ 1'b0 ;
  assign n31946 = n10935 ^ n2445 ^ 1'b0 ;
  assign n31947 = n31946 ^ n13043 ^ 1'b0 ;
  assign n31948 = n14548 & ~n29687 ;
  assign n31949 = n30357 ^ n12218 ^ n5355 ;
  assign n31950 = ~n31948 & n31949 ;
  assign n31951 = n31950 ^ n17247 ^ 1'b0 ;
  assign n31952 = n25722 ^ n563 ^ 1'b0 ;
  assign n31953 = n6964 & n31952 ;
  assign n31954 = n10536 & n31953 ;
  assign n31955 = n3588 & ~n6150 ;
  assign n31956 = n5019 & n31955 ;
  assign n31957 = n16283 ^ n13676 ^ 1'b0 ;
  assign n31958 = ~n31956 & n31957 ;
  assign n31959 = n4867 ^ n1380 ^ 1'b0 ;
  assign n31960 = n31958 & n31959 ;
  assign n31961 = n18461 ^ n8701 ^ 1'b0 ;
  assign n31966 = n12854 ^ x153 ^ 1'b0 ;
  assign n31967 = n15829 & n31966 ;
  assign n31968 = n31967 ^ n8270 ^ 1'b0 ;
  assign n31969 = n21536 | n31968 ;
  assign n31962 = ~n9811 & n22286 ;
  assign n31963 = n12959 & n31962 ;
  assign n31964 = n5372 & ~n31963 ;
  assign n31965 = n31964 ^ n17508 ^ 1'b0 ;
  assign n31970 = n31969 ^ n31965 ^ 1'b0 ;
  assign n31971 = n30089 ^ n12227 ^ 1'b0 ;
  assign n31972 = ~n11505 & n31971 ;
  assign n31973 = ( n14313 & ~n18415 ) | ( n14313 & n31972 ) | ( ~n18415 & n31972 ) ;
  assign n31974 = n4097 ^ n1380 ^ 1'b0 ;
  assign n31975 = ~n998 & n8443 ;
  assign n31976 = ~n9219 & n31975 ;
  assign n31977 = n31976 ^ n1476 ^ 1'b0 ;
  assign n31978 = n17152 & ~n31977 ;
  assign n31979 = ~n15409 & n31877 ;
  assign n31980 = ~n22809 & n31979 ;
  assign n31981 = ~n3624 & n21836 ;
  assign n31982 = n31981 ^ n13077 ^ 1'b0 ;
  assign n31983 = n31982 ^ n27354 ^ 1'b0 ;
  assign n31984 = n31983 ^ n1110 ^ 1'b0 ;
  assign n31985 = n20372 & ~n31984 ;
  assign n31986 = n16628 ^ n16391 ^ 1'b0 ;
  assign n31987 = n14354 | n31986 ;
  assign n31988 = n31987 ^ x214 ^ 1'b0 ;
  assign n31989 = ~n18759 & n31988 ;
  assign n31990 = n5230 & ~n11070 ;
  assign n31991 = n7199 ^ n6810 ^ 1'b0 ;
  assign n31993 = ~n535 & n4532 ;
  assign n31994 = n2712 & n31993 ;
  assign n31992 = n7405 & n17364 ;
  assign n31995 = n31994 ^ n31992 ^ 1'b0 ;
  assign n31996 = n31995 ^ n23161 ^ n16139 ;
  assign n31997 = ~n4789 & n27095 ;
  assign n31998 = n31997 ^ n9164 ^ n849 ;
  assign n31999 = n10066 & ~n31998 ;
  assign n32000 = n31999 ^ n16943 ^ n6322 ;
  assign n32001 = ~n11282 & n13516 ;
  assign n32002 = n7390 ^ n5859 ^ 1'b0 ;
  assign n32003 = n32001 | n32002 ;
  assign n32004 = n7695 ^ n5795 ^ 1'b0 ;
  assign n32005 = ~n3675 & n9844 ;
  assign n32006 = n26961 & n32005 ;
  assign n32007 = n22576 | n32006 ;
  assign n32008 = n32007 ^ n16292 ^ 1'b0 ;
  assign n32009 = n4226 & ~n18288 ;
  assign n32010 = n26616 & n32009 ;
  assign n32011 = ~n15774 & n27699 ;
  assign n32012 = n32011 ^ n4084 ^ 1'b0 ;
  assign n32013 = n32010 | n32012 ;
  assign n32014 = n32008 & ~n32013 ;
  assign n32015 = n13553 | n27635 ;
  assign n32016 = n32015 ^ n20622 ^ 1'b0 ;
  assign n32017 = n10749 | n10990 ;
  assign n32018 = n11316 | n32017 ;
  assign n32019 = ~n5986 & n7016 ;
  assign n32020 = n32019 ^ n24643 ^ 1'b0 ;
  assign n32021 = n32018 & ~n32020 ;
  assign n32022 = n24833 ^ n20624 ^ n11942 ;
  assign n32023 = n32022 ^ n13321 ^ 1'b0 ;
  assign n32024 = ( ~n29084 & n30417 ) | ( ~n29084 & n32023 ) | ( n30417 & n32023 ) ;
  assign n32025 = n5772 | n8899 ;
  assign n32026 = n7007 | n25343 ;
  assign n32027 = n32025 | n32026 ;
  assign n32028 = n32027 ^ n12113 ^ n3752 ;
  assign n32029 = n1524 | n22619 ;
  assign n32030 = n16709 ^ n6360 ^ 1'b0 ;
  assign n32031 = n6123 ^ n2484 ^ 1'b0 ;
  assign n32032 = ~n12268 & n32031 ;
  assign n32033 = ( n271 & n3692 ) | ( n271 & ~n32032 ) | ( n3692 & ~n32032 ) ;
  assign n32034 = n6221 | n11755 ;
  assign n32035 = n1543 & n13243 ;
  assign n32036 = n32035 ^ n30604 ^ 1'b0 ;
  assign n32037 = n32034 & n32036 ;
  assign n32038 = ~n3350 & n5477 ;
  assign n32039 = ~n3272 & n9987 ;
  assign n32040 = n15671 & n32039 ;
  assign n32041 = ~n32038 & n32040 ;
  assign n32042 = n29290 ^ n10111 ^ 1'b0 ;
  assign n32046 = n25913 ^ n2543 ^ 1'b0 ;
  assign n32047 = ( n1200 & n10093 ) | ( n1200 & ~n32046 ) | ( n10093 & ~n32046 ) ;
  assign n32048 = n18577 & n32047 ;
  assign n32049 = n32048 ^ n7293 ^ 1'b0 ;
  assign n32050 = ~n7399 & n13754 ;
  assign n32051 = ~n4729 & n32050 ;
  assign n32052 = n32049 & n32051 ;
  assign n32043 = n7675 ^ n3183 ^ 1'b0 ;
  assign n32044 = n3501 | n32043 ;
  assign n32045 = n32044 ^ n15200 ^ n9249 ;
  assign n32053 = n32052 ^ n32045 ^ 1'b0 ;
  assign n32054 = n5978 & n32053 ;
  assign n32055 = ~n8887 & n32054 ;
  assign n32056 = n29332 ^ n2763 ^ 1'b0 ;
  assign n32057 = n10444 ^ n9418 ^ 1'b0 ;
  assign n32058 = ( n2284 & n7093 ) | ( n2284 & n32057 ) | ( n7093 & n32057 ) ;
  assign n32059 = n24825 ^ n12762 ^ 1'b0 ;
  assign n32060 = n32058 | n32059 ;
  assign n32061 = n15834 & n32060 ;
  assign n32062 = n4123 | n6874 ;
  assign n32063 = n32062 ^ n2337 ^ 1'b0 ;
  assign n32064 = n18718 & ~n32063 ;
  assign n32065 = n2752 ^ n349 ^ 1'b0 ;
  assign n32066 = n5996 & n32065 ;
  assign n32067 = n10870 ^ n3597 ^ 1'b0 ;
  assign n32068 = n32066 & ~n32067 ;
  assign n32069 = n8544 ^ n1234 ^ 1'b0 ;
  assign n32070 = n2519 & n32069 ;
  assign n32071 = n27527 & n32070 ;
  assign n32072 = n15091 ^ n11908 ^ n10568 ;
  assign n32073 = n32072 ^ n16146 ^ 1'b0 ;
  assign n32074 = n5901 & n6683 ;
  assign n32075 = n32073 & n32074 ;
  assign n32076 = ~n16021 & n23560 ;
  assign n32077 = ~n905 & n32076 ;
  assign n32078 = ( ~n5780 & n6330 ) | ( ~n5780 & n22133 ) | ( n6330 & n22133 ) ;
  assign n32079 = n15307 ^ n10434 ^ n9670 ;
  assign n32080 = ~n26851 & n32079 ;
  assign n32081 = n32080 ^ n15609 ^ 1'b0 ;
  assign n32082 = n32081 ^ n3523 ^ 1'b0 ;
  assign n32083 = n25593 | n28480 ;
  assign n32084 = n3921 | n7881 ;
  assign n32085 = n32084 ^ n31061 ^ 1'b0 ;
  assign n32086 = n32085 ^ n22140 ^ 1'b0 ;
  assign n32087 = ~n12970 & n26035 ;
  assign n32088 = n21377 & n32087 ;
  assign n32089 = n17755 | n32088 ;
  assign n32090 = n12199 ^ n1795 ^ 1'b0 ;
  assign n32091 = ~n6649 & n29296 ;
  assign n32092 = n19887 ^ n8170 ^ n6409 ;
  assign n32093 = n6430 | n32092 ;
  assign n32094 = ~n5805 & n18042 ;
  assign n32095 = n18114 ^ n5677 ^ 1'b0 ;
  assign n32096 = n10631 | n32095 ;
  assign n32097 = n8809 & ~n32096 ;
  assign n32100 = n1916 ^ n1249 ^ n502 ;
  assign n32098 = n15034 ^ n3528 ^ 1'b0 ;
  assign n32099 = ~n7831 & n32098 ;
  assign n32101 = n32100 ^ n32099 ^ 1'b0 ;
  assign n32102 = ( n12162 & n26191 ) | ( n12162 & n29076 ) | ( n26191 & n29076 ) ;
  assign n32103 = n17599 & ~n32102 ;
  assign n32104 = n32103 ^ n10396 ^ n3438 ;
  assign n32105 = n32104 ^ n8362 ^ 1'b0 ;
  assign n32106 = n17257 & ~n32105 ;
  assign n32107 = n6235 ^ n735 ^ 1'b0 ;
  assign n32108 = n1099 | n32107 ;
  assign n32109 = n14639 ^ n1285 ^ 1'b0 ;
  assign n32110 = n32109 ^ n25487 ^ 1'b0 ;
  assign n32111 = ~n32108 & n32110 ;
  assign n32112 = ~n9835 & n32111 ;
  assign n32113 = n21316 ^ n17767 ^ n8938 ;
  assign n32114 = n14203 ^ n1995 ^ 1'b0 ;
  assign n32115 = n32113 & ~n32114 ;
  assign n32117 = n7880 ^ n4754 ^ n2913 ;
  assign n32116 = n11818 ^ n387 ^ 1'b0 ;
  assign n32118 = n32117 ^ n32116 ^ 1'b0 ;
  assign n32119 = n3734 & n32118 ;
  assign n32120 = n11934 & ~n12408 ;
  assign n32121 = n6327 & ~n10272 ;
  assign n32122 = n12554 ^ n10782 ^ 1'b0 ;
  assign n32123 = ~n1541 & n9215 ;
  assign n32124 = ~n4724 & n32123 ;
  assign n32125 = n32124 ^ n20822 ^ n4552 ;
  assign n32126 = n15902 & n32125 ;
  assign n32127 = n20058 & n32126 ;
  assign n32128 = ~n579 & n23400 ;
  assign n32129 = n32128 ^ n2915 ^ 1'b0 ;
  assign n32133 = n9221 & ~n11418 ;
  assign n32131 = ~n2732 & n21056 ;
  assign n32132 = ~n11425 & n32131 ;
  assign n32130 = n23049 ^ n8458 ^ 1'b0 ;
  assign n32134 = n32133 ^ n32132 ^ n32130 ;
  assign n32135 = ~x254 & n4787 ;
  assign n32136 = n32135 ^ n8493 ^ 1'b0 ;
  assign n32137 = ~n7785 & n32136 ;
  assign n32138 = n773 & n18586 ;
  assign n32139 = n32138 ^ n17845 ^ n11666 ;
  assign n32140 = n9819 & ~n10138 ;
  assign n32141 = n4026 & n32140 ;
  assign n32142 = n1323 | n32141 ;
  assign n32143 = n32142 ^ n7339 ^ 1'b0 ;
  assign n32144 = n6049 ^ n5568 ^ 1'b0 ;
  assign n32145 = x28 | n5844 ;
  assign n32146 = ( n6298 & ~n8112 ) | ( n6298 & n10571 ) | ( ~n8112 & n10571 ) ;
  assign n32147 = n11536 & ~n15502 ;
  assign n32148 = ( n3723 & n32146 ) | ( n3723 & ~n32147 ) | ( n32146 & ~n32147 ) ;
  assign n32149 = ~n7087 & n29249 ;
  assign n32150 = n32149 ^ x170 ^ 1'b0 ;
  assign n32151 = n32150 ^ n28698 ^ 1'b0 ;
  assign n32152 = ( ~n12282 & n13977 ) | ( ~n12282 & n15053 ) | ( n13977 & n15053 ) ;
  assign n32153 = n4193 & ~n12485 ;
  assign n32154 = n13612 & n32153 ;
  assign n32155 = n17046 & ~n32154 ;
  assign n32156 = n6363 & n21121 ;
  assign n32157 = n18857 & n32156 ;
  assign n32158 = n32157 ^ n2950 ^ 1'b0 ;
  assign n32159 = n16071 | n19056 ;
  assign n32160 = n32159 ^ n6010 ^ 1'b0 ;
  assign n32161 = ~n5588 & n32160 ;
  assign n32162 = n14429 | n32161 ;
  assign n32163 = n10261 ^ n5256 ^ 1'b0 ;
  assign n32164 = n29645 & ~n32163 ;
  assign n32165 = n5546 & n8236 ;
  assign n32166 = ~n32164 & n32165 ;
  assign n32167 = ~n7809 & n25108 ;
  assign n32168 = n21508 ^ n11710 ^ n1021 ;
  assign n32169 = x88 & n913 ;
  assign n32170 = ~n913 & n32169 ;
  assign n32171 = n5338 & ~n32170 ;
  assign n32172 = n32171 ^ n11210 ^ n2519 ;
  assign n32173 = ( ~n1155 & n23894 ) | ( ~n1155 & n25771 ) | ( n23894 & n25771 ) ;
  assign n32174 = n32172 | n32173 ;
  assign n32175 = n5274 & ~n6728 ;
  assign n32176 = ~n30945 & n32175 ;
  assign n32177 = n32176 ^ n22999 ^ 1'b0 ;
  assign n32178 = n32177 ^ n19447 ^ 1'b0 ;
  assign n32179 = n24078 ^ n2638 ^ 1'b0 ;
  assign n32180 = ~n7556 & n32179 ;
  assign n32181 = n9561 & n27807 ;
  assign n32182 = n2431 | n25018 ;
  assign n32183 = n13406 ^ n3093 ^ 1'b0 ;
  assign n32184 = ~n759 & n32183 ;
  assign n32185 = ( ~n1263 & n4436 ) | ( ~n1263 & n18205 ) | ( n4436 & n18205 ) ;
  assign n32186 = n32185 ^ n17884 ^ n2881 ;
  assign n32187 = ~n9960 & n29231 ;
  assign n32188 = n17830 & n32187 ;
  assign n32189 = n13904 ^ n1136 ^ 1'b0 ;
  assign n32190 = n32188 | n32189 ;
  assign n32191 = n14531 & ~n29834 ;
  assign n32192 = n32190 & n32191 ;
  assign n32193 = n32192 ^ n4172 ^ 1'b0 ;
  assign n32194 = n32186 & n32193 ;
  assign n32195 = n17456 ^ n11448 ^ 1'b0 ;
  assign n32196 = ~n4402 & n29886 ;
  assign n32197 = n32196 ^ n20166 ^ 1'b0 ;
  assign n32198 = n26127 | n32197 ;
  assign n32199 = n32198 ^ n24117 ^ 1'b0 ;
  assign n32200 = n8390 & n8478 ;
  assign n32202 = n5733 ^ n2960 ^ 1'b0 ;
  assign n32201 = n3706 & ~n14557 ;
  assign n32203 = n32202 ^ n32201 ^ 1'b0 ;
  assign n32204 = n27787 ^ n12485 ^ 1'b0 ;
  assign n32205 = n9121 & ~n21732 ;
  assign n32206 = n32205 ^ n20284 ^ 1'b0 ;
  assign n32207 = ~n13801 & n14571 ;
  assign n32208 = ~n4242 & n32207 ;
  assign n32209 = n353 | n32208 ;
  assign n32210 = n1483 & n32209 ;
  assign n32211 = n32210 ^ n2558 ^ 1'b0 ;
  assign n32212 = n32206 | n32211 ;
  assign n32213 = n20600 & ~n32212 ;
  assign n32214 = ( x169 & n25319 ) | ( x169 & ~n32213 ) | ( n25319 & ~n32213 ) ;
  assign n32215 = n19686 ^ n522 ^ 1'b0 ;
  assign n32216 = n16846 | n32215 ;
  assign n32220 = n9544 ^ n4463 ^ 1'b0 ;
  assign n32217 = n26308 ^ n6338 ^ 1'b0 ;
  assign n32218 = ~n17110 & n32217 ;
  assign n32219 = ~n2463 & n32218 ;
  assign n32221 = n32220 ^ n32219 ^ 1'b0 ;
  assign n32222 = n18876 & ~n32221 ;
  assign n32223 = n32216 & n32222 ;
  assign n32224 = n7593 | n11468 ;
  assign n32225 = n32224 ^ n21615 ^ 1'b0 ;
  assign n32226 = ~n8865 & n32225 ;
  assign n32227 = n32226 ^ n4294 ^ 1'b0 ;
  assign n32228 = n2278 & n11764 ;
  assign n32229 = n10155 & n32228 ;
  assign n32230 = n28305 & ~n32229 ;
  assign n32231 = n32230 ^ n3294 ^ 1'b0 ;
  assign n32232 = n22742 ^ n13462 ^ 1'b0 ;
  assign n32233 = n8809 & ~n32232 ;
  assign n32237 = n2518 & ~n4402 ;
  assign n32234 = n1166 & n18759 ;
  assign n32235 = ~n8577 & n32234 ;
  assign n32236 = ( n23579 & ~n28536 ) | ( n23579 & n32235 ) | ( ~n28536 & n32235 ) ;
  assign n32238 = n32237 ^ n32236 ^ 1'b0 ;
  assign n32241 = n28129 ^ n12876 ^ n5988 ;
  assign n32239 = ~n20463 & n23430 ;
  assign n32240 = ~n4757 & n32239 ;
  assign n32242 = n32241 ^ n32240 ^ n6128 ;
  assign n32243 = n2500 & n10530 ;
  assign n32244 = n20658 | n28101 ;
  assign n32245 = n10258 & n32244 ;
  assign n32246 = n7367 ^ n6279 ^ n2002 ;
  assign n32247 = n2320 & n3119 ;
  assign n32248 = n32247 ^ n23773 ^ n19604 ;
  assign n32249 = ~n572 & n3127 ;
  assign n32250 = n32249 ^ n15670 ^ n6683 ;
  assign n32251 = n19754 | n32250 ;
  assign n32252 = n32251 ^ n27170 ^ 1'b0 ;
  assign n32253 = n21140 ^ n8531 ^ n6811 ;
  assign n32254 = n32252 & n32253 ;
  assign n32255 = ~n16261 & n27605 ;
  assign n32256 = n18099 | n28426 ;
  assign n32257 = n13230 | n32256 ;
  assign n32258 = ~n3340 & n32257 ;
  assign n32259 = ~n2431 & n12429 ;
  assign n32260 = n10411 & n32259 ;
  assign n32261 = n32260 ^ n9343 ^ n9106 ;
  assign n32262 = n21851 ^ n12118 ^ 1'b0 ;
  assign n32263 = n15644 & n32262 ;
  assign n32264 = n32263 ^ n20335 ^ 1'b0 ;
  assign n32265 = n10258 | n32264 ;
  assign n32266 = n12942 ^ n4575 ^ 1'b0 ;
  assign n32267 = ~n29290 & n32266 ;
  assign n32269 = ~n7458 & n12640 ;
  assign n32270 = ~n3305 & n32269 ;
  assign n32268 = ~n15541 & n22486 ;
  assign n32271 = n32270 ^ n32268 ^ 1'b0 ;
  assign n32272 = ( n3929 & n5259 ) | ( n3929 & ~n16124 ) | ( n5259 & ~n16124 ) ;
  assign n32273 = n31603 ^ n31042 ^ 1'b0 ;
  assign n32274 = ( ~n438 & n15440 ) | ( ~n438 & n25806 ) | ( n15440 & n25806 ) ;
  assign n32275 = n9649 & ~n10416 ;
  assign n32276 = n32274 & n32275 ;
  assign n32277 = n10311 ^ n8488 ^ 1'b0 ;
  assign n32278 = ~n14261 & n32277 ;
  assign n32279 = ~n8315 & n8494 ;
  assign n32280 = n23203 ^ n2311 ^ n397 ;
  assign n32281 = ( x232 & n2924 ) | ( x232 & ~n32280 ) | ( n2924 & ~n32280 ) ;
  assign n32282 = n20879 & n32281 ;
  assign n32283 = ~n32279 & n32282 ;
  assign n32284 = n729 | n26115 ;
  assign n32285 = n13623 & ~n32284 ;
  assign n32286 = n24635 ^ n19639 ^ 1'b0 ;
  assign n32287 = n24374 ^ n17817 ^ n645 ;
  assign n32288 = n12193 ^ n11249 ^ 1'b0 ;
  assign n32289 = n8648 | n32288 ;
  assign n32290 = n15932 | n18388 ;
  assign n32291 = n32290 ^ n24318 ^ 1'b0 ;
  assign n32293 = n32108 ^ n2794 ^ 1'b0 ;
  assign n32292 = n14259 & ~n21234 ;
  assign n32294 = n32293 ^ n32292 ^ 1'b0 ;
  assign n32295 = n719 | n32294 ;
  assign n32296 = n20914 | n29245 ;
  assign n32297 = n14412 & ~n32296 ;
  assign n32298 = n8252 & ~n15117 ;
  assign n32299 = ~n22442 & n32298 ;
  assign n32300 = n20692 ^ n1703 ^ 1'b0 ;
  assign n32301 = n24833 ^ n11827 ^ n642 ;
  assign n32302 = n32301 ^ n30036 ^ n7097 ;
  assign n32303 = n14256 ^ n4510 ^ 1'b0 ;
  assign n32304 = ( ~n13004 & n20309 ) | ( ~n13004 & n32303 ) | ( n20309 & n32303 ) ;
  assign n32305 = n16510 ^ n14105 ^ 1'b0 ;
  assign n32306 = n7303 | n32305 ;
  assign n32307 = n32304 & ~n32306 ;
  assign n32308 = n12059 ^ n5653 ^ n3201 ;
  assign n32309 = n32308 ^ n15408 ^ 1'b0 ;
  assign n32310 = n11234 & n32309 ;
  assign n32311 = n18481 & n32310 ;
  assign n32312 = n13868 & n32311 ;
  assign n32313 = n4055 | n32312 ;
  assign n32314 = n14648 & ~n32313 ;
  assign n32315 = n11203 | n32314 ;
  assign n32316 = ~n2843 & n6177 ;
  assign n32317 = n32316 ^ n31341 ^ 1'b0 ;
  assign n32318 = n32317 ^ n9105 ^ 1'b0 ;
  assign n32319 = n11614 & n32318 ;
  assign n32320 = ( n1486 & ~n8229 ) | ( n1486 & n15302 ) | ( ~n8229 & n15302 ) ;
  assign n32321 = n32320 ^ n2024 ^ 1'b0 ;
  assign n32322 = n2329 & n16435 ;
  assign n32323 = n32322 ^ n9170 ^ 1'b0 ;
  assign n32324 = ~n21732 & n32323 ;
  assign n32325 = n9440 & ~n30124 ;
  assign n32326 = ( ~n7786 & n23305 ) | ( ~n7786 & n32325 ) | ( n23305 & n32325 ) ;
  assign n32329 = n7407 ^ n4208 ^ n3138 ;
  assign n32327 = n26091 ^ n6539 ^ 1'b0 ;
  assign n32328 = n26893 | n32327 ;
  assign n32330 = n32329 ^ n32328 ^ 1'b0 ;
  assign n32331 = n7321 & n17243 ;
  assign n32332 = n9280 & n32331 ;
  assign n32333 = n9482 & ~n32332 ;
  assign n32334 = n18003 & ~n26066 ;
  assign n32335 = n26112 ^ n2744 ^ 1'b0 ;
  assign n32336 = n15998 ^ n3193 ^ 1'b0 ;
  assign n32337 = n23924 ^ n5944 ^ x104 ;
  assign n32338 = n3791 ^ n1970 ^ 1'b0 ;
  assign n32339 = n30463 & ~n32338 ;
  assign n32340 = n32339 ^ n3814 ^ 1'b0 ;
  assign n32341 = ( n3912 & ~n7130 ) | ( n3912 & n22945 ) | ( ~n7130 & n22945 ) ;
  assign n32342 = n13988 | n32341 ;
  assign n32343 = n32342 ^ n10775 ^ 1'b0 ;
  assign n32344 = n27615 & ~n32343 ;
  assign n32345 = n17810 ^ n15408 ^ 1'b0 ;
  assign n32346 = n30349 & ~n32345 ;
  assign n32350 = ( ~n3825 & n4464 ) | ( ~n3825 & n10757 ) | ( n4464 & n10757 ) ;
  assign n32347 = n1281 & ~n4128 ;
  assign n32348 = n32347 ^ n2419 ^ 1'b0 ;
  assign n32349 = ~n8149 & n32348 ;
  assign n32351 = n32350 ^ n32349 ^ 1'b0 ;
  assign n32352 = n24847 ^ n14113 ^ 1'b0 ;
  assign n32353 = n32351 | n32352 ;
  assign n32354 = x155 | n10221 ;
  assign n32355 = ~n15168 & n32354 ;
  assign n32356 = n27852 ^ n12760 ^ 1'b0 ;
  assign n32357 = n24644 ^ n10066 ^ n1365 ;
  assign n32358 = n23164 ^ n14992 ^ 1'b0 ;
  assign n32359 = ~n12841 & n32358 ;
  assign n32360 = ~n29376 & n32359 ;
  assign n32361 = n31342 ^ n12608 ^ 1'b0 ;
  assign n32362 = n4694 & n15589 ;
  assign n32363 = ~n11134 & n32362 ;
  assign n32364 = n18140 & n32363 ;
  assign n32365 = n2946 ^ n2345 ^ 1'b0 ;
  assign n32366 = n32365 ^ n1253 ^ 1'b0 ;
  assign n32367 = n7358 & n9529 ;
  assign n32368 = n32367 ^ n29856 ^ 1'b0 ;
  assign n32369 = n23495 ^ n6149 ^ 1'b0 ;
  assign n32370 = n23763 & ~n32369 ;
  assign n32372 = ~n3498 & n4144 ;
  assign n32373 = n32372 ^ n4832 ^ 1'b0 ;
  assign n32371 = n15757 & n30689 ;
  assign n32374 = n32373 ^ n32371 ^ 1'b0 ;
  assign n32375 = n18099 ^ n12774 ^ 1'b0 ;
  assign n32376 = n21484 & n32375 ;
  assign n32377 = n20082 | n27296 ;
  assign n32378 = n9761 | n16563 ;
  assign n32379 = n32378 ^ n24833 ^ n2732 ;
  assign n32380 = n21051 ^ n11812 ^ 1'b0 ;
  assign n32381 = n1665 | n30490 ;
  assign n32382 = n10095 ^ n8619 ^ n747 ;
  assign n32383 = n7099 | n32382 ;
  assign n32384 = x173 & n24416 ;
  assign n32385 = n7930 ^ n5134 ^ 1'b0 ;
  assign n32386 = ~n32384 & n32385 ;
  assign n32388 = n3204 ^ n2313 ^ 1'b0 ;
  assign n32389 = n4417 & ~n32388 ;
  assign n32387 = n8445 | n12342 ;
  assign n32390 = n32389 ^ n32387 ^ 1'b0 ;
  assign n32391 = ~n3511 & n32390 ;
  assign n32393 = n29071 ^ n14357 ^ x22 ;
  assign n32392 = n3700 & n4031 ;
  assign n32394 = n32393 ^ n32392 ^ 1'b0 ;
  assign n32395 = n32391 & n32394 ;
  assign n32396 = n32395 ^ n11660 ^ n1293 ;
  assign n32397 = n985 | n6937 ;
  assign n32398 = n2804 & n32397 ;
  assign n32399 = n32398 ^ n11175 ^ n5735 ;
  assign n32400 = ~n15085 & n32399 ;
  assign n32401 = n2553 & n22593 ;
  assign n32402 = n19536 & ~n32401 ;
  assign n32403 = n994 & ~n16558 ;
  assign n32404 = ( n2481 & n21573 ) | ( n2481 & n32403 ) | ( n21573 & n32403 ) ;
  assign n32405 = n22999 ^ n16824 ^ n10593 ;
  assign n32406 = n10552 | n32405 ;
  assign n32407 = n5884 & ~n32406 ;
  assign n32408 = ( n5099 & ~n23229 ) | ( n5099 & n32407 ) | ( ~n23229 & n32407 ) ;
  assign n32409 = n3198 | n5433 ;
  assign n32410 = n20073 & ~n32409 ;
  assign n32411 = n2733 | n8287 ;
  assign n32413 = n1411 & n2294 ;
  assign n32412 = ~n5292 & n10017 ;
  assign n32414 = n32413 ^ n32412 ^ 1'b0 ;
  assign n32415 = n5839 & n32414 ;
  assign n32416 = n12199 ^ n5853 ^ 1'b0 ;
  assign n32417 = n19494 ^ n2459 ^ 1'b0 ;
  assign n32418 = ~n25455 & n32417 ;
  assign n32419 = n32418 ^ n9591 ^ n4902 ;
  assign n32421 = n17374 ^ n1155 ^ 1'b0 ;
  assign n32422 = ( n3371 & n5298 ) | ( n3371 & n32421 ) | ( n5298 & n32421 ) ;
  assign n32420 = ~n4073 & n15458 ;
  assign n32423 = n32422 ^ n32420 ^ 1'b0 ;
  assign n32424 = n10589 ^ n5583 ^ 1'b0 ;
  assign n32425 = n11087 | n32424 ;
  assign n32426 = ~n17827 & n27534 ;
  assign n32427 = n32426 ^ n32029 ^ 1'b0 ;
  assign n32428 = n9350 | n28847 ;
  assign n32429 = n4549 & ~n31095 ;
  assign n32431 = ~n329 & n5836 ;
  assign n32432 = ~n2302 & n32431 ;
  assign n32433 = n3095 | n32432 ;
  assign n32434 = n14218 & ~n32433 ;
  assign n32435 = n32434 ^ n23251 ^ 1'b0 ;
  assign n32436 = n8308 & ~n32435 ;
  assign n32430 = n24311 ^ n19126 ^ n18742 ;
  assign n32437 = n32436 ^ n32430 ^ 1'b0 ;
  assign n32438 = n8334 | n32057 ;
  assign n32439 = ~n27354 & n32438 ;
  assign n32440 = n25851 ^ n1129 ^ 1'b0 ;
  assign n32441 = n11204 & ~n32440 ;
  assign n32442 = n32441 ^ n21808 ^ 1'b0 ;
  assign n32443 = ~n3366 & n4059 ;
  assign n32444 = n11657 & n32443 ;
  assign n32445 = n9299 & n22081 ;
  assign n32446 = n13313 & ~n31913 ;
  assign n32447 = ~n32445 & n32446 ;
  assign n32448 = n22078 ^ n4558 ^ 1'b0 ;
  assign n32449 = ~n18009 & n28208 ;
  assign n32450 = n5218 & n32449 ;
  assign n32451 = n1666 | n21460 ;
  assign n32452 = ( ~n18205 & n25599 ) | ( ~n18205 & n32451 ) | ( n25599 & n32451 ) ;
  assign n32453 = n25996 ^ n1033 ^ 1'b0 ;
  assign n32454 = n3388 | n13943 ;
  assign n32455 = n32454 ^ n17219 ^ 1'b0 ;
  assign n32456 = n10842 | n32455 ;
  assign n32457 = n6359 & n8813 ;
  assign n32458 = n32457 ^ n15440 ^ 1'b0 ;
  assign n32459 = n32458 ^ n8686 ^ 1'b0 ;
  assign n32460 = n24614 | n32459 ;
  assign n32461 = n3325 & n16718 ;
  assign n32462 = n32461 ^ n6975 ^ 1'b0 ;
  assign n32463 = n9201 & ~n17322 ;
  assign n32464 = ~n32462 & n32463 ;
  assign n32465 = n2580 | n27222 ;
  assign n32466 = n32465 ^ n27508 ^ 1'b0 ;
  assign n32467 = ~x182 & n16060 ;
  assign n32468 = ~n3860 & n5954 ;
  assign n32469 = ( n12901 & ~n32467 ) | ( n12901 & n32468 ) | ( ~n32467 & n32468 ) ;
  assign n32470 = ~n15378 & n16251 ;
  assign n32471 = ~n18070 & n20522 ;
  assign n32472 = ~n13697 & n32471 ;
  assign n32474 = ~n8073 & n21151 ;
  assign n32473 = ~n9873 & n18657 ;
  assign n32475 = n32474 ^ n32473 ^ 1'b0 ;
  assign n32476 = ( n1546 & ~n8011 ) | ( n1546 & n23485 ) | ( ~n8011 & n23485 ) ;
  assign n32477 = n7521 | n19137 ;
  assign n32478 = n32477 ^ n20370 ^ 1'b0 ;
  assign n32479 = ~n32476 & n32478 ;
  assign n32480 = n3493 | n12044 ;
  assign n32481 = n32480 ^ n10882 ^ 1'b0 ;
  assign n32484 = ~n8324 & n9542 ;
  assign n32482 = n755 | n1279 ;
  assign n32483 = n25257 & n32482 ;
  assign n32485 = n32484 ^ n32483 ^ 1'b0 ;
  assign n32486 = n308 | n7629 ;
  assign n32487 = ( n6698 & ~n16429 ) | ( n6698 & n32486 ) | ( ~n16429 & n32486 ) ;
  assign n32488 = n2743 & ~n32487 ;
  assign n32489 = n2120 & n32488 ;
  assign n32490 = n8212 & ~n11014 ;
  assign n32491 = n16964 ^ n753 ^ 1'b0 ;
  assign n32492 = n32490 | n32491 ;
  assign n32493 = n16606 & ~n32492 ;
  assign n32494 = n25673 ^ n1321 ^ 1'b0 ;
  assign n32495 = n14262 & ~n32494 ;
  assign n32501 = ( n5010 & n18152 ) | ( n5010 & ~n21603 ) | ( n18152 & ~n21603 ) ;
  assign n32496 = ( n5223 & n13506 ) | ( n5223 & n20382 ) | ( n13506 & n20382 ) ;
  assign n32497 = x188 & n16629 ;
  assign n32498 = n32496 & n32497 ;
  assign n32499 = n32498 ^ n4031 ^ n3693 ;
  assign n32500 = n12827 & n32499 ;
  assign n32502 = n32501 ^ n32500 ^ 1'b0 ;
  assign n32503 = ( n3034 & n32495 ) | ( n3034 & ~n32502 ) | ( n32495 & ~n32502 ) ;
  assign n32504 = n7617 & ~n10534 ;
  assign n32505 = ~n8780 & n32504 ;
  assign n32507 = n30788 ^ n25229 ^ 1'b0 ;
  assign n32508 = n11927 & n32507 ;
  assign n32506 = ~n2509 & n4867 ;
  assign n32509 = n32508 ^ n32506 ^ 1'b0 ;
  assign n32510 = n32112 ^ n3382 ^ 1'b0 ;
  assign n32511 = n7325 & ~n32510 ;
  assign n32512 = n1493 | n8260 ;
  assign n32513 = n420 & ~n32512 ;
  assign n32514 = ( n952 & n6053 ) | ( n952 & n8098 ) | ( n6053 & n8098 ) ;
  assign n32515 = n7405 | n32514 ;
  assign n32516 = ( n579 & n3411 ) | ( n579 & n28160 ) | ( n3411 & n28160 ) ;
  assign n32518 = n9642 & ~n15746 ;
  assign n32517 = ~n1036 & n23087 ;
  assign n32519 = n32518 ^ n32517 ^ 1'b0 ;
  assign n32520 = n1362 & ~n32519 ;
  assign n32523 = x56 & ~n3013 ;
  assign n32524 = n32523 ^ n3010 ^ 1'b0 ;
  assign n32521 = ~n2810 & n21330 ;
  assign n32522 = n32521 ^ x111 ^ 1'b0 ;
  assign n32525 = n32524 ^ n32522 ^ n11908 ;
  assign n32526 = n10134 ^ n4553 ^ n2563 ;
  assign n32527 = n32525 & ~n32526 ;
  assign n32528 = n32527 ^ n10723 ^ 1'b0 ;
  assign n32529 = n20205 & ~n28094 ;
  assign n32530 = ~n279 & n22902 ;
  assign n32531 = n32530 ^ n5311 ^ 1'b0 ;
  assign n32532 = ~n5772 & n5895 ;
  assign n32534 = ( ~n2577 & n7146 ) | ( ~n2577 & n15049 ) | ( n7146 & n15049 ) ;
  assign n32533 = n28138 ^ n1571 ^ n531 ;
  assign n32535 = n32534 ^ n32533 ^ 1'b0 ;
  assign n32536 = n5388 | n19259 ;
  assign n32537 = n29210 & ~n32536 ;
  assign n32538 = n11976 & n22947 ;
  assign n32539 = n32538 ^ n7196 ^ 1'b0 ;
  assign n32540 = n14302 ^ n3812 ^ 1'b0 ;
  assign n32541 = n677 & n749 ;
  assign n32542 = n23232 & n32541 ;
  assign n32546 = ( n4957 & n13613 ) | ( n4957 & ~n26158 ) | ( n13613 & ~n26158 ) ;
  assign n32547 = ( n1499 & n8635 ) | ( n1499 & ~n18759 ) | ( n8635 & ~n18759 ) ;
  assign n32548 = n32547 ^ n15986 ^ 1'b0 ;
  assign n32549 = n32546 & n32548 ;
  assign n32543 = ~n7869 & n22072 ;
  assign n32544 = ~n7346 & n10675 ;
  assign n32545 = ~n32543 & n32544 ;
  assign n32550 = n32549 ^ n32545 ^ 1'b0 ;
  assign n32551 = n9273 & ~n32550 ;
  assign n32552 = n3773 & ~n16348 ;
  assign n32553 = ~n13048 & n24825 ;
  assign n32554 = n1975 & n2219 ;
  assign n32555 = n32554 ^ n20111 ^ 1'b0 ;
  assign n32556 = n32555 ^ n2100 ^ 1'b0 ;
  assign n32557 = n12244 & ~n29287 ;
  assign n32558 = n30543 ^ n12435 ^ 1'b0 ;
  assign n32559 = n21393 | n32558 ;
  assign n32560 = ~n734 & n11351 ;
  assign n32561 = n12313 & ~n18905 ;
  assign n32562 = n8829 & n18143 ;
  assign n32563 = n32562 ^ n20239 ^ 1'b0 ;
  assign n32564 = ( n10292 & n18050 ) | ( n10292 & ~n32563 ) | ( n18050 & ~n32563 ) ;
  assign n32565 = n32564 ^ n28802 ^ 1'b0 ;
  assign n32566 = n17311 ^ n11000 ^ n6888 ;
  assign n32568 = ~n13753 & n27558 ;
  assign n32569 = n32568 ^ n6362 ^ 1'b0 ;
  assign n32567 = n1813 | n5228 ;
  assign n32570 = n32569 ^ n32567 ^ 1'b0 ;
  assign n32571 = n8774 & n32570 ;
  assign n32572 = n32571 ^ n6516 ^ 1'b0 ;
  assign n32573 = n28979 ^ n22934 ^ 1'b0 ;
  assign n32574 = n9436 ^ n3362 ^ 1'b0 ;
  assign n32575 = n7437 | n28951 ;
  assign n32576 = n13715 & ~n32575 ;
  assign n32577 = n13332 | n32576 ;
  assign n32578 = n781 & ~n32577 ;
  assign n32579 = n20254 | n32578 ;
  assign n32580 = n10258 | n13477 ;
  assign n32581 = n32580 ^ n24066 ^ 1'b0 ;
  assign n32582 = ~n369 & n28874 ;
  assign n32583 = n3497 | n15095 ;
  assign n32584 = n32583 ^ n3326 ^ 1'b0 ;
  assign n32589 = n25697 ^ n11837 ^ 1'b0 ;
  assign n32585 = n32472 ^ n5680 ^ 1'b0 ;
  assign n32586 = n21214 & n32585 ;
  assign n32587 = ~n4026 & n32586 ;
  assign n32588 = n32587 ^ n10835 ^ 1'b0 ;
  assign n32590 = n32589 ^ n32588 ^ n31935 ;
  assign n32591 = n23297 ^ n8325 ^ 1'b0 ;
  assign n32592 = n26659 ^ x139 ^ 1'b0 ;
  assign n32593 = ~n14416 & n32592 ;
  assign n32594 = ( n4746 & ~n13338 ) | ( n4746 & n13921 ) | ( ~n13338 & n13921 ) ;
  assign n32595 = n32594 ^ n17127 ^ n1826 ;
  assign n32596 = n32595 ^ n20989 ^ 1'b0 ;
  assign n32597 = n6227 & n32596 ;
  assign n32598 = n13832 & n27402 ;
  assign n32599 = n6563 | n12660 ;
  assign n32600 = n28160 & ~n32599 ;
  assign n32601 = n7639 & ~n15075 ;
  assign n32602 = n13623 ^ n8239 ^ 1'b0 ;
  assign n32603 = n9871 & n32602 ;
  assign n32604 = ( n3204 & n10692 ) | ( n3204 & ~n25374 ) | ( n10692 & ~n25374 ) ;
  assign n32605 = ( ~n12692 & n25771 ) | ( ~n12692 & n32604 ) | ( n25771 & n32604 ) ;
  assign n32606 = n10338 & ~n21771 ;
  assign n32607 = n6766 & n10502 ;
  assign n32608 = n32607 ^ n20007 ^ 1'b0 ;
  assign n32610 = ( n7255 & n16644 ) | ( n7255 & ~n18098 ) | ( n16644 & ~n18098 ) ;
  assign n32609 = ~n1038 & n20829 ;
  assign n32611 = n32610 ^ n32609 ^ 1'b0 ;
  assign n32612 = ~n8293 & n32611 ;
  assign n32613 = n20112 ^ n13212 ^ 1'b0 ;
  assign n32614 = ( n1949 & n9175 ) | ( n1949 & ~n23732 ) | ( n9175 & ~n23732 ) ;
  assign n32615 = n28861 ^ n17780 ^ 1'b0 ;
  assign n32616 = n345 & n5511 ;
  assign n32617 = n32615 & n32616 ;
  assign n32618 = n6383 ^ n4560 ^ 1'b0 ;
  assign n32619 = n5419 & n32618 ;
  assign n32620 = n32619 ^ n8152 ^ 1'b0 ;
  assign n32621 = n27478 & ~n30034 ;
  assign n32622 = n32620 & n32621 ;
  assign n32623 = ~n5740 & n32622 ;
  assign n32624 = n6917 & ~n8009 ;
  assign n32628 = n22486 & ~n31622 ;
  assign n32625 = n1467 | n30192 ;
  assign n32626 = n32625 ^ n12101 ^ n2952 ;
  assign n32627 = n19992 & ~n32626 ;
  assign n32629 = n32628 ^ n32627 ^ 1'b0 ;
  assign n32630 = n7377 | n20429 ;
  assign n32631 = n4323 ^ n4024 ^ 1'b0 ;
  assign n32632 = n18386 & ~n32631 ;
  assign n32633 = ~n21411 & n32632 ;
  assign n32634 = n12952 ^ n7421 ^ n6334 ;
  assign n32635 = n32634 ^ n17146 ^ 1'b0 ;
  assign n32636 = n18406 & ~n23474 ;
  assign n32637 = n26876 ^ n21663 ^ 1'b0 ;
  assign n32638 = ~n770 & n32637 ;
  assign n32639 = x39 & ~n31927 ;
  assign n32640 = n32639 ^ n31845 ^ 1'b0 ;
  assign n32641 = n17772 & ~n19235 ;
  assign n32642 = n11268 & n31422 ;
  assign n32643 = n32642 ^ n7474 ^ n3894 ;
  assign n32644 = n11440 | n25456 ;
  assign n32645 = n2418 | n18313 ;
  assign n32646 = n32645 ^ x184 ^ 1'b0 ;
  assign n32647 = n909 & ~n32646 ;
  assign n32648 = n32647 ^ n13744 ^ 1'b0 ;
  assign n32649 = ~n1339 & n32648 ;
  assign n32650 = n2201 & n4542 ;
  assign n32651 = n2991 | n4895 ;
  assign n32652 = x248 & n11017 ;
  assign n32653 = n32652 ^ n19105 ^ 1'b0 ;
  assign n32654 = ( n1468 & ~n31715 ) | ( n1468 & n32653 ) | ( ~n31715 & n32653 ) ;
  assign n32655 = n15055 ^ n13356 ^ n8103 ;
  assign n32658 = ~n4528 & n9891 ;
  assign n32659 = ~n3447 & n32658 ;
  assign n32660 = ( n5473 & n9678 ) | ( n5473 & n32659 ) | ( n9678 & n32659 ) ;
  assign n32661 = n7928 & ~n32660 ;
  assign n32656 = n20214 ^ n16729 ^ n8855 ;
  assign n32657 = n1425 | n32656 ;
  assign n32662 = n32661 ^ n32657 ^ 1'b0 ;
  assign n32664 = n6411 | n15938 ;
  assign n32665 = n21878 ^ n5190 ^ 1'b0 ;
  assign n32666 = ~n32664 & n32665 ;
  assign n32663 = n4493 & n18754 ;
  assign n32667 = n32666 ^ n32663 ^ 1'b0 ;
  assign n32668 = n6119 | n7655 ;
  assign n32669 = n32668 ^ n14003 ^ 1'b0 ;
  assign n32670 = n32669 ^ n22207 ^ 1'b0 ;
  assign n32674 = ( ~n13419 & n16392 ) | ( ~n13419 & n26243 ) | ( n16392 & n26243 ) ;
  assign n32675 = n32674 ^ n20833 ^ n8823 ;
  assign n32671 = ( n2696 & ~n6529 ) | ( n2696 & n8451 ) | ( ~n6529 & n8451 ) ;
  assign n32672 = ( n2795 & n6516 ) | ( n2795 & ~n7632 ) | ( n6516 & ~n7632 ) ;
  assign n32673 = ~n32671 & n32672 ;
  assign n32676 = n32675 ^ n32673 ^ 1'b0 ;
  assign n32677 = n6867 | n16965 ;
  assign n32678 = n10133 ^ n1180 ^ 1'b0 ;
  assign n32679 = n32678 ^ n31407 ^ 1'b0 ;
  assign n32680 = n10166 & ~n32679 ;
  assign n32681 = x245 & n4339 ;
  assign n32682 = n32681 ^ n8120 ^ n3949 ;
  assign n32683 = ~n13925 & n32682 ;
  assign n32684 = n11298 ^ n7184 ^ 1'b0 ;
  assign n32685 = n10334 & ~n32684 ;
  assign n32686 = n12699 | n13327 ;
  assign n32687 = n2823 & ~n32686 ;
  assign n32688 = n21501 & n32687 ;
  assign n32689 = ~n8630 & n16485 ;
  assign n32690 = n17529 ^ n7602 ^ n407 ;
  assign n32691 = n23540 | n32690 ;
  assign n32692 = n32691 ^ n3369 ^ 1'b0 ;
  assign n32693 = ( n6121 & n10801 ) | ( n6121 & ~n32692 ) | ( n10801 & ~n32692 ) ;
  assign n32694 = n1969 | n4835 ;
  assign n32695 = ~n11849 & n20517 ;
  assign n32696 = n32695 ^ n27072 ^ n18083 ;
  assign n32697 = n10274 ^ n2353 ^ n994 ;
  assign n32698 = x87 & n10964 ;
  assign n32699 = ~n32697 & n32698 ;
  assign n32700 = n32699 ^ n6749 ^ 1'b0 ;
  assign n32701 = ~n32696 & n32700 ;
  assign n32702 = n15862 & n23902 ;
  assign n32703 = x101 & n32702 ;
  assign n32704 = n11872 ^ n5430 ^ 1'b0 ;
  assign n32705 = n8756 & ~n32704 ;
  assign n32706 = n8639 & ~n8914 ;
  assign n32707 = n32706 ^ n18935 ^ 1'b0 ;
  assign n32708 = n14667 | n32707 ;
  assign n32709 = n10051 | n32708 ;
  assign n32710 = n32705 & ~n32709 ;
  assign n32711 = ( n13746 & ~n19292 ) | ( n13746 & n31671 ) | ( ~n19292 & n31671 ) ;
  assign n32712 = n1746 & ~n10779 ;
  assign n32713 = n32712 ^ n25269 ^ 1'b0 ;
  assign n32714 = ~n23084 & n32713 ;
  assign n32715 = n32714 ^ n20251 ^ 1'b0 ;
  assign n32716 = ~n1688 & n32715 ;
  assign n32717 = ~n6563 & n7859 ;
  assign n32718 = n32717 ^ n3749 ^ 1'b0 ;
  assign n32719 = n32718 ^ n20152 ^ 1'b0 ;
  assign n32720 = ( n908 & n998 ) | ( n908 & n21000 ) | ( n998 & n21000 ) ;
  assign n32721 = ( n4358 & ~n4599 ) | ( n4358 & n9986 ) | ( ~n4599 & n9986 ) ;
  assign n32722 = n32721 ^ n10204 ^ n9820 ;
  assign n32723 = n27026 ^ n9213 ^ 1'b0 ;
  assign n32724 = n28157 ^ n1963 ^ 1'b0 ;
  assign n32725 = n24772 & ~n29714 ;
  assign n32726 = n29202 ^ n5783 ^ 1'b0 ;
  assign n32727 = ~n27365 & n29574 ;
  assign n32728 = n6197 ^ n1153 ^ 1'b0 ;
  assign n32729 = ~n1665 & n11112 ;
  assign n32730 = ~n26643 & n32729 ;
  assign n32731 = ( n9632 & n21229 ) | ( n9632 & ~n21252 ) | ( n21229 & ~n21252 ) ;
  assign n32732 = ( n3909 & ~n7973 ) | ( n3909 & n32731 ) | ( ~n7973 & n32731 ) ;
  assign n32733 = n2846 | n32732 ;
  assign n32734 = n18673 ^ n7888 ^ 1'b0 ;
  assign n32735 = ~n11718 & n32734 ;
  assign n32736 = n4478 & n32735 ;
  assign n32737 = ~n16709 & n18832 ;
  assign n32738 = n32737 ^ n1070 ^ 1'b0 ;
  assign n32739 = n8594 & ~n32738 ;
  assign n32740 = n32736 & n32739 ;
  assign n32741 = n13466 | n26869 ;
  assign n32742 = n18427 | n32741 ;
  assign n32743 = ~n3505 & n8586 ;
  assign n32744 = n13404 | n24204 ;
  assign n32745 = n32744 ^ n3683 ^ 1'b0 ;
  assign n32746 = n32745 ^ n24906 ^ n6274 ;
  assign n32747 = n3988 ^ n2514 ^ 1'b0 ;
  assign n32748 = n15233 ^ n3497 ^ 1'b0 ;
  assign n32749 = n16651 & ~n32748 ;
  assign n32750 = n32749 ^ n28643 ^ n9595 ;
  assign n32751 = n20684 ^ n11933 ^ n9331 ;
  assign n32752 = x64 | n17714 ;
  assign n32753 = n6114 & n32752 ;
  assign n32754 = n17187 & n32753 ;
  assign n32755 = n26405 ^ n681 ^ n553 ;
  assign n32756 = n32755 ^ n22878 ^ n15746 ;
  assign n32757 = ~n29324 & n32756 ;
  assign n32758 = n12815 & n29106 ;
  assign n32759 = n32758 ^ n9779 ^ 1'b0 ;
  assign n32760 = ~n5888 & n32759 ;
  assign n32761 = n3506 & n18600 ;
  assign n32762 = n32761 ^ n17766 ^ 1'b0 ;
  assign n32763 = n32762 ^ n9761 ^ 1'b0 ;
  assign n32764 = n5768 | n26373 ;
  assign n32765 = n19510 | n31259 ;
  assign n32766 = ~n26993 & n27111 ;
  assign n32767 = n32766 ^ n14046 ^ 1'b0 ;
  assign n32768 = ( n13803 & n20922 ) | ( n13803 & ~n28676 ) | ( n20922 & ~n28676 ) ;
  assign n32769 = ~n25501 & n32768 ;
  assign n32770 = n14368 & ~n20015 ;
  assign n32771 = n32770 ^ n2888 ^ 1'b0 ;
  assign n32772 = n5923 & ~n6034 ;
  assign n32773 = ( n10319 & ~n15950 ) | ( n10319 & n32772 ) | ( ~n15950 & n32772 ) ;
  assign n32774 = n14268 ^ x111 ^ 1'b0 ;
  assign n32775 = ( n1880 & ~n18181 ) | ( n1880 & n27819 ) | ( ~n18181 & n27819 ) ;
  assign n32776 = n13040 ^ n8931 ^ 1'b0 ;
  assign n32777 = n4628 & ~n20369 ;
  assign n32778 = ( n2034 & n19295 ) | ( n2034 & n32777 ) | ( n19295 & n32777 ) ;
  assign n32779 = n19627 ^ n5373 ^ 1'b0 ;
  assign n32780 = n6647 & n32779 ;
  assign n32781 = n25171 ^ n17049 ^ x201 ;
  assign n32782 = n311 & n32781 ;
  assign n32783 = n3918 & n18292 ;
  assign n32784 = ~n5872 & n32783 ;
  assign n32785 = n20453 ^ n14631 ^ 1'b0 ;
  assign n32786 = x46 & ~n27266 ;
  assign n32787 = n32786 ^ n7469 ^ 1'b0 ;
  assign n32788 = n15121 | n16343 ;
  assign n32789 = n32788 ^ n20232 ^ n8167 ;
  assign n32790 = n28669 ^ n3172 ^ 1'b0 ;
  assign n32791 = ~n10839 & n28885 ;
  assign n32792 = n11645 | n32791 ;
  assign n32793 = n32790 & ~n32792 ;
  assign n32794 = n7077 ^ n1876 ^ 1'b0 ;
  assign n32795 = n7804 & n32794 ;
  assign n32796 = n32795 ^ n4346 ^ 1'b0 ;
  assign n32797 = n516 | n780 ;
  assign n32798 = ~n605 & n16464 ;
  assign n32799 = ~n6585 & n32798 ;
  assign n32800 = n11351 & n32799 ;
  assign n32801 = n24796 ^ n2483 ^ 1'b0 ;
  assign n32802 = n32801 ^ n19269 ^ 1'b0 ;
  assign n32803 = n538 & ~n16094 ;
  assign n32805 = x212 & ~n12882 ;
  assign n32804 = ( n12347 & ~n19849 ) | ( n12347 & n24156 ) | ( ~n19849 & n24156 ) ;
  assign n32806 = n32805 ^ n32804 ^ n27932 ;
  assign n32807 = ~n4622 & n18114 ;
  assign n32808 = ~n22307 & n32807 ;
  assign n32809 = n32808 ^ n9978 ^ 1'b0 ;
  assign n32810 = ( n4828 & n24995 ) | ( n4828 & ~n32809 ) | ( n24995 & ~n32809 ) ;
  assign n32811 = ~n11869 & n24917 ;
  assign n32812 = n32811 ^ n5302 ^ 1'b0 ;
  assign n32813 = n31834 ^ n1489 ^ 1'b0 ;
  assign n32814 = x155 & ~n32813 ;
  assign n32815 = n32814 ^ n29744 ^ 1'b0 ;
  assign n32816 = n6655 | n22863 ;
  assign n32817 = n32816 ^ n1755 ^ 1'b0 ;
  assign n32818 = n18238 | n32817 ;
  assign n32819 = n10621 & n32818 ;
  assign n32820 = n1358 & n32819 ;
  assign n32821 = n3777 ^ n3617 ^ n3129 ;
  assign n32822 = n32821 ^ n24546 ^ n2165 ;
  assign n32823 = n4266 & n10522 ;
  assign n32824 = ~n18256 & n27951 ;
  assign n32825 = n30593 & ~n32758 ;
  assign n32826 = n32825 ^ n14465 ^ 1'b0 ;
  assign n32827 = ( ~n15230 & n32824 ) | ( ~n15230 & n32826 ) | ( n32824 & n32826 ) ;
  assign n32828 = ~n21487 & n27860 ;
  assign n32829 = n9840 & n32828 ;
  assign n32830 = n23865 & ~n23940 ;
  assign n32833 = ( ~n12723 & n19178 ) | ( ~n12723 & n26614 ) | ( n19178 & n26614 ) ;
  assign n32831 = n5916 ^ n4657 ^ 1'b0 ;
  assign n32832 = n23857 | n32831 ;
  assign n32834 = n32833 ^ n32832 ^ n6122 ;
  assign n32835 = ~n2337 & n5758 ;
  assign n32836 = n19587 ^ n11314 ^ 1'b0 ;
  assign n32837 = n32835 & ~n32836 ;
  assign n32838 = ~n19185 & n20030 ;
  assign n32839 = n32837 & ~n32838 ;
  assign n32840 = n10198 & ~n15111 ;
  assign n32841 = n32840 ^ n23005 ^ 1'b0 ;
  assign n32842 = n22142 ^ n9069 ^ n2896 ;
  assign n32843 = n23887 & n32842 ;
  assign n32844 = n400 & ~n19880 ;
  assign n32845 = n2332 | n15181 ;
  assign n32846 = n32845 ^ n27946 ^ n7267 ;
  assign n32847 = n5802 & n32451 ;
  assign n32848 = n5544 & n32847 ;
  assign n32849 = ~n5129 & n7621 ;
  assign n32850 = n11284 & ~n32849 ;
  assign n32851 = n2749 & ~n11064 ;
  assign n32852 = n32851 ^ n7593 ^ 1'b0 ;
  assign n32853 = n12018 | n15026 ;
  assign n32854 = n1987 | n32853 ;
  assign n32855 = n17936 ^ n3504 ^ 1'b0 ;
  assign n32856 = ~n15629 & n32855 ;
  assign n32857 = n7443 & n29721 ;
  assign n32858 = n4498 & n32857 ;
  assign n32859 = n25927 ^ n19116 ^ 1'b0 ;
  assign n32860 = ~n32858 & n32859 ;
  assign n32861 = n11449 & n32860 ;
  assign n32862 = ~n25994 & n32861 ;
  assign n32863 = ~n23966 & n32862 ;
  assign n32864 = n7404 & n12379 ;
  assign n32866 = n4473 | n13823 ;
  assign n32865 = n10490 | n18534 ;
  assign n32867 = n32866 ^ n32865 ^ 1'b0 ;
  assign n32868 = n21392 & n23970 ;
  assign n32869 = n32868 ^ n26323 ^ 1'b0 ;
  assign n32870 = n23463 ^ n9551 ^ 1'b0 ;
  assign n32871 = n6093 & n32870 ;
  assign n32872 = n32871 ^ x38 ^ 1'b0 ;
  assign n32873 = ~n718 & n26594 ;
  assign n32874 = ~n32872 & n32873 ;
  assign n32875 = ( n3322 & n3374 ) | ( n3322 & n3474 ) | ( n3374 & n3474 ) ;
  assign n32876 = n22909 & n32875 ;
  assign n32877 = ~n4418 & n32876 ;
  assign n32878 = n9865 & ~n32877 ;
  assign n32879 = n32878 ^ n28296 ^ 1'b0 ;
  assign n32880 = n32874 | n32879 ;
  assign n32881 = ( n8375 & n9447 ) | ( n8375 & n31249 ) | ( n9447 & n31249 ) ;
  assign n32882 = n32881 ^ n9937 ^ 1'b0 ;
  assign n32883 = n1618 ^ x125 ^ 1'b0 ;
  assign n32884 = n1272 | n4592 ;
  assign n32885 = n32883 | n32884 ;
  assign n32886 = ~n7745 & n13575 ;
  assign n32888 = n11706 ^ n8415 ^ 1'b0 ;
  assign n32889 = ~n1274 & n32888 ;
  assign n32887 = n7795 | n13687 ;
  assign n32890 = n32889 ^ n32887 ^ 1'b0 ;
  assign n32891 = n4207 & n8520 ;
  assign n32892 = n12781 & n32891 ;
  assign n32893 = ( n4689 & n14000 ) | ( n4689 & n27706 ) | ( n14000 & n27706 ) ;
  assign n32894 = n27296 | n32893 ;
  assign n32895 = n18335 ^ n16925 ^ 1'b0 ;
  assign n32896 = n19138 & ~n32895 ;
  assign n32897 = ~n5033 & n5296 ;
  assign n32898 = n1113 & ~n2289 ;
  assign n32899 = ~n25056 & n32898 ;
  assign n32900 = n32899 ^ n14817 ^ x200 ;
  assign n32901 = n5975 & ~n17091 ;
  assign n32902 = ~n4615 & n15205 ;
  assign n32903 = n2504 & n32902 ;
  assign n32904 = x155 & ~n32903 ;
  assign n32905 = n32904 ^ n1394 ^ 1'b0 ;
  assign n32906 = n27551 & n32905 ;
  assign n32907 = n17523 & n32906 ;
  assign n32908 = n14776 | n24498 ;
  assign n32909 = n20159 | n32908 ;
  assign n32910 = ~n7378 & n11353 ;
  assign n32911 = ( n3415 & n7221 ) | ( n3415 & n32910 ) | ( n7221 & n32910 ) ;
  assign n32912 = n14550 & n25576 ;
  assign n32913 = n32912 ^ n5800 ^ 1'b0 ;
  assign n32914 = n19494 ^ n8220 ^ 1'b0 ;
  assign n32915 = n13789 | n32914 ;
  assign n32916 = ~n19832 & n23810 ;
  assign n32917 = ~n2759 & n5227 ;
  assign n32918 = ~n13707 & n32917 ;
  assign n32919 = n11135 & n20388 ;
  assign n32920 = n32919 ^ n6415 ^ 1'b0 ;
  assign n32921 = n1327 & ~n19511 ;
  assign n32922 = n1674 & n32921 ;
  assign n32923 = n7696 & ~n32922 ;
  assign n32924 = n2502 & n32923 ;
  assign n32925 = ( n3465 & ~n5279 ) | ( n3465 & n5976 ) | ( ~n5279 & n5976 ) ;
  assign n32926 = n16346 ^ n15455 ^ 1'b0 ;
  assign n32927 = n32925 & ~n32926 ;
  assign n32928 = n32924 | n32927 ;
  assign n32929 = ( ~n1166 & n3972 ) | ( ~n1166 & n18399 ) | ( n3972 & n18399 ) ;
  assign n32930 = ~n5768 & n32929 ;
  assign n32931 = n18534 ^ n2981 ^ 1'b0 ;
  assign n32932 = n1494 | n2524 ;
  assign n32933 = n19591 & ~n32932 ;
  assign n32934 = n31471 | n32933 ;
  assign n32935 = n15555 & ~n24647 ;
  assign n32936 = n9175 ^ n4068 ^ 1'b0 ;
  assign n32937 = n20293 & n32936 ;
  assign n32938 = n32937 ^ n7004 ^ 1'b0 ;
  assign n32939 = n1036 & n9661 ;
  assign n32940 = n32939 ^ n1697 ^ 1'b0 ;
  assign n32941 = n3336 & n12408 ;
  assign n32942 = n32941 ^ n2661 ^ 1'b0 ;
  assign n32943 = ~n6357 & n13007 ;
  assign n32944 = n32943 ^ n30032 ^ 1'b0 ;
  assign n32945 = ~n9952 & n15258 ;
  assign n32946 = n20980 & ~n32945 ;
  assign n32947 = ( ~n5446 & n13400 ) | ( ~n5446 & n32946 ) | ( n13400 & n32946 ) ;
  assign n32948 = n10567 & n27736 ;
  assign n32949 = n22666 ^ n3783 ^ n768 ;
  assign n32950 = n32949 ^ n5043 ^ 1'b0 ;
  assign n32951 = n19704 ^ n16575 ^ 1'b0 ;
  assign n32952 = n12938 & n32951 ;
  assign n32953 = ~n4672 & n17689 ;
  assign n32954 = n32953 ^ n19799 ^ n2821 ;
  assign n32955 = n8029 | n11349 ;
  assign n32956 = n3505 & ~n10534 ;
  assign n32957 = n32956 ^ n5843 ^ 1'b0 ;
  assign n32958 = ~n4630 & n11080 ;
  assign n32959 = n32958 ^ n612 ^ 1'b0 ;
  assign n32960 = n13897 ^ n12887 ^ 1'b0 ;
  assign n32961 = n32959 & n32960 ;
  assign n32962 = ( n6645 & n32957 ) | ( n6645 & ~n32961 ) | ( n32957 & ~n32961 ) ;
  assign n32963 = n32962 ^ n12503 ^ n6388 ;
  assign n32964 = ( n8901 & ~n16180 ) | ( n8901 & n18161 ) | ( ~n16180 & n18161 ) ;
  assign n32965 = ~n6363 & n20438 ;
  assign n32966 = n2991 & ~n6309 ;
  assign n32967 = n18183 & n32966 ;
  assign n32968 = n32967 ^ n22516 ^ 1'b0 ;
  assign n32969 = n24663 ^ n8029 ^ 1'b0 ;
  assign n32970 = n32968 & n32969 ;
  assign n32971 = ~n1036 & n15473 ;
  assign n32972 = ~n20013 & n32971 ;
  assign n32974 = n13676 ^ n895 ^ 1'b0 ;
  assign n32975 = n790 & ~n32974 ;
  assign n32973 = n972 | n16996 ;
  assign n32976 = n32975 ^ n32973 ^ 1'b0 ;
  assign n32978 = n18431 ^ n4153 ^ 1'b0 ;
  assign n32979 = n16605 & ~n32978 ;
  assign n32980 = n17882 & n32979 ;
  assign n32981 = n32980 ^ n14086 ^ 1'b0 ;
  assign n32977 = n7570 & n26086 ;
  assign n32982 = n32981 ^ n32977 ^ 1'b0 ;
  assign n32983 = n26906 ^ n25615 ^ n24681 ;
  assign n32984 = n1046 & n8752 ;
  assign n32985 = n20279 & n32984 ;
  assign n32986 = n9287 | n32985 ;
  assign n32987 = ~n3430 & n21053 ;
  assign n32988 = n23016 ^ n12802 ^ 1'b0 ;
  assign n32989 = n17420 & n32988 ;
  assign n32990 = n4600 & n12683 ;
  assign n32991 = n32990 ^ n5366 ^ 1'b0 ;
  assign n32992 = ~n2814 & n15423 ;
  assign n32993 = n22928 ^ n1093 ^ 1'b0 ;
  assign n32994 = n17150 & ~n21941 ;
  assign n32995 = n8052 ^ n559 ^ 1'b0 ;
  assign n32996 = n22787 & ~n32995 ;
  assign n32997 = n10830 & n32996 ;
  assign n32998 = n21988 ^ n9897 ^ 1'b0 ;
  assign n32999 = n27145 ^ n20192 ^ 1'b0 ;
  assign n33000 = n32096 ^ n18214 ^ n3505 ;
  assign n33001 = n17650 & n21572 ;
  assign n33002 = n33000 & n33001 ;
  assign n33003 = ~n13372 & n25238 ;
  assign n33004 = n33003 ^ n5549 ^ 1'b0 ;
  assign n33005 = n25705 ^ n24242 ^ 1'b0 ;
  assign n33006 = n6151 & n6242 ;
  assign n33007 = n2577 & n33006 ;
  assign n33008 = n911 & ~n8453 ;
  assign n33009 = ~n11153 & n33008 ;
  assign n33010 = n33007 | n33009 ;
  assign n33013 = n9583 & ~n16465 ;
  assign n33012 = n19501 ^ n12865 ^ 1'b0 ;
  assign n33011 = n4119 & n7901 ;
  assign n33014 = n33013 ^ n33012 ^ n33011 ;
  assign n33015 = n18410 ^ n650 ^ 1'b0 ;
  assign n33016 = n8882 & n33015 ;
  assign n33017 = ( n1506 & ~n12134 ) | ( n1506 & n33016 ) | ( ~n12134 & n33016 ) ;
  assign n33018 = ~n10692 & n20273 ;
  assign n33019 = n33018 ^ n1022 ^ 1'b0 ;
  assign n33020 = n15993 & ~n22293 ;
  assign n33021 = n24500 ^ n14571 ^ n9123 ;
  assign n33022 = ( n1049 & n19866 ) | ( n1049 & ~n27040 ) | ( n19866 & ~n27040 ) ;
  assign n33023 = ~n3124 & n3196 ;
  assign n33024 = n33023 ^ n3709 ^ 1'b0 ;
  assign n33025 = n2810 & n26646 ;
  assign n33026 = n33025 ^ n23815 ^ 1'b0 ;
  assign n33027 = n20301 | n33026 ;
  assign n33028 = n20887 ^ n6196 ^ 1'b0 ;
  assign n33029 = n13017 | n33028 ;
  assign n33030 = n13183 & n17025 ;
  assign n33031 = n33029 & n33030 ;
  assign n33032 = n12025 ^ n11201 ^ 1'b0 ;
  assign n33033 = n20061 | n33032 ;
  assign n33034 = n11048 & ~n33033 ;
  assign n33035 = n29787 & ~n33034 ;
  assign n33036 = n3922 & n33035 ;
  assign n33037 = ( n1892 & n28724 ) | ( n1892 & n32177 ) | ( n28724 & n32177 ) ;
  assign n33039 = n11866 ^ n7255 ^ 1'b0 ;
  assign n33040 = ~n11646 & n33039 ;
  assign n33041 = n33040 ^ n1850 ^ 1'b0 ;
  assign n33038 = n32247 ^ n30899 ^ n1254 ;
  assign n33042 = n33041 ^ n33038 ^ n26779 ;
  assign n33043 = n22836 & n24914 ;
  assign n33044 = ~n21121 & n33043 ;
  assign n33045 = n10206 & ~n33044 ;
  assign n33046 = ~n19793 & n33045 ;
  assign n33047 = n978 & n28757 ;
  assign n33048 = n6895 ^ n1360 ^ 1'b0 ;
  assign n33049 = n27207 ^ n16709 ^ 1'b0 ;
  assign n33050 = n33048 & n33049 ;
  assign n33051 = n4063 & ~n12083 ;
  assign n33052 = n33051 ^ n28140 ^ n24191 ;
  assign n33053 = ~n1433 & n11073 ;
  assign n33058 = ~n4518 & n6161 ;
  assign n33059 = ~n10004 & n33058 ;
  assign n33054 = ~n5181 & n10825 ;
  assign n33055 = n25317 ^ n9769 ^ 1'b0 ;
  assign n33056 = ( n1435 & ~n19905 ) | ( n1435 & n33055 ) | ( ~n19905 & n33055 ) ;
  assign n33057 = ~n33054 & n33056 ;
  assign n33060 = n33059 ^ n33057 ^ 1'b0 ;
  assign n33061 = n14989 ^ n2279 ^ 1'b0 ;
  assign n33062 = n25219 | n33061 ;
  assign n33063 = n16916 & ~n33062 ;
  assign n33064 = n33063 ^ n27967 ^ 1'b0 ;
  assign n33065 = n24441 ^ n15126 ^ n14862 ;
  assign n33066 = n405 & n18889 ;
  assign n33067 = n29937 & n33066 ;
  assign n33068 = n33065 | n33067 ;
  assign n33069 = n29937 ^ n26846 ^ 1'b0 ;
  assign n33070 = n32837 ^ n30516 ^ 1'b0 ;
  assign n33073 = ( ~n6572 & n7321 ) | ( ~n6572 & n23506 ) | ( n7321 & n23506 ) ;
  assign n33072 = n32641 ^ n5267 ^ n1870 ;
  assign n33071 = ( n365 & n6766 ) | ( n365 & ~n7087 ) | ( n6766 & ~n7087 ) ;
  assign n33074 = n33073 ^ n33072 ^ n33071 ;
  assign n33075 = n33074 ^ n27270 ^ n15095 ;
  assign n33076 = n17809 ^ n9343 ^ n1884 ;
  assign n33077 = n33076 ^ n11505 ^ 1'b0 ;
  assign n33078 = n3048 | n4446 ;
  assign n33079 = n33078 ^ n3108 ^ 1'b0 ;
  assign n33080 = ( n11951 & n27319 ) | ( n11951 & n33079 ) | ( n27319 & n33079 ) ;
  assign n33081 = ~n6136 & n28083 ;
  assign n33082 = ~n8977 & n33081 ;
  assign n33083 = n33082 ^ n3405 ^ 1'b0 ;
  assign n33084 = ~n5731 & n33083 ;
  assign n33085 = n33084 ^ n16324 ^ 1'b0 ;
  assign n33086 = ( n30656 & ~n33080 ) | ( n30656 & n33085 ) | ( ~n33080 & n33085 ) ;
  assign n33087 = n19821 ^ n6574 ^ 1'b0 ;
  assign n33088 = ( n7056 & n16524 ) | ( n7056 & n33087 ) | ( n16524 & n33087 ) ;
  assign n33089 = n12273 ^ n3712 ^ 1'b0 ;
  assign n33090 = n12494 ^ n4192 ^ 1'b0 ;
  assign n33091 = ~n21550 & n33090 ;
  assign n33092 = n33091 ^ n29158 ^ 1'b0 ;
  assign n33093 = n7804 & ~n29100 ;
  assign n33094 = n6607 & n33093 ;
  assign n33095 = n1393 & ~n6064 ;
  assign n33096 = n33095 ^ n4029 ^ 1'b0 ;
  assign n33097 = n10771 ^ n7160 ^ 1'b0 ;
  assign n33098 = n20753 | n33097 ;
  assign n33099 = n4578 | n15074 ;
  assign n33100 = n13530 | n33099 ;
  assign n33101 = n33100 ^ n9295 ^ n3848 ;
  assign n33102 = n574 & n5208 ;
  assign n33103 = n21057 ^ x41 ^ 1'b0 ;
  assign n33104 = n8405 ^ n6409 ^ 1'b0 ;
  assign n33109 = ~n6844 & n33012 ;
  assign n33110 = n8554 & ~n33109 ;
  assign n33111 = n33110 ^ n2561 ^ 1'b0 ;
  assign n33105 = ~n4246 & n6930 ;
  assign n33106 = n18380 & n33105 ;
  assign n33107 = ~n19694 & n33106 ;
  assign n33108 = n23430 & n33107 ;
  assign n33112 = n33111 ^ n33108 ^ 1'b0 ;
  assign n33113 = n2055 | n16118 ;
  assign n33114 = n33113 ^ n31019 ^ 1'b0 ;
  assign n33115 = n20823 ^ n5295 ^ 1'b0 ;
  assign n33116 = ( n15930 & n20197 ) | ( n15930 & n33115 ) | ( n20197 & n33115 ) ;
  assign n33117 = n18055 & n33116 ;
  assign n33118 = n33117 ^ n28458 ^ 1'b0 ;
  assign n33119 = n15601 ^ n14071 ^ 1'b0 ;
  assign n33120 = n26441 ^ n7452 ^ 1'b0 ;
  assign n33121 = n33119 | n33120 ;
  assign n33123 = ( ~n1255 & n7293 ) | ( ~n1255 & n19019 ) | ( n7293 & n19019 ) ;
  assign n33122 = n11458 & ~n11941 ;
  assign n33124 = n33123 ^ n33122 ^ 1'b0 ;
  assign n33125 = n20447 & n23685 ;
  assign n33126 = ~n1228 & n8088 ;
  assign n33127 = n2701 & n12021 ;
  assign n33128 = n33127 ^ n16103 ^ 1'b0 ;
  assign n33129 = n28395 ^ n8585 ^ 1'b0 ;
  assign n33130 = n4117 & ~n27663 ;
  assign n33133 = n6594 & n14631 ;
  assign n33134 = n29381 & n33133 ;
  assign n33131 = n24192 ^ n18413 ^ 1'b0 ;
  assign n33132 = n8716 & n33131 ;
  assign n33135 = n33134 ^ n33132 ^ 1'b0 ;
  assign n33136 = n32862 ^ n17866 ^ 1'b0 ;
  assign n33137 = n33136 ^ n12551 ^ 1'b0 ;
  assign n33138 = ( n1106 & n10336 ) | ( n1106 & n17822 ) | ( n10336 & n17822 ) ;
  assign n33139 = n33138 ^ n22361 ^ 1'b0 ;
  assign n33140 = n32104 ^ n15040 ^ 1'b0 ;
  assign n33141 = n17875 ^ n11109 ^ 1'b0 ;
  assign n33142 = n24001 ^ n1655 ^ 1'b0 ;
  assign n33143 = ~n12923 & n33142 ;
  assign n33144 = ( n4415 & ~n7157 ) | ( n4415 & n33143 ) | ( ~n7157 & n33143 ) ;
  assign n33145 = n2203 | n33144 ;
  assign n33146 = n33141 & ~n33145 ;
  assign n33147 = ~n6779 & n15387 ;
  assign n33148 = n33147 ^ n2399 ^ 1'b0 ;
  assign n33149 = n3301 ^ n1010 ^ x248 ;
  assign n33150 = ( n16024 & ~n33148 ) | ( n16024 & n33149 ) | ( ~n33148 & n33149 ) ;
  assign n33151 = n13542 ^ x130 ^ 1'b0 ;
  assign n33152 = ~n13603 & n22134 ;
  assign n33153 = n15941 & n26834 ;
  assign n33154 = n10699 ^ n3641 ^ 1'b0 ;
  assign n33155 = ( n14272 & n16555 ) | ( n14272 & ~n32569 ) | ( n16555 & ~n32569 ) ;
  assign n33156 = n3273 & n5947 ;
  assign n33157 = ( ~n8325 & n17055 ) | ( ~n8325 & n33156 ) | ( n17055 & n33156 ) ;
  assign n33158 = n7053 ^ n5054 ^ 1'b0 ;
  assign n33159 = n12802 & ~n33158 ;
  assign n33160 = ~n8672 & n33159 ;
  assign n33161 = n26821 ^ n4547 ^ 1'b0 ;
  assign n33162 = n8356 & n33161 ;
  assign n33163 = n5124 & ~n14482 ;
  assign n33164 = n29120 ^ n16681 ^ 1'b0 ;
  assign n33165 = ~n33163 & n33164 ;
  assign n33166 = ( n25900 & n33162 ) | ( n25900 & ~n33165 ) | ( n33162 & ~n33165 ) ;
  assign n33167 = n9319 & ~n23341 ;
  assign n33168 = n15247 | n25650 ;
  assign n33169 = n7756 & ~n33168 ;
  assign n33170 = n33169 ^ n5061 ^ 1'b0 ;
  assign n33171 = ~n32671 & n33170 ;
  assign n33172 = n16558 ^ n2225 ^ 1'b0 ;
  assign n33173 = n29042 ^ n6986 ^ 1'b0 ;
  assign n33174 = ~n20285 & n33173 ;
  assign n33179 = n14843 ^ n2849 ^ 1'b0 ;
  assign n33175 = n7273 & n17339 ;
  assign n33176 = n16510 & n33175 ;
  assign n33177 = n11932 & n33176 ;
  assign n33178 = n33177 ^ n19887 ^ n2026 ;
  assign n33180 = n33179 ^ n33178 ^ n27056 ;
  assign n33184 = n10726 ^ n7341 ^ 1'b0 ;
  assign n33181 = n6869 ^ n2416 ^ 1'b0 ;
  assign n33182 = n11511 | n33181 ;
  assign n33183 = n12843 | n33182 ;
  assign n33185 = n33184 ^ n33183 ^ n23401 ;
  assign n33186 = n11024 & n23390 ;
  assign n33187 = n2434 ^ n723 ^ 1'b0 ;
  assign n33188 = ~n5997 & n33187 ;
  assign n33189 = ~n33186 & n33188 ;
  assign n33190 = n1097 & n4723 ;
  assign n33191 = n33190 ^ n16330 ^ 1'b0 ;
  assign n33192 = ~n16929 & n18176 ;
  assign n33193 = n33192 ^ n6971 ^ 1'b0 ;
  assign n33194 = n28117 ^ n4312 ^ 1'b0 ;
  assign n33195 = n3326 | n33194 ;
  assign n33196 = n21675 ^ n18963 ^ n5338 ;
  assign n33197 = n10468 ^ n8673 ^ 1'b0 ;
  assign n33198 = n4137 & n33197 ;
  assign n33199 = ~n33196 & n33198 ;
  assign n33202 = n6513 & ~n16185 ;
  assign n33203 = n33202 ^ n30077 ^ 1'b0 ;
  assign n33200 = n18124 ^ n8951 ^ 1'b0 ;
  assign n33201 = n23055 | n33200 ;
  assign n33204 = n33203 ^ n33201 ^ 1'b0 ;
  assign n33205 = n12170 ^ n6119 ^ 1'b0 ;
  assign n33206 = n10137 & n12636 ;
  assign n33207 = n17171 & n33206 ;
  assign n33208 = n33207 ^ n7217 ^ n432 ;
  assign n33209 = n33208 ^ n32880 ^ 1'b0 ;
  assign n33210 = n33205 & n33209 ;
  assign n33211 = ~n8329 & n21464 ;
  assign n33212 = ~n397 & n7857 ;
  assign n33213 = ( ~n1063 & n1989 ) | ( ~n1063 & n5219 ) | ( n1989 & n5219 ) ;
  assign n33214 = n17766 ^ x203 ^ 1'b0 ;
  assign n33215 = n33213 & ~n33214 ;
  assign n33216 = ( n8211 & ~n24988 ) | ( n8211 & n33215 ) | ( ~n24988 & n33215 ) ;
  assign n33217 = n24882 ^ n9447 ^ 1'b0 ;
  assign n33218 = ( n26541 & n27300 ) | ( n26541 & ~n33217 ) | ( n27300 & ~n33217 ) ;
  assign n33219 = n19893 ^ n12406 ^ n7244 ;
  assign n33220 = ~n7220 & n10518 ;
  assign n33221 = n33220 ^ n360 ^ 1'b0 ;
  assign n33222 = n10338 ^ n5839 ^ 1'b0 ;
  assign n33223 = n12180 | n33222 ;
  assign n33224 = n10886 & ~n33223 ;
  assign n33225 = n33224 ^ n20411 ^ 1'b0 ;
  assign n33226 = n15353 ^ n4207 ^ 1'b0 ;
  assign n33227 = n13837 ^ n5805 ^ 1'b0 ;
  assign n33228 = n33226 & ~n33227 ;
  assign n33229 = n17892 ^ n12843 ^ 1'b0 ;
  assign n33230 = ~n1430 & n33229 ;
  assign n33231 = n30188 ^ n2130 ^ 1'b0 ;
  assign n33232 = n30768 | n33231 ;
  assign n33233 = ( n3918 & n20524 ) | ( n3918 & n26281 ) | ( n20524 & n26281 ) ;
  assign n33235 = ( n4165 & n5063 ) | ( n4165 & ~n11649 ) | ( n5063 & ~n11649 ) ;
  assign n33234 = ~n6501 & n9267 ;
  assign n33236 = n33235 ^ n33234 ^ 1'b0 ;
  assign n33237 = n19566 & ~n33236 ;
  assign n33238 = n1323 & n5542 ;
  assign n33239 = n2801 & n30357 ;
  assign n33240 = n11108 ^ x214 ^ 1'b0 ;
  assign n33241 = n33239 & n33240 ;
  assign n33242 = n7454 & n13608 ;
  assign n33243 = n3879 | n12899 ;
  assign n33244 = n33242 & ~n33243 ;
  assign n33252 = n7916 & n9899 ;
  assign n33253 = ~n9899 & n33252 ;
  assign n33254 = n5312 & ~n11866 ;
  assign n33255 = n11866 & n33254 ;
  assign n33256 = ~n5157 & n8808 ;
  assign n33257 = n33255 & n33256 ;
  assign n33258 = n33257 ^ n3898 ^ 1'b0 ;
  assign n33259 = n33253 | n33258 ;
  assign n33260 = n33259 ^ x114 ^ 1'b0 ;
  assign n33249 = n9177 | n14476 ;
  assign n33250 = n14795 | n33249 ;
  assign n33245 = n27992 ^ n3413 ^ 1'b0 ;
  assign n33246 = n4425 | n33245 ;
  assign n33247 = n11844 ^ n4396 ^ 1'b0 ;
  assign n33248 = ~n33246 & n33247 ;
  assign n33251 = n33250 ^ n33248 ^ n11836 ;
  assign n33261 = n33260 ^ n33251 ^ n27498 ;
  assign n33262 = n14935 ^ n12339 ^ 1'b0 ;
  assign n33263 = ( n11706 & n20715 ) | ( n11706 & ~n26630 ) | ( n20715 & ~n26630 ) ;
  assign n33264 = n4765 & n14070 ;
  assign n33265 = n33263 & n33264 ;
  assign n33266 = n13703 | n28895 ;
  assign n33267 = n33266 ^ n11872 ^ 1'b0 ;
  assign n33268 = n271 & ~n3380 ;
  assign n33269 = n33268 ^ n20453 ^ 1'b0 ;
  assign n33270 = ~n13903 & n33269 ;
  assign n33271 = n33270 ^ n8270 ^ 1'b0 ;
  assign n33272 = n12772 & n19398 ;
  assign n33273 = n33272 ^ n22870 ^ 1'b0 ;
  assign n33274 = n21705 ^ n6851 ^ 1'b0 ;
  assign n33275 = ( ~n5521 & n6027 ) | ( ~n5521 & n33274 ) | ( n6027 & n33274 ) ;
  assign n33276 = n27660 ^ n26876 ^ 1'b0 ;
  assign n33277 = n7680 ^ n6762 ^ 1'b0 ;
  assign n33278 = n30206 ^ n2232 ^ 1'b0 ;
  assign n33279 = n29566 | n33278 ;
  assign n33280 = n14093 & ~n33279 ;
  assign n33281 = n18583 ^ n6079 ^ 1'b0 ;
  assign n33282 = n18529 ^ n4091 ^ 1'b0 ;
  assign n33283 = n33282 ^ n10420 ^ 1'b0 ;
  assign n33284 = n33281 | n33283 ;
  assign n33285 = ( n6907 & ~n9467 ) | ( n6907 & n10536 ) | ( ~n9467 & n10536 ) ;
  assign n33286 = n33285 ^ n20920 ^ 1'b0 ;
  assign n33287 = ( ~n12691 & n28565 ) | ( ~n12691 & n33286 ) | ( n28565 & n33286 ) ;
  assign n33288 = n1587 & n2281 ;
  assign n33289 = n6153 & n33288 ;
  assign n33290 = n4790 & ~n15946 ;
  assign n33291 = n33289 & n33290 ;
  assign n33292 = n33291 ^ n5190 ^ 1'b0 ;
  assign n33293 = n19118 & n33292 ;
  assign n33294 = n4778 & n19462 ;
  assign n33295 = n1097 & n15047 ;
  assign n33296 = n9126 & n33295 ;
  assign n33297 = ( n12760 & ~n19586 ) | ( n12760 & n33296 ) | ( ~n19586 & n33296 ) ;
  assign n33298 = n27604 ^ n8103 ^ 1'b0 ;
  assign n33299 = n22278 ^ n17259 ^ 1'b0 ;
  assign n33300 = ~n6504 & n8893 ;
  assign n33301 = n33300 ^ n9247 ^ n7033 ;
  assign n33302 = ~x199 & n33301 ;
  assign n33303 = n6762 & n22307 ;
  assign n33304 = n9952 | n10840 ;
  assign n33305 = n5134 & n33304 ;
  assign n33306 = n13240 & n26395 ;
  assign n33307 = n6101 & n33306 ;
  assign n33308 = n33305 | n33307 ;
  assign n33309 = ~n5177 & n10441 ;
  assign n33310 = ( n7624 & ~n14314 ) | ( n7624 & n18896 ) | ( ~n14314 & n18896 ) ;
  assign n33311 = n15392 | n25041 ;
  assign n33312 = n33310 & ~n33311 ;
  assign n33313 = n9986 ^ n2882 ^ 1'b0 ;
  assign n33314 = ~n15179 & n33313 ;
  assign n33315 = ( n7215 & n19874 ) | ( n7215 & n22753 ) | ( n19874 & n22753 ) ;
  assign n33316 = n14065 & ~n33315 ;
  assign n33317 = n16480 & n33316 ;
  assign n33318 = n11482 & ~n32554 ;
  assign n33319 = ~n27556 & n33318 ;
  assign n33320 = ~n29346 & n33319 ;
  assign n33321 = ~n4117 & n8999 ;
  assign n33322 = n2271 & ~n33321 ;
  assign n33323 = ~n3230 & n33322 ;
  assign n33324 = n25702 & ~n33323 ;
  assign n33325 = n31364 ^ n27629 ^ 1'b0 ;
  assign n33326 = n16006 & ~n25656 ;
  assign n33327 = n33326 ^ n22080 ^ 1'b0 ;
  assign n33328 = n5945 & n11918 ;
  assign n33329 = n26513 ^ n6790 ^ 1'b0 ;
  assign n33330 = ~n33328 & n33329 ;
  assign n33331 = n4287 ^ n1952 ^ 1'b0 ;
  assign n33332 = n930 | n15284 ;
  assign n33333 = n33331 | n33332 ;
  assign n33334 = n11088 ^ n7755 ^ 1'b0 ;
  assign n33335 = n8105 & ~n33334 ;
  assign n33336 = n33335 ^ n817 ^ 1'b0 ;
  assign n33337 = n33336 ^ n31317 ^ 1'b0 ;
  assign n33338 = ( ~n6272 & n14574 ) | ( ~n6272 & n33337 ) | ( n14574 & n33337 ) ;
  assign n33340 = n6644 | n13453 ;
  assign n33341 = n33340 ^ n9411 ^ 1'b0 ;
  assign n33342 = n10746 | n33341 ;
  assign n33339 = n2484 & ~n7040 ;
  assign n33343 = n33342 ^ n33339 ^ n7708 ;
  assign n33346 = n7593 | n21713 ;
  assign n33347 = n4994 & ~n33346 ;
  assign n33344 = ~n19489 & n26741 ;
  assign n33345 = n33344 ^ n1646 ^ 1'b0 ;
  assign n33348 = n33347 ^ n33345 ^ n22022 ;
  assign n33349 = n5051 ^ n1287 ^ 1'b0 ;
  assign n33350 = n33349 ^ n23024 ^ 1'b0 ;
  assign n33351 = n33348 & n33350 ;
  assign n33352 = n23472 & n33351 ;
  assign n33353 = ~n21209 & n24926 ;
  assign n33354 = ~n5294 & n33353 ;
  assign n33355 = n26614 & n33354 ;
  assign n33356 = n4379 ^ n2600 ^ 1'b0 ;
  assign n33357 = n2376 & ~n33356 ;
  assign n33358 = n1879 & n33357 ;
  assign n33359 = n33358 ^ n7064 ^ 1'b0 ;
  assign n33360 = ~n14975 & n33359 ;
  assign n33361 = n33360 ^ n13175 ^ 1'b0 ;
  assign n33362 = n428 | n33361 ;
  assign n33363 = n27499 & ~n33362 ;
  assign n33364 = n13741 | n19587 ;
  assign n33365 = n26158 & ~n33364 ;
  assign n33367 = n3278 | n19471 ;
  assign n33368 = n33367 ^ n28249 ^ n2797 ;
  assign n33366 = n12415 & n30859 ;
  assign n33369 = n33368 ^ n33366 ^ n23221 ;
  assign n33370 = n18653 & n27626 ;
  assign n33371 = n16252 & n33370 ;
  assign n33372 = n8632 & ~n21707 ;
  assign n33373 = n385 & n3254 ;
  assign n33374 = n33373 ^ n10322 ^ 1'b0 ;
  assign n33375 = ~n8096 & n31261 ;
  assign n33376 = n33374 | n33375 ;
  assign n33377 = n33376 ^ n20561 ^ 1'b0 ;
  assign n33378 = ( n23642 & n33372 ) | ( n23642 & ~n33377 ) | ( n33372 & ~n33377 ) ;
  assign n33379 = ( x85 & n556 ) | ( x85 & ~n1692 ) | ( n556 & ~n1692 ) ;
  assign n33380 = n14397 ^ n2544 ^ 1'b0 ;
  assign n33381 = n8296 & ~n33380 ;
  assign n33382 = n33381 ^ n19001 ^ 1'b0 ;
  assign n33383 = n33379 & ~n33382 ;
  assign n33384 = ~n18344 & n23114 ;
  assign n33385 = n33384 ^ n2669 ^ 1'b0 ;
  assign n33386 = ( ~n6290 & n33383 ) | ( ~n6290 & n33385 ) | ( n33383 & n33385 ) ;
  assign n33387 = n14881 & n17113 ;
  assign n33388 = n33387 ^ n8310 ^ 1'b0 ;
  assign n33389 = ~n11416 & n11427 ;
  assign n33390 = n26227 ^ n16908 ^ n3697 ;
  assign n33392 = n4542 & n8886 ;
  assign n33391 = ~n9653 & n11372 ;
  assign n33393 = n33392 ^ n33391 ^ n29901 ;
  assign n33394 = n33390 & ~n33393 ;
  assign n33395 = n18673 | n28528 ;
  assign n33396 = n33395 ^ n22246 ^ 1'b0 ;
  assign n33397 = n33396 ^ n20469 ^ n16026 ;
  assign n33398 = n7677 & n33397 ;
  assign n33399 = ~n6731 & n33398 ;
  assign n33400 = n9901 & n29143 ;
  assign n33401 = ~n553 & n33400 ;
  assign n33402 = n27423 ^ n23520 ^ n931 ;
  assign n33403 = ~n6589 & n14406 ;
  assign n33404 = n11004 ^ n6114 ^ x156 ;
  assign n33405 = n33404 ^ n25993 ^ 1'b0 ;
  assign n33406 = ( ~n7969 & n9746 ) | ( ~n7969 & n33405 ) | ( n9746 & n33405 ) ;
  assign n33407 = n33406 ^ n26906 ^ 1'b0 ;
  assign n33408 = n33403 | n33407 ;
  assign n33409 = ( x83 & n17480 ) | ( x83 & n30516 ) | ( n17480 & n30516 ) ;
  assign n33410 = n33409 ^ n4832 ^ 1'b0 ;
  assign n33411 = n9054 & n33410 ;
  assign n33412 = n14566 & ~n29373 ;
  assign n33413 = ~n18797 & n33412 ;
  assign n33414 = n33413 ^ n12493 ^ 1'b0 ;
  assign n33415 = ~n1791 & n33414 ;
  assign n33416 = n7853 ^ n1225 ^ 1'b0 ;
  assign n33417 = n33416 ^ n3122 ^ 1'b0 ;
  assign n33418 = n3333 & ~n33417 ;
  assign n33419 = n33418 ^ n27757 ^ 1'b0 ;
  assign n33420 = n19763 ^ n19471 ^ n7892 ;
  assign n33421 = n24394 ^ n17627 ^ 1'b0 ;
  assign n33422 = n3648 & n12339 ;
  assign n33423 = n33422 ^ n1686 ^ 1'b0 ;
  assign n33431 = ( n15468 & n16077 ) | ( n15468 & n29371 ) | ( n16077 & n29371 ) ;
  assign n33426 = n13146 ^ n3029 ^ 1'b0 ;
  assign n33425 = n2959 | n31004 ;
  assign n33427 = n33426 ^ n33425 ^ n3201 ;
  assign n33428 = n5725 | n33427 ;
  assign n33429 = n25522 | n33428 ;
  assign n33424 = n1115 | n20623 ;
  assign n33430 = n33429 ^ n33424 ^ 1'b0 ;
  assign n33432 = n33431 ^ n33430 ^ 1'b0 ;
  assign n33433 = n33423 & ~n33432 ;
  assign n33434 = n19370 & n22639 ;
  assign n33435 = n33434 ^ n8395 ^ 1'b0 ;
  assign n33436 = n33435 ^ n28734 ^ 1'b0 ;
  assign n33437 = n33436 ^ n17548 ^ n13563 ;
  assign n33438 = n33437 ^ n21229 ^ n3158 ;
  assign n33439 = ~n7423 & n19050 ;
  assign n33440 = n33438 & n33439 ;
  assign n33441 = n33440 ^ n14285 ^ 1'b0 ;
  assign n33442 = n13481 ^ n10943 ^ 1'b0 ;
  assign n33443 = n21358 & n33442 ;
  assign n33444 = n33443 ^ n21581 ^ 1'b0 ;
  assign n33445 = ( n3222 & n25554 ) | ( n3222 & ~n33444 ) | ( n25554 & ~n33444 ) ;
  assign n33446 = n3445 & ~n4445 ;
  assign n33447 = n33446 ^ n15433 ^ 1'b0 ;
  assign n33448 = x164 & n33447 ;
  assign n33449 = ( n829 & n3567 ) | ( n829 & ~n25406 ) | ( n3567 & ~n25406 ) ;
  assign n33450 = n33449 ^ n7603 ^ 1'b0 ;
  assign n33451 = n28157 ^ n26525 ^ n11847 ;
  assign n33452 = n481 & ~n10995 ;
  assign n33453 = ( ~n2781 & n10566 ) | ( ~n2781 & n33452 ) | ( n10566 & n33452 ) ;
  assign n33455 = n16657 & ~n32398 ;
  assign n33456 = ~n18189 & n33455 ;
  assign n33454 = ~n4580 & n14446 ;
  assign n33457 = n33456 ^ n33454 ^ 1'b0 ;
  assign n33458 = n3895 ^ x151 ^ 1'b0 ;
  assign n33459 = n570 & ~n33458 ;
  assign n33460 = n1996 & ~n4984 ;
  assign n33461 = n16391 & ~n33460 ;
  assign n33462 = n18987 ^ n12421 ^ 1'b0 ;
  assign n33463 = n7812 & ~n33462 ;
  assign n33464 = n33463 ^ n7112 ^ 1'b0 ;
  assign n33465 = n6163 & n7004 ;
  assign n33466 = ( n14285 & ~n14816 ) | ( n14285 & n33465 ) | ( ~n14816 & n33465 ) ;
  assign n33467 = n11601 & n15194 ;
  assign n33468 = n3785 & n33467 ;
  assign n33469 = ~n1246 & n31236 ;
  assign n33470 = n2180 | n27222 ;
  assign n33471 = n33470 ^ n26488 ^ 1'b0 ;
  assign n33472 = n33471 ^ n25747 ^ 1'b0 ;
  assign n33473 = ( n33468 & n33469 ) | ( n33468 & ~n33472 ) | ( n33469 & ~n33472 ) ;
  assign n33474 = n22574 ^ n6164 ^ 1'b0 ;
  assign n33475 = n33474 ^ n13784 ^ 1'b0 ;
  assign n33476 = ~n1965 & n3831 ;
  assign n33477 = ( n11718 & ~n17572 ) | ( n11718 & n33476 ) | ( ~n17572 & n33476 ) ;
  assign n33478 = n8440 & ~n33477 ;
  assign n33479 = ~n5131 & n24905 ;
  assign n33480 = ~n4550 & n33479 ;
  assign n33481 = n14451 ^ n11414 ^ n9522 ;
  assign n33482 = ( n27198 & n33480 ) | ( n27198 & ~n33481 ) | ( n33480 & ~n33481 ) ;
  assign n33483 = ( n5485 & ~n5635 ) | ( n5485 & n27814 ) | ( ~n5635 & n27814 ) ;
  assign n33484 = ~n5398 & n21341 ;
  assign n33485 = n31775 & n33484 ;
  assign n33486 = ( n10087 & ~n12335 ) | ( n10087 & n33485 ) | ( ~n12335 & n33485 ) ;
  assign n33487 = n15994 ^ n4114 ^ 1'b0 ;
  assign n33488 = ~n27981 & n33487 ;
  assign n33489 = ~n23865 & n33488 ;
  assign n33490 = ~n6141 & n23871 ;
  assign n33491 = ( n7411 & n9439 ) | ( n7411 & ~n15140 ) | ( n9439 & ~n15140 ) ;
  assign n33492 = n8173 & n12903 ;
  assign n33493 = n33491 & n33492 ;
  assign n33494 = n10279 | n18279 ;
  assign n33495 = n10431 ^ n462 ^ 1'b0 ;
  assign n33496 = ~n29502 & n33495 ;
  assign n33497 = n10596 ^ n2040 ^ n1814 ;
  assign n33498 = n5439 & ~n16299 ;
  assign n33499 = n1690 & n5934 ;
  assign n33500 = ~n15583 & n33499 ;
  assign n33501 = n33500 ^ n7675 ^ 1'b0 ;
  assign n33502 = n33498 & ~n33501 ;
  assign n33503 = ~n5760 & n22827 ;
  assign n33504 = n8887 & ~n33503 ;
  assign n33505 = n8720 & n9068 ;
  assign n33506 = ( n2481 & n10637 ) | ( n2481 & n17300 ) | ( n10637 & n17300 ) ;
  assign n33507 = ~n20784 & n33506 ;
  assign n33508 = n14715 & n33507 ;
  assign n33509 = n16662 ^ n14957 ^ 1'b0 ;
  assign n33510 = n20591 ^ n18072 ^ 1'b0 ;
  assign n33511 = x147 & ~n8013 ;
  assign n33512 = n7418 & n33511 ;
  assign n33513 = n33512 ^ x46 ^ 1'b0 ;
  assign n33514 = n16466 & ~n33513 ;
  assign n33515 = n10658 ^ n5590 ^ 1'b0 ;
  assign n33516 = n18015 | n33515 ;
  assign n33517 = n15450 ^ n5241 ^ 1'b0 ;
  assign n33518 = ~n1944 & n8276 ;
  assign n33519 = n10893 & n33518 ;
  assign n33520 = n33519 ^ n20750 ^ 1'b0 ;
  assign n33521 = n33517 & ~n33520 ;
  assign n33522 = n1126 | n3365 ;
  assign n33523 = n33522 ^ n4824 ^ 1'b0 ;
  assign n33524 = n33523 ^ n30866 ^ n18140 ;
  assign n33525 = n12187 | n33524 ;
  assign n33526 = n14609 ^ n13500 ^ 1'b0 ;
  assign n33527 = n28432 ^ n19052 ^ 1'b0 ;
  assign n33528 = n28640 & n33527 ;
  assign n33529 = n9199 & ~n15428 ;
  assign n33530 = n33529 ^ n21548 ^ 1'b0 ;
  assign n33531 = n28461 & ~n33530 ;
  assign n33532 = n33531 ^ n8836 ^ 1'b0 ;
  assign n33533 = n25211 | n33532 ;
  assign n33534 = ~n9561 & n30257 ;
  assign n33535 = n33534 ^ n27083 ^ 1'b0 ;
  assign n33536 = ( n481 & n950 ) | ( n481 & n33535 ) | ( n950 & n33535 ) ;
  assign n33537 = ( ~n15194 & n24609 ) | ( ~n15194 & n33536 ) | ( n24609 & n33536 ) ;
  assign n33538 = n7196 & n30551 ;
  assign n33539 = n33538 ^ n706 ^ 1'b0 ;
  assign n33540 = n16939 ^ n10949 ^ 1'b0 ;
  assign n33541 = n23902 & n33540 ;
  assign n33542 = n33539 & ~n33541 ;
  assign n33543 = ( n6189 & n17150 ) | ( n6189 & n32569 ) | ( n17150 & n32569 ) ;
  assign n33544 = ~n2791 & n8839 ;
  assign n33545 = n33543 & n33544 ;
  assign n33546 = ~n5091 & n7608 ;
  assign n33547 = n33545 & n33546 ;
  assign n33548 = n7585 ^ n1506 ^ 1'b0 ;
  assign n33549 = n981 & ~n8453 ;
  assign n33550 = ~n5770 & n33549 ;
  assign n33551 = n790 & ~n26937 ;
  assign n33552 = ( x22 & n10348 ) | ( x22 & ~n15675 ) | ( n10348 & ~n15675 ) ;
  assign n33553 = n2080 & n3344 ;
  assign n33554 = ~n11577 & n33553 ;
  assign n33555 = n5355 | n15079 ;
  assign n33556 = n8846 & ~n16047 ;
  assign n33557 = n14589 & ~n33556 ;
  assign n33558 = n3025 & n33557 ;
  assign n33561 = n5797 & ~n33054 ;
  assign n33559 = n6964 & ~n12745 ;
  assign n33560 = n33559 ^ n15840 ^ 1'b0 ;
  assign n33562 = n33561 ^ n33560 ^ 1'b0 ;
  assign n33563 = n10382 | n12973 ;
  assign n33568 = n13480 ^ n7683 ^ 1'b0 ;
  assign n33564 = n7997 ^ n4184 ^ n2527 ;
  assign n33565 = n20723 ^ n14490 ^ 1'b0 ;
  assign n33566 = ~n6824 & n33565 ;
  assign n33567 = ~n33564 & n33566 ;
  assign n33569 = n33568 ^ n33567 ^ 1'b0 ;
  assign n33570 = n21184 & ~n22709 ;
  assign n33571 = n33570 ^ n11616 ^ 1'b0 ;
  assign n33572 = n33571 ^ n27627 ^ 1'b0 ;
  assign n33573 = n3483 & ~n33572 ;
  assign n33574 = ~x52 & n1626 ;
  assign n33575 = n33574 ^ n24129 ^ 1'b0 ;
  assign n33576 = ~n2149 & n33575 ;
  assign n33577 = n33576 ^ n19783 ^ 1'b0 ;
  assign n33578 = n15618 ^ n4160 ^ n4038 ;
  assign n33579 = ~n17085 & n33578 ;
  assign n33580 = n27591 ^ n24327 ^ 1'b0 ;
  assign n33581 = n11262 & ~n33580 ;
  assign n33582 = ( n2129 & ~n33579 ) | ( n2129 & n33581 ) | ( ~n33579 & n33581 ) ;
  assign n33583 = n11718 ^ n9534 ^ 1'b0 ;
  assign n33584 = ~n27678 & n33583 ;
  assign n33585 = n21750 ^ n4998 ^ 1'b0 ;
  assign n33586 = n11692 ^ n5465 ^ 1'b0 ;
  assign n33587 = n26893 | n33586 ;
  assign n33588 = ~n5075 & n17522 ;
  assign n33589 = n33588 ^ n2581 ^ 1'b0 ;
  assign n33590 = ~n2879 & n27339 ;
  assign n33591 = n16244 ^ n15281 ^ 1'b0 ;
  assign n33592 = n3407 & n33591 ;
  assign n33593 = ~n17272 & n18390 ;
  assign n33594 = n11046 & n33593 ;
  assign n33595 = n33594 ^ n527 ^ 1'b0 ;
  assign n33596 = ~n981 & n2882 ;
  assign n33597 = n8516 & n33596 ;
  assign n33598 = n33597 ^ n3369 ^ 1'b0 ;
  assign n33599 = x70 & n33598 ;
  assign n33600 = n1110 & n4899 ;
  assign n33601 = n33600 ^ n9902 ^ n749 ;
  assign n33602 = n650 & ~n12835 ;
  assign n33603 = ( n7890 & n18601 ) | ( n7890 & n33602 ) | ( n18601 & n33602 ) ;
  assign n33604 = n3359 ^ n490 ^ 1'b0 ;
  assign n33605 = ( n4722 & ~n4802 ) | ( n4722 & n33604 ) | ( ~n4802 & n33604 ) ;
  assign n33606 = n24977 ^ n11145 ^ 1'b0 ;
  assign n33607 = ~n17194 & n29337 ;
  assign n33608 = n33607 ^ n26629 ^ 1'b0 ;
  assign n33609 = n15784 ^ n884 ^ 1'b0 ;
  assign n33610 = ~n3009 & n33609 ;
  assign n33611 = n32742 & ~n33610 ;
  assign n33612 = ~n1314 & n5137 ;
  assign n33613 = ~x187 & n33612 ;
  assign n33614 = n19369 ^ n12886 ^ n12353 ;
  assign n33615 = n9971 ^ n6369 ^ 1'b0 ;
  assign n33616 = n14636 ^ n5693 ^ 1'b0 ;
  assign n33617 = n3336 & n11464 ;
  assign n33618 = n2033 ^ n909 ^ 1'b0 ;
  assign n33619 = n13902 & ~n33618 ;
  assign n33620 = n33619 ^ n11643 ^ 1'b0 ;
  assign n33621 = n22497 ^ n14040 ^ n8905 ;
  assign n33622 = n33621 ^ n31919 ^ 1'b0 ;
  assign n33623 = n20511 | n33622 ;
  assign n33624 = n21499 | n33623 ;
  assign n33625 = n31806 | n33624 ;
  assign n33626 = n18337 ^ n2810 ^ 1'b0 ;
  assign n33627 = n7317 | n33626 ;
  assign n33628 = n13052 ^ n10023 ^ 1'b0 ;
  assign n33629 = n33627 | n33628 ;
  assign n33630 = n20777 ^ n7958 ^ 1'b0 ;
  assign n33631 = n22885 & n33630 ;
  assign n33632 = n2118 & ~n4382 ;
  assign n33633 = n653 | n3415 ;
  assign n33634 = n33633 ^ n6462 ^ 1'b0 ;
  assign n33635 = ( n2702 & n8618 ) | ( n2702 & n30401 ) | ( n8618 & n30401 ) ;
  assign n33636 = n20670 ^ n1890 ^ 1'b0 ;
  assign n33637 = n6613 ^ n5806 ^ 1'b0 ;
  assign n33638 = n5200 & n33637 ;
  assign n33639 = n1191 | n33638 ;
  assign n33640 = ( n26319 & ~n33636 ) | ( n26319 & n33639 ) | ( ~n33636 & n33639 ) ;
  assign n33641 = n19570 ^ n16129 ^ 1'b0 ;
  assign n33642 = n2144 | n33641 ;
  assign n33643 = n29573 & ~n33642 ;
  assign n33644 = ~n21796 & n33643 ;
  assign n33645 = ~n18695 & n28779 ;
  assign n33646 = n13635 & n33645 ;
  assign n33647 = n33646 ^ n30995 ^ 1'b0 ;
  assign n33648 = n3261 ^ n1646 ^ 1'b0 ;
  assign n33649 = ~n4039 & n33648 ;
  assign n33650 = n22659 ^ n4391 ^ 1'b0 ;
  assign n33651 = n739 & ~n33650 ;
  assign n33652 = ~n8828 & n33651 ;
  assign n33653 = ~n22027 & n33652 ;
  assign n33654 = n19225 | n33653 ;
  assign n33655 = n33649 | n33654 ;
  assign n33656 = n7048 & ~n7871 ;
  assign n33657 = n671 & n33656 ;
  assign n33658 = n33657 ^ n8666 ^ 1'b0 ;
  assign n33659 = n15347 ^ n7354 ^ 1'b0 ;
  assign n33660 = ~n3620 & n14229 ;
  assign n33661 = n5461 | n33660 ;
  assign n33662 = n33659 & ~n33661 ;
  assign n33663 = n20511 ^ n4292 ^ 1'b0 ;
  assign n33664 = ~n14344 & n33663 ;
  assign n33665 = ~n10598 & n13774 ;
  assign n33666 = n6727 & n13621 ;
  assign n33667 = n16186 ^ n12271 ^ 1'b0 ;
  assign n33668 = n16026 | n17013 ;
  assign n33669 = n16351 | n33668 ;
  assign n33670 = n17644 ^ n12839 ^ 1'b0 ;
  assign n33671 = n33669 & n33670 ;
  assign n33672 = n33667 & n33671 ;
  assign n33673 = n33666 | n33672 ;
  assign n33674 = n30330 ^ n17200 ^ 1'b0 ;
  assign n33675 = n28394 & ~n30535 ;
  assign n33676 = n9456 & n33675 ;
  assign n33677 = n28150 ^ n5376 ^ 1'b0 ;
  assign n33678 = n11719 | n33677 ;
  assign n33679 = n15710 ^ n4154 ^ 1'b0 ;
  assign n33680 = n12500 | n33679 ;
  assign n33681 = n23133 | n33680 ;
  assign n33682 = n33678 & ~n33681 ;
  assign n33683 = n12572 & n25875 ;
  assign n33684 = n33683 ^ n10539 ^ 1'b0 ;
  assign n33685 = ~n1687 & n5976 ;
  assign n33686 = n1323 & n27232 ;
  assign n33687 = n33685 & n33686 ;
  assign n33688 = n1558 & n3988 ;
  assign n33689 = n22079 & ~n33688 ;
  assign n33690 = ~n22079 & n33689 ;
  assign n33691 = n33690 ^ n17071 ^ 1'b0 ;
  assign n33692 = n5359 & ~n26961 ;
  assign n33693 = n33692 ^ n16485 ^ 1'b0 ;
  assign n33694 = ~n6851 & n8229 ;
  assign n33695 = n10943 & n33694 ;
  assign n33696 = n1297 | n4207 ;
  assign n33697 = n32554 & ~n33696 ;
  assign n33698 = n33697 ^ n5306 ^ 1'b0 ;
  assign n33699 = ( n26515 & n33695 ) | ( n26515 & ~n33698 ) | ( n33695 & ~n33698 ) ;
  assign n33700 = n31163 ^ n8948 ^ 1'b0 ;
  assign n33701 = n3451 | n33700 ;
  assign n33702 = n33699 | n33701 ;
  assign n33703 = n16392 ^ n8428 ^ 1'b0 ;
  assign n33704 = n3445 & n33703 ;
  assign n33705 = n2017 & n33704 ;
  assign n33706 = n33705 ^ n12637 ^ 1'b0 ;
  assign n33707 = n33706 ^ n21506 ^ n10160 ;
  assign n33708 = n12917 ^ n702 ^ 1'b0 ;
  assign n33709 = n4892 & n33708 ;
  assign n33710 = n10051 & n33709 ;
  assign n33711 = n33710 ^ n8739 ^ 1'b0 ;
  assign n33712 = n33711 ^ n7382 ^ 1'b0 ;
  assign n33713 = ( n9783 & ~n20950 ) | ( n9783 & n33712 ) | ( ~n20950 & n33712 ) ;
  assign n33714 = n33379 ^ n16911 ^ 1'b0 ;
  assign n33715 = ~n5971 & n13835 ;
  assign n33716 = n5497 | n33715 ;
  assign n33717 = n27563 | n33716 ;
  assign n33718 = n33119 ^ n4370 ^ n2793 ;
  assign n33721 = n10774 ^ n5513 ^ 1'b0 ;
  assign n33722 = ~n15362 & n33721 ;
  assign n33719 = ~n2354 & n4749 ;
  assign n33720 = n1046 & ~n33719 ;
  assign n33723 = n33722 ^ n33720 ^ 1'b0 ;
  assign n33724 = n33723 ^ n25505 ^ n5549 ;
  assign n33725 = n33724 ^ n21783 ^ n11123 ;
  assign n33726 = ~n16179 & n23717 ;
  assign n33727 = n5592 | n27133 ;
  assign n33728 = n33727 ^ n4026 ^ 1'b0 ;
  assign n33729 = n33728 ^ n6805 ^ 1'b0 ;
  assign n33730 = n7627 & ~n23971 ;
  assign n33732 = ~n13584 & n15322 ;
  assign n33731 = ~n16384 & n19008 ;
  assign n33733 = n33732 ^ n33731 ^ 1'b0 ;
  assign n33734 = n26559 & ~n33733 ;
  assign n33735 = ~x207 & n10575 ;
  assign n33736 = ( n8782 & n22517 ) | ( n8782 & n33735 ) | ( n22517 & n33735 ) ;
  assign n33737 = n9342 ^ n4413 ^ 1'b0 ;
  assign n33738 = ~n33736 & n33737 ;
  assign n33739 = n12603 ^ n9242 ^ 1'b0 ;
  assign n33740 = n3332 & n33739 ;
  assign n33741 = n33740 ^ n3953 ^ 1'b0 ;
  assign n33742 = ( ~n23700 & n33738 ) | ( ~n23700 & n33741 ) | ( n33738 & n33741 ) ;
  assign n33744 = n8463 & ~n24151 ;
  assign n33743 = n10759 | n20321 ;
  assign n33745 = n33744 ^ n33743 ^ 1'b0 ;
  assign n33746 = n6825 & n10253 ;
  assign n33747 = ~x107 & n33746 ;
  assign n33748 = n33747 ^ n6808 ^ 1'b0 ;
  assign n33749 = n25221 & n33748 ;
  assign n33750 = n4724 ^ n2824 ^ 1'b0 ;
  assign n33751 = x120 & n33750 ;
  assign n33752 = n33751 ^ n5560 ^ 1'b0 ;
  assign n33753 = n28658 & ~n33752 ;
  assign n33754 = ~n7559 & n25318 ;
  assign n33755 = ~n25318 & n33754 ;
  assign n33756 = n7812 ^ n4775 ^ 1'b0 ;
  assign n33757 = n6901 | n33756 ;
  assign n33758 = n33757 ^ n13896 ^ 1'b0 ;
  assign n33759 = n25773 ^ n8554 ^ n4174 ;
  assign n33760 = ~n16444 & n28035 ;
  assign n33761 = n15098 & ~n23814 ;
  assign n33762 = n33761 ^ n436 ^ 1'b0 ;
  assign n33763 = n875 | n33762 ;
  assign n33764 = n4369 ^ n3000 ^ 1'b0 ;
  assign n33765 = x7 & n5196 ;
  assign n33766 = n33765 ^ n24246 ^ 1'b0 ;
  assign n33767 = ~n3664 & n32134 ;
  assign n33768 = ~n516 & n12068 ;
  assign n33769 = ~n10114 & n33768 ;
  assign n33770 = n33769 ^ n24347 ^ n9653 ;
  assign n33772 = n18903 ^ n9451 ^ n3506 ;
  assign n33773 = n8929 | n33772 ;
  assign n33771 = n27914 ^ n10333 ^ n5051 ;
  assign n33774 = n33773 ^ n33771 ^ n1495 ;
  assign n33777 = ~n7975 & n28798 ;
  assign n33778 = ~n28798 & n33777 ;
  assign n33775 = n13021 ^ n1843 ^ 1'b0 ;
  assign n33776 = n1199 | n33775 ;
  assign n33779 = n33778 ^ n33776 ^ n10068 ;
  assign n33780 = n23121 & ~n25776 ;
  assign n33781 = n2286 & n33780 ;
  assign n33782 = n8557 ^ n2692 ^ 1'b0 ;
  assign n33783 = n17489 & ~n33782 ;
  assign n33784 = ~n8819 & n15027 ;
  assign n33785 = n931 & ~n18323 ;
  assign n33786 = ~n18296 & n33785 ;
  assign n33787 = ~n11649 & n33786 ;
  assign n33788 = n1713 | n9431 ;
  assign n33789 = n17766 | n33788 ;
  assign n33790 = n3809 & ~n33789 ;
  assign n33791 = n5681 & ~n30025 ;
  assign n33792 = n5446 & ~n9881 ;
  assign n33793 = n27055 ^ n23230 ^ n7115 ;
  assign n33794 = ( ~n5006 & n10331 ) | ( ~n5006 & n10846 ) | ( n10331 & n10846 ) ;
  assign n33795 = n33794 ^ n13201 ^ n11009 ;
  assign n33798 = n23637 ^ n5740 ^ 1'b0 ;
  assign n33797 = n1860 & n11888 ;
  assign n33799 = n33798 ^ n33797 ^ 1'b0 ;
  assign n33796 = n2930 & n30144 ;
  assign n33800 = n33799 ^ n33796 ^ 1'b0 ;
  assign n33807 = n7154 ^ n3757 ^ 1'b0 ;
  assign n33801 = n9054 | n29093 ;
  assign n33802 = ( ~n11504 & n12934 ) | ( ~n11504 & n33801 ) | ( n12934 & n33801 ) ;
  assign n33803 = x67 | n33802 ;
  assign n33804 = n3574 | n33803 ;
  assign n33805 = ~x222 & n15204 ;
  assign n33806 = ~n33804 & n33805 ;
  assign n33808 = n33807 ^ n33806 ^ n21685 ;
  assign n33809 = n20071 ^ n14314 ^ 1'b0 ;
  assign n33810 = n33808 & n33809 ;
  assign n33811 = ~n19406 & n23071 ;
  assign n33812 = ~n1374 & n33811 ;
  assign n33813 = n24018 ^ n18367 ^ n7348 ;
  assign n33814 = n4476 & n16735 ;
  assign n33815 = n18561 ^ n6382 ^ 1'b0 ;
  assign n33816 = n2073 | n11754 ;
  assign n33817 = n25290 & ~n33816 ;
  assign n33818 = n11335 & ~n33817 ;
  assign n33819 = n1489 & ~n15241 ;
  assign n33820 = n17882 ^ n16519 ^ 1'b0 ;
  assign n33821 = x8 & n33820 ;
  assign n33822 = ~n5666 & n33821 ;
  assign n33823 = n2443 & ~n31555 ;
  assign n33824 = ~n28452 & n33823 ;
  assign n33825 = ~n6555 & n15268 ;
  assign n33826 = n2203 ^ n936 ^ n883 ;
  assign n33827 = ~n19117 & n33826 ;
  assign n33828 = n33827 ^ n16098 ^ 1'b0 ;
  assign n33829 = ( ~n18451 & n32910 ) | ( ~n18451 & n33828 ) | ( n32910 & n33828 ) ;
  assign n33830 = ~n4590 & n8520 ;
  assign n33831 = n33830 ^ n15350 ^ 1'b0 ;
  assign n33832 = n24376 ^ n19948 ^ n13279 ;
  assign n33833 = n12102 ^ n2057 ^ 1'b0 ;
  assign n33834 = n33832 & n33833 ;
  assign n33835 = ( x71 & n645 ) | ( x71 & ~n10985 ) | ( n645 & ~n10985 ) ;
  assign n33836 = n33835 ^ n18364 ^ 1'b0 ;
  assign n33837 = n25420 ^ n21393 ^ n8715 ;
  assign n33838 = ( x161 & n11109 ) | ( x161 & ~n33837 ) | ( n11109 & ~n33837 ) ;
  assign n33839 = n7037 ^ n1401 ^ 1'b0 ;
  assign n33840 = n24085 & n33839 ;
  assign n33841 = ~n2522 & n33840 ;
  assign n33842 = n2853 & ~n33841 ;
  assign n33843 = n4826 & ~n5830 ;
  assign n33844 = n22666 ^ n1340 ^ 1'b0 ;
  assign n33845 = n790 & ~n11241 ;
  assign n33846 = n12773 ^ n12291 ^ 1'b0 ;
  assign n33847 = n33845 & n33846 ;
  assign n33848 = ~n6045 & n16836 ;
  assign n33849 = n33848 ^ n3822 ^ 1'b0 ;
  assign n33850 = ~n631 & n33849 ;
  assign n33851 = n26866 ^ n24320 ^ 1'b0 ;
  assign n33852 = n33850 & ~n33851 ;
  assign n33854 = n7119 ^ n3848 ^ 1'b0 ;
  assign n33855 = n18503 & ~n33854 ;
  assign n33853 = n2955 | n3752 ;
  assign n33856 = n33855 ^ n33853 ^ 1'b0 ;
  assign n33857 = ( n3879 & n33150 ) | ( n3879 & ~n33856 ) | ( n33150 & ~n33856 ) ;
  assign n33858 = n32929 ^ n23978 ^ 1'b0 ;
  assign n33859 = ~n19276 & n33858 ;
  assign n33860 = n11168 & ~n21940 ;
  assign n33861 = n1090 & n33436 ;
  assign n33862 = ~n31609 & n33861 ;
  assign n33863 = n17557 ^ x15 ^ 1'b0 ;
  assign n33864 = n5805 & n33863 ;
  assign n33865 = ~n3320 & n6232 ;
  assign n33866 = ~n1669 & n33865 ;
  assign n33867 = n24275 & ~n33866 ;
  assign n33868 = n33867 ^ n10600 ^ 1'b0 ;
  assign n33869 = ~n9496 & n33868 ;
  assign n33870 = n15932 ^ n3666 ^ 1'b0 ;
  assign n33871 = ( n4194 & n18618 ) | ( n4194 & ~n33870 ) | ( n18618 & ~n33870 ) ;
  assign n33872 = n33869 & n33871 ;
  assign n33873 = ( ~n7002 & n9500 ) | ( ~n7002 & n23797 ) | ( n9500 & n23797 ) ;
  assign n33874 = ~n5348 & n16307 ;
  assign n33875 = ~n12169 & n33874 ;
  assign n33876 = n12572 & ~n33875 ;
  assign n33877 = ~n7012 & n29033 ;
  assign n33878 = n16012 ^ n10626 ^ 1'b0 ;
  assign n33879 = n33878 ^ n7380 ^ 1'b0 ;
  assign n33880 = n19079 | n33879 ;
  assign n33881 = n256 & ~n263 ;
  assign n33882 = ~n14584 & n33881 ;
  assign n33883 = n23513 ^ n8747 ^ 1'b0 ;
  assign n33884 = n33882 | n33883 ;
  assign n33885 = n15692 ^ n5740 ^ 1'b0 ;
  assign n33888 = n18839 ^ n10653 ^ 1'b0 ;
  assign n33889 = ~n10736 & n33888 ;
  assign n33890 = n32824 ^ n11297 ^ 1'b0 ;
  assign n33891 = n33889 & ~n33890 ;
  assign n33886 = n23469 ^ n1768 ^ 1'b0 ;
  assign n33887 = n5139 & ~n33886 ;
  assign n33892 = n33891 ^ n33887 ^ 1'b0 ;
  assign n33893 = n14328 ^ n2149 ^ 1'b0 ;
  assign n33894 = n31322 | n33893 ;
  assign n33895 = ~n20493 & n25723 ;
  assign n33896 = n33894 & n33895 ;
  assign n33897 = n27627 ^ n6333 ^ 1'b0 ;
  assign n33898 = n25552 ^ n1019 ^ 1'b0 ;
  assign n33899 = n26099 & ~n33898 ;
  assign n33900 = n26989 & n33899 ;
  assign n33901 = ( ~n9530 & n17993 ) | ( ~n9530 & n33900 ) | ( n17993 & n33900 ) ;
  assign n33902 = n1381 ^ x63 ^ 1'b0 ;
  assign n33903 = n33902 ^ n3043 ^ n1941 ;
  assign n33904 = n32641 & ~n33903 ;
  assign n33905 = ~n8237 & n33904 ;
  assign n33906 = n6768 | n8484 ;
  assign n33907 = n393 & ~n4921 ;
  assign n33908 = ( ~n3111 & n18096 ) | ( ~n3111 & n33907 ) | ( n18096 & n33907 ) ;
  assign n33909 = n1448 & n9699 ;
  assign n33910 = n28895 ^ n9073 ^ 1'b0 ;
  assign n33923 = n677 & ~n24748 ;
  assign n33924 = n33923 ^ n4493 ^ 1'b0 ;
  assign n33925 = n2765 | n33924 ;
  assign n33926 = n33925 ^ n3326 ^ 1'b0 ;
  assign n33927 = n33926 ^ n14251 ^ 1'b0 ;
  assign n33918 = n10377 & n14603 ;
  assign n33912 = n22438 ^ n10787 ^ n1036 ;
  assign n33913 = n31294 ^ n835 ^ 1'b0 ;
  assign n33914 = n33913 ^ n1122 ^ n681 ;
  assign n33915 = n33914 ^ n6808 ^ 1'b0 ;
  assign n33916 = ~n33912 & n33915 ;
  assign n33917 = n23591 & n33916 ;
  assign n33919 = n33918 ^ n33917 ^ 1'b0 ;
  assign n33920 = ( n1930 & ~n4359 ) | ( n1930 & n11573 ) | ( ~n4359 & n11573 ) ;
  assign n33921 = n12256 & n33920 ;
  assign n33922 = n33919 & n33921 ;
  assign n33911 = n23157 ^ n6802 ^ n723 ;
  assign n33928 = n33927 ^ n33922 ^ n33911 ;
  assign n33929 = n7673 & ~n16596 ;
  assign n33930 = n7726 & n33929 ;
  assign n33931 = n33930 ^ n7233 ^ n5302 ;
  assign n33932 = n5920 & ~n11503 ;
  assign n33933 = n15806 & n33932 ;
  assign n33934 = n30082 & ~n33933 ;
  assign n33935 = n33934 ^ n5484 ^ 1'b0 ;
  assign n33936 = n12836 ^ n704 ^ 1'b0 ;
  assign n33938 = n1348 & n19363 ;
  assign n33939 = n33938 ^ n24221 ^ 1'b0 ;
  assign n33937 = n24926 ^ n15819 ^ n10625 ;
  assign n33940 = n33939 ^ n33937 ^ 1'b0 ;
  assign n33941 = ~n33936 & n33940 ;
  assign n33942 = n8681 ^ n1473 ^ 1'b0 ;
  assign n33943 = n15741 & ~n33942 ;
  assign n33944 = n33943 ^ n5657 ^ 1'b0 ;
  assign n33945 = n8527 ^ n7431 ^ 1'b0 ;
  assign n33946 = n21638 & n33945 ;
  assign n33947 = n17150 ^ n3254 ^ 1'b0 ;
  assign n33948 = n26593 | n32126 ;
  assign n33949 = n33948 ^ n2158 ^ 1'b0 ;
  assign n33950 = n33947 & ~n33949 ;
  assign n33953 = n12986 & n19138 ;
  assign n33951 = ~n11722 & n29815 ;
  assign n33952 = ~n11571 & n33951 ;
  assign n33954 = n33953 ^ n33952 ^ 1'b0 ;
  assign n33955 = ~n15347 & n33954 ;
  assign n33956 = n24781 ^ n21556 ^ n12603 ;
  assign n33957 = n7178 ^ n2423 ^ 1'b0 ;
  assign n33958 = n5538 & ~n33957 ;
  assign n33959 = n9998 ^ n5898 ^ n3633 ;
  assign n33960 = n33958 & n33959 ;
  assign n33961 = n31213 ^ n5934 ^ 1'b0 ;
  assign n33962 = ~n669 & n16147 ;
  assign n33963 = n23400 ^ n2093 ^ 1'b0 ;
  assign n33964 = n19526 & ~n33963 ;
  assign n33965 = n33964 ^ n17352 ^ 1'b0 ;
  assign n33966 = ( n1215 & ~n6764 ) | ( n1215 & n33965 ) | ( ~n6764 & n33965 ) ;
  assign n33967 = n15462 & n33966 ;
  assign n33968 = ~n11350 & n19456 ;
  assign n33969 = ~n9336 & n33968 ;
  assign n33970 = n2839 & ~n7839 ;
  assign n33971 = n10275 | n33970 ;
  assign n33972 = n33017 ^ n1289 ^ 1'b0 ;
  assign n33973 = n33971 & n33972 ;
  assign n33974 = n2120 & n27881 ;
  assign n33975 = n30437 & ~n33974 ;
  assign n33976 = n33975 ^ n14655 ^ 1'b0 ;
  assign n33977 = n6440 | n12198 ;
  assign n33978 = n33977 ^ n13264 ^ 1'b0 ;
  assign n33979 = n9345 & n33978 ;
  assign n33980 = n11861 & ~n33979 ;
  assign n33981 = n33980 ^ n11267 ^ 1'b0 ;
  assign n33982 = n33981 ^ n33822 ^ n31540 ;
  assign n33983 = ~n3050 & n32713 ;
  assign n33984 = n33983 ^ n19602 ^ 1'b0 ;
  assign n33985 = n33984 ^ n14828 ^ n10325 ;
  assign n33986 = n19753 ^ n12233 ^ 1'b0 ;
  assign n33987 = n13186 & n33986 ;
  assign n33988 = n15516 | n16237 ;
  assign n33989 = n24834 | n33988 ;
  assign n33990 = n33989 ^ n18773 ^ 1'b0 ;
  assign n33991 = ~n18725 & n19787 ;
  assign n33992 = ~n11263 & n33991 ;
  assign n33993 = ( n18784 & n25636 ) | ( n18784 & ~n33992 ) | ( n25636 & ~n33992 ) ;
  assign n33994 = n29886 ^ n21750 ^ n1442 ;
  assign n33995 = n5642 | n10779 ;
  assign n33996 = n14267 & ~n33995 ;
  assign n33997 = n22888 ^ n11842 ^ 1'b0 ;
  assign n33998 = x84 & n33997 ;
  assign n33999 = n1069 & n4030 ;
  assign n34000 = n20976 ^ n11301 ^ 1'b0 ;
  assign n34001 = ~n10586 & n34000 ;
  assign n34002 = n13693 ^ n11474 ^ 1'b0 ;
  assign n34003 = n34001 & n34002 ;
  assign n34004 = n6384 | n16633 ;
  assign n34005 = n24705 ^ n17131 ^ n10385 ;
  assign n34006 = n16971 ^ n15561 ^ n1029 ;
  assign n34007 = n15975 & ~n24585 ;
  assign n34008 = n34007 ^ n21004 ^ 1'b0 ;
  assign n34009 = ~n5725 & n13533 ;
  assign n34010 = n34009 ^ n27947 ^ 1'b0 ;
  assign n34011 = n10049 ^ n8725 ^ 1'b0 ;
  assign n34012 = n22704 & ~n34011 ;
  assign n34013 = n12943 ^ n4741 ^ 1'b0 ;
  assign n34016 = ~n2739 & n7000 ;
  assign n34017 = n34016 ^ n983 ^ 1'b0 ;
  assign n34018 = n10122 | n34017 ;
  assign n34014 = n9890 ^ n2339 ^ 1'b0 ;
  assign n34015 = n3263 & n34014 ;
  assign n34019 = n34018 ^ n34015 ^ 1'b0 ;
  assign n34020 = n3053 & n34019 ;
  assign n34021 = n13749 & n34020 ;
  assign n34023 = n7788 | n29392 ;
  assign n34024 = n12419 | n34023 ;
  assign n34022 = n15093 ^ n10302 ^ 1'b0 ;
  assign n34025 = n34024 ^ n34022 ^ n26508 ;
  assign n34026 = n13936 & n22070 ;
  assign n34027 = ~n24337 & n34026 ;
  assign n34028 = n5099 ^ n2806 ^ 1'b0 ;
  assign n34029 = n25963 & ~n34028 ;
  assign n34036 = n6432 ^ n3178 ^ 1'b0 ;
  assign n34037 = n9952 & n34036 ;
  assign n34030 = n18879 ^ n1669 ^ 1'b0 ;
  assign n34031 = n6808 | n34030 ;
  assign n34032 = ( n838 & ~n11831 ) | ( n838 & n34031 ) | ( ~n11831 & n34031 ) ;
  assign n34033 = n12800 & ~n34032 ;
  assign n34034 = n34033 ^ n12187 ^ 1'b0 ;
  assign n34035 = ( ~n2525 & n10334 ) | ( ~n2525 & n34034 ) | ( n10334 & n34034 ) ;
  assign n34038 = n34037 ^ n34035 ^ n5766 ;
  assign n34039 = n12175 & n20015 ;
  assign n34040 = n34038 & n34039 ;
  assign n34041 = ~n7710 & n33866 ;
  assign n34042 = n34040 | n34041 ;
  assign n34043 = n1489 & ~n34042 ;
  assign n34044 = n33866 ^ n14862 ^ 1'b0 ;
  assign n34045 = ~n1930 & n9157 ;
  assign n34046 = n34045 ^ n23066 ^ 1'b0 ;
  assign n34047 = n34044 | n34046 ;
  assign n34048 = n10696 & ~n34047 ;
  assign n34049 = n20743 & n21605 ;
  assign n34050 = n20695 ^ n6044 ^ 1'b0 ;
  assign n34051 = x185 & n34050 ;
  assign n34052 = n22709 ^ n4657 ^ 1'b0 ;
  assign n34053 = ( n5678 & ~n34051 ) | ( n5678 & n34052 ) | ( ~n34051 & n34052 ) ;
  assign n34054 = ~n3847 & n14062 ;
  assign n34055 = ~n24945 & n34054 ;
  assign n34056 = ~n824 & n5740 ;
  assign n34057 = ( n7867 & ~n34055 ) | ( n7867 & n34056 ) | ( ~n34055 & n34056 ) ;
  assign n34058 = n28937 ^ n17178 ^ 1'b0 ;
  assign n34059 = n591 & n13936 ;
  assign n34060 = n34059 ^ n6188 ^ 1'b0 ;
  assign n34061 = n26642 ^ n12762 ^ 1'b0 ;
  assign n34062 = n20392 | n34061 ;
  assign n34063 = n12917 | n18906 ;
  assign n34064 = n34062 & ~n34063 ;
  assign n34065 = n26192 ^ n4622 ^ 1'b0 ;
  assign n34066 = n7916 ^ n7035 ^ x107 ;
  assign n34067 = n21334 | n34066 ;
  assign n34068 = n17026 ^ n14383 ^ 1'b0 ;
  assign n34069 = n7608 & n34068 ;
  assign n34070 = n20723 & ~n34069 ;
  assign n34071 = n1387 | n6152 ;
  assign n34072 = n13981 ^ n2728 ^ 1'b0 ;
  assign n34073 = n3877 & n34072 ;
  assign n34074 = ~n2166 & n34073 ;
  assign n34075 = n12072 & n30851 ;
  assign n34076 = n26045 & n34075 ;
  assign n34077 = n26777 ^ n1088 ^ 1'b0 ;
  assign n34078 = n13830 & n34077 ;
  assign n34079 = ( ~n5967 & n9127 ) | ( ~n5967 & n13386 ) | ( n9127 & n13386 ) ;
  assign n34080 = n19470 ^ n19298 ^ n2257 ;
  assign n34081 = n23175 | n34080 ;
  assign n34082 = n34079 & ~n34081 ;
  assign n34083 = n32586 ^ n24317 ^ 1'b0 ;
  assign n34084 = n12443 ^ n3359 ^ 1'b0 ;
  assign n34085 = n34083 | n34084 ;
  assign n34086 = n32549 | n34085 ;
  assign n34087 = n707 & ~n813 ;
  assign n34088 = ~n4541 & n34087 ;
  assign n34089 = n34088 ^ n3104 ^ n2812 ;
  assign n34090 = n34089 ^ n17891 ^ 1'b0 ;
  assign n34091 = n34090 ^ n26020 ^ n25732 ;
  assign n34092 = ~n9988 & n13516 ;
  assign n34093 = n22120 ^ n10046 ^ 1'b0 ;
  assign n34094 = n34092 & n34093 ;
  assign n34095 = ~n11047 & n27239 ;
  assign n34096 = ~n9784 & n34095 ;
  assign n34100 = ( n2267 & ~n7542 ) | ( n2267 & n10368 ) | ( ~n7542 & n10368 ) ;
  assign n34101 = n34100 ^ n6528 ^ 1'b0 ;
  assign n34102 = n10935 & ~n34101 ;
  assign n34103 = n15692 ^ n10172 ^ 1'b0 ;
  assign n34104 = n34102 & ~n34103 ;
  assign n34097 = n527 | n711 ;
  assign n34098 = n24269 & ~n34097 ;
  assign n34099 = n11624 | n34098 ;
  assign n34105 = n34104 ^ n34099 ^ 1'b0 ;
  assign n34106 = n9581 & n28456 ;
  assign n34107 = n34106 ^ n1878 ^ 1'b0 ;
  assign n34108 = n34107 ^ n6013 ^ 1'b0 ;
  assign n34109 = n13757 ^ n11857 ^ 1'b0 ;
  assign n34110 = n32030 | n34109 ;
  assign n34111 = n3363 | n34110 ;
  assign n34112 = n34111 ^ n29076 ^ 1'b0 ;
  assign n34113 = n25244 ^ n24818 ^ n8828 ;
  assign n34114 = n13712 & n34113 ;
  assign n34115 = n34114 ^ n27163 ^ 1'b0 ;
  assign n34116 = n32955 ^ n16090 ^ 1'b0 ;
  assign n34117 = n4049 ^ n472 ^ 1'b0 ;
  assign n34118 = n34117 ^ n14555 ^ 1'b0 ;
  assign n34119 = n22566 ^ n1255 ^ n305 ;
  assign n34120 = ( n10206 & n19486 ) | ( n10206 & n34119 ) | ( n19486 & n34119 ) ;
  assign n34121 = ( n13764 & n24306 ) | ( n13764 & ~n27706 ) | ( n24306 & ~n27706 ) ;
  assign n34122 = ( n12576 & n28432 ) | ( n12576 & n34121 ) | ( n28432 & n34121 ) ;
  assign n34123 = n8375 | n33415 ;
  assign n34124 = n14586 ^ n11914 ^ 1'b0 ;
  assign n34125 = ( n24258 & ~n25464 ) | ( n24258 & n29428 ) | ( ~n25464 & n29428 ) ;
  assign n34126 = n16752 ^ n8474 ^ 1'b0 ;
  assign n34131 = n8570 | n22680 ;
  assign n34132 = n34131 ^ n1488 ^ 1'b0 ;
  assign n34127 = n4542 ^ n2816 ^ 1'b0 ;
  assign n34128 = ~n11941 & n34127 ;
  assign n34129 = n8179 ^ n7626 ^ n3391 ;
  assign n34130 = n34128 & ~n34129 ;
  assign n34133 = n34132 ^ n34130 ^ 1'b0 ;
  assign n34134 = n29354 & ~n34133 ;
  assign n34135 = ~n12080 & n31769 ;
  assign n34136 = ~n3281 & n34135 ;
  assign n34137 = n34136 ^ n20605 ^ n858 ;
  assign n34138 = ~n7027 & n8119 ;
  assign n34139 = ( ~n8025 & n34137 ) | ( ~n8025 & n34138 ) | ( n34137 & n34138 ) ;
  assign n34140 = n28932 ^ n26637 ^ 1'b0 ;
  assign n34142 = n3016 ^ n2955 ^ 1'b0 ;
  assign n34143 = n26035 & n34142 ;
  assign n34141 = ~n4160 & n23089 ;
  assign n34144 = n34143 ^ n34141 ^ 1'b0 ;
  assign n34145 = n12940 & ~n25845 ;
  assign n34146 = n34145 ^ n20193 ^ 1'b0 ;
  assign n34147 = n33007 ^ n15449 ^ n9326 ;
  assign n34148 = ~n11813 & n34147 ;
  assign n34152 = n1595 | n20009 ;
  assign n34149 = n538 & ~n7559 ;
  assign n34150 = n18449 | n34149 ;
  assign n34151 = n24872 | n34150 ;
  assign n34153 = n34152 ^ n34151 ^ n9477 ;
  assign n34154 = n17231 ^ n8025 ^ 1'b0 ;
  assign n34155 = n34154 ^ n17007 ^ 1'b0 ;
  assign n34156 = n19649 & n32159 ;
  assign n34157 = n34156 ^ n14086 ^ 1'b0 ;
  assign n34158 = n8725 & n34157 ;
  assign n34159 = n26463 ^ n19729 ^ 1'b0 ;
  assign n34160 = n24526 & ~n34159 ;
  assign n34161 = n345 & ~n535 ;
  assign n34162 = ~n345 & n34161 ;
  assign n34163 = n1833 | n3903 ;
  assign n34164 = n3903 & ~n34163 ;
  assign n34165 = n1289 & ~n2441 ;
  assign n34166 = ~n1289 & n34165 ;
  assign n34167 = n34164 | n34166 ;
  assign n34168 = n34164 & ~n34167 ;
  assign n34169 = n34162 & ~n34168 ;
  assign n34170 = ~n23276 & n34169 ;
  assign n34171 = ~n1763 & n5584 ;
  assign n34172 = ~n5584 & n34171 ;
  assign n34173 = n1733 & n34172 ;
  assign n34174 = ~n26187 & n34173 ;
  assign n34175 = ~n15996 & n34174 ;
  assign n34176 = n6246 | n34175 ;
  assign n34177 = n11222 & ~n34176 ;
  assign n34178 = n6459 | n34177 ;
  assign n34179 = n34177 & ~n34178 ;
  assign n34180 = n8411 & ~n34179 ;
  assign n34181 = n34170 & n34180 ;
  assign n34182 = n8004 & ~n34181 ;
  assign n34183 = n34182 ^ n16403 ^ 1'b0 ;
  assign n34184 = n1132 | n1702 ;
  assign n34185 = n1702 & ~n34184 ;
  assign n34186 = n1281 & ~n1514 ;
  assign n34187 = n1514 & n34186 ;
  assign n34188 = n1395 | n34187 ;
  assign n34189 = n34187 & ~n34188 ;
  assign n34190 = n4100 & ~n34189 ;
  assign n34191 = ~n1244 & n34190 ;
  assign n34192 = n34185 & n34191 ;
  assign n34193 = n14982 | n34192 ;
  assign n34194 = n34183 & ~n34193 ;
  assign n34196 = n26909 ^ n13473 ^ 1'b0 ;
  assign n34197 = ( n13223 & n16004 ) | ( n13223 & ~n34196 ) | ( n16004 & ~n34196 ) ;
  assign n34195 = ~n12518 & n20555 ;
  assign n34198 = n34197 ^ n34195 ^ 1'b0 ;
  assign n34199 = n34198 ^ n19178 ^ 1'b0 ;
  assign n34200 = n3786 & ~n11337 ;
  assign n34201 = n29123 | n34200 ;
  assign n34202 = n34201 ^ n26210 ^ 1'b0 ;
  assign n34203 = ( n6005 & n10237 ) | ( n6005 & n34202 ) | ( n10237 & n34202 ) ;
  assign n34204 = n18294 ^ n6844 ^ 1'b0 ;
  assign n34205 = ~n3320 & n34204 ;
  assign n34206 = n20975 ^ n279 ^ 1'b0 ;
  assign n34207 = n3384 | n34206 ;
  assign n34208 = n30201 | n34207 ;
  assign n34209 = n7101 ^ n4779 ^ 1'b0 ;
  assign n34210 = n32690 ^ n5177 ^ 1'b0 ;
  assign n34211 = ~n9502 & n19543 ;
  assign n34212 = n6388 | n13046 ;
  assign n34213 = n7154 & ~n34212 ;
  assign n34214 = n16933 & ~n34213 ;
  assign n34215 = n34211 & n34214 ;
  assign n34216 = n5404 & n34215 ;
  assign n34217 = ~n18322 & n33772 ;
  assign n34218 = n21452 & n34217 ;
  assign n34219 = n34218 ^ x124 ^ 1'b0 ;
  assign n34220 = n6565 | n23895 ;
  assign n34221 = n26671 & ~n34220 ;
  assign n34222 = n33452 ^ n18123 ^ 1'b0 ;
  assign n34223 = n17451 ^ n11721 ^ 1'b0 ;
  assign n34224 = n1281 & ~n34223 ;
  assign n34225 = n7418 | n10049 ;
  assign n34226 = n34225 ^ n3316 ^ 1'b0 ;
  assign n34227 = n33339 ^ n6096 ^ n2272 ;
  assign n34228 = n34227 ^ n2860 ^ 1'b0 ;
  assign n34229 = ~n6145 & n34228 ;
  assign n34230 = n26431 ^ n6818 ^ 1'b0 ;
  assign n34231 = n3334 | n6445 ;
  assign n34232 = n4872 & ~n34231 ;
  assign n34233 = ~n13685 & n34232 ;
  assign n34234 = n30945 ^ n5102 ^ n1666 ;
  assign n34235 = n18294 ^ n17963 ^ 1'b0 ;
  assign n34236 = ( ~n1943 & n2727 ) | ( ~n1943 & n6930 ) | ( n2727 & n6930 ) ;
  assign n34237 = n34236 ^ n25519 ^ 1'b0 ;
  assign n34238 = n3096 & ~n23924 ;
  assign n34239 = n7769 & n34238 ;
  assign n34240 = n18917 ^ n17459 ^ 1'b0 ;
  assign n34243 = n31926 ^ n2733 ^ 1'b0 ;
  assign n34244 = n15264 | n34243 ;
  assign n34241 = ~n4246 & n23151 ;
  assign n34242 = n10842 & n34241 ;
  assign n34245 = n34244 ^ n34242 ^ 1'b0 ;
  assign n34246 = n34240 & n34245 ;
  assign n34247 = n3581 & n7559 ;
  assign n34248 = n1453 & n34247 ;
  assign n34249 = n2727 | n34248 ;
  assign n34250 = n34249 ^ n6703 ^ 1'b0 ;
  assign n34251 = n17013 | n34250 ;
  assign n34252 = n34251 ^ n12707 ^ 1'b0 ;
  assign n34253 = n21817 | n34252 ;
  assign n34254 = n34253 ^ n18696 ^ 1'b0 ;
  assign n34255 = n12208 ^ n8317 ^ 1'b0 ;
  assign n34256 = n13117 & ~n34255 ;
  assign n34257 = ~x174 & n18171 ;
  assign n34258 = n25905 ^ n19601 ^ n14995 ;
  assign n34259 = n34257 & n34258 ;
  assign n34260 = ( n4894 & ~n5720 ) | ( n4894 & n12720 ) | ( ~n5720 & n12720 ) ;
  assign n34261 = n14077 ^ n6151 ^ 1'b0 ;
  assign n34262 = n3122 | n34261 ;
  assign n34263 = ~n21286 & n34262 ;
  assign n34264 = n25909 & n34263 ;
  assign n34265 = n34260 | n34264 ;
  assign n34266 = n13640 | n28996 ;
  assign n34267 = n17300 & ~n34266 ;
  assign n34268 = ~n20448 & n30871 ;
  assign n34269 = ( ~n704 & n2073 ) | ( ~n704 & n24124 ) | ( n2073 & n24124 ) ;
  assign n34270 = n506 & n34269 ;
  assign n34271 = n34270 ^ n4734 ^ 1'b0 ;
  assign n34272 = ( n6590 & ~n29207 ) | ( n6590 & n32045 ) | ( ~n29207 & n32045 ) ;
  assign n34273 = n34272 ^ n28553 ^ 1'b0 ;
  assign n34274 = n25609 | n34273 ;
  assign n34275 = n31901 | n33347 ;
  assign n34276 = n3330 ^ x73 ^ 1'b0 ;
  assign n34277 = n34276 ^ n32339 ^ n4330 ;
  assign n34278 = n24151 ^ n14918 ^ n10794 ;
  assign n34279 = n16283 & n32363 ;
  assign n34280 = n33506 & n34279 ;
  assign n34281 = n3088 & n34280 ;
  assign n34282 = n12070 & n27777 ;
  assign n34283 = n24661 ^ n17226 ^ 1'b0 ;
  assign n34284 = n16373 & n34283 ;
  assign n34285 = ~n33878 & n34284 ;
  assign n34286 = n20523 ^ n9771 ^ 1'b0 ;
  assign n34287 = n34286 ^ n15468 ^ 1'b0 ;
  assign n34288 = n2243 & n34287 ;
  assign n34290 = n2107 & ~n5671 ;
  assign n34291 = n7306 ^ n2922 ^ n1147 ;
  assign n34292 = ~n34290 & n34291 ;
  assign n34289 = n4555 | n25124 ;
  assign n34293 = n34292 ^ n34289 ^ 1'b0 ;
  assign n34294 = n10785 & ~n28891 ;
  assign n34295 = ~n31724 & n33639 ;
  assign n34296 = n34295 ^ n33720 ^ 1'b0 ;
  assign n34297 = ~n34294 & n34296 ;
  assign n34298 = ( n1382 & n7908 ) | ( n1382 & ~n28107 ) | ( n7908 & ~n28107 ) ;
  assign n34299 = ( n3783 & n15629 ) | ( n3783 & n23628 ) | ( n15629 & n23628 ) ;
  assign n34300 = n11813 | n11893 ;
  assign n34301 = n13785 | n34300 ;
  assign n34302 = ( n363 & n29534 ) | ( n363 & n34301 ) | ( n29534 & n34301 ) ;
  assign n34303 = n34302 ^ n33129 ^ 1'b0 ;
  assign n34304 = n23877 & ~n34303 ;
  assign n34305 = n6075 & n6419 ;
  assign n34306 = n8949 & n32442 ;
  assign n34307 = n34306 ^ n7559 ^ 1'b0 ;
  assign n34308 = n9268 ^ n8038 ^ 1'b0 ;
  assign n34309 = n16931 ^ n3396 ^ 1'b0 ;
  assign n34310 = ( n961 & ~n8963 ) | ( n961 & n27296 ) | ( ~n8963 & n27296 ) ;
  assign n34312 = ~n271 & n1158 ;
  assign n34311 = n21964 ^ n20293 ^ 1'b0 ;
  assign n34313 = n34312 ^ n34311 ^ n7118 ;
  assign n34314 = n441 & n34313 ;
  assign n34315 = ~n34310 & n34314 ;
  assign n34316 = n8509 & ~n14576 ;
  assign n34317 = n34316 ^ n29257 ^ 1'b0 ;
  assign n34318 = n15578 ^ n9978 ^ n9694 ;
  assign n34320 = ~n13464 & n34069 ;
  assign n34319 = n23307 | n25063 ;
  assign n34321 = n34320 ^ n34319 ^ 1'b0 ;
  assign n34322 = n21390 ^ n16808 ^ 1'b0 ;
  assign n34323 = n8237 & n34322 ;
  assign n34324 = n19150 ^ n16492 ^ 1'b0 ;
  assign n34325 = n8894 & n24020 ;
  assign n34326 = ~n23490 & n34325 ;
  assign n34327 = ~n11672 & n24856 ;
  assign n34329 = n546 | n17640 ;
  assign n34330 = n34329 ^ n4694 ^ 1'b0 ;
  assign n34328 = ~n2548 & n21938 ;
  assign n34331 = n34330 ^ n34328 ^ 1'b0 ;
  assign n34332 = n34331 ^ n16977 ^ 1'b0 ;
  assign n34333 = n31740 ^ n27198 ^ n6142 ;
  assign n34334 = n14112 & ~n34333 ;
  assign n34335 = n20455 ^ n7762 ^ n3642 ;
  assign n34336 = n34335 ^ n12045 ^ 1'b0 ;
  assign n34337 = n32216 & ~n34079 ;
  assign n34338 = n15351 & ~n34337 ;
  assign n34339 = n6607 & ~n34338 ;
  assign n34340 = n5905 & n14951 ;
  assign n34341 = n11507 & n34340 ;
  assign n34342 = ( n10352 & n12435 ) | ( n10352 & ~n16227 ) | ( n12435 & ~n16227 ) ;
  assign n34343 = n34342 ^ n21489 ^ 1'b0 ;
  assign n34344 = ~n25676 & n34343 ;
  assign n34345 = ~n33185 & n34260 ;
  assign n34346 = n34345 ^ n9338 ^ 1'b0 ;
  assign n34347 = n6510 & ~n13391 ;
  assign n34348 = n9774 | n34347 ;
  assign n34349 = n23660 & n34348 ;
  assign n34350 = ~n7727 & n34349 ;
  assign n34351 = n34350 ^ n22824 ^ n3826 ;
  assign n34354 = ~n8930 & n13258 ;
  assign n34355 = n34354 ^ n30274 ^ 1'b0 ;
  assign n34352 = n7852 ^ n6284 ^ 1'b0 ;
  assign n34353 = n34352 ^ n19019 ^ n8572 ;
  assign n34356 = n34355 ^ n34353 ^ 1'b0 ;
  assign n34357 = n2425 ^ n1618 ^ 1'b0 ;
  assign n34358 = n6170 & ~n34357 ;
  assign n34359 = n17601 | n34358 ;
  assign n34360 = n34356 & ~n34359 ;
  assign n34361 = ~n4081 & n7627 ;
  assign n34366 = ( n15677 & ~n17127 ) | ( n15677 & n31949 ) | ( ~n17127 & n31949 ) ;
  assign n34362 = n6218 ^ n2305 ^ 1'b0 ;
  assign n34363 = n14016 & ~n34362 ;
  assign n34364 = n7805 & n20561 ;
  assign n34365 = ~n34363 & n34364 ;
  assign n34367 = n34366 ^ n34365 ^ 1'b0 ;
  assign n34368 = ( n8179 & n34361 ) | ( n8179 & ~n34367 ) | ( n34361 & ~n34367 ) ;
  assign n34370 = n3078 | n8707 ;
  assign n34371 = n34370 ^ n11167 ^ 1'b0 ;
  assign n34369 = n2587 & ~n28388 ;
  assign n34372 = n34371 ^ n34369 ^ 1'b0 ;
  assign n34373 = ~n21702 & n31611 ;
  assign n34374 = n34373 ^ n7844 ^ 1'b0 ;
  assign n34375 = n20685 ^ n734 ^ 1'b0 ;
  assign n34376 = n34375 ^ n17798 ^ n2146 ;
  assign n34377 = n1186 & n19895 ;
  assign n34378 = n34377 ^ n25343 ^ n23199 ;
  assign n34379 = n11203 ^ n5330 ^ n1081 ;
  assign n34380 = ~n2296 & n34379 ;
  assign n34381 = n12845 & ~n33002 ;
  assign n34382 = n34381 ^ n20960 ^ 1'b0 ;
  assign n34383 = n6493 & n8573 ;
  assign n34384 = ~n3216 & n7745 ;
  assign n34385 = n31386 & n34384 ;
  assign n34386 = n34383 & n34385 ;
  assign n34387 = n5477 ^ n4774 ^ n608 ;
  assign n34388 = ( n11729 & n25203 ) | ( n11729 & ~n34387 ) | ( n25203 & ~n34387 ) ;
  assign n34389 = n15758 ^ n8777 ^ 1'b0 ;
  assign n34390 = ( n11314 & ~n29901 ) | ( n11314 & n34389 ) | ( ~n29901 & n34389 ) ;
  assign n34391 = n8787 & n23783 ;
  assign n34392 = n5300 & n34391 ;
  assign n34393 = n29673 ^ n3967 ^ 1'b0 ;
  assign n34394 = n30870 & n34393 ;
  assign n34395 = n22067 ^ n14382 ^ 1'b0 ;
  assign n34396 = ~n34394 & n34395 ;
  assign n34397 = n2971 & ~n5103 ;
  assign n34398 = n12845 ^ n7315 ^ n2727 ;
  assign n34399 = n34397 & ~n34398 ;
  assign n34400 = n13002 ^ n6607 ^ 1'b0 ;
  assign n34401 = n29202 & ~n34400 ;
  assign n34402 = n8998 ^ n2925 ^ 1'b0 ;
  assign n34403 = n22062 ^ n8829 ^ 1'b0 ;
  assign n34404 = n8655 & ~n34403 ;
  assign n34405 = n34404 ^ n31753 ^ n4137 ;
  assign n34406 = ~n5568 & n18140 ;
  assign n34407 = ~n2905 & n34406 ;
  assign n34408 = n26362 ^ n13764 ^ 1'b0 ;
  assign n34409 = n14394 & n34408 ;
  assign n34410 = n5481 | n7952 ;
  assign n34411 = n14961 | n34410 ;
  assign n34412 = n5233 & ~n34411 ;
  assign n34413 = n21467 ^ n17891 ^ 1'b0 ;
  assign n34414 = ~n13873 & n18254 ;
  assign n34415 = n12756 | n34414 ;
  assign n34416 = ( ~n2843 & n17477 ) | ( ~n2843 & n34138 ) | ( n17477 & n34138 ) ;
  assign n34417 = n11258 | n26545 ;
  assign n34418 = n1024 & ~n10565 ;
  assign n34419 = n22092 ^ n16653 ^ n9371 ;
  assign n34420 = n18061 & ~n34419 ;
  assign n34421 = n34420 ^ n13608 ^ 1'b0 ;
  assign n34422 = n34421 ^ n7184 ^ 1'b0 ;
  assign n34423 = n28713 | n34422 ;
  assign n34424 = ( n2950 & n13404 ) | ( n2950 & ~n29493 ) | ( n13404 & ~n29493 ) ;
  assign n34425 = n2630 & n6556 ;
  assign n34426 = ~n6298 & n18694 ;
  assign n34427 = n34426 ^ n15378 ^ 1'b0 ;
  assign n34428 = n18516 ^ n13019 ^ n6440 ;
  assign n34429 = n9706 ^ n5740 ^ 1'b0 ;
  assign n34430 = n34428 & n34429 ;
  assign n34431 = n12629 & n32860 ;
  assign n34432 = n33803 & n34431 ;
  assign n34433 = ~n8688 & n28548 ;
  assign n34434 = n22166 ^ n17853 ^ 1'b0 ;
  assign n34435 = n20185 ^ n3257 ^ 1'b0 ;
  assign n34436 = n530 & ~n34435 ;
  assign n34437 = n16005 ^ n2608 ^ 1'b0 ;
  assign n34438 = n15851 | n34437 ;
  assign n34439 = ~n20269 & n34438 ;
  assign n34440 = n34439 ^ n24858 ^ 1'b0 ;
  assign n34441 = n17694 & n34440 ;
  assign n34442 = ~n20876 & n34441 ;
  assign n34444 = n13723 ^ n11335 ^ 1'b0 ;
  assign n34445 = n6448 & ~n34444 ;
  assign n34443 = n4711 & n12790 ;
  assign n34446 = n34445 ^ n34443 ^ 1'b0 ;
  assign n34447 = n3675 | n9932 ;
  assign n34448 = n34447 ^ n3600 ^ 1'b0 ;
  assign n34449 = n10035 & n25193 ;
  assign n34450 = ~n559 & n34449 ;
  assign n34451 = n5532 ^ n790 ^ 1'b0 ;
  assign n34452 = n259 & ~n10707 ;
  assign n34453 = n34452 ^ n6724 ^ 1'b0 ;
  assign n34454 = ~n34451 & n34453 ;
  assign n34455 = ~n11641 & n34454 ;
  assign n34456 = ~n261 & n427 ;
  assign n34457 = n34456 ^ n1920 ^ 1'b0 ;
  assign n34458 = n3448 & ~n34457 ;
  assign n34459 = n9382 & n17530 ;
  assign n34460 = ~n12528 & n34459 ;
  assign n34461 = n7915 & ~n32130 ;
  assign n34462 = n24176 ^ n18415 ^ n702 ;
  assign n34463 = n5716 | n16553 ;
  assign n34464 = n34463 ^ n8978 ^ 1'b0 ;
  assign n34465 = ~x187 & n33741 ;
  assign n34466 = ( n5399 & n16749 ) | ( n5399 & n23617 ) | ( n16749 & n23617 ) ;
  assign n34467 = x2 & n34466 ;
  assign n34468 = ~n8848 & n34467 ;
  assign n34469 = n12903 ^ n1271 ^ 1'b0 ;
  assign n34470 = n15922 | n34469 ;
  assign n34471 = n2543 & ~n16706 ;
  assign n34472 = n34471 ^ n16338 ^ 1'b0 ;
  assign n34473 = n34472 ^ n16680 ^ n10360 ;
  assign n34474 = n12546 | n34473 ;
  assign n34475 = ( ~n1925 & n26986 ) | ( ~n1925 & n34474 ) | ( n26986 & n34474 ) ;
  assign n34476 = n4991 & ~n20877 ;
  assign n34477 = n34476 ^ n13668 ^ 1'b0 ;
  assign n34478 = n294 | n20203 ;
  assign n34479 = n33724 & ~n34478 ;
  assign n34480 = n16777 ^ n12950 ^ 1'b0 ;
  assign n34482 = n2557 & ~n15378 ;
  assign n34483 = ~n13948 & n34482 ;
  assign n34481 = n7200 | n14607 ;
  assign n34484 = n34483 ^ n34481 ^ 1'b0 ;
  assign n34485 = n5150 & n9880 ;
  assign n34486 = n34485 ^ n20921 ^ 1'b0 ;
  assign n34487 = n3938 & n26792 ;
  assign n34488 = n34487 ^ n30516 ^ 1'b0 ;
  assign n34489 = n20004 ^ n12547 ^ 1'b0 ;
  assign n34490 = n12359 & ~n21286 ;
  assign n34492 = n1493 & ~n10601 ;
  assign n34491 = ( ~n1232 & n9416 ) | ( ~n1232 & n33974 ) | ( n9416 & n33974 ) ;
  assign n34493 = n34492 ^ n34491 ^ n23413 ;
  assign n34495 = n21643 ^ n19019 ^ 1'b0 ;
  assign n34494 = n10974 & n15398 ;
  assign n34496 = n34495 ^ n34494 ^ 1'b0 ;
  assign n34497 = n24855 ^ n20463 ^ n4074 ;
  assign n34498 = n33361 ^ n14636 ^ 1'b0 ;
  assign n34499 = n34497 & n34498 ;
  assign n34500 = n15508 ^ n12178 ^ 1'b0 ;
  assign n34501 = n12002 & ~n34500 ;
  assign n34502 = n9334 ^ n8232 ^ n1473 ;
  assign n34503 = n1824 & n10158 ;
  assign n34504 = n34152 ^ n2704 ^ 1'b0 ;
  assign n34505 = n34503 & n34504 ;
  assign n34506 = n34505 ^ n18999 ^ 1'b0 ;
  assign n34507 = n34502 | n34506 ;
  assign n34508 = n1342 | n13172 ;
  assign n34509 = n446 & ~n29982 ;
  assign n34510 = n34509 ^ n13355 ^ 1'b0 ;
  assign n34512 = n10243 | n12591 ;
  assign n34511 = ~n10870 & n29837 ;
  assign n34513 = n34512 ^ n34511 ^ 1'b0 ;
  assign n34514 = n7047 & n8859 ;
  assign n34515 = ~n2682 & n34514 ;
  assign n34516 = n34515 ^ n30434 ^ 1'b0 ;
  assign n34517 = n8375 | n31552 ;
  assign n34518 = n34517 ^ n21381 ^ 1'b0 ;
  assign n34520 = n3778 | n6795 ;
  assign n34521 = n11519 | n34520 ;
  assign n34519 = n12805 & n19759 ;
  assign n34522 = n34521 ^ n34519 ^ 1'b0 ;
  assign n34523 = n34522 ^ n17366 ^ n10594 ;
  assign n34524 = n4015 | n16363 ;
  assign n34525 = x102 | n34524 ;
  assign n34526 = n26137 ^ n17772 ^ n991 ;
  assign n34527 = n34526 ^ x42 ^ 1'b0 ;
  assign n34528 = ( n23307 & n34525 ) | ( n23307 & ~n34527 ) | ( n34525 & ~n34527 ) ;
  assign n34529 = ( n3257 & n4895 ) | ( n3257 & ~n25989 ) | ( n4895 & ~n25989 ) ;
  assign n34530 = ( n9249 & ~n34389 ) | ( n9249 & n34529 ) | ( ~n34389 & n34529 ) ;
  assign n34531 = ( n1259 & n2652 ) | ( n1259 & n12685 ) | ( n2652 & n12685 ) ;
  assign n34532 = ~n642 & n34531 ;
  assign n34533 = n24911 ^ n16570 ^ 1'b0 ;
  assign n34534 = n5129 ^ n3456 ^ 1'b0 ;
  assign n34535 = n13453 | n30679 ;
  assign n34536 = n31214 ^ n12041 ^ 1'b0 ;
  assign n34537 = n29322 | n34536 ;
  assign n34538 = n7411 ^ n1450 ^ 1'b0 ;
  assign n34539 = n28107 | n34538 ;
  assign n34540 = n34539 ^ n773 ^ 1'b0 ;
  assign n34541 = n12379 & n34540 ;
  assign n34542 = ~n27852 & n34541 ;
  assign n34543 = ~n2351 & n34542 ;
  assign n34544 = n10757 & n15588 ;
  assign n34545 = ~n2081 & n34544 ;
  assign n34546 = n34545 ^ n25821 ^ 1'b0 ;
  assign n34547 = n18562 & n34546 ;
  assign n34548 = n22855 ^ n18997 ^ 1'b0 ;
  assign n34553 = n8294 | n10434 ;
  assign n34554 = n18213 & ~n34553 ;
  assign n34549 = n11230 | n21124 ;
  assign n34550 = n4364 | n34549 ;
  assign n34551 = n2488 & n34550 ;
  assign n34552 = n34551 ^ n10344 ^ 1'b0 ;
  assign n34555 = n34554 ^ n34552 ^ 1'b0 ;
  assign n34556 = ( n1362 & n4876 ) | ( n1362 & n23390 ) | ( n4876 & n23390 ) ;
  assign n34557 = n16324 & n34556 ;
  assign n34558 = n27185 & ~n34557 ;
  assign n34559 = n15657 ^ n5145 ^ 1'b0 ;
  assign n34560 = n8118 | n9442 ;
  assign n34561 = n34560 ^ n5115 ^ 1'b0 ;
  assign n34562 = ~n15679 & n34561 ;
  assign n34563 = n2386 & n34562 ;
  assign n34564 = n11300 ^ n5869 ^ 1'b0 ;
  assign n34565 = ~n34563 & n34564 ;
  assign n34566 = n15441 & ~n21941 ;
  assign n34567 = n34566 ^ n4967 ^ 1'b0 ;
  assign n34568 = ~n3668 & n7245 ;
  assign n34569 = n5896 & ~n13787 ;
  assign n34570 = n12530 ^ n8588 ^ 1'b0 ;
  assign n34571 = n2034 ^ n555 ^ 1'b0 ;
  assign n34572 = ~n18413 & n34571 ;
  assign n34573 = n34572 ^ n4900 ^ 1'b0 ;
  assign n34574 = n27642 ^ n17091 ^ 1'b0 ;
  assign n34575 = n3473 & ~n34574 ;
  assign n34576 = ~n7660 & n34575 ;
  assign n34577 = n12660 ^ n5043 ^ 1'b0 ;
  assign n34578 = n2704 & ~n34577 ;
  assign n34579 = n21988 ^ n13573 ^ 1'b0 ;
  assign n34580 = n34578 | n34579 ;
  assign n34581 = n34580 ^ n24458 ^ 1'b0 ;
  assign n34582 = n23053 ^ n6704 ^ 1'b0 ;
  assign n34583 = ( n1753 & n32901 ) | ( n1753 & ~n34582 ) | ( n32901 & ~n34582 ) ;
  assign n34584 = n31662 ^ n7721 ^ 1'b0 ;
  assign n34585 = n34584 ^ n10123 ^ n2507 ;
  assign n34586 = n8352 & n14113 ;
  assign n34587 = n34585 & n34586 ;
  assign n34588 = n3248 ^ n2659 ^ 1'b0 ;
  assign n34589 = ~n11804 & n34588 ;
  assign n34590 = ~n16285 & n34589 ;
  assign n34591 = n5422 & ~n17523 ;
  assign n34592 = ( ~n1071 & n10828 ) | ( ~n1071 & n34591 ) | ( n10828 & n34591 ) ;
  assign n34593 = ( n12810 & ~n12869 ) | ( n12810 & n34592 ) | ( ~n12869 & n34592 ) ;
  assign n34594 = ~n17669 & n20508 ;
  assign n34595 = n34594 ^ n28480 ^ 1'b0 ;
  assign n34596 = n30690 ^ n11732 ^ n7627 ;
  assign n34597 = n34596 ^ n18327 ^ n3027 ;
  assign n34598 = n13677 & ~n20623 ;
  assign n34599 = n26886 & n34598 ;
  assign n34600 = ( n7372 & ~n20625 ) | ( n7372 & n32758 ) | ( ~n20625 & n32758 ) ;
  assign n34601 = n30809 ^ n300 ^ 1'b0 ;
  assign n34602 = n34600 | n34601 ;
  assign n34603 = n7429 | n13134 ;
  assign n34604 = n34603 ^ n671 ^ 1'b0 ;
  assign n34605 = n12788 ^ n8776 ^ n1674 ;
  assign n34606 = n18034 | n34605 ;
  assign n34608 = n1875 ^ n1395 ^ 1'b0 ;
  assign n34609 = n9048 & ~n34608 ;
  assign n34610 = ~n25598 & n34609 ;
  assign n34607 = n32081 ^ n2726 ^ 1'b0 ;
  assign n34611 = n34610 ^ n34607 ^ 1'b0 ;
  assign n34612 = n12265 ^ n11726 ^ n5073 ;
  assign n34615 = n22666 ^ n9484 ^ 1'b0 ;
  assign n34613 = n11028 ^ x31 ^ 1'b0 ;
  assign n34614 = n30859 & n34613 ;
  assign n34616 = n34615 ^ n34614 ^ 1'b0 ;
  assign n34617 = n5163 | n18559 ;
  assign n34618 = n34617 ^ n5418 ^ 1'b0 ;
  assign n34619 = n3018 | n21147 ;
  assign n34620 = ~n28310 & n34619 ;
  assign n34621 = n18464 ^ n9442 ^ 1'b0 ;
  assign n34622 = n22214 & ~n34621 ;
  assign n34623 = n3968 ^ n558 ^ 1'b0 ;
  assign n34624 = n34623 ^ n16889 ^ n13744 ;
  assign n34625 = n31261 ^ n6214 ^ n3056 ;
  assign n34626 = n16783 ^ n6670 ^ 1'b0 ;
  assign n34627 = n32804 ^ n32543 ^ 1'b0 ;
  assign n34628 = ~n10215 & n27127 ;
  assign n34629 = n34628 ^ n21626 ^ 1'b0 ;
  assign n34631 = n2504 | n15774 ;
  assign n34632 = n34631 ^ n2632 ^ 1'b0 ;
  assign n34630 = n17184 & ~n28585 ;
  assign n34633 = n34632 ^ n34630 ^ 1'b0 ;
  assign n34634 = n12937 ^ n5477 ^ 1'b0 ;
  assign n34635 = n1102 & ~n34634 ;
  assign n34636 = n34635 ^ n15911 ^ 1'b0 ;
  assign n34637 = n28057 ^ n11282 ^ 1'b0 ;
  assign n34638 = n22692 ^ n17979 ^ n9556 ;
  assign n34639 = n21660 | n25911 ;
  assign n34640 = ( ~n15027 & n22020 ) | ( ~n15027 & n34639 ) | ( n22020 & n34639 ) ;
  assign n34641 = n34640 ^ n3116 ^ 1'b0 ;
  assign n34642 = n14709 ^ n7593 ^ 1'b0 ;
  assign n34643 = n12981 | n34642 ;
  assign n34644 = n7297 ^ n3332 ^ 1'b0 ;
  assign n34645 = ~n10473 & n34644 ;
  assign n34646 = n7914 & n34645 ;
  assign n34647 = n34646 ^ n25795 ^ 1'b0 ;
  assign n34648 = n14294 & n15430 ;
  assign n34649 = n34648 ^ n8612 ^ 1'b0 ;
  assign n34650 = n22636 & ~n33232 ;
  assign n34651 = n34649 & n34650 ;
  assign n34652 = n10648 & ~n34651 ;
  assign n34654 = n8115 | n13423 ;
  assign n34655 = n591 & n34654 ;
  assign n34653 = x80 & n14801 ;
  assign n34656 = n34655 ^ n34653 ^ 1'b0 ;
  assign n34657 = n6251 & ~n29753 ;
  assign n34658 = n34656 & n34657 ;
  assign n34659 = n9159 & ~n12384 ;
  assign n34660 = n34659 ^ n16772 ^ 1'b0 ;
  assign n34661 = n5776 & n34660 ;
  assign n34662 = n9545 | n15551 ;
  assign n34665 = ~n18404 & n19209 ;
  assign n34664 = n19635 ^ x71 ^ 1'b0 ;
  assign n34663 = ~n12651 & n27109 ;
  assign n34666 = n34665 ^ n34664 ^ n34663 ;
  assign n34667 = n6705 & n7122 ;
  assign n34668 = n28256 ^ n17178 ^ 1'b0 ;
  assign n34669 = n34667 & ~n34668 ;
  assign n34670 = n3453 | n13126 ;
  assign n34671 = n34670 ^ n552 ^ 1'b0 ;
  assign n34672 = n23360 ^ n5968 ^ n915 ;
  assign n34673 = ( ~n6023 & n8496 ) | ( ~n6023 & n32260 ) | ( n8496 & n32260 ) ;
  assign n34674 = n18429 & ~n18802 ;
  assign n34675 = n34674 ^ n24234 ^ n21743 ;
  assign n34676 = ( n23373 & n34673 ) | ( n23373 & n34675 ) | ( n34673 & n34675 ) ;
  assign n34677 = ( n3445 & n6060 ) | ( n3445 & n15582 ) | ( n6060 & n15582 ) ;
  assign n34678 = n18277 & n19719 ;
  assign n34679 = ~n5807 & n34678 ;
  assign n34680 = n34679 ^ n29261 ^ 1'b0 ;
  assign n34681 = n485 & ~n34680 ;
  assign n34682 = n19255 & n34681 ;
  assign n34683 = n34682 ^ n6642 ^ 1'b0 ;
  assign n34684 = ( n3061 & n34677 ) | ( n3061 & ~n34683 ) | ( n34677 & ~n34683 ) ;
  assign n34685 = ~n22680 & n34684 ;
  assign n34686 = n9831 ^ n5797 ^ n1540 ;
  assign n34687 = ( n13705 & n15585 ) | ( n13705 & ~n34686 ) | ( n15585 & ~n34686 ) ;
  assign n34688 = x61 | n3884 ;
  assign n34689 = n8404 & n34688 ;
  assign n34690 = n14858 ^ n6541 ^ 1'b0 ;
  assign n34691 = n7294 & ~n30922 ;
  assign n34692 = n34691 ^ n14028 ^ 1'b0 ;
  assign n34693 = n6290 & n34692 ;
  assign n34694 = n34693 ^ n30213 ^ 1'b0 ;
  assign n34695 = ~n14396 & n34694 ;
  assign n34696 = ~n2438 & n14329 ;
  assign n34697 = n5255 & n34696 ;
  assign n34698 = ( n867 & ~n34695 ) | ( n867 & n34697 ) | ( ~n34695 & n34697 ) ;
  assign n34699 = n34698 ^ n28789 ^ 1'b0 ;
  assign n34700 = n34045 ^ n5514 ^ 1'b0 ;
  assign n34701 = n9658 ^ n5103 ^ 1'b0 ;
  assign n34702 = n3480 & ~n34701 ;
  assign n34703 = ( ~n3554 & n11597 ) | ( ~n3554 & n34702 ) | ( n11597 & n34702 ) ;
  assign n34704 = n5373 & n31256 ;
  assign n34705 = n34703 | n34704 ;
  assign n34706 = n8039 | n11870 ;
  assign n34707 = n10558 | n34706 ;
  assign n34708 = n34707 ^ n28648 ^ 1'b0 ;
  assign n34709 = n9222 & ~n11499 ;
  assign n34710 = ( n11261 & n28677 ) | ( n11261 & n34709 ) | ( n28677 & n34709 ) ;
  assign n34712 = n13750 ^ n11011 ^ 1'b0 ;
  assign n34713 = n10123 & n34712 ;
  assign n34711 = n12368 & n24298 ;
  assign n34714 = n34713 ^ n34711 ^ n29567 ;
  assign n34715 = n20119 ^ n16764 ^ 1'b0 ;
  assign n34716 = n26524 ^ n8440 ^ 1'b0 ;
  assign n34717 = n8119 | n30845 ;
  assign n34718 = n14092 | n34717 ;
  assign n34719 = n34718 ^ n27167 ^ n10258 ;
  assign n34720 = n1701 ^ n933 ^ 1'b0 ;
  assign n34721 = n12845 & ~n34720 ;
  assign n34722 = n34719 & n34721 ;
  assign n34723 = n14732 ^ x9 ^ 1'b0 ;
  assign n34724 = n17290 | n34723 ;
  assign n34725 = n14976 & ~n19937 ;
  assign n34726 = n10261 | n12162 ;
  assign n34727 = n34725 & ~n34726 ;
  assign n34728 = n2826 | n34727 ;
  assign n34729 = n10206 | n34728 ;
  assign n34730 = n2223 & ~n5685 ;
  assign n34731 = n20979 | n31797 ;
  assign n34732 = ~n2751 & n34731 ;
  assign n34738 = n2973 ^ n1671 ^ 1'b0 ;
  assign n34734 = n9817 & ~n10977 ;
  assign n34735 = n15244 & n34734 ;
  assign n34733 = n17143 ^ n16953 ^ 1'b0 ;
  assign n34736 = n34735 ^ n34733 ^ n22340 ;
  assign n34737 = ~n14371 & n34736 ;
  assign n34739 = n34738 ^ n34737 ^ 1'b0 ;
  assign n34740 = n17680 ^ n1210 ^ 1'b0 ;
  assign n34741 = n12981 & n14359 ;
  assign n34742 = n34741 ^ n18612 ^ 1'b0 ;
  assign n34743 = n15178 & n34742 ;
  assign n34744 = n11742 & ~n14487 ;
  assign n34745 = n6379 | n12290 ;
  assign n34746 = n10777 | n34745 ;
  assign n34747 = x48 | n29842 ;
  assign n34748 = n34746 & ~n34747 ;
  assign n34753 = n13883 ^ n1569 ^ 1'b0 ;
  assign n34754 = n8673 & ~n34753 ;
  assign n34750 = n12830 & ~n16307 ;
  assign n34751 = n34750 ^ n9331 ^ 1'b0 ;
  assign n34749 = n9692 & n29702 ;
  assign n34752 = n34751 ^ n34749 ^ 1'b0 ;
  assign n34755 = n34754 ^ n34752 ^ n25531 ;
  assign n34756 = n13671 & n20420 ;
  assign n34757 = n432 & n34756 ;
  assign n34758 = n26195 | n34757 ;
  assign n34759 = n34758 ^ n20080 ^ 1'b0 ;
  assign n34760 = ( n4278 & n7554 ) | ( n4278 & ~n13313 ) | ( n7554 & ~n13313 ) ;
  assign n34761 = n19609 ^ n2993 ^ 1'b0 ;
  assign n34762 = n34760 | n34761 ;
  assign n34763 = n11117 & ~n34762 ;
  assign n34764 = n29170 ^ n8590 ^ 1'b0 ;
  assign n34765 = n674 & n7398 ;
  assign n34766 = n34765 ^ n23902 ^ 1'b0 ;
  assign n34767 = n34764 & n34766 ;
  assign n34768 = n34763 & ~n34767 ;
  assign n34769 = n24196 ^ n2414 ^ 1'b0 ;
  assign n34770 = n7161 ^ n5220 ^ n5040 ;
  assign n34771 = ( n21603 & n33761 ) | ( n21603 & n34770 ) | ( n33761 & n34770 ) ;
  assign n34772 = n24860 ^ n1570 ^ 1'b0 ;
  assign n34773 = n10244 | n22067 ;
  assign n34774 = n34773 ^ n21977 ^ 1'b0 ;
  assign n34775 = ( ~n10411 & n13673 ) | ( ~n10411 & n34774 ) | ( n13673 & n34774 ) ;
  assign n34776 = n15271 | n30113 ;
  assign n34777 = ~x17 & n1709 ;
  assign n34778 = n28920 ^ n19323 ^ 1'b0 ;
  assign n34779 = n429 & ~n1103 ;
  assign n34780 = n31557 & n34779 ;
  assign n34781 = n15390 | n29251 ;
  assign n34782 = n27793 ^ n13992 ^ n12372 ;
  assign n34783 = ~n1989 & n29482 ;
  assign n34784 = n9745 & ~n25890 ;
  assign n34785 = n34784 ^ n13246 ^ n4287 ;
  assign n34786 = n1663 | n28772 ;
  assign n34787 = n34786 ^ n1878 ^ 1'b0 ;
  assign n34788 = ( x205 & n8343 ) | ( x205 & ~n18205 ) | ( n8343 & ~n18205 ) ;
  assign n34789 = n13574 ^ n2979 ^ 1'b0 ;
  assign n34790 = n34789 ^ n12905 ^ n4917 ;
  assign n34791 = n34788 & n34790 ;
  assign n34792 = x16 & n4764 ;
  assign n34793 = n5411 & n34792 ;
  assign n34794 = n12160 | n34793 ;
  assign n34795 = n14080 | n34794 ;
  assign n34796 = n12069 & ~n23147 ;
  assign n34797 = n34796 ^ n3588 ^ 1'b0 ;
  assign n34798 = ~n19548 & n26704 ;
  assign n34799 = n34797 & n34798 ;
  assign n34800 = n34799 ^ n11026 ^ 1'b0 ;
  assign n34801 = n3668 ^ n2618 ^ n1919 ;
  assign n34802 = n8077 | n34801 ;
  assign n34803 = n4137 | n34802 ;
  assign n34804 = n34803 ^ n24713 ^ 1'b0 ;
  assign n34806 = n766 | n16498 ;
  assign n34807 = n30810 & ~n34806 ;
  assign n34805 = n13928 & ~n19067 ;
  assign n34808 = n34807 ^ n34805 ^ 1'b0 ;
  assign n34809 = n16966 ^ n9934 ^ 1'b0 ;
  assign n34810 = n11312 | n34809 ;
  assign n34811 = n18122 & n26375 ;
  assign n34812 = n23337 & n34811 ;
  assign n34813 = ~n24828 & n34812 ;
  assign n34814 = n3683 & ~n26454 ;
  assign n34815 = ( n1517 & n15569 ) | ( n1517 & ~n19055 ) | ( n15569 & ~n19055 ) ;
  assign n34816 = ~n14992 & n34815 ;
  assign n34817 = n4797 & ~n15668 ;
  assign n34818 = n34817 ^ n2690 ^ 1'b0 ;
  assign n34819 = n34818 ^ n16180 ^ 1'b0 ;
  assign n34820 = n744 & ~n34819 ;
  assign n34821 = n5465 & n34820 ;
  assign n34822 = n1925 & n27723 ;
  assign n34823 = n34822 ^ n759 ^ 1'b0 ;
  assign n34826 = n3175 & ~n3451 ;
  assign n34827 = ~n3175 & n34826 ;
  assign n34824 = n471 & ~n1477 ;
  assign n34825 = n34824 ^ n4470 ^ 1'b0 ;
  assign n34828 = n34827 ^ n34825 ^ n6865 ;
  assign n34829 = n6805 ^ n3126 ^ 1'b0 ;
  assign n34830 = n28358 ^ n9317 ^ n6994 ;
  assign n34831 = n34830 ^ n7895 ^ 1'b0 ;
  assign n34832 = n13212 & n34831 ;
  assign n34833 = ( ~n655 & n8033 ) | ( ~n655 & n8848 ) | ( n8033 & n8848 ) ;
  assign n34834 = n17328 ^ n7852 ^ n1590 ;
  assign n34835 = n34833 & n34834 ;
  assign n34836 = n12453 & ~n17967 ;
  assign n34837 = ~n937 & n34836 ;
  assign n34838 = n13572 ^ n10186 ^ 1'b0 ;
  assign n34839 = n16400 & ~n34838 ;
  assign n34840 = n33491 ^ n29737 ^ 1'b0 ;
  assign n34841 = n19157 ^ n18802 ^ 1'b0 ;
  assign n34842 = n23248 & ~n34841 ;
  assign n34843 = n31800 ^ n2276 ^ 1'b0 ;
  assign n34844 = n17917 & n34843 ;
  assign n34845 = n15302 ^ n4035 ^ 1'b0 ;
  assign n34846 = n34844 & ~n34845 ;
  assign n34847 = ( n5288 & ~n12895 ) | ( n5288 & n27278 ) | ( ~n12895 & n27278 ) ;
  assign n34848 = n4977 & n34847 ;
  assign n34849 = n583 ^ n327 ^ 1'b0 ;
  assign n34850 = n18283 ^ n6846 ^ 1'b0 ;
  assign n34851 = n3433 & ~n34850 ;
  assign n34852 = ~n34849 & n34851 ;
  assign n34853 = ~n34848 & n34852 ;
  assign n34854 = n24560 ^ n12089 ^ n5341 ;
  assign n34855 = n34854 ^ n18082 ^ n9891 ;
  assign n34856 = ~n436 & n7714 ;
  assign n34857 = n16895 & n34856 ;
  assign n34858 = n34857 ^ n33370 ^ n27547 ;
  assign n34859 = n34605 ^ n11123 ^ 1'b0 ;
  assign n34860 = ~n3409 & n12718 ;
  assign n34861 = ~n5115 & n34860 ;
  assign n34862 = n8171 & n8438 ;
  assign n34863 = ( ~n7567 & n11805 ) | ( ~n7567 & n28072 ) | ( n11805 & n28072 ) ;
  assign n34864 = n34863 ^ n22653 ^ n10432 ;
  assign n34865 = x168 & n7151 ;
  assign n34866 = n12711 & ~n13706 ;
  assign n34867 = n34866 ^ n13727 ^ 1'b0 ;
  assign n34868 = ( n3907 & n13353 ) | ( n3907 & n34867 ) | ( n13353 & n34867 ) ;
  assign n34869 = ~n6096 & n21032 ;
  assign n34870 = n34869 ^ n7603 ^ 1'b0 ;
  assign n34871 = n19642 | n34870 ;
  assign n34872 = ~n18514 & n21468 ;
  assign n34873 = n34871 & n34872 ;
  assign n34874 = n5223 ^ n894 ^ 1'b0 ;
  assign n34875 = n34873 | n34874 ;
  assign n34876 = n2199 | n26207 ;
  assign n34877 = n34876 ^ n7231 ^ 1'b0 ;
  assign n34878 = n34877 ^ n21144 ^ 1'b0 ;
  assign n34879 = n23387 | n34878 ;
  assign n34881 = n4565 ^ n1013 ^ 1'b0 ;
  assign n34882 = n34881 ^ n18592 ^ n8821 ;
  assign n34880 = n22985 | n29786 ;
  assign n34883 = n34882 ^ n34880 ^ 1'b0 ;
  assign n34884 = n4058 & ~n32634 ;
  assign n34885 = n24994 ^ n5918 ^ 1'b0 ;
  assign n34886 = n10117 & n34885 ;
  assign n34887 = ~n15833 & n34886 ;
  assign n34888 = n15178 & n34887 ;
  assign n34889 = n608 & ~n13132 ;
  assign n34890 = ~n25631 & n34889 ;
  assign n34891 = n13995 & n19735 ;
  assign n34892 = ( n3692 & ~n10709 ) | ( n3692 & n30565 ) | ( ~n10709 & n30565 ) ;
  assign n34893 = ~n34891 & n34892 ;
  assign n34894 = ~n16723 & n34893 ;
  assign n34895 = ~n11608 & n33339 ;
  assign n34896 = ~n34894 & n34895 ;
  assign n34897 = ( n329 & n981 ) | ( n329 & n13362 ) | ( n981 & n13362 ) ;
  assign n34898 = ~n6035 & n34897 ;
  assign n34899 = n34898 ^ n14854 ^ 1'b0 ;
  assign n34900 = x23 & ~n34899 ;
  assign n34901 = ( n1260 & n7408 ) | ( n1260 & ~n18645 ) | ( n7408 & ~n18645 ) ;
  assign n34902 = n34901 ^ n22453 ^ n21509 ;
  assign n34903 = n29132 ^ n13752 ^ 1'b0 ;
  assign n34904 = n22914 ^ n2937 ^ 1'b0 ;
  assign n34905 = n34903 & ~n34904 ;
  assign n34906 = n3283 ^ n1535 ^ 1'b0 ;
  assign n34907 = n22541 | n23350 ;
  assign n34908 = n23861 | n34907 ;
  assign n34909 = n23474 & ~n34908 ;
  assign n34910 = n21000 ^ n5836 ^ 1'b0 ;
  assign n34911 = n742 & ~n14738 ;
  assign n34912 = ~n31119 & n34911 ;
  assign n34913 = n14581 & ~n23623 ;
  assign n34914 = n34913 ^ n14306 ^ 1'b0 ;
  assign n34915 = n16516 ^ n12678 ^ 1'b0 ;
  assign n34916 = ( n7807 & n22194 ) | ( n7807 & n33493 ) | ( n22194 & n33493 ) ;
  assign n34917 = n7633 & ~n20730 ;
  assign n34918 = ~n836 & n34917 ;
  assign n34919 = n34918 ^ n28728 ^ 1'b0 ;
  assign n34920 = n20511 & ~n21705 ;
  assign n34921 = n34244 ^ n23678 ^ n12834 ;
  assign n34922 = n28138 ^ n17283 ^ n12788 ;
  assign n34923 = n2582 | n9001 ;
  assign n34924 = n34923 ^ n8102 ^ 1'b0 ;
  assign n34925 = n5946 | n10686 ;
  assign n34930 = n2966 & n7977 ;
  assign n34926 = n4750 & ~n6469 ;
  assign n34927 = n34926 ^ n14736 ^ n289 ;
  assign n34928 = n27442 & n34927 ;
  assign n34929 = n34928 ^ n930 ^ 1'b0 ;
  assign n34931 = n34930 ^ n34929 ^ n15939 ;
  assign n34932 = n24403 ^ n11446 ^ 1'b0 ;
  assign n34934 = n5430 & ~n21089 ;
  assign n34935 = n34934 ^ n10973 ^ 1'b0 ;
  assign n34936 = n1476 & n12760 ;
  assign n34937 = ~n8913 & n34936 ;
  assign n34938 = n34937 ^ n24456 ^ n23542 ;
  assign n34939 = n34935 & n34938 ;
  assign n34940 = n18289 & n34939 ;
  assign n34941 = n34940 ^ n9686 ^ 1'b0 ;
  assign n34933 = n8501 & n25757 ;
  assign n34942 = n34941 ^ n34933 ^ 1'b0 ;
  assign n34943 = n24884 ^ n22690 ^ 1'b0 ;
  assign n34944 = n19557 ^ n2344 ^ 1'b0 ;
  assign n34945 = n16491 & n34944 ;
  assign n34946 = ( n11401 & n23068 ) | ( n11401 & ~n34945 ) | ( n23068 & ~n34945 ) ;
  assign n34947 = ~n1253 & n4494 ;
  assign n34948 = n4097 & ~n5031 ;
  assign n34949 = n7112 & ~n26903 ;
  assign n34950 = n25990 ^ n2318 ^ 1'b0 ;
  assign n34951 = n34950 ^ n20182 ^ n3111 ;
  assign n34952 = n22096 & n34951 ;
  assign n34953 = n34952 ^ n14227 ^ 1'b0 ;
  assign n34954 = n27801 | n32858 ;
  assign n34955 = n34954 ^ n18636 ^ 1'b0 ;
  assign n34956 = n20496 | n34955 ;
  assign n34957 = n34956 ^ n12947 ^ 1'b0 ;
  assign n34958 = n34957 ^ n6481 ^ 1'b0 ;
  assign n34959 = n7607 & ~n11885 ;
  assign n34960 = n33826 ^ n10733 ^ 1'b0 ;
  assign n34961 = ~n1453 & n15760 ;
  assign n34962 = ~n14715 & n25944 ;
  assign n34963 = n24081 & n34962 ;
  assign n34964 = ( n1635 & n14057 ) | ( n1635 & n27423 ) | ( n14057 & n27423 ) ;
  assign n34965 = n24123 ^ n14886 ^ n11914 ;
  assign n34966 = ~n34964 & n34965 ;
  assign n34967 = n14673 & n26625 ;
  assign n34968 = n34967 ^ n6354 ^ 1'b0 ;
  assign n34969 = ~n21903 & n25920 ;
  assign n34970 = n7663 & n19671 ;
  assign n34971 = n2217 & ~n34970 ;
  assign n34972 = n34971 ^ n20293 ^ 1'b0 ;
  assign n34973 = n34972 ^ n7377 ^ 1'b0 ;
  assign n34974 = n34973 ^ n9707 ^ 1'b0 ;
  assign n34975 = n681 | n29159 ;
  assign n34976 = n2722 | n4698 ;
  assign n34977 = n34976 ^ n4975 ^ 1'b0 ;
  assign n34978 = ( n6661 & n24175 ) | ( n6661 & ~n34977 ) | ( n24175 & ~n34977 ) ;
  assign n34983 = n14375 & n19953 ;
  assign n34984 = n34983 ^ n28358 ^ 1'b0 ;
  assign n34979 = n692 & ~n14697 ;
  assign n34980 = ~n5701 & n34979 ;
  assign n34981 = n34980 ^ n28117 ^ n13272 ;
  assign n34982 = n7696 & ~n34981 ;
  assign n34985 = n34984 ^ n34982 ^ 1'b0 ;
  assign n34986 = n1983 & ~n16802 ;
  assign n34987 = n34986 ^ n6940 ^ 1'b0 ;
  assign n34988 = n8246 & n15814 ;
  assign n34989 = n34988 ^ n4043 ^ 1'b0 ;
  assign n34990 = n5247 ^ n400 ^ 1'b0 ;
  assign n34991 = n10026 & ~n34990 ;
  assign n34992 = x11 & n22150 ;
  assign n34993 = ~n7705 & n34992 ;
  assign n34995 = n16018 ^ n5719 ^ 1'b0 ;
  assign n34996 = n21608 ^ n1127 ^ 1'b0 ;
  assign n34997 = n34995 & ~n34996 ;
  assign n34994 = n275 & ~n16491 ;
  assign n34998 = n34997 ^ n34994 ^ 1'b0 ;
  assign n34999 = n2044 & n31364 ;
  assign n35000 = n20599 ^ n2686 ^ 1'b0 ;
  assign n35001 = n35000 ^ n30977 ^ 1'b0 ;
  assign n35003 = ~n2549 & n15170 ;
  assign n35004 = n35003 ^ n536 ^ 1'b0 ;
  assign n35002 = n10028 & n22658 ;
  assign n35005 = n35004 ^ n35002 ^ n13386 ;
  assign n35006 = n21464 & n35005 ;
  assign n35007 = ~n24116 & n35006 ;
  assign n35008 = n35007 ^ n2856 ^ 1'b0 ;
  assign n35009 = n2437 | n6971 ;
  assign n35010 = n2186 & n11091 ;
  assign n35011 = ~n35009 & n35010 ;
  assign n35012 = n3756 & ~n26261 ;
  assign n35013 = n8262 & n15945 ;
  assign n35014 = n16143 & n35013 ;
  assign n35015 = n18490 | n32204 ;
  assign n35016 = ~n1339 & n18076 ;
  assign n35017 = n26674 & n35016 ;
  assign n35018 = n22056 | n35017 ;
  assign n35019 = n2991 & n11709 ;
  assign n35020 = n35019 ^ n4184 ^ 1'b0 ;
  assign n35021 = ~n2726 & n8367 ;
  assign n35022 = n35021 ^ n18733 ^ 1'b0 ;
  assign n35023 = n35020 | n35022 ;
  assign n35025 = n2033 & ~n13475 ;
  assign n35026 = ~n16245 & n35025 ;
  assign n35024 = n7636 & n34493 ;
  assign n35027 = n35026 ^ n35024 ^ 1'b0 ;
  assign n35028 = n12437 ^ n2965 ^ 1'b0 ;
  assign n35029 = ~n22832 & n35028 ;
  assign n35030 = n6018 | n7027 ;
  assign n35031 = n35030 ^ n23538 ^ 1'b0 ;
  assign n35033 = n21361 ^ n13149 ^ 1'b0 ;
  assign n35034 = n13915 & n35033 ;
  assign n35032 = n3830 & ~n32439 ;
  assign n35035 = n35034 ^ n35032 ^ 1'b0 ;
  assign n35036 = n30041 ^ n25033 ^ 1'b0 ;
  assign n35037 = n1102 & n22497 ;
  assign n35038 = n28181 ^ n3528 ^ 1'b0 ;
  assign n35039 = n26893 & n35038 ;
  assign n35040 = n6572 | n17758 ;
  assign n35041 = n14604 ^ n5675 ^ 1'b0 ;
  assign n35042 = n26119 ^ n16490 ^ 1'b0 ;
  assign n35043 = n10389 & ~n35042 ;
  assign n35044 = n35043 ^ n26899 ^ 1'b0 ;
  assign n35045 = n1594 & ~n7469 ;
  assign n35046 = ~n7846 & n24165 ;
  assign n35047 = n2868 | n35046 ;
  assign n35048 = ~n6692 & n22873 ;
  assign n35049 = ~n7033 & n35048 ;
  assign n35050 = n16288 ^ n1543 ^ 1'b0 ;
  assign n35051 = n20538 & n35050 ;
  assign n35052 = ~n28287 & n35051 ;
  assign n35053 = n3036 | n14816 ;
  assign n35054 = n34980 & ~n35053 ;
  assign n35055 = n31916 ^ n3765 ^ 1'b0 ;
  assign n35056 = n4631 & n35055 ;
  assign n35060 = n6382 & ~n9259 ;
  assign n35061 = n15155 | n35060 ;
  assign n35062 = n35061 ^ n29285 ^ 1'b0 ;
  assign n35063 = n35062 ^ n1897 ^ 1'b0 ;
  assign n35064 = ~n8372 & n35063 ;
  assign n35057 = n4093 | n14563 ;
  assign n35058 = n20574 & ~n35057 ;
  assign n35059 = n13972 & ~n35058 ;
  assign n35065 = n35064 ^ n35059 ^ 1'b0 ;
  assign n35066 = n2875 & n17838 ;
  assign n35067 = n35066 ^ n6364 ^ 1'b0 ;
  assign n35068 = n15265 ^ n13266 ^ n2839 ;
  assign n35069 = n1281 & n1619 ;
  assign n35070 = ~n35068 & n35069 ;
  assign n35071 = n8274 ^ n5927 ^ n2320 ;
  assign n35072 = n28752 ^ n7821 ^ 1'b0 ;
  assign n35073 = n35071 & n35072 ;
  assign n35074 = ~n267 & n11724 ;
  assign n35075 = ~n21834 & n30310 ;
  assign n35076 = n9133 ^ n6198 ^ x216 ;
  assign n35077 = n35076 ^ n22503 ^ 1'b0 ;
  assign n35078 = n1044 | n35077 ;
  assign n35079 = n2173 & ~n26422 ;
  assign n35080 = n7073 ^ n6594 ^ 1'b0 ;
  assign n35081 = n7760 & n35080 ;
  assign n35082 = n26744 | n35081 ;
  assign n35083 = n20783 ^ n5857 ^ 1'b0 ;
  assign n35084 = n4844 | n35083 ;
  assign n35085 = n22340 ^ x139 ^ 1'b0 ;
  assign n35086 = n16106 & ~n35085 ;
  assign n35087 = ~n35084 & n35086 ;
  assign n35088 = n35087 ^ n28510 ^ 1'b0 ;
  assign n35089 = n2490 & ~n21343 ;
  assign n35090 = n35089 ^ n33123 ^ n6227 ;
  assign n35091 = n677 & ~n12701 ;
  assign n35092 = ~n20878 & n35091 ;
  assign n35093 = n35090 & n35092 ;
  assign n35094 = ~n4590 & n17640 ;
  assign n35095 = n35094 ^ n31949 ^ 1'b0 ;
  assign n35096 = n25945 ^ n21060 ^ 1'b0 ;
  assign n35097 = ~n9423 & n18560 ;
  assign n35098 = n35096 & n35097 ;
  assign n35099 = ~n19467 & n28410 ;
  assign n35100 = n35099 ^ n24374 ^ 1'b0 ;
  assign n35101 = ( n6373 & n7636 ) | ( n6373 & ~n23242 ) | ( n7636 & ~n23242 ) ;
  assign n35102 = n10039 ^ n3604 ^ 1'b0 ;
  assign n35103 = x42 & n35102 ;
  assign n35104 = ~n11405 & n35103 ;
  assign n35105 = n35104 ^ n26318 ^ 1'b0 ;
  assign n35106 = ~n2723 & n35105 ;
  assign n35107 = n4047 & n35106 ;
  assign n35108 = n1173 & n20424 ;
  assign n35109 = n35108 ^ n11070 ^ 1'b0 ;
  assign n35113 = n9819 & ~n26057 ;
  assign n35114 = n985 & n35113 ;
  assign n35110 = n27702 ^ n832 ^ 1'b0 ;
  assign n35111 = n4139 | n35110 ;
  assign n35112 = n21361 | n35111 ;
  assign n35115 = n35114 ^ n35112 ^ 1'b0 ;
  assign n35116 = n22261 ^ n17917 ^ 1'b0 ;
  assign n35117 = n6684 & n17657 ;
  assign n35118 = ~n28680 & n35117 ;
  assign n35119 = n35118 ^ n22245 ^ n6692 ;
  assign n35120 = n18264 | n35119 ;
  assign n35121 = n21048 ^ n19257 ^ 1'b0 ;
  assign n35122 = n13860 & n35121 ;
  assign n35123 = n35122 ^ n18714 ^ 1'b0 ;
  assign n35124 = ( x190 & ~n17830 ) | ( x190 & n26616 ) | ( ~n17830 & n26616 ) ;
  assign n35125 = n35117 ^ n24776 ^ n8663 ;
  assign n35126 = n4658 & ~n6207 ;
  assign n35127 = n35126 ^ n22936 ^ n5182 ;
  assign n35128 = ( ~n6518 & n26595 ) | ( ~n6518 & n29295 ) | ( n26595 & n29295 ) ;
  assign n35129 = n26328 | n35128 ;
  assign n35130 = n1471 & ~n13327 ;
  assign n35131 = n35130 ^ n27444 ^ 1'b0 ;
  assign n35132 = n32746 ^ n9056 ^ 1'b0 ;
  assign n35133 = n5200 & n16827 ;
  assign n35134 = ~n35132 & n35133 ;
  assign n35135 = ( n674 & n11183 ) | ( n674 & n27456 ) | ( n11183 & n27456 ) ;
  assign n35136 = n10513 | n21216 ;
  assign n35137 = n21377 & ~n35136 ;
  assign n35138 = n20263 ^ n841 ^ 1'b0 ;
  assign n35139 = n35137 & ~n35138 ;
  assign n35140 = n35139 ^ n34102 ^ 1'b0 ;
  assign n35141 = n14179 & n35140 ;
  assign n35142 = n500 & n32955 ;
  assign n35143 = n12251 & n22214 ;
  assign n35144 = n35143 ^ n8121 ^ 1'b0 ;
  assign n35145 = ~n33907 & n35073 ;
  assign n35146 = n25257 ^ n12715 ^ 1'b0 ;
  assign n35147 = n9170 ^ n6929 ^ n3716 ;
  assign n35148 = n14858 ^ n2664 ^ 1'b0 ;
  assign n35149 = n8519 ^ n3864 ^ 1'b0 ;
  assign n35150 = ~n5373 & n20643 ;
  assign n35151 = n35150 ^ n18860 ^ 1'b0 ;
  assign n35152 = n35149 & n35151 ;
  assign n35153 = n30814 ^ n27997 ^ 1'b0 ;
  assign n35154 = ~n7251 & n35153 ;
  assign n35155 = ~n18442 & n35154 ;
  assign n35156 = n35155 ^ n16574 ^ 1'b0 ;
  assign n35157 = n23625 & ~n35156 ;
  assign n35158 = ~n3597 & n35157 ;
  assign n35164 = n2277 & ~n8554 ;
  assign n35165 = ~n2277 & n35164 ;
  assign n35166 = n35165 ^ n2497 ^ 1'b0 ;
  assign n35159 = n1213 | n3490 ;
  assign n35160 = n3490 & ~n35159 ;
  assign n35161 = n12961 ^ n8612 ^ 1'b0 ;
  assign n35162 = ~n35160 & n35161 ;
  assign n35163 = ( n11710 & n21756 ) | ( n11710 & n35162 ) | ( n21756 & n35162 ) ;
  assign n35167 = n35166 ^ n35163 ^ n21490 ;
  assign n35168 = n6781 ^ n2723 ^ n1177 ;
  assign n35169 = n2253 | n35168 ;
  assign n35170 = n19821 & ~n35169 ;
  assign n35171 = n35167 | n35170 ;
  assign n35183 = n28165 ^ n12480 ^ 1'b0 ;
  assign n35184 = n26768 ^ n16709 ^ 1'b0 ;
  assign n35185 = ~n35183 & n35184 ;
  assign n35186 = n35185 ^ n19736 ^ n14967 ;
  assign n35172 = n16291 ^ n9531 ^ 1'b0 ;
  assign n35173 = n35172 ^ n10045 ^ 1'b0 ;
  assign n35174 = ~n11651 & n35173 ;
  assign n35175 = n25142 ^ n6756 ^ 1'b0 ;
  assign n35176 = n35174 & n35175 ;
  assign n35177 = n704 | n1957 ;
  assign n35178 = n8271 & ~n35177 ;
  assign n35179 = n35178 ^ n8366 ^ 1'b0 ;
  assign n35180 = ~n5033 & n35179 ;
  assign n35181 = n25290 & n35180 ;
  assign n35182 = n35176 & ~n35181 ;
  assign n35187 = n35186 ^ n35182 ^ 1'b0 ;
  assign n35188 = n18615 ^ n17891 ^ 1'b0 ;
  assign n35189 = ~n8001 & n35188 ;
  assign n35190 = ~n10733 & n15723 ;
  assign n35191 = n22572 & n35190 ;
  assign n35192 = n20759 & ~n35191 ;
  assign n35193 = n35192 ^ n26213 ^ 1'b0 ;
  assign n35194 = ( n3347 & ~n13941 ) | ( n3347 & n15074 ) | ( ~n13941 & n15074 ) ;
  assign n35195 = x111 & n35194 ;
  assign n35196 = n35195 ^ n2623 ^ 1'b0 ;
  assign n35197 = n27591 ^ n25506 ^ 1'b0 ;
  assign n35198 = n8281 & n14894 ;
  assign n35199 = n27255 ^ n15931 ^ 1'b0 ;
  assign n35200 = ( n4991 & n7068 ) | ( n4991 & ~n9045 ) | ( n7068 & ~n9045 ) ;
  assign n35201 = n21275 & ~n35200 ;
  assign n35202 = n2480 & n35201 ;
  assign n35203 = n735 | n35202 ;
  assign n35204 = n35199 & ~n35203 ;
  assign n35205 = n28829 ^ n1865 ^ n780 ;
  assign n35206 = n2260 | n8268 ;
  assign n35207 = n12238 & n35206 ;
  assign n35208 = n26137 ^ n11818 ^ 1'b0 ;
  assign n35209 = n3497 | n3749 ;
  assign n35210 = n1797 & ~n35209 ;
  assign n35211 = n17731 & ~n33413 ;
  assign n35212 = n35211 ^ n21109 ^ 1'b0 ;
  assign n35213 = n15188 & n35212 ;
  assign n35214 = n35213 ^ n7682 ^ 1'b0 ;
  assign n35215 = ~n35210 & n35214 ;
  assign n35218 = ( n3746 & ~n17655 ) | ( n3746 & n22985 ) | ( ~n17655 & n22985 ) ;
  assign n35216 = n3898 & ~n12275 ;
  assign n35217 = n25357 & n35216 ;
  assign n35219 = n35218 ^ n35217 ^ n16186 ;
  assign n35220 = n16482 ^ n10026 ^ 1'b0 ;
  assign n35221 = n1009 & ~n35220 ;
  assign n35222 = ~n14422 & n35221 ;
  assign n35223 = n3877 & n35222 ;
  assign n35224 = n35219 & n35223 ;
  assign n35225 = n27545 ^ n26234 ^ 1'b0 ;
  assign n35226 = n9885 | n35225 ;
  assign n35227 = n3556 | n35226 ;
  assign n35228 = n9247 | n23764 ;
  assign n35229 = n35227 | n35228 ;
  assign n35230 = n15951 ^ n7632 ^ 1'b0 ;
  assign n35231 = n3647 & n35230 ;
  assign n35232 = ( n14576 & ~n20503 ) | ( n14576 & n35231 ) | ( ~n20503 & n35231 ) ;
  assign n35233 = ~n1310 & n1688 ;
  assign n35234 = n35233 ^ n14668 ^ n5238 ;
  assign n35235 = ( n843 & ~n27334 ) | ( n843 & n29876 ) | ( ~n27334 & n29876 ) ;
  assign n35236 = ( ~n7709 & n8785 ) | ( ~n7709 & n35235 ) | ( n8785 & n35235 ) ;
  assign n35237 = ~n5471 & n13994 ;
  assign n35238 = ~n14482 & n35237 ;
  assign n35239 = ( n14579 & ~n16702 ) | ( n14579 & n35238 ) | ( ~n16702 & n35238 ) ;
  assign n35240 = n13535 | n24333 ;
  assign n35241 = n5988 ^ n3919 ^ 1'b0 ;
  assign n35242 = ~n6131 & n35241 ;
  assign n35243 = ~n6567 & n19220 ;
  assign n35244 = n14570 ^ n8393 ^ 1'b0 ;
  assign n35245 = n27831 | n35244 ;
  assign n35246 = n13527 ^ n3352 ^ 1'b0 ;
  assign n35247 = ( n8342 & n14410 ) | ( n8342 & n25320 ) | ( n14410 & n25320 ) ;
  assign n35248 = n35247 ^ n13920 ^ n283 ;
  assign n35249 = n2300 & ~n8823 ;
  assign n35250 = n8823 & n35249 ;
  assign n35251 = n35250 ^ n15440 ^ 1'b0 ;
  assign n35252 = ~n3882 & n5306 ;
  assign n35253 = ~n5306 & n35252 ;
  assign n35254 = ~n7644 & n35253 ;
  assign n35255 = ~n3523 & n35254 ;
  assign n35256 = n35255 ^ n6747 ^ 1'b0 ;
  assign n35257 = n35251 & ~n35256 ;
  assign n35258 = ( n11633 & n27083 ) | ( n11633 & ~n35257 ) | ( n27083 & ~n35257 ) ;
  assign n35259 = n28276 ^ n24348 ^ 1'b0 ;
  assign n35260 = n3714 | n35259 ;
  assign n35261 = n21242 ^ n12805 ^ 1'b0 ;
  assign n35262 = n512 | n7685 ;
  assign n35263 = ~n6801 & n23647 ;
  assign n35264 = n4415 & ~n15516 ;
  assign n35265 = ( n17829 & ~n23773 ) | ( n17829 & n35264 ) | ( ~n23773 & n35264 ) ;
  assign n35266 = n17515 & ~n35265 ;
  assign n35267 = n15519 ^ n2623 ^ 1'b0 ;
  assign n35268 = ~n1991 & n7801 ;
  assign n35269 = ~n7999 & n35268 ;
  assign n35270 = n10191 & ~n14268 ;
  assign n35271 = n35270 ^ n22225 ^ 1'b0 ;
  assign n35272 = n8007 | n35271 ;
  assign n35274 = n4797 & n9804 ;
  assign n35275 = n35274 ^ n4533 ^ 1'b0 ;
  assign n35276 = n10881 | n35275 ;
  assign n35277 = n3475 | n35276 ;
  assign n35278 = n11191 & n35277 ;
  assign n35273 = ~n681 & n12606 ;
  assign n35279 = n35278 ^ n35273 ^ 1'b0 ;
  assign n35280 = n1122 & ~n9070 ;
  assign n35281 = n516 & n35280 ;
  assign n35282 = n8776 ^ n292 ^ 1'b0 ;
  assign n35283 = x82 & ~n605 ;
  assign n35284 = n605 & n35283 ;
  assign n35285 = n3434 | n35284 ;
  assign n35286 = n9077 ^ n8941 ^ n6995 ;
  assign n35287 = ~n11001 & n35286 ;
  assign n35288 = n35287 ^ n30859 ^ 1'b0 ;
  assign n35289 = n35288 ^ n25958 ^ 1'b0 ;
  assign n35290 = n35285 | n35289 ;
  assign n35291 = n23228 ^ n9456 ^ 1'b0 ;
  assign n35292 = ( n8288 & ~n9402 ) | ( n8288 & n20516 ) | ( ~n9402 & n20516 ) ;
  assign n35293 = n10334 & n35292 ;
  assign n35294 = n5569 ^ n1170 ^ 1'b0 ;
  assign n35295 = n35294 ^ n13982 ^ 1'b0 ;
  assign n35296 = n20686 ^ n11898 ^ 1'b0 ;
  assign n35297 = ~n35295 & n35296 ;
  assign n35298 = n4534 & ~n27296 ;
  assign n35299 = n5260 ^ n4062 ^ 1'b0 ;
  assign n35300 = n5967 & n22713 ;
  assign n35301 = n34445 & n35300 ;
  assign n35302 = n26431 & ~n35301 ;
  assign n35303 = n24129 & n35302 ;
  assign n35304 = ( n6272 & ~n12557 ) | ( n6272 & n19412 ) | ( ~n12557 & n19412 ) ;
  assign n35305 = ~n7679 & n35304 ;
  assign n35306 = n14206 & n35305 ;
  assign n35307 = ~n18394 & n35306 ;
  assign n35308 = n9977 | n21034 ;
  assign n35309 = n15381 & n25895 ;
  assign n35310 = n35309 ^ n23470 ^ 1'b0 ;
  assign n35311 = n12128 ^ n7569 ^ 1'b0 ;
  assign n35312 = n30565 & ~n35311 ;
  assign n35313 = ( n27481 & n30483 ) | ( n27481 & ~n35312 ) | ( n30483 & ~n35312 ) ;
  assign n35314 = n6936 & n25587 ;
  assign n35315 = n16122 & n35314 ;
  assign n35316 = n21606 | n32127 ;
  assign n35317 = n35316 ^ n31542 ^ 1'b0 ;
  assign n35318 = ~n11532 & n32070 ;
  assign n35319 = ~n9875 & n35318 ;
  assign n35320 = n22895 ^ n21061 ^ n8780 ;
  assign n35321 = n29921 ^ n21575 ^ 1'b0 ;
  assign n35322 = n35320 | n35321 ;
  assign n35323 = ~n5758 & n9255 ;
  assign n35324 = n16405 & ~n26402 ;
  assign n35325 = ~n35323 & n35324 ;
  assign n35326 = ~n10504 & n14054 ;
  assign n35327 = n35325 & n35326 ;
  assign n35328 = n31084 ^ n18431 ^ n9783 ;
  assign n35329 = n26029 & ~n35328 ;
  assign n35331 = n29612 ^ n5616 ^ 1'b0 ;
  assign n35332 = n33903 ^ n27626 ^ 1'b0 ;
  assign n35333 = n35331 | n35332 ;
  assign n35330 = n15493 & n25094 ;
  assign n35334 = n35333 ^ n35330 ^ 1'b0 ;
  assign n35335 = n2096 | n11857 ;
  assign n35336 = n34040 ^ n5728 ^ n3278 ;
  assign n35337 = n15966 ^ n14469 ^ 1'b0 ;
  assign n35338 = n33282 | n35337 ;
  assign n35339 = n15990 ^ n9385 ^ 1'b0 ;
  assign n35340 = n32253 & n35339 ;
  assign n35341 = n4731 & n35017 ;
  assign n35342 = n5085 & n35341 ;
  assign n35343 = n4366 ^ n4282 ^ 1'b0 ;
  assign n35344 = n9188 & n11572 ;
  assign n35345 = n9525 & n35344 ;
  assign n35346 = ( ~n6714 & n35343 ) | ( ~n6714 & n35345 ) | ( n35343 & n35345 ) ;
  assign n35347 = ~n26130 & n35346 ;
  assign n35348 = ~n1730 & n35347 ;
  assign n35349 = ( n6182 & n6896 ) | ( n6182 & ~n29172 ) | ( n6896 & ~n29172 ) ;
  assign n35351 = n16599 & ~n20707 ;
  assign n35350 = n9106 ^ n5411 ^ 1'b0 ;
  assign n35352 = n35351 ^ n35350 ^ n31696 ;
  assign n35353 = n18440 ^ n449 ^ 1'b0 ;
  assign n35354 = n7301 & n15246 ;
  assign n35355 = n33856 ^ n20753 ^ 1'b0 ;
  assign n35356 = n28583 | n35355 ;
  assign n35357 = n4326 & n33953 ;
  assign n35358 = ( n17218 & n22040 ) | ( n17218 & n35357 ) | ( n22040 & n35357 ) ;
  assign n35359 = n19609 ^ n12955 ^ 1'b0 ;
  assign n35360 = n842 & n35359 ;
  assign n35361 = n35360 ^ n28658 ^ n18592 ;
  assign n35362 = ( n14876 & n30407 ) | ( n14876 & n34999 ) | ( n30407 & n34999 ) ;
  assign n35363 = n756 | n4241 ;
  assign n35364 = n30478 & ~n35363 ;
  assign n35365 = ~n23533 & n35364 ;
  assign n35366 = n17534 & n34148 ;
  assign n35367 = n35366 ^ n9332 ^ 1'b0 ;
  assign n35368 = n20757 ^ n388 ^ 1'b0 ;
  assign n35369 = n35368 ^ x239 ^ 1'b0 ;
  assign n35370 = n9897 & ~n35369 ;
  assign n35371 = n17802 ^ n1836 ^ 1'b0 ;
  assign n35372 = n30052 ^ n19887 ^ 1'b0 ;
  assign n35373 = n35371 | n35372 ;
  assign n35374 = n3617 & ~n7908 ;
  assign n35375 = ( ~n5330 & n21265 ) | ( ~n5330 & n35374 ) | ( n21265 & n35374 ) ;
  assign n35376 = n35375 ^ n25527 ^ n10078 ;
  assign n35377 = n11389 & ~n30032 ;
  assign n35378 = n924 | n1365 ;
  assign n35379 = n1365 & ~n35378 ;
  assign n35380 = n5885 | n35379 ;
  assign n35381 = n35379 & ~n35380 ;
  assign n35382 = n4860 | n35381 ;
  assign n35383 = n35381 & ~n35382 ;
  assign n35384 = ~n2797 & n4194 ;
  assign n35385 = n35384 ^ n8406 ^ 1'b0 ;
  assign n35386 = n35385 ^ n17282 ^ 1'b0 ;
  assign n35387 = n24234 & ~n35386 ;
  assign n35388 = n35387 ^ n9033 ^ 1'b0 ;
  assign n35389 = ~n35383 & n35388 ;
  assign n35390 = n33305 ^ n13584 ^ 1'b0 ;
  assign n35391 = ~n13749 & n35390 ;
  assign n35392 = ~n9359 & n35391 ;
  assign n35393 = x187 & n35392 ;
  assign n35394 = n1464 & ~n9695 ;
  assign n35395 = ( n1829 & ~n15843 ) | ( n1829 & n20753 ) | ( ~n15843 & n20753 ) ;
  assign n35396 = ( ~n22655 & n35394 ) | ( ~n22655 & n35395 ) | ( n35394 & n35395 ) ;
  assign n35397 = ( n4726 & n5558 ) | ( n4726 & ~n22140 ) | ( n5558 & ~n22140 ) ;
  assign n35398 = n25908 & ~n34871 ;
  assign n35399 = ~n17942 & n35398 ;
  assign n35400 = ~n12172 & n26883 ;
  assign n35401 = n9020 & n15522 ;
  assign n35402 = n35400 & n35401 ;
  assign n35403 = n7565 | n35402 ;
  assign n35404 = n7033 | n13513 ;
  assign n35405 = n9173 & ~n35404 ;
  assign n35406 = n35405 ^ n3920 ^ 1'b0 ;
  assign n35407 = n35406 ^ n6233 ^ 1'b0 ;
  assign n35408 = n8917 & ~n35407 ;
  assign n35409 = ~n9971 & n10204 ;
  assign n35410 = n10201 & n35409 ;
  assign n35411 = n12625 | n35410 ;
  assign n35412 = n35411 ^ n7843 ^ 1'b0 ;
  assign n35413 = ~n3003 & n6450 ;
  assign n35414 = n17128 | n34318 ;
  assign n35415 = n35414 ^ n5521 ^ 1'b0 ;
  assign n35416 = n366 & n15533 ;
  assign n35417 = n7265 | n27205 ;
  assign n35418 = n35417 ^ n26618 ^ 1'b0 ;
  assign n35419 = ~n919 & n35418 ;
  assign n35420 = ~n35416 & n35419 ;
  assign n35421 = n16904 & n24210 ;
  assign n35422 = n35421 ^ n10962 ^ 1'b0 ;
  assign n35423 = n26527 ^ n14368 ^ 1'b0 ;
  assign n35424 = ~n7074 & n35423 ;
  assign n35425 = n35424 ^ n14028 ^ 1'b0 ;
  assign n35426 = n5514 ^ n4587 ^ 1'b0 ;
  assign n35428 = n13131 ^ n9133 ^ 1'b0 ;
  assign n35429 = n9375 & n35428 ;
  assign n35427 = n1536 & ~n5813 ;
  assign n35430 = n35429 ^ n35427 ^ 1'b0 ;
  assign n35431 = n5361 & ~n17128 ;
  assign n35433 = n25455 ^ n23614 ^ 1'b0 ;
  assign n35434 = n6481 & n35433 ;
  assign n35435 = ~n32053 & n35434 ;
  assign n35432 = ~n5720 & n31238 ;
  assign n35436 = n35435 ^ n35432 ^ 1'b0 ;
  assign n35437 = n28589 ^ n3272 ^ 1'b0 ;
  assign n35438 = n10102 | n15406 ;
  assign n35439 = n17666 ^ n17302 ^ n4618 ;
  assign n35440 = n34805 ^ n29811 ^ n26193 ;
  assign n35441 = ( ~n15851 & n19746 ) | ( ~n15851 & n30634 ) | ( n19746 & n30634 ) ;
  assign n35442 = n9074 | n35441 ;
  assign n35443 = n35442 ^ n23706 ^ 1'b0 ;
  assign n35454 = n2528 | n2550 ;
  assign n35455 = n2550 & ~n35454 ;
  assign n35444 = x239 & ~n536 ;
  assign n35445 = n536 & n35444 ;
  assign n35446 = x61 & ~n1510 ;
  assign n35447 = n1510 & n35446 ;
  assign n35448 = n320 | n35447 ;
  assign n35449 = n320 & ~n35448 ;
  assign n35450 = x35 & ~n35449 ;
  assign n35451 = n35445 & n35450 ;
  assign n35452 = n10033 & ~n35451 ;
  assign n35453 = n35451 & n35452 ;
  assign n35456 = n35455 ^ n35453 ^ 1'b0 ;
  assign n35457 = ~n20730 & n35456 ;
  assign n35458 = n27150 & ~n30491 ;
  assign n35459 = n28158 ^ n22123 ^ 1'b0 ;
  assign n35460 = ( n2327 & ~n8813 ) | ( n2327 & n10835 ) | ( ~n8813 & n10835 ) ;
  assign n35461 = n18536 & n32673 ;
  assign n35462 = n16846 ^ n15118 ^ 1'b0 ;
  assign n35463 = ~n16848 & n35462 ;
  assign n35464 = n35463 ^ n4960 ^ 1'b0 ;
  assign n35465 = n9219 & ~n35464 ;
  assign n35466 = n2991 & ~n19085 ;
  assign n35469 = n8854 ^ n2327 ^ n2204 ;
  assign n35467 = n5907 ^ n1460 ^ n1073 ;
  assign n35468 = n35467 ^ n21370 ^ n6077 ;
  assign n35470 = n35469 ^ n35468 ^ n4135 ;
  assign n35471 = n16793 ^ n15778 ^ 1'b0 ;
  assign n35472 = n27591 & n35471 ;
  assign n35473 = n32790 ^ n1809 ^ 1'b0 ;
  assign n35474 = n3245 & ~n35473 ;
  assign n35475 = n8083 & ~n35294 ;
  assign n35476 = n35475 ^ n7593 ^ 1'b0 ;
  assign n35477 = n6232 & n35476 ;
  assign n35478 = n35477 ^ n13768 ^ 1'b0 ;
  assign n35479 = ( n5642 & ~n9877 ) | ( n5642 & n15282 ) | ( ~n9877 & n15282 ) ;
  assign n35480 = n35479 ^ n24214 ^ 1'b0 ;
  assign n35481 = n8246 & n35480 ;
  assign n35482 = n27019 ^ n22909 ^ n2518 ;
  assign n35483 = n5230 | n23199 ;
  assign n35484 = n7841 & n28480 ;
  assign n35485 = n35484 ^ n28801 ^ 1'b0 ;
  assign n35486 = n30978 ^ n13932 ^ 1'b0 ;
  assign n35487 = ~n35485 & n35486 ;
  assign n35488 = n9524 ^ n3551 ^ 1'b0 ;
  assign n35489 = n7600 & n35488 ;
  assign n35490 = n35489 ^ n11596 ^ 1'b0 ;
  assign n35491 = n29497 | n35490 ;
  assign n35492 = ( n635 & n23518 ) | ( n635 & n35491 ) | ( n23518 & n35491 ) ;
  assign n35493 = ( n2183 & n18675 ) | ( n2183 & n22960 ) | ( n18675 & n22960 ) ;
  assign n35494 = n11292 & ~n25069 ;
  assign n35495 = n35494 ^ n14020 ^ 1'b0 ;
  assign n35496 = n25137 & ~n35495 ;
  assign n35497 = n6701 & n26923 ;
  assign n35498 = n35497 ^ n28083 ^ 1'b0 ;
  assign n35499 = n30622 ^ x167 ^ 1'b0 ;
  assign n35500 = n21945 & ~n35499 ;
  assign n35501 = n2413 & ~n7794 ;
  assign n35502 = ~n20984 & n35501 ;
  assign n35503 = n21761 | n35502 ;
  assign n35504 = n35503 ^ n6624 ^ 1'b0 ;
  assign n35505 = ~n31379 & n35504 ;
  assign n35507 = n9713 ^ n4518 ^ 1'b0 ;
  assign n35508 = n8820 & n35507 ;
  assign n35506 = n14489 | n17731 ;
  assign n35509 = n35508 ^ n35506 ^ n30233 ;
  assign n35510 = n15231 | n21194 ;
  assign n35511 = n35510 ^ n17982 ^ 1'b0 ;
  assign n35512 = n30739 ^ n6455 ^ 1'b0 ;
  assign n35513 = n35511 | n35512 ;
  assign n35514 = n5868 ^ n5598 ^ 1'b0 ;
  assign n35515 = n35514 ^ n27530 ^ 1'b0 ;
  assign n35517 = n2728 | n5685 ;
  assign n35518 = n9083 & ~n35517 ;
  assign n35519 = ~n13080 & n35518 ;
  assign n35516 = n6945 & n19149 ;
  assign n35520 = n35519 ^ n35516 ^ 1'b0 ;
  assign n35521 = n19827 ^ n13077 ^ 1'b0 ;
  assign n35522 = n1000 ^ n686 ^ 1'b0 ;
  assign n35523 = n7756 | n27102 ;
  assign n35524 = n35523 ^ n14704 ^ 1'b0 ;
  assign n35525 = n8610 ^ n8120 ^ 1'b0 ;
  assign n35526 = n30001 & ~n35525 ;
  assign n35527 = n14531 ^ x121 ^ 1'b0 ;
  assign n35528 = ~n2160 & n35527 ;
  assign n35529 = n33124 ^ n8389 ^ 1'b0 ;
  assign n35530 = n11489 & ~n33310 ;
  assign n35531 = ~n4656 & n35530 ;
  assign n35532 = n30229 | n35531 ;
  assign n35533 = n35532 ^ n21611 ^ 1'b0 ;
  assign n35534 = ~n2839 & n26124 ;
  assign n35535 = n9055 ^ n7401 ^ 1'b0 ;
  assign n35536 = n29586 ^ n6579 ^ n1419 ;
  assign n35537 = n25659 | n35536 ;
  assign n35538 = n2539 & ~n33926 ;
  assign n35539 = n22897 & n35538 ;
  assign n35540 = ~n2098 & n6674 ;
  assign n35541 = n35540 ^ n5829 ^ 1'b0 ;
  assign n35542 = n4912 | n6331 ;
  assign n35543 = n16373 | n35542 ;
  assign n35544 = n35543 ^ n12001 ^ 1'b0 ;
  assign n35545 = ~n861 & n35544 ;
  assign n35546 = n35545 ^ n30465 ^ 1'b0 ;
  assign n35547 = n5892 ^ n5624 ^ 1'b0 ;
  assign n35548 = n27346 ^ n26666 ^ 1'b0 ;
  assign n35549 = n7443 & ~n35548 ;
  assign n35550 = n29421 ^ n9678 ^ 1'b0 ;
  assign n35551 = n27724 ^ n23690 ^ 1'b0 ;
  assign n35552 = ( n1024 & n12665 ) | ( n1024 & ~n35551 ) | ( n12665 & ~n35551 ) ;
  assign n35553 = n35552 ^ n10120 ^ 1'b0 ;
  assign n35554 = ( n1546 & n17716 ) | ( n1546 & ~n23764 ) | ( n17716 & ~n23764 ) ;
  assign n35555 = ( n14057 & n16939 ) | ( n14057 & n35554 ) | ( n16939 & n35554 ) ;
  assign n35556 = n7201 | n9849 ;
  assign n35557 = n24849 | n35556 ;
  assign n35558 = n35557 ^ n33474 ^ n3658 ;
  assign n35559 = n26550 ^ n21467 ^ 1'b0 ;
  assign n35560 = n22665 ^ n2949 ^ 1'b0 ;
  assign n35561 = n10331 | n35560 ;
  assign n35565 = ( n2355 & n4253 ) | ( n2355 & ~n20038 ) | ( n4253 & ~n20038 ) ;
  assign n35562 = ~n7233 & n28284 ;
  assign n35563 = n19671 & n35562 ;
  assign n35564 = n10102 & n35563 ;
  assign n35566 = n35565 ^ n35564 ^ n508 ;
  assign n35567 = n23369 ^ n4973 ^ 1'b0 ;
  assign n35568 = ~n9981 & n21462 ;
  assign n35569 = n33947 ^ n9128 ^ 1'b0 ;
  assign n35570 = n24340 & ~n35569 ;
  assign n35571 = n30520 ^ n18923 ^ 1'b0 ;
  assign n35572 = n7318 & ~n35571 ;
  assign n35573 = n19857 & n35572 ;
  assign n35574 = ( ~n19269 & n25622 ) | ( ~n19269 & n34895 ) | ( n25622 & n34895 ) ;
  assign n35575 = n30235 | n35574 ;
  assign n35576 = n35575 ^ n2608 ^ 1'b0 ;
  assign n35577 = ~n3804 & n6276 ;
  assign n35578 = ~n6182 & n35577 ;
  assign n35579 = n35578 ^ n9233 ^ 1'b0 ;
  assign n35580 = n27974 & ~n31322 ;
  assign n35581 = n6461 & n35580 ;
  assign n35582 = n10770 ^ n7630 ^ 1'b0 ;
  assign n35583 = n443 & ~n35582 ;
  assign n35584 = ~n1524 & n35583 ;
  assign n35585 = ( n31167 & n35581 ) | ( n31167 & ~n35584 ) | ( n35581 & ~n35584 ) ;
  assign n35586 = n12523 & ~n28340 ;
  assign n35587 = n35586 ^ n10720 ^ 1'b0 ;
  assign n35588 = n35587 ^ n2441 ^ 1'b0 ;
  assign n35589 = n1097 & n35588 ;
  assign n35590 = n17339 ^ n5116 ^ 1'b0 ;
  assign n35591 = n21789 & n35590 ;
  assign n35592 = ~n23413 & n35591 ;
  assign n35593 = n30084 ^ n15437 ^ 1'b0 ;
  assign n35594 = n34955 ^ n12698 ^ 1'b0 ;
  assign n35595 = n35594 ^ n9697 ^ x202 ;
  assign n35596 = ~n23172 & n24083 ;
  assign n35597 = n14548 ^ n2910 ^ 1'b0 ;
  assign n35598 = ~n7344 & n35597 ;
  assign n35599 = ~n9471 & n35598 ;
  assign n35600 = n22336 ^ n11007 ^ 1'b0 ;
  assign n35601 = n28169 & n35600 ;
  assign n35602 = n5418 ^ n1553 ^ 1'b0 ;
  assign n35603 = n21344 | n35602 ;
  assign n35604 = n35603 ^ n5177 ^ 1'b0 ;
  assign n35605 = ~n10252 & n35604 ;
  assign n35606 = n11781 ^ n2372 ^ 1'b0 ;
  assign n35607 = n6761 & n35606 ;
  assign n35608 = n7070 & ~n26404 ;
  assign n35609 = ~n1415 & n17263 ;
  assign n35610 = n14306 ^ n3647 ^ 1'b0 ;
  assign n35611 = ~n14533 & n24095 ;
  assign n35612 = ~n8555 & n35611 ;
  assign n35613 = ( ~n8864 & n13992 ) | ( ~n8864 & n35612 ) | ( n13992 & n35612 ) ;
  assign n35614 = n22164 & ~n35613 ;
  assign n35615 = n23978 ^ n6727 ^ 1'b0 ;
  assign n35616 = n2107 | n35615 ;
  assign n35617 = n5719 & n33303 ;
  assign n35618 = n35617 ^ n12440 ^ 1'b0 ;
  assign n35619 = ~n6045 & n26409 ;
  assign n35620 = n35619 ^ n7141 ^ 1'b0 ;
  assign n35621 = n5843 & ~n15933 ;
  assign n35622 = n25291 & n35621 ;
  assign n35623 = n4808 | n35622 ;
  assign n35624 = ~n6153 & n9651 ;
  assign n35625 = n3316 | n18642 ;
  assign n35626 = n15426 & ~n35625 ;
  assign n35627 = n35624 & ~n35626 ;
  assign n35628 = n14102 | n35627 ;
  assign n35629 = ~n6271 & n18057 ;
  assign n35630 = n35629 ^ n15128 ^ 1'b0 ;
  assign n35631 = n35076 ^ n4226 ^ n1098 ;
  assign n35632 = n11861 & ~n15276 ;
  assign n35633 = n26194 ^ n13640 ^ 1'b0 ;
  assign n35634 = n8223 & n35633 ;
  assign n35636 = ( n456 & n1855 ) | ( n456 & n9472 ) | ( n1855 & n9472 ) ;
  assign n35637 = n35636 ^ n13793 ^ n1665 ;
  assign n35638 = ( ~n2855 & n9355 ) | ( ~n2855 & n35637 ) | ( n9355 & n35637 ) ;
  assign n35635 = n7572 & ~n24661 ;
  assign n35639 = n35638 ^ n35635 ^ 1'b0 ;
  assign n35640 = ( x73 & n33226 ) | ( x73 & ~n34292 ) | ( n33226 & ~n34292 ) ;
  assign n35641 = ( ~x206 & n7842 ) | ( ~x206 & n18058 ) | ( n7842 & n18058 ) ;
  assign n35642 = n1798 & ~n13464 ;
  assign n35643 = ~n34276 & n35642 ;
  assign n35644 = n1533 | n27290 ;
  assign n35645 = n21117 & ~n35644 ;
  assign n35646 = n35645 ^ n16138 ^ 1'b0 ;
  assign n35647 = n18805 ^ n18776 ^ n15585 ;
  assign n35648 = n28917 ^ n20935 ^ 1'b0 ;
  assign n35649 = n5129 & n6276 ;
  assign n35650 = n35649 ^ n10614 ^ 1'b0 ;
  assign n35651 = n35650 ^ n6302 ^ 1'b0 ;
  assign n35652 = n10111 & n35651 ;
  assign n35653 = n6444 | n13894 ;
  assign n35654 = n35653 ^ n14842 ^ 1'b0 ;
  assign n35655 = n2151 & n20397 ;
  assign n35656 = n35655 ^ n24084 ^ 1'b0 ;
  assign n35657 = n1618 ^ n681 ^ x125 ;
  assign n35658 = n3824 | n12778 ;
  assign n35659 = n3824 & ~n35658 ;
  assign n35660 = n27085 ^ n1048 ^ 1'b0 ;
  assign n35661 = n25849 ^ n17109 ^ 1'b0 ;
  assign n35662 = n12325 ^ n9525 ^ 1'b0 ;
  assign n35663 = n10255 & n35662 ;
  assign n35664 = n3624 ^ n915 ^ 1'b0 ;
  assign n35665 = n21139 ^ n17167 ^ 1'b0 ;
  assign n35666 = n25743 ^ n13640 ^ n4599 ;
  assign n35667 = n7861 & ~n23049 ;
  assign n35668 = ( n35048 & ~n35666 ) | ( n35048 & n35667 ) | ( ~n35666 & n35667 ) ;
  assign n35669 = ( n15063 & n21899 ) | ( n15063 & ~n35168 ) | ( n21899 & ~n35168 ) ;
  assign n35670 = ( ~n1666 & n14679 ) | ( ~n1666 & n35669 ) | ( n14679 & n35669 ) ;
  assign n35671 = ~n32304 & n35670 ;
  assign n35672 = n33941 & ~n35671 ;
  assign n35673 = n25390 ^ n24972 ^ 1'b0 ;
  assign n35674 = n35673 ^ n27623 ^ 1'b0 ;
  assign n35675 = n22220 | n35674 ;
  assign n35676 = ~x233 & n33916 ;
  assign n35677 = n34750 ^ n22764 ^ n7518 ;
  assign n35678 = n35677 ^ x142 ^ 1'b0 ;
  assign n35679 = n31562 & ~n35678 ;
  assign n35680 = n35676 & n35679 ;
  assign n35682 = n4545 ^ n2085 ^ 1'b0 ;
  assign n35681 = n30548 ^ n11312 ^ n4831 ;
  assign n35683 = n35682 ^ n35681 ^ 1'b0 ;
  assign n35684 = n747 & ~n26323 ;
  assign n35685 = n10752 ^ n5052 ^ 1'b0 ;
  assign n35686 = ~n27793 & n35685 ;
  assign n35689 = n24620 ^ n4662 ^ 1'b0 ;
  assign n35690 = ( ~n18716 & n33123 ) | ( ~n18716 & n35689 ) | ( n33123 & n35689 ) ;
  assign n35687 = n5865 | n34073 ;
  assign n35688 = ~n2495 & n35687 ;
  assign n35691 = n35690 ^ n35688 ^ 1'b0 ;
  assign n35692 = ( n5549 & n7213 ) | ( n5549 & ~n18161 ) | ( n7213 & ~n18161 ) ;
  assign n35693 = n25534 | n35692 ;
  assign n35694 = ( n4899 & n12873 ) | ( n4899 & n12915 ) | ( n12873 & n12915 ) ;
  assign n35695 = n1775 & n35694 ;
  assign n35696 = ~n7812 & n17613 ;
  assign n35697 = n20439 & n27572 ;
  assign n35698 = n2384 | n8746 ;
  assign n35699 = n19113 ^ n512 ^ 1'b0 ;
  assign n35700 = n35698 | n35699 ;
  assign n35701 = n1837 & ~n2253 ;
  assign n35702 = n8011 & n17625 ;
  assign n35703 = n35702 ^ n16631 ^ 1'b0 ;
  assign n35704 = n35703 ^ n15018 ^ n11763 ;
  assign n35705 = n35704 ^ n3947 ^ 1'b0 ;
  assign n35706 = n4973 | n35705 ;
  assign n35707 = ( n9055 & ~n16435 ) | ( n9055 & n21750 ) | ( ~n16435 & n21750 ) ;
  assign n35708 = n15672 & n25593 ;
  assign n35709 = n35708 ^ n22639 ^ 1'b0 ;
  assign n35710 = ( n5812 & ~n35707 ) | ( n5812 & n35709 ) | ( ~n35707 & n35709 ) ;
  assign n35711 = n19769 ^ n6232 ^ 1'b0 ;
  assign n35712 = n5043 & n27494 ;
  assign n35713 = n35712 ^ n20165 ^ 1'b0 ;
  assign n35714 = n25186 ^ n23444 ^ 1'b0 ;
  assign n35715 = ~n18925 & n31920 ;
  assign n35716 = n4509 | n21902 ;
  assign n35717 = n3389 & ~n35716 ;
  assign n35718 = ( x160 & n32363 ) | ( x160 & n35717 ) | ( n32363 & n35717 ) ;
  assign n35719 = n16577 ^ n9598 ^ 1'b0 ;
  assign n35720 = n12774 | n35719 ;
  assign n35721 = n23024 ^ n5648 ^ 1'b0 ;
  assign n35722 = n24160 ^ n10512 ^ 1'b0 ;
  assign n35723 = n6871 | n22429 ;
  assign n35724 = n14992 & ~n35723 ;
  assign n35725 = n34857 ^ n3448 ^ 1'b0 ;
  assign n35726 = n35724 | n35725 ;
  assign n35728 = n19785 ^ n18425 ^ 1'b0 ;
  assign n35729 = ~n2274 & n35728 ;
  assign n35727 = ~n3675 & n25105 ;
  assign n35730 = n35729 ^ n35727 ^ 1'b0 ;
  assign n35731 = ( n6992 & n13155 ) | ( n6992 & n17178 ) | ( n13155 & n17178 ) ;
  assign n35732 = n16466 ^ x21 ^ 1'b0 ;
  assign n35733 = ~n9997 & n13471 ;
  assign n35734 = ~n35732 & n35733 ;
  assign n35735 = n35734 ^ n23252 ^ 1'b0 ;
  assign n35736 = n35735 ^ n20314 ^ n13877 ;
  assign n35738 = n14036 & n14181 ;
  assign n35739 = n7632 & n35738 ;
  assign n35737 = n29270 | n31817 ;
  assign n35740 = n35739 ^ n35737 ^ 1'b0 ;
  assign n35741 = x11 & n8899 ;
  assign n35742 = n35741 ^ n2826 ^ 1'b0 ;
  assign n35743 = n7748 ^ n2852 ^ 1'b0 ;
  assign n35744 = n32910 ^ n8554 ^ 1'b0 ;
  assign n35745 = n9103 | n35744 ;
  assign n35746 = n21265 | n35745 ;
  assign n35747 = n18593 | n35746 ;
  assign n35748 = n9044 & ~n14356 ;
  assign n35749 = n35748 ^ n34423 ^ 1'b0 ;
  assign n35750 = n10443 ^ n3834 ^ 1'b0 ;
  assign n35751 = n34579 & n35750 ;
  assign n35752 = n604 & n35751 ;
  assign n35753 = ~n2134 & n10780 ;
  assign n35754 = n35753 ^ n7194 ^ 1'b0 ;
  assign n35755 = ~n8560 & n35754 ;
  assign n35756 = n31948 ^ n21209 ^ n18723 ;
  assign n35757 = ( x254 & ~n634 ) | ( x254 & n4796 ) | ( ~n634 & n4796 ) ;
  assign n35758 = n27779 ^ n7512 ^ 1'b0 ;
  assign n35759 = n35758 ^ n14760 ^ 1'b0 ;
  assign n35760 = n2324 & n35759 ;
  assign n35761 = n15589 & n30225 ;
  assign n35762 = n3897 & n35761 ;
  assign n35763 = n27623 ^ n3278 ^ 1'b0 ;
  assign n35764 = n35762 | n35763 ;
  assign n35765 = n21029 & n27989 ;
  assign n35766 = n35765 ^ n6762 ^ 1'b0 ;
  assign n35767 = n35396 ^ n20605 ^ 1'b0 ;
  assign n35768 = n2164 | n19596 ;
  assign n35769 = n8903 & ~n12182 ;
  assign n35770 = n35769 ^ n25494 ^ 1'b0 ;
  assign n35771 = n35770 ^ n9508 ^ 1'b0 ;
  assign n35772 = x247 & n5065 ;
  assign n35773 = ~n671 & n35772 ;
  assign n35774 = ( ~n7824 & n34833 ) | ( ~n7824 & n35773 ) | ( n34833 & n35773 ) ;
  assign n35775 = n19606 | n26296 ;
  assign n35776 = n26600 | n35775 ;
  assign n35777 = n1653 & ~n35663 ;
  assign n35778 = n32057 ^ n6822 ^ 1'b0 ;
  assign n35779 = n13372 | n33680 ;
  assign n35780 = n35779 ^ n639 ^ 1'b0 ;
  assign n35781 = ~n22641 & n23408 ;
  assign n35782 = n35781 ^ n12344 ^ 1'b0 ;
  assign n35783 = n15389 & ~n16769 ;
  assign n35784 = n35782 & n35783 ;
  assign n35785 = n28859 ^ n23110 ^ 1'b0 ;
  assign n35786 = ~n18434 & n35785 ;
  assign n35787 = n8131 & ~n11061 ;
  assign n35788 = n22936 ^ n957 ^ x130 ;
  assign n35791 = n10068 ^ n861 ^ 1'b0 ;
  assign n35792 = ~n18975 & n35791 ;
  assign n35789 = n25105 & ~n29138 ;
  assign n35790 = n30357 & n35789 ;
  assign n35793 = n35792 ^ n35790 ^ 1'b0 ;
  assign n35794 = ( n5277 & n10272 ) | ( n5277 & n26308 ) | ( n10272 & n26308 ) ;
  assign n35795 = ( ~n13453 & n24253 ) | ( ~n13453 & n35794 ) | ( n24253 & n35794 ) ;
  assign n35796 = ~n22895 & n27207 ;
  assign n35797 = n22564 ^ n6911 ^ 1'b0 ;
  assign n35798 = n24594 & n35797 ;
  assign n35799 = n28691 | n33386 ;
  assign n35800 = n35799 ^ n5160 ^ 1'b0 ;
  assign n35801 = n21241 ^ n10322 ^ 1'b0 ;
  assign n35802 = ~n27142 & n35801 ;
  assign n35803 = n33196 ^ n25061 ^ n5323 ;
  assign n35804 = n16970 & ~n27264 ;
  assign n35805 = n35804 ^ n21383 ^ n5961 ;
  assign n35806 = ~n5552 & n17442 ;
  assign n35807 = n35806 ^ n10186 ^ 1'b0 ;
  assign n35808 = ~n2783 & n2975 ;
  assign n35809 = ~n15096 & n35808 ;
  assign n35810 = ~n11344 & n16598 ;
  assign n35811 = n3094 & n35810 ;
  assign n35812 = n12528 ^ n360 ^ 1'b0 ;
  assign n35813 = n32237 ^ n7683 ^ 1'b0 ;
  assign n35814 = ~n6884 & n28514 ;
  assign n35815 = n7758 | n20009 ;
  assign n35816 = n17402 | n35815 ;
  assign n35817 = n35816 ^ n31055 ^ n9542 ;
  assign n35818 = n3248 & ~n8728 ;
  assign n35819 = n16391 & ~n20839 ;
  assign n35820 = n14750 | n35819 ;
  assign n35821 = n35820 ^ n3136 ^ 1'b0 ;
  assign n35823 = n1667 & n29530 ;
  assign n35822 = n5876 & n15816 ;
  assign n35824 = n35823 ^ n35822 ^ 1'b0 ;
  assign n35825 = n1947 | n35824 ;
  assign n35827 = n28058 ^ n17873 ^ 1'b0 ;
  assign n35826 = n26087 ^ n18114 ^ n404 ;
  assign n35828 = n35827 ^ n35826 ^ 1'b0 ;
  assign n35829 = n21718 ^ n16142 ^ 1'b0 ;
  assign n35830 = n3490 | n8578 ;
  assign n35831 = n35830 ^ n29246 ^ 1'b0 ;
  assign n35832 = n20895 & ~n35831 ;
  assign n35833 = n27546 ^ n23147 ^ n10882 ;
  assign n35834 = n9213 & n18555 ;
  assign n35835 = n35834 ^ n5861 ^ 1'b0 ;
  assign n35836 = n14913 & n14981 ;
  assign n35837 = n35836 ^ n8989 ^ 1'b0 ;
  assign n35838 = n4806 & ~n32006 ;
  assign n35839 = n35838 ^ n3305 ^ 1'b0 ;
  assign n35840 = n26724 ^ n14530 ^ 1'b0 ;
  assign n35841 = n32697 & ~n35840 ;
  assign n35842 = n35841 ^ n25193 ^ n9559 ;
  assign n35843 = n22665 ^ n14960 ^ n5330 ;
  assign n35844 = n2207 | n35843 ;
  assign n35845 = ~n4413 & n20007 ;
  assign n35846 = n3698 & n35845 ;
  assign n35847 = n19642 & n35846 ;
  assign n35848 = n4544 & ~n35847 ;
  assign n35849 = ~n14851 & n35848 ;
  assign n35850 = n8651 ^ n7072 ^ 1'b0 ;
  assign n35851 = n610 & ~n2950 ;
  assign n35852 = ~n1233 & n35851 ;
  assign n35853 = n35852 ^ n342 ^ 1'b0 ;
  assign n35854 = n4192 | n35853 ;
  assign n35855 = n31881 & ~n35854 ;
  assign n35856 = ~n9366 & n35855 ;
  assign n35857 = n20643 ^ n4507 ^ 1'b0 ;
  assign n35858 = n8790 & ~n35857 ;
  assign n35859 = n35858 ^ n32791 ^ 1'b0 ;
  assign n35860 = n14818 ^ n11447 ^ 1'b0 ;
  assign n35861 = ( ~n27570 & n27891 ) | ( ~n27570 & n35860 ) | ( n27891 & n35860 ) ;
  assign n35862 = n2190 ^ x133 ^ 1'b0 ;
  assign n35863 = n13475 ^ n9688 ^ 1'b0 ;
  assign n35864 = n14231 ^ n1567 ^ 1'b0 ;
  assign n35865 = n15500 ^ n6206 ^ 1'b0 ;
  assign n35866 = n22789 & ~n35865 ;
  assign n35867 = n35866 ^ n1042 ^ 1'b0 ;
  assign n35868 = ~n35864 & n35867 ;
  assign n35869 = n6665 & ~n18994 ;
  assign n35870 = ~n12845 & n35869 ;
  assign n35871 = n35870 ^ n8002 ^ 1'b0 ;
  assign n35872 = n12720 ^ n10013 ^ n2033 ;
  assign n35873 = n20648 | n22103 ;
  assign n35874 = x118 & ~n9612 ;
  assign n35875 = n35874 ^ n20095 ^ 1'b0 ;
  assign n35876 = ( ~n35872 & n35873 ) | ( ~n35872 & n35875 ) | ( n35873 & n35875 ) ;
  assign n35877 = n12661 ^ n12429 ^ 1'b0 ;
  assign n35878 = n3536 | n35877 ;
  assign n35879 = ( n11692 & n12001 ) | ( n11692 & n35878 ) | ( n12001 & n35878 ) ;
  assign n35880 = n32508 ^ n8938 ^ 1'b0 ;
  assign n35881 = n26621 ^ n7559 ^ 1'b0 ;
  assign n35882 = n2548 & ~n35881 ;
  assign n35883 = n27418 ^ n19412 ^ n13404 ;
  assign n35884 = n25343 & n35883 ;
  assign n35885 = n34619 ^ n30639 ^ n7805 ;
  assign n35886 = n26779 ^ n2638 ^ 1'b0 ;
  assign n35887 = n19078 ^ n5521 ^ 1'b0 ;
  assign n35888 = n1760 & n35887 ;
  assign n35889 = ~n22753 & n35888 ;
  assign n35890 = n8427 & n35889 ;
  assign n35891 = n21903 | n35890 ;
  assign n35892 = n35891 ^ n10019 ^ 1'b0 ;
  assign n35893 = n17716 ^ n7353 ^ n2667 ;
  assign n35894 = n24153 ^ n20525 ^ 1'b0 ;
  assign n35895 = n35893 | n35894 ;
  assign n35896 = n17878 & ~n35895 ;
  assign n35897 = n2431 & n35896 ;
  assign n35898 = n29109 ^ n8901 ^ 1'b0 ;
  assign n35899 = ( n1389 & n7384 ) | ( n1389 & n15334 ) | ( n7384 & n15334 ) ;
  assign n35900 = n7674 & ~n25589 ;
  assign n35901 = n35900 ^ n10085 ^ 1'b0 ;
  assign n35902 = n12550 ^ n6683 ^ n4686 ;
  assign n35903 = n35901 | n35902 ;
  assign n35904 = n20235 | n20890 ;
  assign n35905 = ~n3954 & n21317 ;
  assign n35906 = n18410 & n35905 ;
  assign n35907 = n31742 ^ n15473 ^ n13151 ;
  assign n35908 = ( n10668 & n14419 ) | ( n10668 & ~n20285 ) | ( n14419 & ~n20285 ) ;
  assign n35909 = n19748 ^ n10612 ^ n3782 ;
  assign n35910 = n35909 ^ n33964 ^ n17557 ;
  assign n35911 = ( n26809 & ~n35908 ) | ( n26809 & n35910 ) | ( ~n35908 & n35910 ) ;
  assign n35912 = ~n315 & n4142 ;
  assign n35913 = n35912 ^ n4038 ^ 1'b0 ;
  assign n35914 = n27780 ^ n7887 ^ n4035 ;
  assign n35915 = n35914 ^ n11374 ^ 1'b0 ;
  assign n35916 = ~n27708 & n31986 ;
  assign n35917 = ( n7859 & ~n24786 ) | ( n7859 & n35916 ) | ( ~n24786 & n35916 ) ;
  assign n35918 = ~n776 & n6202 ;
  assign n35919 = n35918 ^ n5552 ^ n4015 ;
  assign n35920 = ( n7521 & n20332 ) | ( n7521 & n35919 ) | ( n20332 & n35919 ) ;
  assign n35921 = n7710 ^ n1837 ^ 1'b0 ;
  assign n35922 = ( n7152 & n35920 ) | ( n7152 & ~n35921 ) | ( n35920 & ~n35921 ) ;
  assign n35923 = n35922 ^ n23908 ^ 1'b0 ;
  assign n35924 = n34579 & ~n35923 ;
  assign n35925 = n4404 & n35924 ;
  assign n35926 = ~n6300 & n13510 ;
  assign n35927 = n35926 ^ n5915 ^ 1'b0 ;
  assign n35928 = ( n2377 & ~n13870 ) | ( n2377 & n35927 ) | ( ~n13870 & n35927 ) ;
  assign n35929 = n3577 & n3673 ;
  assign n35930 = n16949 ^ n15837 ^ 1'b0 ;
  assign n35931 = ( n529 & n35929 ) | ( n529 & ~n35930 ) | ( n35929 & ~n35930 ) ;
  assign n35932 = n16195 ^ n8311 ^ 1'b0 ;
  assign n35933 = n3123 | n35932 ;
  assign n35934 = n35933 ^ n6853 ^ 1'b0 ;
  assign n35935 = n15434 & n35934 ;
  assign n35936 = n26086 & n35935 ;
  assign n35937 = n28179 ^ n3193 ^ 1'b0 ;
  assign n35938 = n25570 & n35937 ;
  assign n35939 = n3495 & n9167 ;
  assign n35940 = n26367 ^ n24958 ^ 1'b0 ;
  assign n35941 = ( n3439 & ~n13056 ) | ( n3439 & n35940 ) | ( ~n13056 & n35940 ) ;
  assign n35942 = n19188 ^ n19019 ^ n6835 ;
  assign n35943 = ~n23142 & n32032 ;
  assign n35944 = n7457 & n35943 ;
  assign n35945 = n35944 ^ n30318 ^ 1'b0 ;
  assign n35946 = n10935 & n35945 ;
  assign n35947 = n16335 & n17481 ;
  assign n35948 = ~n14736 & n35947 ;
  assign n35949 = n3777 & ~n4751 ;
  assign n35950 = n35949 ^ n482 ^ 1'b0 ;
  assign n35951 = ~n14817 & n32953 ;
  assign n35952 = n13270 & n15813 ;
  assign n35953 = n35952 ^ n27877 ^ 1'b0 ;
  assign n35954 = ( ~n410 & n10012 ) | ( ~n410 & n10498 ) | ( n10012 & n10498 ) ;
  assign n35955 = n5961 & n35954 ;
  assign n35956 = n9946 | n33939 ;
  assign n35957 = n35956 ^ n23059 ^ 1'b0 ;
  assign n35958 = n1903 & ~n3062 ;
  assign n35959 = ~n12572 & n31705 ;
  assign n35960 = n35959 ^ n15703 ^ 1'b0 ;
  assign n35962 = n13939 ^ n7880 ^ n5869 ;
  assign n35961 = n16335 ^ x10 ^ 1'b0 ;
  assign n35963 = n35962 ^ n35961 ^ n27288 ;
  assign n35964 = ( n14969 & n35960 ) | ( n14969 & ~n35963 ) | ( n35960 & ~n35963 ) ;
  assign n35966 = n34719 ^ x188 ^ 1'b0 ;
  assign n35965 = n18462 & n22830 ;
  assign n35967 = n35966 ^ n35965 ^ n18398 ;
  assign n35968 = n14429 ^ n1194 ^ 1'b0 ;
  assign n35969 = n35968 ^ n24343 ^ n9138 ;
  assign n35970 = n31440 & n35969 ;
  assign n35971 = n35970 ^ n23614 ^ 1'b0 ;
  assign n35976 = n8330 ^ n4608 ^ 1'b0 ;
  assign n35972 = n1134 | n17518 ;
  assign n35973 = n9369 & ~n35972 ;
  assign n35974 = n35973 ^ n19758 ^ n4553 ;
  assign n35975 = n1773 & n35974 ;
  assign n35977 = n35976 ^ n35975 ^ 1'b0 ;
  assign n35978 = n6922 & n17440 ;
  assign n35979 = ~n11317 & n35978 ;
  assign n35980 = n9900 & n26843 ;
  assign n35981 = n35980 ^ n10073 ^ 1'b0 ;
  assign n35982 = n6102 & n18687 ;
  assign n35983 = ~n3992 & n35982 ;
  assign n35984 = n1350 | n18269 ;
  assign n35985 = n28724 ^ n25290 ^ n21711 ;
  assign n35986 = n26427 ^ n7796 ^ n5425 ;
  assign n35988 = n6851 & ~n7809 ;
  assign n35987 = ~n1347 & n27597 ;
  assign n35989 = n35988 ^ n35987 ^ n1194 ;
  assign n35990 = n4756 ^ n948 ^ 1'b0 ;
  assign n35991 = ~n10516 & n35990 ;
  assign n35992 = ~n10876 & n21762 ;
  assign n35993 = n35992 ^ n2444 ^ 1'b0 ;
  assign n35994 = n28863 | n35993 ;
  assign n35995 = n13499 ^ n11033 ^ 1'b0 ;
  assign n35996 = ~n2879 & n6428 ;
  assign n35997 = n35996 ^ n19689 ^ 1'b0 ;
  assign n35998 = n10504 | n17574 ;
  assign n35999 = n35997 & ~n35998 ;
  assign n36000 = n35647 | n35999 ;
  assign n36001 = n35995 & ~n36000 ;
  assign n36002 = n20057 | n22927 ;
  assign n36003 = ~n21212 & n36002 ;
  assign n36004 = ~n21041 & n36003 ;
  assign n36005 = ~n6780 & n16205 ;
  assign n36006 = n36005 ^ n33604 ^ n21862 ;
  assign n36007 = n16166 & ~n18024 ;
  assign n36008 = ( n5067 & n14846 ) | ( n5067 & ~n33059 ) | ( n14846 & ~n33059 ) ;
  assign n36009 = n31965 ^ n26319 ^ 1'b0 ;
  assign n36010 = n36008 & n36009 ;
  assign n36011 = n19616 ^ n17959 ^ n872 ;
  assign n36012 = ( n13334 & n13587 ) | ( n13334 & n36011 ) | ( n13587 & n36011 ) ;
  assign n36013 = n36012 ^ n13990 ^ 1'b0 ;
  assign n36014 = n31358 ^ n14855 ^ 1'b0 ;
  assign n36015 = n36014 ^ n2253 ^ 1'b0 ;
  assign n36016 = ~n18881 & n36015 ;
  assign n36017 = ~n16123 & n36016 ;
  assign n36018 = n32975 ^ n14075 ^ 1'b0 ;
  assign n36019 = n34764 & ~n36018 ;
  assign n36020 = n19191 & n36019 ;
  assign n36021 = n36020 ^ n19828 ^ 1'b0 ;
  assign n36022 = n16075 & ~n20797 ;
  assign n36023 = n14176 & n36022 ;
  assign n36024 = ( n23095 & ~n23330 ) | ( n23095 & n36023 ) | ( ~n23330 & n36023 ) ;
  assign n36025 = ~n1806 & n11484 ;
  assign n36026 = n36025 ^ n32405 ^ n25637 ;
  assign n36027 = n31843 ^ n3922 ^ 1'b0 ;
  assign n36028 = n9170 & ~n36027 ;
  assign n36029 = n36028 ^ n8117 ^ n840 ;
  assign n36030 = n25619 & n30236 ;
  assign n36031 = n1266 & n20287 ;
  assign n36032 = n36030 & n36031 ;
  assign n36033 = n14560 ^ n3545 ^ 1'b0 ;
  assign n36034 = ~n6348 & n36033 ;
  assign n36035 = n22614 ^ n11001 ^ 1'b0 ;
  assign n36036 = n31351 | n36035 ;
  assign n36042 = ~n13679 & n15594 ;
  assign n36043 = n36042 ^ n23277 ^ 1'b0 ;
  assign n36037 = ( x96 & n3778 ) | ( x96 & ~n12002 ) | ( n3778 & ~n12002 ) ;
  assign n36038 = n21279 ^ n4244 ^ 1'b0 ;
  assign n36039 = n36037 & n36038 ;
  assign n36040 = n11474 & n36039 ;
  assign n36041 = ~n12947 & n36040 ;
  assign n36044 = n36043 ^ n36041 ^ 1'b0 ;
  assign n36045 = n24265 ^ n22860 ^ 1'b0 ;
  assign n36046 = n7424 & n16562 ;
  assign n36047 = n14016 ^ n6136 ^ n4497 ;
  assign n36048 = n14887 | n22959 ;
  assign n36049 = ( n10506 & n36047 ) | ( n10506 & ~n36048 ) | ( n36047 & ~n36048 ) ;
  assign n36050 = n16836 ^ n6930 ^ n6257 ;
  assign n36051 = n5290 & ~n36050 ;
  assign n36053 = ~n4196 & n5490 ;
  assign n36052 = n26439 & n28704 ;
  assign n36054 = n36053 ^ n36052 ^ 1'b0 ;
  assign n36055 = n24126 ^ n546 ^ 1'b0 ;
  assign n36056 = n11974 ^ n9134 ^ 1'b0 ;
  assign n36057 = n36055 & n36056 ;
  assign n36058 = n13523 ^ n4533 ^ 1'b0 ;
  assign n36059 = ( n15219 & n21379 ) | ( n15219 & n25052 ) | ( n21379 & n25052 ) ;
  assign n36060 = ~n17480 & n33189 ;
  assign n36061 = n36059 & n36060 ;
  assign n36063 = ( n10255 & n14476 ) | ( n10255 & ~n30055 ) | ( n14476 & ~n30055 ) ;
  assign n36062 = n5685 & ~n7477 ;
  assign n36064 = n36063 ^ n36062 ^ 1'b0 ;
  assign n36065 = ( n1795 & ~n6167 ) | ( n1795 & n10970 ) | ( ~n6167 & n10970 ) ;
  assign n36066 = ~n3195 & n4342 ;
  assign n36067 = n36066 ^ n8458 ^ 1'b0 ;
  assign n36068 = ( n4281 & n6189 ) | ( n4281 & ~n36067 ) | ( n6189 & ~n36067 ) ;
  assign n36069 = n10777 & ~n30753 ;
  assign n36070 = ~n12656 & n17748 ;
  assign n36071 = n15403 | n20105 ;
  assign n36072 = ( ~n2916 & n15228 ) | ( ~n2916 & n36071 ) | ( n15228 & n36071 ) ;
  assign n36073 = n13353 | n36072 ;
  assign n36074 = ( n7675 & n10481 ) | ( n7675 & ~n28653 ) | ( n10481 & ~n28653 ) ;
  assign n36075 = ( n6015 & ~n19069 ) | ( n6015 & n33272 ) | ( ~n19069 & n33272 ) ;
  assign n36076 = n2368 & n16170 ;
  assign n36077 = ~n2368 & n36076 ;
  assign n36078 = n1782 | n1890 ;
  assign n36079 = n1890 & ~n36078 ;
  assign n36080 = ~n2921 & n36079 ;
  assign n36081 = n36077 | n36080 ;
  assign n36082 = n36077 & ~n36081 ;
  assign n36083 = n24272 | n36082 ;
  assign n36084 = n26125 & ~n36083 ;
  assign n36085 = n15030 ^ n3462 ^ 1'b0 ;
  assign n36086 = n21983 & ~n36085 ;
  assign n36087 = ~n14110 & n36086 ;
  assign n36088 = n21406 ^ n13902 ^ n4709 ;
  assign n36089 = n34272 ^ n16416 ^ 1'b0 ;
  assign n36090 = n14650 ^ n7180 ^ 1'b0 ;
  assign n36091 = n36090 ^ n3696 ^ 1'b0 ;
  assign n36092 = n25433 & n25637 ;
  assign n36093 = n31037 & ~n33391 ;
  assign n36094 = n2076 | n6818 ;
  assign n36095 = n36094 ^ n10112 ^ 1'b0 ;
  assign n36096 = n10159 & ~n36095 ;
  assign n36097 = n16619 ^ n13873 ^ x117 ;
  assign n36098 = ( ~n2066 & n28951 ) | ( ~n2066 & n36097 ) | ( n28951 & n36097 ) ;
  assign n36099 = n11767 & n15027 ;
  assign n36100 = n28155 & n36099 ;
  assign n36101 = n15486 | n23221 ;
  assign n36102 = n14362 & n33051 ;
  assign n36103 = n15626 & ~n33409 ;
  assign n36104 = n36103 ^ n19438 ^ 1'b0 ;
  assign n36105 = ( ~n4710 & n8860 ) | ( ~n4710 & n9097 ) | ( n8860 & n9097 ) ;
  assign n36106 = ~n5772 & n19889 ;
  assign n36107 = n3030 & n36106 ;
  assign n36108 = n36107 ^ n10614 ^ 1'b0 ;
  assign n36109 = n36105 | n36108 ;
  assign n36110 = ~n13052 & n21411 ;
  assign n36111 = n36110 ^ n8077 ^ n1589 ;
  assign n36112 = n6038 ^ n2782 ^ 1'b0 ;
  assign n36113 = n527 & ~n36112 ;
  assign n36114 = ( n28385 & n30866 ) | ( n28385 & n36113 ) | ( n30866 & n36113 ) ;
  assign n36115 = n10665 ^ n2741 ^ 1'b0 ;
  assign n36116 = n36115 ^ n14868 ^ n5327 ;
  assign n36117 = n21630 ^ n14338 ^ 1'b0 ;
  assign n36118 = n12500 ^ n991 ^ 1'b0 ;
  assign n36119 = n36118 ^ n11032 ^ 1'b0 ;
  assign n36120 = n22856 & ~n36119 ;
  assign n36125 = n25753 ^ n22997 ^ 1'b0 ;
  assign n36121 = n12097 ^ n5542 ^ 1'b0 ;
  assign n36122 = n4282 & ~n36121 ;
  assign n36123 = n36122 ^ n23490 ^ 1'b0 ;
  assign n36124 = n5483 & n36123 ;
  assign n36126 = n36125 ^ n36124 ^ 1'b0 ;
  assign n36127 = ~n2360 & n15807 ;
  assign n36128 = n36127 ^ n19623 ^ 1'b0 ;
  assign n36129 = n36128 ^ n1263 ^ 1'b0 ;
  assign n36130 = n13678 ^ n4905 ^ n4481 ;
  assign n36131 = n13844 | n36130 ;
  assign n36132 = n36131 ^ n14968 ^ 1'b0 ;
  assign n36133 = n1510 & n36132 ;
  assign n36134 = n1501 | n19735 ;
  assign n36135 = n25498 ^ n9798 ^ 1'b0 ;
  assign n36136 = n17504 ^ n11459 ^ 1'b0 ;
  assign n36137 = n5182 & n36136 ;
  assign n36138 = n36137 ^ n17486 ^ 1'b0 ;
  assign n36139 = n9042 ^ n6327 ^ 1'b0 ;
  assign n36140 = n36139 ^ n2507 ^ 1'b0 ;
  assign n36141 = ~n6022 & n36140 ;
  assign n36142 = n12223 & n36141 ;
  assign n36143 = n36142 ^ n25661 ^ 1'b0 ;
  assign n36144 = n5013 & ~n27027 ;
  assign n36145 = ~n27117 & n36144 ;
  assign n36146 = n10412 ^ n4347 ^ 1'b0 ;
  assign n36147 = n8453 | n36146 ;
  assign n36148 = n28653 ^ n3096 ^ 1'b0 ;
  assign n36149 = n9752 & n36148 ;
  assign n36150 = n8408 | n29971 ;
  assign n36151 = n15341 & n36150 ;
  assign n36152 = n36151 ^ n22234 ^ 1'b0 ;
  assign n36153 = n7158 ^ x199 ^ 1'b0 ;
  assign n36154 = ~n2910 & n36153 ;
  assign n36155 = n4503 & n36154 ;
  assign n36156 = n36155 ^ n32213 ^ 1'b0 ;
  assign n36157 = n7843 & n28191 ;
  assign n36158 = n30243 & n36157 ;
  assign n36159 = ( ~x215 & n23510 ) | ( ~x215 & n26158 ) | ( n23510 & n26158 ) ;
  assign n36160 = ( n8167 & n15168 ) | ( n8167 & n36159 ) | ( n15168 & n36159 ) ;
  assign n36161 = n4910 ^ n1802 ^ 1'b0 ;
  assign n36162 = n4582 | n21216 ;
  assign n36163 = n31729 | n36162 ;
  assign n36164 = n11521 ^ n669 ^ 1'b0 ;
  assign n36165 = n34969 ^ n665 ^ 1'b0 ;
  assign n36166 = n36164 | n36165 ;
  assign n36167 = n1767 & ~n12885 ;
  assign n36168 = n36167 ^ n27058 ^ 1'b0 ;
  assign n36169 = n3333 & ~n36168 ;
  assign n36170 = n3666 | n13584 ;
  assign n36171 = ( n795 & ~n21991 ) | ( n795 & n36170 ) | ( ~n21991 & n36170 ) ;
  assign n36172 = n36171 ^ n15031 ^ 1'b0 ;
  assign n36173 = n36169 & ~n36172 ;
  assign n36174 = n16435 ^ n4993 ^ n3752 ;
  assign n36175 = ( n9369 & ~n19689 ) | ( n9369 & n33102 ) | ( ~n19689 & n33102 ) ;
  assign n36176 = n24114 ^ n20297 ^ 1'b0 ;
  assign n36177 = n18694 & ~n36176 ;
  assign n36178 = n35584 & n36177 ;
  assign n36179 = ~n14470 & n36178 ;
  assign n36180 = ~n1969 & n2993 ;
  assign n36181 = n13864 ^ n8944 ^ 1'b0 ;
  assign n36182 = ~n36180 & n36181 ;
  assign n36183 = n27812 ^ n11235 ^ 1'b0 ;
  assign n36184 = ~n28745 & n36183 ;
  assign n36185 = n2096 ^ n1302 ^ 1'b0 ;
  assign n36186 = ~n5725 & n36185 ;
  assign n36187 = n36186 ^ n6827 ^ 1'b0 ;
  assign n36188 = n26571 ^ n9398 ^ n9273 ;
  assign n36189 = n17238 ^ n12754 ^ n9529 ;
  assign n36190 = n36188 & n36189 ;
  assign n36191 = ~n36187 & n36190 ;
  assign n36192 = n17032 & ~n21472 ;
  assign n36193 = n36191 & n36192 ;
  assign n36194 = ~n23088 & n24025 ;
  assign n36195 = n23307 ^ n21316 ^ 1'b0 ;
  assign n36196 = ( n4652 & ~n9014 ) | ( n4652 & n32397 ) | ( ~n9014 & n32397 ) ;
  assign n36197 = n3826 & ~n36196 ;
  assign n36198 = ~x183 & n23747 ;
  assign n36199 = n2701 & ~n3881 ;
  assign n36200 = ~n8663 & n36199 ;
  assign n36201 = n23841 ^ n23706 ^ 1'b0 ;
  assign n36202 = ~n10715 & n36201 ;
  assign n36203 = n3144 & ~n36202 ;
  assign n36204 = n15676 & ~n24131 ;
  assign n36205 = n3328 & n36204 ;
  assign n36207 = n19930 ^ n1191 ^ 1'b0 ;
  assign n36208 = n4758 & n36207 ;
  assign n36206 = n26088 ^ n2155 ^ 1'b0 ;
  assign n36209 = n36208 ^ n36206 ^ 1'b0 ;
  assign n36210 = ~n19364 & n31093 ;
  assign n36211 = n9605 | n32858 ;
  assign n36212 = n10445 & n27245 ;
  assign n36213 = ~n36211 & n36212 ;
  assign n36214 = n29469 ^ n8344 ^ 1'b0 ;
  assign n36215 = n1129 | n29254 ;
  assign n36216 = n36215 ^ n17518 ^ 1'b0 ;
  assign n36217 = ~x58 & n13770 ;
  assign n36218 = n26039 ^ n610 ^ 1'b0 ;
  assign n36219 = n10326 | n36218 ;
  assign n36220 = n25965 ^ n25343 ^ 1'b0 ;
  assign n36221 = n18454 | n33106 ;
  assign n36222 = n19650 & ~n27572 ;
  assign n36223 = n30114 ^ n2144 ^ 1'b0 ;
  assign n36224 = ~n31710 & n36223 ;
  assign n36225 = n11586 ^ n1853 ^ 1'b0 ;
  assign n36226 = n4165 & ~n36225 ;
  assign n36227 = n8225 ^ n1313 ^ 1'b0 ;
  assign n36228 = n17467 & n36227 ;
  assign n36232 = ~n3746 & n11060 ;
  assign n36229 = n10658 & ~n30797 ;
  assign n36230 = n11667 & ~n36229 ;
  assign n36231 = n19562 & n36230 ;
  assign n36233 = n36232 ^ n36231 ^ 1'b0 ;
  assign n36234 = n25123 ^ n20098 ^ 1'b0 ;
  assign n36235 = n10457 | n31289 ;
  assign n36236 = n36235 ^ n9965 ^ 1'b0 ;
  assign n36237 = n17304 & n28614 ;
  assign n36238 = ~x3 & n36237 ;
  assign n36239 = ( ~n5690 & n7377 ) | ( ~n5690 & n8941 ) | ( n7377 & n8941 ) ;
  assign n36240 = n5279 & n23652 ;
  assign n36241 = ~n36239 & n36240 ;
  assign n36242 = n36241 ^ n2925 ^ 1'b0 ;
  assign n36243 = n36238 | n36242 ;
  assign n36244 = n6259 | n32495 ;
  assign n36245 = n31722 ^ n11348 ^ 1'b0 ;
  assign n36246 = ~n20233 & n36245 ;
  assign n36247 = n26899 ^ n14105 ^ 1'b0 ;
  assign n36248 = n16900 & ~n20850 ;
  assign n36249 = n36248 ^ n16420 ^ 1'b0 ;
  assign n36250 = n7113 & ~n36249 ;
  assign n36251 = n36247 & n36250 ;
  assign n36252 = n19419 & ~n36251 ;
  assign n36253 = ~n6849 & n36252 ;
  assign n36254 = n16417 & n28692 ;
  assign n36258 = n12752 | n18835 ;
  assign n36259 = n18498 | n36258 ;
  assign n36256 = n5661 ^ n1388 ^ 1'b0 ;
  assign n36257 = n12661 | n36256 ;
  assign n36260 = n36259 ^ n36257 ^ 1'b0 ;
  assign n36255 = n6022 | n8584 ;
  assign n36261 = n36260 ^ n36255 ^ 1'b0 ;
  assign n36262 = n32801 ^ n6359 ^ 1'b0 ;
  assign n36263 = ( ~n36254 & n36261 ) | ( ~n36254 & n36262 ) | ( n36261 & n36262 ) ;
  assign n36264 = n26425 ^ n1595 ^ 1'b0 ;
  assign n36265 = ~n18272 & n21054 ;
  assign n36266 = ~n3015 & n16902 ;
  assign n36267 = ~n36265 & n36266 ;
  assign n36268 = ~n9493 & n22048 ;
  assign n36269 = n8490 & n36268 ;
  assign n36270 = n19650 | n34000 ;
  assign n36271 = n36269 & ~n36270 ;
  assign n36272 = n2475 | n3574 ;
  assign n36273 = n7870 & n36272 ;
  assign n36274 = n11426 & n36273 ;
  assign n36275 = n28526 | n36274 ;
  assign n36276 = n36275 ^ n10569 ^ 1'b0 ;
  assign n36277 = ~n8356 & n10351 ;
  assign n36278 = n18804 | n34871 ;
  assign n36279 = n36278 ^ n12590 ^ 1'b0 ;
  assign n36280 = ( n933 & n13896 ) | ( n933 & ~n32197 ) | ( n13896 & ~n32197 ) ;
  assign n36282 = n25436 & n27266 ;
  assign n36283 = n36282 ^ n6384 ^ 1'b0 ;
  assign n36281 = n16838 ^ n7745 ^ n7283 ;
  assign n36284 = n36283 ^ n36281 ^ n10419 ;
  assign n36285 = n11145 ^ n698 ^ 1'b0 ;
  assign n36286 = n472 & n12279 ;
  assign n36287 = n24119 ^ n3767 ^ 1'b0 ;
  assign n36288 = n13787 | n36287 ;
  assign n36289 = n14435 ^ n6630 ^ 1'b0 ;
  assign n36290 = ~n36288 & n36289 ;
  assign n36291 = n12902 ^ n10702 ^ n6260 ;
  assign n36292 = n9805 | n11298 ;
  assign n36293 = n36291 | n36292 ;
  assign n36294 = n3453 & n10749 ;
  assign n36295 = ( ~n11438 & n16579 ) | ( ~n11438 & n36294 ) | ( n16579 & n36294 ) ;
  assign n36296 = ( n2523 & n8884 ) | ( n2523 & ~n34793 ) | ( n8884 & ~n34793 ) ;
  assign n36297 = n36296 ^ n30524 ^ n2253 ;
  assign n36298 = n2147 & n22814 ;
  assign n36299 = n13884 & n36298 ;
  assign n36300 = ( n23172 & n36297 ) | ( n23172 & n36299 ) | ( n36297 & n36299 ) ;
  assign n36301 = ( n1279 & n5067 ) | ( n1279 & n29404 ) | ( n5067 & n29404 ) ;
  assign n36302 = ~n4588 & n8794 ;
  assign n36303 = n30812 ^ n919 ^ 1'b0 ;
  assign n36304 = n1666 & ~n7465 ;
  assign n36305 = n36304 ^ n11880 ^ 1'b0 ;
  assign n36306 = ~n704 & n3365 ;
  assign n36307 = ~n36305 & n36306 ;
  assign n36308 = n7101 | n9134 ;
  assign n36309 = ~n11933 & n16405 ;
  assign n36310 = n27056 & n36309 ;
  assign n36313 = n8106 | n13902 ;
  assign n36311 = n13297 & n26083 ;
  assign n36312 = n6108 & n36311 ;
  assign n36314 = n36313 ^ n36312 ^ 1'b0 ;
  assign n36315 = n9731 ^ x183 ^ 1'b0 ;
  assign n36316 = n3175 & n36315 ;
  assign n36317 = n34608 & n36316 ;
  assign n36319 = n18864 & ~n24765 ;
  assign n36320 = ~n12522 & n36319 ;
  assign n36318 = ~n5051 & n21011 ;
  assign n36321 = n36320 ^ n36318 ^ 1'b0 ;
  assign n36322 = ~n6309 & n36321 ;
  assign n36323 = n23032 ^ n4634 ^ 1'b0 ;
  assign n36324 = n8913 & n36323 ;
  assign n36325 = n20673 ^ n13604 ^ 1'b0 ;
  assign n36326 = ~n28890 & n36325 ;
  assign n36327 = n673 & n27110 ;
  assign n36328 = n29476 & n30501 ;
  assign n36329 = n3506 & n36328 ;
  assign n36330 = n28445 | n36329 ;
  assign n36331 = n36330 ^ n10468 ^ 1'b0 ;
  assign n36332 = n3871 ^ x33 ^ 1'b0 ;
  assign n36333 = ~n12034 & n13921 ;
  assign n36334 = n1680 & n36333 ;
  assign n36335 = n35845 ^ n9286 ^ 1'b0 ;
  assign n36336 = ~n3257 & n36335 ;
  assign n36337 = n36336 ^ n16483 ^ n14272 ;
  assign n36338 = ( n3068 & ~n10293 ) | ( n3068 & n36337 ) | ( ~n10293 & n36337 ) ;
  assign n36339 = n36338 ^ n7609 ^ 1'b0 ;
  assign n36340 = n23908 ^ n3604 ^ 1'b0 ;
  assign n36341 = ~n15567 & n20932 ;
  assign n36342 = ~n36340 & n36341 ;
  assign n36343 = n23305 ^ n22191 ^ 1'b0 ;
  assign n36344 = ~n32519 & n36343 ;
  assign n36345 = n36344 ^ n15703 ^ 1'b0 ;
  assign n36346 = n19021 ^ n10126 ^ 1'b0 ;
  assign n36349 = ~n3958 & n20757 ;
  assign n36347 = n9521 & ~n24819 ;
  assign n36348 = ~n7544 & n36347 ;
  assign n36350 = n36349 ^ n36348 ^ 1'b0 ;
  assign n36351 = n14100 & ~n19218 ;
  assign n36352 = n10516 ^ n3630 ^ 1'b0 ;
  assign n36353 = n12704 & n36352 ;
  assign n36354 = n17506 & ~n24293 ;
  assign n36355 = ~n15793 & n36354 ;
  assign n36356 = n6257 | n36355 ;
  assign n36357 = n6102 & ~n6327 ;
  assign n36358 = n360 & n11845 ;
  assign n36359 = n10245 ^ n1783 ^ n527 ;
  assign n36360 = n7629 & ~n31608 ;
  assign n36361 = n36360 ^ n18752 ^ 1'b0 ;
  assign n36362 = ~n36359 & n36361 ;
  assign n36363 = n29534 ^ n5832 ^ 1'b0 ;
  assign n36364 = n1269 & n36363 ;
  assign n36365 = n1911 | n28982 ;
  assign n36366 = n3947 | n29515 ;
  assign n36367 = n22140 | n24833 ;
  assign n36368 = n12074 ^ n1122 ^ 1'b0 ;
  assign n36369 = n22732 ^ n17270 ^ 1'b0 ;
  assign n36370 = ~n2345 & n36369 ;
  assign n36371 = n20392 | n22422 ;
  assign n36372 = n36371 ^ n20075 ^ 1'b0 ;
  assign n36373 = n19639 ^ n19200 ^ n5202 ;
  assign n36374 = n2714 | n32354 ;
  assign n36375 = n13774 & ~n33910 ;
  assign n36376 = n269 & ~n1053 ;
  assign n36377 = n36376 ^ n32310 ^ n14572 ;
  assign n36378 = n30944 | n36377 ;
  assign n36379 = n18303 ^ n18081 ^ n8577 ;
  assign n36381 = ( ~n6365 & n9246 ) | ( ~n6365 & n13780 ) | ( n9246 & n13780 ) ;
  assign n36380 = n19316 ^ n14285 ^ 1'b0 ;
  assign n36382 = n36381 ^ n36380 ^ n1285 ;
  assign n36383 = n12190 & ~n36382 ;
  assign n36384 = n3441 | n11674 ;
  assign n36385 = n20509 ^ n1000 ^ 1'b0 ;
  assign n36386 = n35479 & n36385 ;
  assign n36387 = n27583 ^ n21251 ^ n16702 ;
  assign n36388 = n21903 ^ n19713 ^ 1'b0 ;
  assign n36389 = ~n6993 & n12131 ;
  assign n36390 = n36389 ^ n21253 ^ 1'b0 ;
  assign n36391 = ( n668 & n16445 ) | ( n668 & n36390 ) | ( n16445 & n36390 ) ;
  assign n36392 = n1450 & n18918 ;
  assign n36393 = n31671 ^ n9702 ^ n1033 ;
  assign n36394 = ( n32348 & n32903 ) | ( n32348 & ~n36393 ) | ( n32903 & ~n36393 ) ;
  assign n36395 = ~n35898 & n36394 ;
  assign n36396 = n10686 & n36395 ;
  assign n36401 = n2390 & ~n13939 ;
  assign n36397 = n8246 & ~n28906 ;
  assign n36398 = n12917 & n36397 ;
  assign n36399 = ( n7826 & n28516 ) | ( n7826 & ~n30196 ) | ( n28516 & ~n30196 ) ;
  assign n36400 = n36398 | n36399 ;
  assign n36402 = n36401 ^ n36400 ^ 1'b0 ;
  assign n36403 = n5620 ^ n979 ^ 1'b0 ;
  assign n36404 = n36403 ^ n9867 ^ 1'b0 ;
  assign n36405 = n5404 & n24689 ;
  assign n36406 = ~n15144 & n17974 ;
  assign n36407 = n36406 ^ n8645 ^ 1'b0 ;
  assign n36408 = n15825 ^ n12065 ^ 1'b0 ;
  assign n36409 = n6874 & ~n36408 ;
  assign n36410 = n10334 ^ n9373 ^ 1'b0 ;
  assign n36411 = ~n11809 & n36410 ;
  assign n36412 = x169 & ~n36411 ;
  assign n36413 = n36409 & n36412 ;
  assign n36414 = n32183 ^ n26898 ^ 1'b0 ;
  assign n36415 = n1339 & ~n31299 ;
  assign n36416 = n4222 & ~n7714 ;
  assign n36417 = n6188 & ~n25766 ;
  assign n36418 = n36416 | n36417 ;
  assign n36419 = n3913 & ~n36418 ;
  assign n36420 = n10391 ^ n7781 ^ 1'b0 ;
  assign n36421 = ~n33307 & n36420 ;
  assign n36422 = n488 & ~n18083 ;
  assign n36425 = n18893 | n24647 ;
  assign n36423 = n11631 ^ n8105 ^ 1'b0 ;
  assign n36424 = n12548 & n36423 ;
  assign n36426 = n36425 ^ n36424 ^ 1'b0 ;
  assign n36427 = n28626 ^ n20980 ^ n1489 ;
  assign n36429 = n14100 | n18804 ;
  assign n36430 = ~n23511 & n36429 ;
  assign n36428 = ~n745 & n35161 ;
  assign n36431 = n36430 ^ n36428 ^ 1'b0 ;
  assign n36432 = ~n1304 & n6607 ;
  assign n36433 = n36432 ^ n12119 ^ 1'b0 ;
  assign n36434 = n36433 ^ n30264 ^ 1'b0 ;
  assign n36435 = n13637 & n36434 ;
  assign n36436 = n6491 & ~n21082 ;
  assign n36437 = n34419 ^ n8368 ^ n3960 ;
  assign n36438 = n5415 & n11864 ;
  assign n36439 = n10801 & n36438 ;
  assign n36440 = n36439 ^ n34435 ^ n6961 ;
  assign n36441 = n2466 & n28492 ;
  assign n36442 = n36441 ^ n11537 ^ 1'b0 ;
  assign n36443 = n26886 ^ n3052 ^ 1'b0 ;
  assign n36444 = n4509 & n36443 ;
  assign n36445 = n23845 & n36444 ;
  assign n36446 = n10963 ^ n9207 ^ 1'b0 ;
  assign n36447 = n11236 & n36446 ;
  assign n36448 = n1168 ^ n393 ^ 1'b0 ;
  assign n36449 = n36448 ^ n14740 ^ 1'b0 ;
  assign n36450 = n36447 & n36449 ;
  assign n36451 = n704 & n36450 ;
  assign n36452 = ~n22047 & n36451 ;
  assign n36453 = n5543 ^ x71 ^ 1'b0 ;
  assign n36454 = n32325 | n34133 ;
  assign n36455 = n36454 ^ n24370 ^ 1'b0 ;
  assign n36456 = n26364 ^ n23520 ^ n4816 ;
  assign n36457 = n25944 ^ n8290 ^ 1'b0 ;
  assign n36458 = n21156 ^ n10982 ^ 1'b0 ;
  assign n36459 = n3489 & n14936 ;
  assign n36460 = n29201 & n29375 ;
  assign n36461 = n2253 & n36460 ;
  assign n36462 = n11564 & ~n14489 ;
  assign n36463 = n269 & ~n1384 ;
  assign n36464 = n6153 & ~n36463 ;
  assign n36465 = n18373 ^ n11297 ^ 1'b0 ;
  assign n36466 = n30606 & ~n34283 ;
  assign n36467 = n20684 ^ n16807 ^ 1'b0 ;
  assign n36470 = n4274 & ~n15316 ;
  assign n36471 = n36470 ^ n18728 ^ 1'b0 ;
  assign n36468 = n1168 | n4094 ;
  assign n36469 = n17128 | n36468 ;
  assign n36472 = n36471 ^ n36469 ^ n674 ;
  assign n36473 = ~n31073 & n36472 ;
  assign n36474 = n36473 ^ n15355 ^ 1'b0 ;
  assign n36475 = n14321 ^ n10331 ^ 1'b0 ;
  assign n36476 = n17125 ^ n16508 ^ 1'b0 ;
  assign n36477 = n13423 & ~n36476 ;
  assign n36478 = n4880 | n22671 ;
  assign n36479 = n36477 | n36478 ;
  assign n36480 = n5449 ^ n2532 ^ 1'b0 ;
  assign n36481 = n36480 ^ n17508 ^ 1'b0 ;
  assign n36482 = n12578 | n36481 ;
  assign n36483 = ( n7877 & n18034 ) | ( n7877 & ~n36482 ) | ( n18034 & ~n36482 ) ;
  assign n36484 = n1665 & n9072 ;
  assign n36485 = n36484 ^ n5912 ^ 1'b0 ;
  assign n36486 = n36485 ^ n4738 ^ 1'b0 ;
  assign n36487 = n13475 ^ n9800 ^ 1'b0 ;
  assign n36488 = n17959 | n29937 ;
  assign n36489 = n36488 ^ n14472 ^ 1'b0 ;
  assign n36490 = n28618 & n36489 ;
  assign n36491 = n25651 ^ n10664 ^ 1'b0 ;
  assign n36492 = n29754 ^ n17852 ^ n8171 ;
  assign n36493 = n24169 & n32545 ;
  assign n36494 = ~x4 & n36493 ;
  assign n36495 = n36492 | n36494 ;
  assign n36496 = n36495 ^ n3659 ^ 1'b0 ;
  assign n36498 = n10471 ^ n2418 ^ 1'b0 ;
  assign n36499 = x219 & n36498 ;
  assign n36497 = n30067 ^ n15881 ^ n7010 ;
  assign n36500 = n36499 ^ n36497 ^ 1'b0 ;
  assign n36501 = n32314 ^ n5671 ^ 1'b0 ;
  assign n36502 = n13806 ^ n6141 ^ n3830 ;
  assign n36503 = n36502 ^ n16438 ^ 1'b0 ;
  assign n36504 = ( n7701 & n10088 ) | ( n7701 & ~n28297 ) | ( n10088 & ~n28297 ) ;
  assign n36505 = n36504 ^ n16722 ^ n5830 ;
  assign n36506 = n12180 | n14043 ;
  assign n36507 = n36506 ^ n7048 ^ 1'b0 ;
  assign n36508 = n4383 ^ n3728 ^ 1'b0 ;
  assign n36509 = n36507 | n36508 ;
  assign n36510 = n32848 ^ n30382 ^ 1'b0 ;
  assign n36511 = n8630 & ~n10527 ;
  assign n36512 = n36511 ^ n8667 ^ 1'b0 ;
  assign n36513 = n302 & n1486 ;
  assign n36514 = n14320 & n36513 ;
  assign n36515 = n30601 & n36514 ;
  assign n36516 = n8384 & ~n29490 ;
  assign n36517 = ~n27665 & n36516 ;
  assign n36518 = n947 & ~n21912 ;
  assign n36519 = n36518 ^ n18311 ^ 1'b0 ;
  assign n36520 = ( n4879 & n6548 ) | ( n4879 & n34825 ) | ( n6548 & n34825 ) ;
  assign n36521 = n36520 ^ n31592 ^ 1'b0 ;
  assign n36522 = n32126 & n36521 ;
  assign n36523 = n3979 | n6838 ;
  assign n36524 = n36523 ^ n535 ^ 1'b0 ;
  assign n36525 = n36524 ^ n17964 ^ 1'b0 ;
  assign n36526 = n11338 ^ n4770 ^ 1'b0 ;
  assign n36527 = ~n4915 & n36526 ;
  assign n36528 = n1773 & n36527 ;
  assign n36529 = n20281 & n36528 ;
  assign n36530 = n7070 & ~n8765 ;
  assign n36531 = n36530 ^ n6232 ^ 1'b0 ;
  assign n36532 = n18488 ^ n3325 ^ 1'b0 ;
  assign n36533 = n960 & n12333 ;
  assign n36534 = n36532 & ~n36533 ;
  assign n36535 = n12805 & ~n35637 ;
  assign n36536 = n30092 & ~n31161 ;
  assign n36537 = n16729 ^ n15717 ^ n11122 ;
  assign n36538 = n36537 ^ n35811 ^ 1'b0 ;
  assign n36539 = n8549 | n16731 ;
  assign n36540 = n36539 ^ n33927 ^ n24625 ;
  assign n36541 = n12268 ^ n3920 ^ 1'b0 ;
  assign n36542 = ( ~n8306 & n26509 ) | ( ~n8306 & n36541 ) | ( n26509 & n36541 ) ;
  assign n36543 = n14510 | n28353 ;
  assign n36544 = n36543 ^ n27738 ^ 1'b0 ;
  assign n36545 = n21357 & ~n23050 ;
  assign n36546 = ~n10488 & n18528 ;
  assign n36547 = ~n18506 & n36546 ;
  assign n36548 = n22453 ^ n16100 ^ 1'b0 ;
  assign n36549 = ~n9029 & n11706 ;
  assign n36550 = n36548 & n36549 ;
  assign n36551 = n36550 ^ n18214 ^ 1'b0 ;
  assign n36552 = ~n35300 & n36551 ;
  assign n36553 = n5400 | n26581 ;
  assign n36554 = n5544 & ~n36553 ;
  assign n36555 = n9459 & n15070 ;
  assign n36556 = n24267 ^ n22182 ^ 1'b0 ;
  assign n36557 = n36555 & ~n36556 ;
  assign n36558 = n6539 ^ n5658 ^ 1'b0 ;
  assign n36559 = n5543 & n36558 ;
  assign n36560 = n36559 ^ n3520 ^ n637 ;
  assign n36561 = n23677 & ~n31093 ;
  assign n36562 = ~n571 & n14394 ;
  assign n36563 = n17392 & ~n32555 ;
  assign n36564 = n1564 | n36563 ;
  assign n36565 = n36564 ^ n20067 ^ 1'b0 ;
  assign n36566 = n36565 ^ n14314 ^ 1'b0 ;
  assign n36568 = n17009 & n33688 ;
  assign n36567 = n21053 ^ n4731 ^ 1'b0 ;
  assign n36569 = n36568 ^ n36567 ^ n31123 ;
  assign n36571 = n3635 | n4086 ;
  assign n36572 = n36571 ^ n2158 ^ 1'b0 ;
  assign n36570 = n10091 & n19927 ;
  assign n36573 = n36572 ^ n36570 ^ n29135 ;
  assign n36574 = n16987 & ~n26961 ;
  assign n36575 = n36574 ^ n23716 ^ 1'b0 ;
  assign n36576 = ~n2481 & n8632 ;
  assign n36577 = ~n36575 & n36576 ;
  assign n36578 = n24117 & n29942 ;
  assign n36579 = n36578 ^ n6910 ^ 1'b0 ;
  assign n36580 = n9713 ^ n5142 ^ 1'b0 ;
  assign n36581 = n32070 & n36580 ;
  assign n36582 = n23289 ^ n19210 ^ 1'b0 ;
  assign n36583 = n6110 ^ n5367 ^ n2132 ;
  assign n36584 = ( n1024 & n15388 ) | ( n1024 & n16213 ) | ( n15388 & n16213 ) ;
  assign n36585 = n20233 & ~n29921 ;
  assign n36586 = ( n5817 & ~n36584 ) | ( n5817 & n36585 ) | ( ~n36584 & n36585 ) ;
  assign n36587 = ~n12344 & n19639 ;
  assign n36588 = n36587 ^ n25230 ^ 1'b0 ;
  assign n36589 = n5993 & n36588 ;
  assign n36590 = n5313 ^ n1125 ^ 1'b0 ;
  assign n36591 = ~n27701 & n36590 ;
  assign n36592 = n36591 ^ n1929 ^ 1'b0 ;
  assign n36593 = ~n3164 & n31973 ;
  assign n36594 = n3899 & n18955 ;
  assign n36595 = n2061 & n36594 ;
  assign n36596 = n8813 ^ n1673 ^ n913 ;
  assign n36597 = n14016 ^ n2285 ^ 1'b0 ;
  assign n36598 = n6272 & ~n36597 ;
  assign n36599 = n3976 & ~n28102 ;
  assign n36600 = n36599 ^ n1015 ^ 1'b0 ;
  assign n36601 = ~n660 & n36600 ;
  assign n36602 = n1430 | n8634 ;
  assign n36603 = n340 & n9260 ;
  assign n36604 = n36603 ^ n35682 ^ 1'b0 ;
  assign n36605 = n35418 ^ n18143 ^ 1'b0 ;
  assign n36606 = n14675 ^ n5277 ^ 1'b0 ;
  assign n36607 = n11434 ^ n4812 ^ 1'b0 ;
  assign n36608 = n34660 ^ n12344 ^ 1'b0 ;
  assign n36609 = x241 | n36608 ;
  assign n36610 = ( n32116 & ~n36607 ) | ( n32116 & n36609 ) | ( ~n36607 & n36609 ) ;
  assign n36611 = n8775 | n22945 ;
  assign n36612 = n11043 & ~n36611 ;
  assign n36613 = n31684 ^ n29914 ^ 1'b0 ;
  assign n36614 = n18451 ^ n13679 ^ n8759 ;
  assign n36615 = n4752 ^ n2234 ^ 1'b0 ;
  assign n36616 = ~n13048 & n36615 ;
  assign n36617 = n11842 & ~n22621 ;
  assign n36618 = n3938 & ~n36617 ;
  assign n36619 = n1991 & n3767 ;
  assign n36620 = n36619 ^ n34295 ^ 1'b0 ;
  assign n36621 = n12733 & ~n14495 ;
  assign n36622 = n1258 | n8064 ;
  assign n36623 = ~n21523 & n36622 ;
  assign n36624 = n27444 & n36623 ;
  assign n36625 = n30063 ^ n20165 ^ n6971 ;
  assign n36626 = n24997 ^ n24340 ^ n1212 ;
  assign n36627 = n25986 ^ n17304 ^ n2212 ;
  assign n36629 = n6831 & ~n15724 ;
  assign n36628 = n7641 & ~n12394 ;
  assign n36630 = n36629 ^ n36628 ^ 1'b0 ;
  assign n36631 = x17 | n31747 ;
  assign n36632 = n1380 | n36631 ;
  assign n36633 = ~n2002 & n36632 ;
  assign n36634 = n36633 ^ n22327 ^ 1'b0 ;
  assign n36635 = n7109 ^ n612 ^ 1'b0 ;
  assign n36636 = n3451 | n13322 ;
  assign n36637 = n36636 ^ n12201 ^ 1'b0 ;
  assign n36638 = n36637 ^ n16422 ^ 1'b0 ;
  assign n36640 = n12020 ^ n5276 ^ 1'b0 ;
  assign n36641 = x14 & ~n36640 ;
  assign n36642 = ( n4084 & n19107 ) | ( n4084 & ~n36641 ) | ( n19107 & ~n36641 ) ;
  assign n36639 = n22552 | n30330 ;
  assign n36643 = n36642 ^ n36639 ^ 1'b0 ;
  assign n36644 = n11596 ^ n3833 ^ 1'b0 ;
  assign n36645 = ~n14719 & n36644 ;
  assign n36646 = n17810 & n36645 ;
  assign n36647 = n23194 & n36646 ;
  assign n36648 = n22915 ^ n15012 ^ 1'b0 ;
  assign n36649 = n21385 & ~n26944 ;
  assign n36650 = n5039 & n12978 ;
  assign n36651 = n1848 & n36650 ;
  assign n36652 = ~n17278 & n36296 ;
  assign n36653 = n36651 & ~n36652 ;
  assign n36654 = x97 & ~n1453 ;
  assign n36655 = ~n5150 & n36654 ;
  assign n36656 = n36655 ^ n2195 ^ 1'b0 ;
  assign n36657 = n23013 ^ n7506 ^ 1'b0 ;
  assign n36658 = n15765 ^ n8815 ^ n4339 ;
  assign n36659 = n36657 & n36658 ;
  assign n36660 = n36659 ^ n22723 ^ 1'b0 ;
  assign n36661 = ~n15502 & n36660 ;
  assign n36666 = n2885 & n26531 ;
  assign n36667 = n36666 ^ n16517 ^ 1'b0 ;
  assign n36668 = n6994 | n36667 ;
  assign n36662 = ( ~n14477 & n15829 ) | ( ~n14477 & n22494 ) | ( n15829 & n22494 ) ;
  assign n36663 = n36662 ^ n27475 ^ 1'b0 ;
  assign n36664 = ~n13035 & n36663 ;
  assign n36665 = ~n36488 & n36664 ;
  assign n36669 = n36668 ^ n36665 ^ 1'b0 ;
  assign n36670 = n33138 ^ n16610 ^ n6951 ;
  assign n36671 = n13685 & ~n36670 ;
  assign n36672 = n11827 | n26282 ;
  assign n36673 = n26639 & n36672 ;
  assign n36674 = n36416 ^ n22481 ^ 1'b0 ;
  assign n36675 = n11408 & ~n36674 ;
  assign n36676 = n22956 | n32075 ;
  assign n36677 = n36676 ^ n35582 ^ 1'b0 ;
  assign n36678 = n2384 | n14533 ;
  assign n36679 = n36678 ^ n7756 ^ 1'b0 ;
  assign n36680 = n8704 | n36679 ;
  assign n36681 = n36680 ^ n11822 ^ 1'b0 ;
  assign n36682 = ~n3136 & n6713 ;
  assign n36683 = n9064 ^ n4124 ^ 1'b0 ;
  assign n36684 = ~n36682 & n36683 ;
  assign n36685 = n9074 & ~n18475 ;
  assign n36686 = n36685 ^ n14814 ^ 1'b0 ;
  assign n36687 = ~n1059 & n36686 ;
  assign n36688 = n27295 & n28893 ;
  assign n36689 = n36688 ^ n13906 ^ 1'b0 ;
  assign n36690 = n30254 ^ n26144 ^ 1'b0 ;
  assign n36691 = n8345 & ~n36690 ;
  assign n36692 = n3942 & ~n15693 ;
  assign n36693 = n34286 & n36692 ;
  assign n36694 = n18193 ^ n5678 ^ 1'b0 ;
  assign n36695 = n849 | n36694 ;
  assign n36696 = ( n21024 & ~n22325 ) | ( n21024 & n36695 ) | ( ~n22325 & n36695 ) ;
  assign n36697 = n25758 ^ n10142 ^ 1'b0 ;
  assign n36698 = ( ~n19724 & n21248 ) | ( ~n19724 & n36697 ) | ( n21248 & n36697 ) ;
  assign n36699 = n33500 ^ n14316 ^ 1'b0 ;
  assign n36700 = n9290 & n13765 ;
  assign n36701 = n1034 & n36700 ;
  assign n36702 = n22360 ^ n17830 ^ n2214 ;
  assign n36703 = n16390 | n26359 ;
  assign n36704 = n1951 ^ n1253 ^ 1'b0 ;
  assign n36705 = n24723 ^ n2166 ^ 1'b0 ;
  assign n36706 = ~n28382 & n36705 ;
  assign n36707 = n20855 & n36706 ;
  assign n36708 = n6929 ^ n6831 ^ 1'b0 ;
  assign n36709 = n1415 ^ n1295 ^ x7 ;
  assign n36710 = n36709 ^ n23941 ^ 1'b0 ;
  assign n36711 = n22127 & ~n36710 ;
  assign n36712 = ( n879 & n3885 ) | ( n879 & n8351 ) | ( n3885 & n8351 ) ;
  assign n36713 = n30178 & ~n36712 ;
  assign n36714 = n36713 ^ n2762 ^ n1669 ;
  assign n36715 = n1674 | n33175 ;
  assign n36716 = n34538 & ~n36715 ;
  assign n36717 = n36714 | n36716 ;
  assign n36718 = n2255 | n36717 ;
  assign n36719 = n8239 & ~n20692 ;
  assign n36720 = ~n12867 & n20692 ;
  assign n36721 = n36720 ^ n18734 ^ 1'b0 ;
  assign n36722 = n27909 & n36721 ;
  assign n36723 = n36722 ^ n30922 ^ 1'b0 ;
  assign n36724 = n31892 ^ n2349 ^ 1'b0 ;
  assign n36725 = n7937 ^ n4382 ^ 1'b0 ;
  assign n36726 = n3731 | n13641 ;
  assign n36727 = n36726 ^ n33274 ^ 1'b0 ;
  assign n36728 = n24126 ^ n2558 ^ 1'b0 ;
  assign n36729 = n36728 ^ n17164 ^ n7475 ;
  assign n36730 = n3344 | n13013 ;
  assign n36731 = n672 & ~n15019 ;
  assign n36732 = ~n36730 & n36731 ;
  assign n36733 = n28072 & n36732 ;
  assign n36735 = n6485 ^ n928 ^ 1'b0 ;
  assign n36734 = n10455 & ~n13920 ;
  assign n36736 = n36735 ^ n36734 ^ 1'b0 ;
  assign n36737 = n35663 ^ n1800 ^ 1'b0 ;
  assign n36738 = n36736 | n36737 ;
  assign n36744 = ~n1136 & n13204 ;
  assign n36745 = n21781 & n36744 ;
  assign n36739 = ~n27594 & n27761 ;
  assign n36740 = n36739 ^ n8707 ^ 1'b0 ;
  assign n36741 = n32066 & n36740 ;
  assign n36742 = ~n34805 & n36741 ;
  assign n36743 = n1616 | n36742 ;
  assign n36746 = n36745 ^ n36743 ^ 1'b0 ;
  assign n36747 = n484 & n35275 ;
  assign n36748 = n8485 ^ n6504 ^ 1'b0 ;
  assign n36749 = n36748 ^ n24698 ^ 1'b0 ;
  assign n36750 = n36749 ^ n28238 ^ n14243 ;
  assign n36751 = n27348 ^ n16937 ^ 1'b0 ;
  assign n36752 = n15500 & ~n36751 ;
  assign n36753 = n36752 ^ n31911 ^ n28083 ;
  assign n36754 = n19369 ^ n4587 ^ 1'b0 ;
  assign n36755 = n1202 | n36754 ;
  assign n36758 = n7306 & ~n20144 ;
  assign n36759 = n1731 & n31120 ;
  assign n36760 = ~n36758 & n36759 ;
  assign n36756 = n4137 & n16732 ;
  assign n36757 = n36756 ^ n17942 ^ 1'b0 ;
  assign n36761 = n36760 ^ n36757 ^ n28783 ;
  assign n36762 = n4510 & ~n15500 ;
  assign n36766 = n24114 & n32484 ;
  assign n36767 = n36766 ^ n11421 ^ 1'b0 ;
  assign n36763 = n4194 | n30689 ;
  assign n36764 = n6215 | n36763 ;
  assign n36765 = n26224 | n36764 ;
  assign n36768 = n36767 ^ n36765 ^ 1'b0 ;
  assign n36769 = n11326 | n36645 ;
  assign n36770 = n9480 & ~n11438 ;
  assign n36771 = ~n36769 & n36770 ;
  assign n36772 = n17352 | n21216 ;
  assign n36773 = n32953 | n36772 ;
  assign n36774 = n26673 & n33056 ;
  assign n36775 = n36774 ^ n33150 ^ 1'b0 ;
  assign n36776 = n7007 ^ n6656 ^ 1'b0 ;
  assign n36777 = n2186 ^ n924 ^ 1'b0 ;
  assign n36778 = n18592 ^ n11428 ^ 1'b0 ;
  assign n36779 = n2548 ^ n1160 ^ 1'b0 ;
  assign n36780 = n4278 | n36779 ;
  assign n36781 = n24937 ^ n19675 ^ 1'b0 ;
  assign n36782 = n36780 | n36781 ;
  assign n36783 = ~n7280 & n33138 ;
  assign n36784 = n31194 & n36783 ;
  assign n36785 = n15595 ^ n8369 ^ 1'b0 ;
  assign n36786 = n1377 & ~n36785 ;
  assign n36787 = n23879 & ~n35051 ;
  assign n36788 = n397 & ~n10488 ;
  assign n36789 = ~n20289 & n36788 ;
  assign n36790 = n19518 | n36789 ;
  assign n36791 = n9232 | n36790 ;
  assign n36792 = n683 | n11237 ;
  assign n36793 = n36792 ^ n9800 ^ 1'b0 ;
  assign n36794 = n22723 ^ n3091 ^ 1'b0 ;
  assign n36795 = n5161 | n36794 ;
  assign n36796 = ( n20707 & n27718 ) | ( n20707 & ~n36795 ) | ( n27718 & ~n36795 ) ;
  assign n36797 = n31898 ^ n6021 ^ 1'b0 ;
  assign n36798 = n2380 | n36797 ;
  assign n36799 = n17392 ^ n10394 ^ 1'b0 ;
  assign n36800 = n5433 | n12236 ;
  assign n36801 = x83 & n2260 ;
  assign n36802 = n5025 & n36801 ;
  assign n36803 = n36802 ^ n34513 ^ 1'b0 ;
  assign n36804 = ~n33379 & n36803 ;
  assign n36805 = n5760 ^ n4705 ^ 1'b0 ;
  assign n36806 = n10915 | n36805 ;
  assign n36807 = n7578 & ~n36806 ;
  assign n36808 = n11332 & ~n36807 ;
  assign n36809 = ~n2305 & n36808 ;
  assign n36810 = ( n909 & ~n34484 ) | ( n909 & n36809 ) | ( ~n34484 & n36809 ) ;
  assign n36813 = n8119 | n10425 ;
  assign n36811 = n10637 ^ n8296 ^ n5687 ;
  assign n36812 = n36811 ^ n17071 ^ 1'b0 ;
  assign n36814 = n36813 ^ n36812 ^ n9914 ;
  assign n36815 = n9831 ^ n1836 ^ 1'b0 ;
  assign n36816 = n10177 & n36815 ;
  assign n36818 = n23710 ^ n4936 ^ 1'b0 ;
  assign n36817 = n10711 | n20584 ;
  assign n36819 = n36818 ^ n36817 ^ 1'b0 ;
  assign n36820 = n34257 & ~n36819 ;
  assign n36821 = n29937 ^ n12724 ^ 1'b0 ;
  assign n36822 = n3043 | n36821 ;
  assign n36823 = n3419 | n13303 ;
  assign n36824 = n26396 & ~n26509 ;
  assign n36825 = n14849 ^ n3639 ^ 1'b0 ;
  assign n36826 = n14908 | n36825 ;
  assign n36827 = n17668 ^ n8845 ^ 1'b0 ;
  assign n36828 = ~n24911 & n36827 ;
  assign n36829 = ( ~n3388 & n36789 ) | ( ~n3388 & n36828 ) | ( n36789 & n36828 ) ;
  assign n36830 = n17647 ^ n1909 ^ 1'b0 ;
  assign n36831 = n36829 & ~n36830 ;
  assign n36832 = ~n12350 & n36831 ;
  assign n36833 = n36832 ^ n12872 ^ 1'b0 ;
  assign n36834 = n36492 ^ n22550 ^ 1'b0 ;
  assign n36835 = n26273 & n36834 ;
  assign n36836 = n20921 & n22381 ;
  assign n36837 = n36836 ^ n19196 ^ 1'b0 ;
  assign n36838 = ~n6402 & n36837 ;
  assign n36839 = ~n33366 & n36838 ;
  assign n36840 = n16394 ^ n14605 ^ 1'b0 ;
  assign n36841 = ~n4941 & n36840 ;
  assign n36842 = n6811 & ~n20181 ;
  assign n36843 = ~n36841 & n36842 ;
  assign n36844 = n16428 ^ n12846 ^ 1'b0 ;
  assign n36845 = n31225 | n36844 ;
  assign n36846 = n3297 & n10230 ;
  assign n36847 = n23230 ^ n6643 ^ 1'b0 ;
  assign n36848 = ( n20243 & ~n25390 ) | ( n20243 & n36847 ) | ( ~n25390 & n36847 ) ;
  assign n36849 = ( n323 & n10642 ) | ( n323 & n21245 ) | ( n10642 & n21245 ) ;
  assign n36850 = n5366 & n16085 ;
  assign n36851 = x206 & ~n36850 ;
  assign n36852 = ( n14405 & n30540 ) | ( n14405 & ~n36851 ) | ( n30540 & ~n36851 ) ;
  assign n36853 = n1254 & n16811 ;
  assign n36854 = n5850 & ~n9060 ;
  assign n36855 = n15973 & ~n36854 ;
  assign n36856 = ( n783 & n1259 ) | ( n783 & n3204 ) | ( n1259 & n3204 ) ;
  assign n36857 = n36856 ^ n24565 ^ 1'b0 ;
  assign n36858 = n4900 & n5211 ;
  assign n36859 = n36858 ^ n29147 ^ 1'b0 ;
  assign n36860 = n15383 | n34200 ;
  assign n36861 = ( ~n4896 & n12128 ) | ( ~n4896 & n22419 ) | ( n12128 & n22419 ) ;
  assign n36863 = n23292 ^ n12550 ^ 1'b0 ;
  assign n36864 = n1010 & ~n36863 ;
  assign n36862 = n968 & n18014 ;
  assign n36865 = n36864 ^ n36862 ^ 1'b0 ;
  assign n36866 = n21422 ^ x237 ^ 1'b0 ;
  assign n36867 = n14673 & n25314 ;
  assign n36868 = n36867 ^ n16694 ^ 1'b0 ;
  assign n36869 = n1903 & n36868 ;
  assign n36870 = n36866 & ~n36869 ;
  assign n36871 = n15182 ^ n1963 ^ 1'b0 ;
  assign n36872 = ~n21082 & n36871 ;
  assign n36873 = n14055 | n15075 ;
  assign n36874 = n17181 ^ n16288 ^ 1'b0 ;
  assign n36875 = n28887 & n36874 ;
  assign n36882 = ~n11840 & n18206 ;
  assign n36876 = n24837 ^ n7661 ^ 1'b0 ;
  assign n36877 = n9404 & n21777 ;
  assign n36878 = n12190 | n36877 ;
  assign n36879 = n36876 & ~n36878 ;
  assign n36880 = ~n27899 & n36879 ;
  assign n36881 = ~n12308 & n36880 ;
  assign n36883 = n36882 ^ n36881 ^ n19934 ;
  assign n36884 = n26823 ^ n7116 ^ 1'b0 ;
  assign n36885 = ~n20672 & n36565 ;
  assign n36886 = n13491 ^ n3979 ^ 1'b0 ;
  assign n36887 = n19890 ^ n15010 ^ 1'b0 ;
  assign n36888 = n18841 ^ n15410 ^ 1'b0 ;
  assign n36889 = ~n36887 & n36888 ;
  assign n36890 = n6369 ^ n4406 ^ 1'b0 ;
  assign n36891 = n15551 | n36890 ;
  assign n36892 = n10846 & ~n36891 ;
  assign n36893 = ~n13454 & n36892 ;
  assign n36894 = n36889 & ~n36893 ;
  assign n36895 = ( n9347 & n20127 ) | ( n9347 & ~n33468 ) | ( n20127 & ~n33468 ) ;
  assign n36896 = n12500 | n12527 ;
  assign n36897 = n36896 ^ n11756 ^ 1'b0 ;
  assign n36898 = n16856 & n36897 ;
  assign n36899 = n10985 ^ n867 ^ 1'b0 ;
  assign n36900 = ~n36898 & n36899 ;
  assign n36901 = ( n10810 & n24276 ) | ( n10810 & ~n27499 ) | ( n24276 & ~n27499 ) ;
  assign n36902 = n7714 & ~n36901 ;
  assign n36903 = n1334 & ~n2203 ;
  assign n36904 = n17062 & n36903 ;
  assign n36905 = n22945 & ~n25171 ;
  assign n36906 = ( n3245 & n36904 ) | ( n3245 & n36905 ) | ( n36904 & n36905 ) ;
  assign n36907 = n10017 ^ n3406 ^ 1'b0 ;
  assign n36908 = ~n32197 & n36907 ;
  assign n36909 = n3123 | n28254 ;
  assign n36910 = n36909 ^ n22364 ^ 1'b0 ;
  assign n36911 = n36908 & n36910 ;
  assign n36912 = n2682 | n3493 ;
  assign n36913 = n36912 ^ n4419 ^ 1'b0 ;
  assign n36914 = n36913 ^ n15901 ^ 1'b0 ;
  assign n36915 = n6975 & ~n36914 ;
  assign n36916 = n7945 ^ n1382 ^ n550 ;
  assign n36917 = n9877 | n9889 ;
  assign n36918 = n14973 | n36917 ;
  assign n36919 = ( n23550 & ~n36916 ) | ( n23550 & n36918 ) | ( ~n36916 & n36918 ) ;
  assign n36920 = n31174 ^ n30101 ^ 1'b0 ;
  assign n36921 = n36920 ^ n33034 ^ n24350 ;
  assign n36922 = n12642 ^ n10445 ^ n6045 ;
  assign n36923 = n4497 ^ n4196 ^ 1'b0 ;
  assign n36924 = n19485 & n36923 ;
  assign n36925 = n1469 & n32218 ;
  assign n36926 = n36925 ^ n26168 ^ n20080 ;
  assign n36927 = n36926 ^ n11184 ^ 1'b0 ;
  assign n36928 = n36924 & ~n36927 ;
  assign n36929 = ~n6895 & n16868 ;
  assign n36930 = ~n824 & n13530 ;
  assign n36931 = n36930 ^ n27150 ^ 1'b0 ;
  assign n36932 = ~n31956 & n36931 ;
  assign n36933 = n4878 & n16181 ;
  assign n36934 = n36164 ^ n9347 ^ 1'b0 ;
  assign n36935 = ~n9921 & n36934 ;
  assign n36936 = n12739 ^ n3098 ^ n1075 ;
  assign n36937 = n11660 | n18264 ;
  assign n36938 = n8531 | n36937 ;
  assign n36939 = ( n4920 & n20495 ) | ( n4920 & ~n32490 ) | ( n20495 & ~n32490 ) ;
  assign n36940 = n24183 & ~n36939 ;
  assign n36941 = ~n11416 & n12199 ;
  assign n36942 = x187 & n674 ;
  assign n36943 = ~n12373 & n36942 ;
  assign n36944 = n15734 & ~n24504 ;
  assign n36945 = n16966 ^ n8682 ^ n2103 ;
  assign n36946 = ~n8316 & n36945 ;
  assign n36947 = n36946 ^ n22863 ^ 1'b0 ;
  assign n36948 = n17343 ^ n14603 ^ n3378 ;
  assign n36949 = n36948 ^ n2038 ^ 1'b0 ;
  assign n36950 = n8226 | n36949 ;
  assign n36951 = n36950 ^ n33347 ^ n2882 ;
  assign n36952 = n17182 & n35669 ;
  assign n36953 = n10707 & n13423 ;
  assign n36954 = n3542 | n36953 ;
  assign n36955 = n742 & n13926 ;
  assign n36956 = n1242 & ~n5154 ;
  assign n36957 = n14807 ^ n9582 ^ 1'b0 ;
  assign n36958 = ~n2721 & n25181 ;
  assign n36959 = ( n1396 & n5903 ) | ( n1396 & n36014 ) | ( n5903 & n36014 ) ;
  assign n36960 = n13747 ^ n4705 ^ 1'b0 ;
  assign n36961 = ~n12182 & n36960 ;
  assign n36962 = n780 & n23985 ;
  assign n36963 = ~n36961 & n36962 ;
  assign n36964 = n18520 & n21834 ;
  assign n36965 = n36964 ^ n26989 ^ 1'b0 ;
  assign n36966 = n20144 & ~n28367 ;
  assign n36967 = n2585 | n5724 ;
  assign n36968 = n10582 & ~n36967 ;
  assign n36969 = n36968 ^ n11316 ^ n6001 ;
  assign n36970 = n28382 & ~n36969 ;
  assign n36971 = n627 & ~n17700 ;
  assign n36972 = n36971 ^ n5910 ^ 1'b0 ;
  assign n36973 = n6597 & ~n36972 ;
  assign n36974 = n3540 & ~n8316 ;
  assign n36975 = n36974 ^ n13683 ^ 1'b0 ;
  assign n36976 = n36973 | n36975 ;
  assign n36977 = n31019 ^ n8800 ^ n4686 ;
  assign n36978 = ~n11807 & n12909 ;
  assign n36979 = ( n2080 & n4284 ) | ( n2080 & n9192 ) | ( n4284 & n9192 ) ;
  assign n36980 = n36978 & ~n36979 ;
  assign n36981 = ( n9514 & n15569 ) | ( n9514 & n19039 ) | ( n15569 & n19039 ) ;
  assign n36982 = ( n4925 & n13920 ) | ( n4925 & n31323 ) | ( n13920 & n31323 ) ;
  assign n36983 = n36982 ^ n20337 ^ 1'b0 ;
  assign n36984 = n36981 & n36983 ;
  assign n36985 = n24471 ^ n22665 ^ 1'b0 ;
  assign n36986 = n3668 | n36985 ;
  assign n36987 = n19323 & ~n23207 ;
  assign n36989 = n4964 & n6880 ;
  assign n36990 = ~n6992 & n36989 ;
  assign n36988 = n6232 & n19099 ;
  assign n36991 = n36990 ^ n36988 ^ 1'b0 ;
  assign n36992 = n11844 & ~n36879 ;
  assign n36993 = n36992 ^ n25806 ^ 1'b0 ;
  assign n36994 = n7532 ^ n2096 ^ x235 ;
  assign n36995 = n36994 ^ n5277 ^ 1'b0 ;
  assign n36996 = n32476 ^ n19895 ^ n9275 ;
  assign n36997 = ( n9012 & ~n14760 ) | ( n9012 & n36996 ) | ( ~n14760 & n36996 ) ;
  assign n36998 = n21736 ^ n15694 ^ 1'b0 ;
  assign n36999 = n11273 & n36998 ;
  assign n37000 = n4018 | n34141 ;
  assign n37001 = n2690 | n37000 ;
  assign n37002 = n7569 | n15258 ;
  assign n37003 = n32964 ^ n32709 ^ 1'b0 ;
  assign n37004 = n6811 ^ n1866 ^ n1407 ;
  assign n37005 = n20199 | n30260 ;
  assign n37006 = n28639 & ~n37005 ;
  assign n37007 = n17226 & n37006 ;
  assign n37008 = n18933 | n24341 ;
  assign n37009 = n25304 | n37008 ;
  assign n37010 = n23258 & ~n32538 ;
  assign n37011 = n37010 ^ n2437 ^ 1'b0 ;
  assign n37012 = n504 | n37011 ;
  assign n37013 = n37012 ^ n21655 ^ 1'b0 ;
  assign n37014 = n37013 ^ n17123 ^ n12987 ;
  assign n37015 = n31648 ^ n14482 ^ n7830 ;
  assign n37016 = ~n6278 & n26929 ;
  assign n37017 = n37016 ^ n25160 ^ 1'b0 ;
  assign n37018 = n14110 & ~n35393 ;
  assign n37019 = n37018 ^ n10369 ^ 1'b0 ;
  assign n37020 = n17964 & n26527 ;
  assign n37021 = n32695 & n37020 ;
  assign n37022 = n37021 ^ n7605 ^ n1767 ;
  assign n37023 = n5643 & ~n9244 ;
  assign n37024 = ~n2511 & n10483 ;
  assign n37025 = n404 & n37024 ;
  assign n37026 = n2957 & n12897 ;
  assign n37027 = ~x58 & n37026 ;
  assign n37028 = n5341 & ~n37027 ;
  assign n37029 = ~n10083 & n37028 ;
  assign n37030 = n32394 & ~n37029 ;
  assign n37031 = n37030 ^ n21629 ^ 1'b0 ;
  assign n37032 = n19583 & n37031 ;
  assign n37033 = n828 & n37032 ;
  assign n37034 = n10027 | n27806 ;
  assign n37035 = n37034 ^ n7773 ^ 1'b0 ;
  assign n37036 = n6489 ^ n6041 ^ 1'b0 ;
  assign n37037 = ~n402 & n22536 ;
  assign n37038 = n37037 ^ n9263 ^ n1401 ;
  assign n37039 = ~n37036 & n37038 ;
  assign n37040 = ~n5402 & n25597 ;
  assign n37041 = n19126 | n37040 ;
  assign n37042 = ( n2320 & ~n7911 ) | ( n2320 & n10346 ) | ( ~n7911 & n10346 ) ;
  assign n37043 = n8415 & ~n37042 ;
  assign n37044 = n37043 ^ x141 ^ 1'b0 ;
  assign n37045 = n21570 | n37044 ;
  assign n37046 = n37045 ^ n7831 ^ 1'b0 ;
  assign n37047 = ~n32641 & n37046 ;
  assign n37048 = n5217 & ~n7565 ;
  assign n37049 = n2986 | n25897 ;
  assign n37050 = n28101 ^ n1838 ^ 1'b0 ;
  assign n37051 = n37049 | n37050 ;
  assign n37052 = n5449 & n5698 ;
  assign n37053 = n37052 ^ n23400 ^ 1'b0 ;
  assign n37057 = ~n7758 & n9935 ;
  assign n37058 = ~n26884 & n37057 ;
  assign n37059 = ( n9498 & n11167 ) | ( n9498 & ~n37058 ) | ( n11167 & ~n37058 ) ;
  assign n37054 = ~n3507 & n11586 ;
  assign n37055 = n37054 ^ n5446 ^ 1'b0 ;
  assign n37056 = n37055 ^ n5713 ^ n2372 ;
  assign n37060 = n37059 ^ n37056 ^ 1'b0 ;
  assign n37061 = ~n37053 & n37060 ;
  assign n37062 = n19902 ^ n3401 ^ n369 ;
  assign n37063 = ~n10879 & n32209 ;
  assign n37064 = ~n37062 & n37063 ;
  assign n37065 = n19939 & ~n29438 ;
  assign n37066 = n37065 ^ n10471 ^ 1'b0 ;
  assign n37067 = n12002 ^ n677 ^ 1'b0 ;
  assign n37068 = n37067 ^ n26084 ^ 1'b0 ;
  assign n37069 = n10043 & n37068 ;
  assign n37070 = ~n3981 & n37069 ;
  assign n37071 = n24561 ^ n456 ^ 1'b0 ;
  assign n37072 = n9694 & n20963 ;
  assign n37073 = n37072 ^ n18383 ^ 1'b0 ;
  assign n37074 = n3454 ^ n2481 ^ 1'b0 ;
  assign n37075 = n7157 & n37074 ;
  assign n37076 = n11819 & ~n20375 ;
  assign n37077 = n37076 ^ n9700 ^ 1'b0 ;
  assign n37078 = n31434 | n37077 ;
  assign n37079 = n37075 | n37078 ;
  assign n37080 = n9355 | n11763 ;
  assign n37083 = n7525 | n14696 ;
  assign n37081 = n17570 ^ n6291 ^ 1'b0 ;
  assign n37082 = n7853 & ~n37081 ;
  assign n37084 = n37083 ^ n37082 ^ n30624 ;
  assign n37085 = n13995 ^ n1917 ^ 1'b0 ;
  assign n37086 = n12551 ^ n10900 ^ n593 ;
  assign n37087 = x187 | n34143 ;
  assign n37088 = n37087 ^ n21716 ^ 1'b0 ;
  assign n37089 = n5843 ^ n4721 ^ 1'b0 ;
  assign n37090 = n37088 & n37089 ;
  assign n37091 = ~n14195 & n31136 ;
  assign n37092 = n37091 ^ n16546 ^ n6563 ;
  assign n37093 = n37092 ^ n21004 ^ 1'b0 ;
  assign n37094 = ~n4724 & n5510 ;
  assign n37095 = n2144 & n37094 ;
  assign n37096 = ( x131 & n11072 ) | ( x131 & n37095 ) | ( n11072 & n37095 ) ;
  assign n37097 = n17806 ^ n7844 ^ n2184 ;
  assign n37098 = n30314 ^ n25094 ^ 1'b0 ;
  assign n37099 = ~n5515 & n10085 ;
  assign n37100 = ~n20282 & n37099 ;
  assign n37101 = ~n3294 & n14841 ;
  assign n37102 = ~n27329 & n37101 ;
  assign n37103 = n5864 ^ n5699 ^ 1'b0 ;
  assign n37104 = ~n37102 & n37103 ;
  assign n37105 = ( n1313 & n10372 ) | ( n1313 & ~n29065 ) | ( n10372 & ~n29065 ) ;
  assign n37106 = n14012 & ~n37105 ;
  assign n37107 = n37106 ^ n6980 ^ n3350 ;
  assign n37108 = n37107 ^ n14090 ^ 1'b0 ;
  assign n37109 = n9797 | n37108 ;
  assign n37110 = n37109 ^ n5843 ^ 1'b0 ;
  assign n37111 = n35790 ^ n19205 ^ 1'b0 ;
  assign n37112 = ~n6844 & n10244 ;
  assign n37113 = n37112 ^ n14178 ^ 1'b0 ;
  assign n37114 = n2774 | n37113 ;
  assign n37115 = ( ~n6176 & n11171 ) | ( ~n6176 & n12058 ) | ( n11171 & n12058 ) ;
  assign n37116 = n37115 ^ n4880 ^ 1'b0 ;
  assign n37117 = n1813 & n37116 ;
  assign n37118 = n37117 ^ n31869 ^ n1175 ;
  assign n37119 = n9440 & ~n16557 ;
  assign n37120 = n37119 ^ n30282 ^ n6741 ;
  assign n37121 = n7519 & n23316 ;
  assign n37122 = n2721 & n37121 ;
  assign n37123 = ~n2106 & n37122 ;
  assign n37124 = n4597 & ~n37123 ;
  assign n37125 = n21609 ^ n15010 ^ n5859 ;
  assign n37126 = n9429 | n37125 ;
  assign n37127 = ~n1930 & n21841 ;
  assign n37128 = ~n15597 & n37127 ;
  assign n37129 = ( n4070 & n14390 ) | ( n4070 & n19652 ) | ( n14390 & n19652 ) ;
  assign n37130 = n20829 ^ n13501 ^ 1'b0 ;
  assign n37131 = n16967 & ~n37130 ;
  assign n37132 = n24388 | n31225 ;
  assign n37133 = n26954 ^ n6131 ^ 1'b0 ;
  assign n37134 = ~n29651 & n37133 ;
  assign n37135 = n23307 ^ n19445 ^ 1'b0 ;
  assign n37136 = n31511 | n37135 ;
  assign n37137 = n20770 | n37136 ;
  assign n37138 = n30539 | n37137 ;
  assign n37139 = n5782 & ~n19026 ;
  assign n37140 = n3454 | n10837 ;
  assign n37141 = n37140 ^ n20509 ^ n8212 ;
  assign n37142 = n24052 ^ n4382 ^ 1'b0 ;
  assign n37143 = n13580 & n28810 ;
  assign n37144 = n14469 | n37143 ;
  assign n37145 = n37142 & ~n37144 ;
  assign n37146 = n23152 ^ n5099 ^ 1'b0 ;
  assign n37147 = n4429 & ~n16163 ;
  assign n37148 = n13885 ^ n5331 ^ 1'b0 ;
  assign n37149 = n3777 & ~n37148 ;
  assign n37150 = n9668 & n37149 ;
  assign n37151 = ~n14500 & n32910 ;
  assign n37152 = n37151 ^ n34079 ^ 1'b0 ;
  assign n37153 = n27690 | n37152 ;
  assign n37154 = n37153 ^ n19287 ^ 1'b0 ;
  assign n37155 = ~n6679 & n14698 ;
  assign n37156 = n17366 & ~n26058 ;
  assign n37157 = n20272 & n22037 ;
  assign n37158 = ( n5527 & n37156 ) | ( n5527 & n37157 ) | ( n37156 & n37157 ) ;
  assign n37159 = n6422 & ~n13063 ;
  assign n37160 = n31136 & ~n37159 ;
  assign n37161 = n6103 & n28408 ;
  assign n37162 = n25490 & n32640 ;
  assign n37163 = n37162 ^ n31189 ^ 1'b0 ;
  assign n37164 = n33551 ^ n30384 ^ 1'b0 ;
  assign n37165 = n12080 | n37164 ;
  assign n37166 = ~n2614 & n4703 ;
  assign n37167 = n37166 ^ n10943 ^ 1'b0 ;
  assign n37168 = n6236 & n16073 ;
  assign n37169 = n37167 & n37168 ;
  assign n37170 = x114 & ~n30333 ;
  assign n37171 = n1415 | n9155 ;
  assign n37172 = n37171 ^ n286 ^ 1'b0 ;
  assign n37173 = ~n9425 & n37172 ;
  assign n37174 = n2826 | n37173 ;
  assign n37175 = n9087 & n13835 ;
  assign n37176 = ~n34833 & n37175 ;
  assign n37177 = n2469 & ~n37176 ;
  assign n37178 = n9724 & n25762 ;
  assign n37179 = ~n37177 & n37178 ;
  assign n37180 = n1589 & ~n12778 ;
  assign n37181 = n23284 ^ n7518 ^ 1'b0 ;
  assign n37182 = x40 & ~n37181 ;
  assign n37183 = ~n3490 & n37182 ;
  assign n37184 = n37180 & n37183 ;
  assign n37185 = n22238 ^ n16539 ^ 1'b0 ;
  assign n37186 = n4039 & n37185 ;
  assign n37187 = ~n10979 & n12721 ;
  assign n37188 = n35650 & n37187 ;
  assign n37189 = n29508 ^ n25615 ^ n20935 ;
  assign n37190 = ( ~n10252 & n10265 ) | ( ~n10252 & n30229 ) | ( n10265 & n30229 ) ;
  assign n37191 = n10132 & n18101 ;
  assign n37192 = ( n1102 & n8288 ) | ( n1102 & ~n37191 ) | ( n8288 & ~n37191 ) ;
  assign n37193 = n2654 & ~n23710 ;
  assign n37194 = n37193 ^ n18987 ^ 1'b0 ;
  assign n37195 = n37194 ^ n21000 ^ 1'b0 ;
  assign n37196 = n11210 | n37195 ;
  assign n37197 = ~n1663 & n37196 ;
  assign n37198 = ( n6379 & n18376 ) | ( n6379 & n20651 ) | ( n18376 & n20651 ) ;
  assign n37199 = ~n1400 & n37198 ;
  assign n37200 = n17169 & ~n18997 ;
  assign n37201 = n37199 & n37200 ;
  assign n37202 = n17740 ^ n10001 ^ 1'b0 ;
  assign n37203 = ~n16960 & n37202 ;
  assign n37209 = n8484 & n20795 ;
  assign n37210 = ~n20795 & n37209 ;
  assign n37207 = n2207 | n14310 ;
  assign n37208 = n7977 & ~n37207 ;
  assign n37211 = n37210 ^ n37208 ^ n33051 ;
  assign n37204 = ( n4287 & n8133 ) | ( n4287 & ~n13009 ) | ( n8133 & ~n13009 ) ;
  assign n37205 = n22248 | n37204 ;
  assign n37206 = n22248 & ~n37205 ;
  assign n37212 = n37211 ^ n37206 ^ n15197 ;
  assign n37213 = n32195 ^ n30776 ^ 1'b0 ;
  assign n37214 = n37212 & n37213 ;
  assign n37215 = n3460 ^ x218 ^ 1'b0 ;
  assign n37216 = ~n10771 & n37215 ;
  assign n37217 = n30019 & n37216 ;
  assign n37218 = n11810 ^ n2010 ^ 1'b0 ;
  assign n37219 = n20188 ^ n1577 ^ 1'b0 ;
  assign n37220 = n1362 | n8708 ;
  assign n37221 = n2522 & ~n37220 ;
  assign n37222 = ~n6272 & n37221 ;
  assign n37223 = n23099 & ~n37222 ;
  assign n37224 = n5354 | n27350 ;
  assign n37225 = n591 & ~n12523 ;
  assign n37226 = n2438 | n37225 ;
  assign n37227 = n3515 | n10867 ;
  assign n37228 = n17450 & ~n37227 ;
  assign n37229 = n16485 & ~n19547 ;
  assign n37230 = n37228 & ~n37229 ;
  assign n37231 = ( n11649 & n12255 ) | ( n11649 & n22688 ) | ( n12255 & n22688 ) ;
  assign n37232 = n37231 ^ n2710 ^ 1'b0 ;
  assign n37233 = n2468 & n21584 ;
  assign n37234 = ~n8643 & n29380 ;
  assign n37235 = n37234 ^ n6352 ^ 1'b0 ;
  assign n37236 = n22818 ^ n17980 ^ 1'b0 ;
  assign n37237 = ~n16547 & n26783 ;
  assign n37238 = n25545 | n37237 ;
  assign n37239 = n19242 & ~n31782 ;
  assign n37240 = ~n3264 & n37239 ;
  assign n37242 = ~n1495 & n2939 ;
  assign n37241 = n8564 | n25655 ;
  assign n37243 = n37242 ^ n37241 ^ 1'b0 ;
  assign n37244 = ~n10614 & n19370 ;
  assign n37245 = n31251 ^ n11077 ^ 1'b0 ;
  assign n37246 = ~n15926 & n37245 ;
  assign n37247 = n2692 & ~n37246 ;
  assign n37248 = ~n1430 & n3922 ;
  assign n37249 = n12293 & ~n37248 ;
  assign n37250 = n24062 ^ n22692 ^ n1641 ;
  assign n37251 = n26383 ^ n20038 ^ n12854 ;
  assign n37252 = n11178 ^ n5278 ^ 1'b0 ;
  assign n37253 = n4638 & ~n37252 ;
  assign n37254 = ~n1111 & n32682 ;
  assign n37255 = n12004 & n37254 ;
  assign n37256 = n3729 & ~n4368 ;
  assign n37257 = n6548 & n37256 ;
  assign n37258 = x7 | n13651 ;
  assign n37259 = n11341 & ~n37258 ;
  assign n37260 = n17983 & ~n37259 ;
  assign n37261 = ~n26950 & n37260 ;
  assign n37262 = x234 | n26675 ;
  assign n37263 = n14406 ^ n2836 ^ 1'b0 ;
  assign n37264 = n10228 ^ n3317 ^ 1'b0 ;
  assign n37265 = n9249 | n37264 ;
  assign n37266 = ~n32484 & n37265 ;
  assign n37267 = n5967 & ~n10808 ;
  assign n37268 = n3926 & n4721 ;
  assign n37269 = n37268 ^ n9099 ^ 1'b0 ;
  assign n37270 = n9518 ^ n7544 ^ 1'b0 ;
  assign n37271 = n8029 ^ n8013 ^ 1'b0 ;
  assign n37272 = n37270 | n37271 ;
  assign n37273 = n37272 ^ n9369 ^ 1'b0 ;
  assign n37274 = n20968 ^ n1532 ^ 1'b0 ;
  assign n37275 = ~n18805 & n37274 ;
  assign n37276 = n5224 | n14227 ;
  assign n37277 = n26177 | n37276 ;
  assign n37278 = ( n8712 & n12674 ) | ( n8712 & ~n19566 ) | ( n12674 & ~n19566 ) ;
  assign n37279 = n14299 | n37278 ;
  assign n37280 = n37279 ^ n22066 ^ 1'b0 ;
  assign n37281 = n33566 ^ n26695 ^ 1'b0 ;
  assign n37282 = n29593 & ~n37281 ;
  assign n37283 = x239 & n7926 ;
  assign n37284 = n37283 ^ n12917 ^ 1'b0 ;
  assign n37285 = n34886 | n35118 ;
  assign n37286 = n8343 ^ n713 ^ 1'b0 ;
  assign n37287 = n8851 | n24444 ;
  assign n37288 = n37286 | n37287 ;
  assign n37289 = n37288 ^ n33993 ^ 1'b0 ;
  assign n37290 = ~n27296 & n37289 ;
  assign n37291 = n28327 ^ n4977 ^ 1'b0 ;
  assign n37292 = n4895 & ~n17069 ;
  assign n37293 = n37292 ^ n860 ^ 1'b0 ;
  assign n37294 = n37293 ^ n24614 ^ 1'b0 ;
  assign n37295 = ~n7650 & n25594 ;
  assign n37296 = ~n22814 & n37295 ;
  assign n37297 = n35234 ^ n15996 ^ 1'b0 ;
  assign n37298 = ~n37296 & n37297 ;
  assign n37299 = n33493 ^ n20497 ^ n7115 ;
  assign n37300 = n26934 ^ n7995 ^ 1'b0 ;
  assign n37301 = n37299 & n37300 ;
  assign n37302 = n22469 ^ n9710 ^ n7337 ;
  assign n37303 = n28075 ^ n26456 ^ n8167 ;
  assign n37304 = n8924 | n11137 ;
  assign n37305 = n1029 & ~n37304 ;
  assign n37306 = n37303 & n37305 ;
  assign n37307 = n28737 & ~n37306 ;
  assign n37308 = n12112 & n21421 ;
  assign n37309 = ~n1145 & n37308 ;
  assign n37310 = n15469 ^ n6770 ^ 1'b0 ;
  assign n37311 = n19281 | n37310 ;
  assign n37312 = n20983 ^ n5888 ^ n3144 ;
  assign n37313 = n36347 & ~n37312 ;
  assign n37314 = n3401 & n6381 ;
  assign n37315 = ~n2806 & n12576 ;
  assign n37316 = n37315 ^ n12525 ^ 1'b0 ;
  assign n37317 = n21223 & n37316 ;
  assign n37318 = n28752 | n37317 ;
  assign n37319 = n37318 ^ n10372 ^ 1'b0 ;
  assign n37320 = n8772 & ~n24271 ;
  assign n37321 = n25698 ^ n15240 ^ 1'b0 ;
  assign n37322 = ~n34333 & n37321 ;
  assign n37328 = n12008 ^ n10032 ^ 1'b0 ;
  assign n37323 = n9771 & ~n15655 ;
  assign n37324 = n37323 ^ n7101 ^ 1'b0 ;
  assign n37325 = n37324 ^ n2930 ^ 1'b0 ;
  assign n37326 = n24997 & n37325 ;
  assign n37327 = n1559 & n37326 ;
  assign n37329 = n37328 ^ n37327 ^ 1'b0 ;
  assign n37330 = n20128 ^ n11938 ^ n10151 ;
  assign n37331 = n37330 ^ n683 ^ 1'b0 ;
  assign n37332 = n13977 & ~n37331 ;
  assign n37333 = ( n4962 & n13656 ) | ( n4962 & ~n19070 ) | ( n13656 & ~n19070 ) ;
  assign n37334 = ~n10709 & n17806 ;
  assign n37335 = n17368 ^ n2264 ^ 1'b0 ;
  assign n37336 = ~n18222 & n37335 ;
  assign n37337 = n37336 ^ n4072 ^ 1'b0 ;
  assign n37338 = n2561 & n10649 ;
  assign n37339 = ~n11248 & n37338 ;
  assign n37340 = n11359 ^ n1858 ^ 1'b0 ;
  assign n37341 = n24392 ^ n14489 ^ n9463 ;
  assign n37342 = n9716 ^ n5765 ^ 1'b0 ;
  assign n37343 = n1120 | n37342 ;
  assign n37344 = ~n4366 & n37149 ;
  assign n37345 = ~n8805 & n37344 ;
  assign n37346 = n24669 ^ n18424 ^ n2176 ;
  assign n37347 = n37345 | n37346 ;
  assign n37348 = ( n28282 & ~n37343 ) | ( n28282 & n37347 ) | ( ~n37343 & n37347 ) ;
  assign n37349 = n17411 & ~n32363 ;
  assign n37350 = ~n17003 & n37349 ;
  assign n37351 = n26846 & ~n33500 ;
  assign n37353 = n4867 ^ n2871 ^ 1'b0 ;
  assign n37352 = ~n1026 & n33474 ;
  assign n37354 = n37353 ^ n37352 ^ 1'b0 ;
  assign n37355 = n15179 ^ n8800 ^ 1'b0 ;
  assign n37356 = n16596 | n37355 ;
  assign n37357 = n5986 ^ n5932 ^ 1'b0 ;
  assign n37358 = n24136 & n37357 ;
  assign n37359 = ~n1550 & n37358 ;
  assign n37360 = n31601 | n37359 ;
  assign n37361 = n37356 & ~n37360 ;
  assign n37362 = n7406 ^ n7145 ^ n6788 ;
  assign n37363 = n1618 & ~n4150 ;
  assign n37364 = n37362 & n37363 ;
  assign n37365 = n4342 & n18757 ;
  assign n37366 = n1510 ^ x32 ^ 1'b0 ;
  assign n37367 = n37366 ^ n21701 ^ n18193 ;
  assign n37368 = n37367 ^ n24225 ^ n18713 ;
  assign n37369 = ~n30807 & n37368 ;
  assign n37370 = n1250 | n3342 ;
  assign n37371 = n26140 & ~n37370 ;
  assign n37372 = n2746 & ~n4021 ;
  assign n37373 = ~n21608 & n37372 ;
  assign n37374 = ( n13750 & n18839 ) | ( n13750 & n37373 ) | ( n18839 & n37373 ) ;
  assign n37375 = n11173 & n37374 ;
  assign n37376 = n29460 ^ n27759 ^ n2972 ;
  assign n37377 = n17532 | n31069 ;
  assign n37378 = n12221 & ~n28741 ;
  assign n37379 = n8533 & ~n23465 ;
  assign n37380 = n10191 | n37379 ;
  assign n37381 = n24392 | n37380 ;
  assign n37382 = ( n4957 & n21951 ) | ( n4957 & n37381 ) | ( n21951 & n37381 ) ;
  assign n37383 = n10064 & ~n37382 ;
  assign n37384 = n11078 & n37383 ;
  assign n37385 = n34938 ^ n24599 ^ 1'b0 ;
  assign n37386 = n36208 & ~n37385 ;
  assign n37387 = ~n12613 & n24110 ;
  assign n37388 = n6363 & ~n37387 ;
  assign n37389 = n2706 & ~n31097 ;
  assign n37392 = n3477 & ~n6808 ;
  assign n37393 = n37392 ^ n21600 ^ 1'b0 ;
  assign n37394 = ~n8409 & n37393 ;
  assign n37395 = n37394 ^ n11142 ^ 1'b0 ;
  assign n37396 = n37395 ^ n20272 ^ n455 ;
  assign n37390 = n9603 | n14618 ;
  assign n37391 = n10490 & ~n37390 ;
  assign n37397 = n37396 ^ n37391 ^ n18994 ;
  assign n37398 = n19194 ^ n18403 ^ 1'b0 ;
  assign n37399 = n5196 | n37398 ;
  assign n37400 = ( ~n15440 & n17769 ) | ( ~n15440 & n37399 ) | ( n17769 & n37399 ) ;
  assign n37401 = n28103 ^ n13723 ^ 1'b0 ;
  assign n37402 = n30387 & n37401 ;
  assign n37403 = ~n5499 & n32966 ;
  assign n37404 = n27779 & n37403 ;
  assign n37405 = n21508 & ~n37404 ;
  assign n37406 = ~n3905 & n8945 ;
  assign n37407 = n7246 & n37406 ;
  assign n37408 = n31588 & n37407 ;
  assign n37409 = n17023 ^ n6937 ^ 1'b0 ;
  assign n37410 = n34107 & ~n37409 ;
  assign n37411 = n319 & ~n17574 ;
  assign n37412 = ( ~n12718 & n18334 ) | ( ~n12718 & n23532 ) | ( n18334 & n23532 ) ;
  assign n37413 = n9788 | n37412 ;
  assign n37414 = n33487 ^ n14020 ^ n12099 ;
  assign n37415 = n4489 & ~n10068 ;
  assign n37416 = n37415 ^ n13917 ^ 1'b0 ;
  assign n37417 = n30709 ^ n19375 ^ 1'b0 ;
  assign n37418 = n37416 & n37417 ;
  assign n37419 = n29351 ^ n11808 ^ 1'b0 ;
  assign n37420 = ~n3059 & n37419 ;
  assign n37421 = n37420 ^ n18193 ^ n5683 ;
  assign n37422 = ( ~n6296 & n8748 ) | ( ~n6296 & n13632 ) | ( n8748 & n13632 ) ;
  assign n37423 = ~n20476 & n37422 ;
  assign n37424 = n22392 ^ n12291 ^ 1'b0 ;
  assign n37425 = ~n21941 & n37424 ;
  assign n37426 = n37425 ^ n21763 ^ 1'b0 ;
  assign n37431 = n18004 ^ n6906 ^ 1'b0 ;
  assign n37427 = n13033 ^ n12895 ^ 1'b0 ;
  assign n37428 = n27159 & n37427 ;
  assign n37429 = n37428 ^ n1308 ^ 1'b0 ;
  assign n37430 = n21248 & ~n37429 ;
  assign n37432 = n37431 ^ n37430 ^ 1'b0 ;
  assign n37433 = n21592 ^ n10128 ^ 1'b0 ;
  assign n37434 = n25599 ^ n15381 ^ n12126 ;
  assign n37435 = ~n5406 & n37434 ;
  assign n37436 = n37435 ^ n4294 ^ 1'b0 ;
  assign n37437 = ~n3088 & n7049 ;
  assign n37438 = ( n1111 & n7849 ) | ( n1111 & n37437 ) | ( n7849 & n37437 ) ;
  assign n37439 = n17359 ^ n271 ^ 1'b0 ;
  assign n37440 = n3968 ^ x27 ^ 1'b0 ;
  assign n37441 = ~n37439 & n37440 ;
  assign n37442 = n37438 & n37441 ;
  assign n37443 = n463 & n13324 ;
  assign n37444 = n15962 & n20103 ;
  assign n37445 = ~n4562 & n24039 ;
  assign n37446 = ( n11227 & n21062 ) | ( n11227 & n37445 ) | ( n21062 & n37445 ) ;
  assign n37447 = n21106 & ~n34926 ;
  assign n37448 = ~n5361 & n12327 ;
  assign n37449 = n37448 ^ n27243 ^ 1'b0 ;
  assign n37450 = n29795 ^ n21067 ^ 1'b0 ;
  assign n37451 = n6895 & n37450 ;
  assign n37452 = n37451 ^ n23978 ^ 1'b0 ;
  assign n37453 = n4789 ^ n4418 ^ 1'b0 ;
  assign n37454 = n37452 | n37453 ;
  assign n37455 = n19882 | n35129 ;
  assign n37456 = n37455 ^ n22200 ^ 1'b0 ;
  assign n37457 = ( n6833 & n11345 ) | ( n6833 & n27011 ) | ( n11345 & n27011 ) ;
  assign n37458 = n19390 ^ n18610 ^ 1'b0 ;
  assign n37459 = ( ~n7070 & n37457 ) | ( ~n7070 & n37458 ) | ( n37457 & n37458 ) ;
  assign n37460 = ~n30194 & n37459 ;
  assign n37462 = n6476 & n16595 ;
  assign n37463 = n37462 ^ n5770 ^ 1'b0 ;
  assign n37461 = n2744 | n13103 ;
  assign n37464 = n37463 ^ n37461 ^ 1'b0 ;
  assign n37465 = ( n19743 & n20346 ) | ( n19743 & n20879 ) | ( n20346 & n20879 ) ;
  assign n37466 = n12253 ^ n7051 ^ x128 ;
  assign n37467 = n11915 | n37466 ;
  assign n37468 = n33530 ^ n7306 ^ 1'b0 ;
  assign n37469 = n16278 & n21761 ;
  assign n37470 = ~x222 & n27726 ;
  assign n37471 = n34196 | n37470 ;
  assign n37475 = ~n2284 & n2976 ;
  assign n37476 = n37475 ^ n2966 ^ 1'b0 ;
  assign n37472 = ~n1998 & n8826 ;
  assign n37473 = n6572 & n37472 ;
  assign n37474 = n2028 & ~n37473 ;
  assign n37477 = n37476 ^ n37474 ^ 1'b0 ;
  assign n37478 = n37477 ^ n1982 ^ n328 ;
  assign n37479 = n13780 & ~n20706 ;
  assign n37480 = n11227 | n12138 ;
  assign n37481 = n5972 ^ n2359 ^ n1206 ;
  assign n37482 = n33181 | n37481 ;
  assign n37483 = n37482 ^ n34578 ^ 1'b0 ;
  assign n37484 = n37483 ^ n23536 ^ 1'b0 ;
  assign n37485 = n15181 ^ n13538 ^ 1'b0 ;
  assign n37486 = n37485 ^ n10657 ^ 1'b0 ;
  assign n37487 = ~n13868 & n37486 ;
  assign n37488 = n13851 ^ n13214 ^ 1'b0 ;
  assign n37489 = ~n3077 & n12095 ;
  assign n37490 = n37489 ^ n3907 ^ n3126 ;
  assign n37491 = n24623 & n32403 ;
  assign n37492 = n37491 ^ x175 ^ 1'b0 ;
  assign n37493 = ~n2610 & n30689 ;
  assign n37494 = ~n37492 & n37493 ;
  assign n37495 = n20152 ^ n14043 ^ 1'b0 ;
  assign n37496 = n1206 & ~n2830 ;
  assign n37497 = n35408 ^ n29398 ^ 1'b0 ;
  assign n37498 = n27594 | n37497 ;
  assign n37499 = n32393 ^ n27155 ^ 1'b0 ;
  assign n37500 = n360 & ~n10969 ;
  assign n37501 = n10694 ^ n5939 ^ 1'b0 ;
  assign n37502 = x101 | n5620 ;
  assign n37503 = n4436 | n37502 ;
  assign n37504 = n37501 | n37503 ;
  assign n37505 = n37504 ^ n25909 ^ n19759 ;
  assign n37506 = n2875 & ~n6462 ;
  assign n37507 = n34334 ^ n19230 ^ 1'b0 ;
  assign n37508 = n8562 | n37507 ;
  assign n37509 = n23349 ^ n4593 ^ 1'b0 ;
  assign n37510 = n21663 & ~n37509 ;
  assign n37511 = n37510 ^ n5141 ^ 1'b0 ;
  assign n37512 = ~n1657 & n13195 ;
  assign n37513 = n10791 & ~n14110 ;
  assign n37514 = n3955 & n13426 ;
  assign n37515 = ~n13574 & n37514 ;
  assign n37516 = n4361 ^ n1697 ^ n617 ;
  assign n37517 = n13230 & n14858 ;
  assign n37518 = ~n37516 & n37517 ;
  assign n37519 = n20781 ^ n11567 ^ 1'b0 ;
  assign n37521 = n7225 ^ n1239 ^ 1'b0 ;
  assign n37522 = n13744 & n37521 ;
  assign n37523 = ~n3277 & n37522 ;
  assign n37520 = n791 | n6681 ;
  assign n37524 = n37523 ^ n37520 ^ 1'b0 ;
  assign n37525 = ~n4758 & n31097 ;
  assign n37526 = n37525 ^ n11408 ^ 1'b0 ;
  assign n37527 = n7686 & n18409 ;
  assign n37528 = ~n692 & n9853 ;
  assign n37529 = n14562 & ~n14911 ;
  assign n37530 = n5895 | n37529 ;
  assign n37531 = n972 & ~n37530 ;
  assign n37532 = n1188 | n30123 ;
  assign n37533 = n3947 & ~n37532 ;
  assign n37534 = n5452 & n17597 ;
  assign n37535 = n37534 ^ n7203 ^ 1'b0 ;
  assign n37536 = n1195 & n4007 ;
  assign n37537 = n37536 ^ n20010 ^ n3294 ;
  assign n37538 = ~n29066 & n37537 ;
  assign n37539 = ~n37535 & n37538 ;
  assign n37540 = n37539 ^ n5326 ^ 1'b0 ;
  assign n37541 = n35670 ^ n8112 ^ 1'b0 ;
  assign n37542 = ~n11396 & n37541 ;
  assign n37543 = ~n11607 & n20531 ;
  assign n37544 = n37543 ^ n13442 ^ 1'b0 ;
  assign n37545 = n19686 & n27695 ;
  assign n37546 = ~n24691 & n37545 ;
  assign n37547 = n12604 & ~n37546 ;
  assign n37548 = ( n5875 & n18053 ) | ( n5875 & ~n21560 ) | ( n18053 & ~n21560 ) ;
  assign n37549 = n37548 ^ n13528 ^ 1'b0 ;
  assign n37550 = n5411 | n37549 ;
  assign n37551 = n2431 | n13189 ;
  assign n37552 = n37551 ^ n20809 ^ 1'b0 ;
  assign n37553 = n20476 & n37552 ;
  assign n37554 = n37553 ^ n3967 ^ 1'b0 ;
  assign n37555 = n16443 & n29780 ;
  assign n37556 = n37555 ^ n1432 ^ 1'b0 ;
  assign n37557 = ~n790 & n23706 ;
  assign n37558 = n37556 | n37557 ;
  assign n37559 = n37558 ^ n11983 ^ 1'b0 ;
  assign n37560 = n19860 & ~n28632 ;
  assign n37561 = n37560 ^ n594 ^ 1'b0 ;
  assign n37562 = n14359 & n29144 ;
  assign n37563 = n18971 & n37562 ;
  assign n37564 = n17282 ^ n11516 ^ 1'b0 ;
  assign n37565 = ( ~n4721 & n10020 ) | ( ~n4721 & n20309 ) | ( n10020 & n20309 ) ;
  assign n37566 = n27295 ^ n6887 ^ n4137 ;
  assign n37567 = n37566 ^ n30032 ^ 1'b0 ;
  assign n37568 = n37567 ^ n23286 ^ n23111 ;
  assign n37569 = n13343 ^ n12542 ^ 1'b0 ;
  assign n37570 = n9483 | n34018 ;
  assign n37571 = ~n4027 & n16832 ;
  assign n37572 = n5252 & ~n37571 ;
  assign n37573 = x64 & n37572 ;
  assign n37574 = n1010 | n37573 ;
  assign n37575 = n6770 | n37574 ;
  assign n37576 = n37575 ^ n8212 ^ 1'b0 ;
  assign n37577 = n20123 ^ n5226 ^ 1'b0 ;
  assign n37578 = n1669 & ~n33296 ;
  assign n37579 = ~n30101 & n37578 ;
  assign n37580 = n6121 ^ n1380 ^ 1'b0 ;
  assign n37581 = n1453 & ~n32100 ;
  assign n37582 = n37581 ^ n10378 ^ 1'b0 ;
  assign n37583 = ( n1056 & n26715 ) | ( n1056 & n37582 ) | ( n26715 & n37582 ) ;
  assign n37584 = ~n1856 & n37583 ;
  assign n37585 = ( n2448 & n37580 ) | ( n2448 & n37584 ) | ( n37580 & n37584 ) ;
  assign n37587 = n28217 ^ n8101 ^ 1'b0 ;
  assign n37586 = n17817 & n20483 ;
  assign n37588 = n37587 ^ n37586 ^ n7206 ;
  assign n37589 = n23436 ^ n9241 ^ 1'b0 ;
  assign n37590 = ~n2097 & n27703 ;
  assign n37591 = ~n18337 & n37590 ;
  assign n37592 = n12024 ^ n1124 ^ 1'b0 ;
  assign n37593 = x94 & n32532 ;
  assign n37594 = ~n37592 & n37593 ;
  assign n37595 = n23946 & n36752 ;
  assign n37596 = n37595 ^ n37429 ^ 1'b0 ;
  assign n37597 = n18524 | n35081 ;
  assign n37598 = n19121 ^ n8159 ^ 1'b0 ;
  assign n37599 = ~n9068 & n20845 ;
  assign n37600 = n37599 ^ n14990 ^ 1'b0 ;
  assign n37601 = n37598 & ~n37600 ;
  assign n37602 = ( n17375 & ~n19100 ) | ( n17375 & n37036 ) | ( ~n19100 & n37036 ) ;
  assign n37603 = n23592 & ~n27295 ;
  assign n37604 = ~n10296 & n20493 ;
  assign n37605 = n7066 ^ n4180 ^ 1'b0 ;
  assign n37612 = n4727 ^ n1824 ^ 1'b0 ;
  assign n37606 = n8129 & ~n8461 ;
  assign n37607 = n991 | n37606 ;
  assign n37608 = n37607 ^ n31175 ^ 1'b0 ;
  assign n37609 = n25486 ^ n21383 ^ 1'b0 ;
  assign n37610 = n37608 | n37609 ;
  assign n37611 = n905 & ~n37610 ;
  assign n37613 = n37612 ^ n37611 ^ 1'b0 ;
  assign n37614 = n8330 & ~n13103 ;
  assign n37615 = ~n13757 & n37614 ;
  assign n37616 = n23110 ^ n12469 ^ 1'b0 ;
  assign n37617 = n37615 | n37616 ;
  assign n37618 = n21749 | n37617 ;
  assign n37619 = n26416 | n37618 ;
  assign n37620 = n37619 ^ n9722 ^ 1'b0 ;
  assign n37625 = n17128 ^ n9500 ^ n329 ;
  assign n37621 = n24071 ^ n7624 ^ 1'b0 ;
  assign n37622 = n4142 & ~n37621 ;
  assign n37623 = n37622 ^ n31919 ^ 1'b0 ;
  assign n37624 = n10757 & ~n37623 ;
  assign n37626 = n37625 ^ n37624 ^ 1'b0 ;
  assign n37627 = n1620 & n37626 ;
  assign n37628 = ~n17596 & n37627 ;
  assign n37629 = ~n13644 & n37628 ;
  assign n37630 = n3643 & n37629 ;
  assign n37631 = n23048 ^ n18514 ^ 1'b0 ;
  assign n37633 = ~n2663 & n25129 ;
  assign n37632 = ~n2774 & n16240 ;
  assign n37634 = n37633 ^ n37632 ^ 1'b0 ;
  assign n37635 = n2687 & n31759 ;
  assign n37636 = ~n30183 & n36502 ;
  assign n37637 = n26856 ^ n2664 ^ 1'b0 ;
  assign n37638 = n34693 & ~n37637 ;
  assign n37639 = n6295 & n21746 ;
  assign n37640 = ( n679 & n2789 ) | ( n679 & ~n17013 ) | ( n2789 & ~n17013 ) ;
  assign n37641 = ~n6505 & n7303 ;
  assign n37642 = ( n5958 & n12917 ) | ( n5958 & n20712 ) | ( n12917 & n20712 ) ;
  assign n37643 = n20757 & ~n37642 ;
  assign n37644 = ( n15960 & n18277 ) | ( n15960 & n26579 ) | ( n18277 & n26579 ) ;
  assign n37648 = n15275 & n21035 ;
  assign n37645 = ~n3196 & n9694 ;
  assign n37646 = n21411 & ~n37645 ;
  assign n37647 = n37646 ^ x139 ^ 1'b0 ;
  assign n37649 = n37648 ^ n37647 ^ n32044 ;
  assign n37650 = n3641 & n18238 ;
  assign n37651 = ( n4137 & n37649 ) | ( n4137 & n37650 ) | ( n37649 & n37650 ) ;
  assign n37653 = n18987 | n25921 ;
  assign n37652 = n5923 & ~n16841 ;
  assign n37654 = n37653 ^ n37652 ^ 1'b0 ;
  assign n37655 = ~n982 & n8154 ;
  assign n37656 = n4201 & n37655 ;
  assign n37657 = n5067 | n5469 ;
  assign n37658 = n15500 | n37657 ;
  assign n37659 = n27940 ^ n2609 ^ 1'b0 ;
  assign n37660 = n11053 ^ n3499 ^ 1'b0 ;
  assign n37661 = n37659 | n37660 ;
  assign n37662 = n26035 & ~n37661 ;
  assign n37663 = n37662 ^ n32088 ^ n9598 ;
  assign n37664 = ~n21005 & n37663 ;
  assign n37665 = n15642 ^ n1981 ^ 1'b0 ;
  assign n37666 = n37665 ^ n6842 ^ n5465 ;
  assign n37667 = n3598 ^ n3523 ^ 1'b0 ;
  assign n37668 = n3718 | n37667 ;
  assign n37669 = ( n27292 & ~n32957 ) | ( n27292 & n37668 ) | ( ~n32957 & n37668 ) ;
  assign n37670 = n10628 | n15802 ;
  assign n37671 = n32012 ^ n12518 ^ n10550 ;
  assign n37672 = n37671 ^ n20320 ^ n17823 ;
  assign n37673 = n19147 ^ n8340 ^ 1'b0 ;
  assign n37674 = n37672 & ~n37673 ;
  assign n37675 = n5843 & n7415 ;
  assign n37676 = n37675 ^ n21190 ^ 1'b0 ;
  assign n37677 = n5027 | n9537 ;
  assign n37678 = n37676 | n37677 ;
  assign n37679 = n12812 & n37678 ;
  assign n37680 = n18587 & n27726 ;
  assign n37681 = ~n37679 & n37680 ;
  assign n37682 = ( n4836 & n15234 ) | ( n4836 & n25519 ) | ( n15234 & n25519 ) ;
  assign n37683 = n1594 | n20883 ;
  assign n37684 = n37682 | n37683 ;
  assign n37685 = n2237 & ~n37684 ;
  assign n37686 = ~n7002 & n37685 ;
  assign n37687 = n6235 | n6667 ;
  assign n37688 = ( n5232 & n15829 ) | ( n5232 & ~n37687 ) | ( n15829 & ~n37687 ) ;
  assign n37689 = n37112 & n37688 ;
  assign n37690 = n37099 ^ n5939 ^ 1'b0 ;
  assign n37691 = n22836 & ~n37690 ;
  assign n37692 = n37689 & n37691 ;
  assign n37693 = n33101 ^ n26934 ^ 1'b0 ;
  assign n37694 = n32547 ^ n4352 ^ 1'b0 ;
  assign n37695 = n18270 & n23252 ;
  assign n37696 = n17124 ^ n3757 ^ n1733 ;
  assign n37697 = n37695 | n37696 ;
  assign n37698 = n27501 ^ n18225 ^ 1'b0 ;
  assign n37699 = n15489 & ~n17518 ;
  assign n37700 = n37699 ^ n35304 ^ 1'b0 ;
  assign n37701 = n15453 & n16054 ;
  assign n37702 = ~n35816 & n37701 ;
  assign n37703 = n13322 ^ n4440 ^ 1'b0 ;
  assign n37704 = n26060 ^ n5849 ^ n2311 ;
  assign n37705 = n6656 & n37704 ;
  assign n37706 = n21498 & n37705 ;
  assign n37707 = n18645 & n32762 ;
  assign n37708 = ~n30751 & n37707 ;
  assign n37709 = ~n16169 & n21879 ;
  assign n37710 = n23533 ^ n4368 ^ n3111 ;
  assign n37711 = n37710 ^ n9286 ^ 1'b0 ;
  assign n37712 = n25640 & ~n32117 ;
  assign n37714 = n2022 | n6869 ;
  assign n37715 = n37714 ^ n21177 ^ 1'b0 ;
  assign n37713 = n16126 | n29505 ;
  assign n37716 = n37715 ^ n37713 ^ 1'b0 ;
  assign n37717 = n13673 & ~n24263 ;
  assign n37718 = n37717 ^ n6811 ^ 1'b0 ;
  assign n37719 = n17788 & n22006 ;
  assign n37720 = n37719 ^ n2038 ^ 1'b0 ;
  assign n37721 = n24134 & n37720 ;
  assign n37722 = n37721 ^ n15178 ^ 1'b0 ;
  assign n37723 = ~n37718 & n37722 ;
  assign n37724 = n7883 & ~n8551 ;
  assign n37725 = n23798 & n33818 ;
  assign n37726 = n23619 & n37725 ;
  assign n37727 = n32910 ^ n5162 ^ n3533 ;
  assign n37728 = n37727 ^ n15722 ^ 1'b0 ;
  assign n37729 = n24833 ^ n3464 ^ n1023 ;
  assign n37730 = ~n23222 & n37729 ;
  assign n37733 = ~n7776 & n37115 ;
  assign n37731 = n26060 ^ n4026 ^ 1'b0 ;
  assign n37732 = ~n32738 & n37731 ;
  assign n37734 = n37733 ^ n37732 ^ 1'b0 ;
  assign n37735 = n12798 & ~n13937 ;
  assign n37736 = n37735 ^ n16836 ^ 1'b0 ;
  assign n37737 = ~n7791 & n33468 ;
  assign n37738 = n15005 ^ n3972 ^ 1'b0 ;
  assign n37739 = n23776 & ~n37738 ;
  assign n37740 = ( n14848 & n31915 ) | ( n14848 & ~n37739 ) | ( n31915 & ~n37739 ) ;
  assign n37741 = n3104 | n10398 ;
  assign n37742 = n37740 & ~n37741 ;
  assign n37743 = ( n12693 & ~n32899 ) | ( n12693 & n37742 ) | ( ~n32899 & n37742 ) ;
  assign n37744 = n3588 | n23978 ;
  assign n37745 = ~n10237 & n12515 ;
  assign n37746 = n24200 ^ n14513 ^ 1'b0 ;
  assign n37747 = n19540 ^ n17124 ^ 1'b0 ;
  assign n37748 = n37746 & n37747 ;
  assign n37749 = ~n1894 & n37748 ;
  assign n37750 = n37749 ^ n4145 ^ 1'b0 ;
  assign n37751 = n6950 ^ n3381 ^ 1'b0 ;
  assign n37752 = n6027 & ~n37751 ;
  assign n37753 = n18989 & n37752 ;
  assign n37754 = n37753 ^ n26895 ^ 1'b0 ;
  assign n37755 = ~n11827 & n18136 ;
  assign n37756 = n37755 ^ n23962 ^ 1'b0 ;
  assign n37757 = n37756 ^ n23860 ^ 1'b0 ;
  assign n37758 = n17411 & n37757 ;
  assign n37759 = n2578 ^ n1287 ^ 1'b0 ;
  assign n37760 = x225 & ~n37759 ;
  assign n37761 = n33964 ^ n11050 ^ 1'b0 ;
  assign n37762 = n22593 | n37761 ;
  assign n37763 = n37762 ^ n16296 ^ 1'b0 ;
  assign n37764 = n3769 ^ n482 ^ 1'b0 ;
  assign n37765 = ~n9826 & n9881 ;
  assign n37766 = ~n31290 & n37765 ;
  assign n37767 = n3983 | n24204 ;
  assign n37768 = n5119 | n37767 ;
  assign n37769 = n37768 ^ n29985 ^ 1'b0 ;
  assign n37770 = n5678 & ~n13167 ;
  assign n37771 = ~n32117 & n37770 ;
  assign n37772 = n18276 | n26178 ;
  assign n37776 = x177 & n15322 ;
  assign n37777 = n37776 ^ n3002 ^ 1'b0 ;
  assign n37773 = n880 & n2850 ;
  assign n37774 = ~n18893 & n28453 ;
  assign n37775 = n37773 & n37774 ;
  assign n37778 = n37777 ^ n37775 ^ n12184 ;
  assign n37779 = n12710 & ~n37359 ;
  assign n37780 = n37779 ^ n5474 ^ 1'b0 ;
  assign n37781 = n1782 | n35362 ;
  assign n37782 = n20964 ^ n2082 ^ 1'b0 ;
  assign n37783 = n12476 & ~n12998 ;
  assign n37784 = n17567 & n37783 ;
  assign n37785 = ~n9861 & n37784 ;
  assign n37786 = n37744 ^ n20292 ^ 1'b0 ;
  assign n37787 = n6131 ^ n6069 ^ n5221 ;
  assign n37788 = n17724 ^ n791 ^ 1'b0 ;
  assign n37789 = ~n18179 & n37788 ;
  assign n37790 = n2761 & n37789 ;
  assign n37791 = n13921 ^ n9388 ^ 1'b0 ;
  assign n37792 = n950 & ~n33799 ;
  assign n37793 = n12914 ^ n6366 ^ 1'b0 ;
  assign n37794 = n28628 & ~n37793 ;
  assign n37795 = n10552 | n32966 ;
  assign n37796 = n37794 | n37795 ;
  assign n37797 = n28706 ^ n13081 ^ n9103 ;
  assign n37798 = ( n6660 & n23172 ) | ( n6660 & ~n37797 ) | ( n23172 & ~n37797 ) ;
  assign n37799 = n37798 ^ n37676 ^ 1'b0 ;
  assign n37800 = n25340 ^ n8848 ^ 1'b0 ;
  assign n37801 = n37800 ^ n25897 ^ 1'b0 ;
  assign n37802 = n14027 ^ n11703 ^ 1'b0 ;
  assign n37803 = n17685 | n37802 ;
  assign n37804 = n2407 & n20771 ;
  assign n37805 = n10548 ^ n5200 ^ 1'b0 ;
  assign n37806 = n6313 & n37805 ;
  assign n37807 = n11901 & n37806 ;
  assign n37808 = n37807 ^ x133 ^ 1'b0 ;
  assign n37809 = n1442 | n37808 ;
  assign n37810 = n25673 | n37809 ;
  assign n37811 = n1164 & n19602 ;
  assign n37812 = n1613 | n37811 ;
  assign n37813 = n37812 ^ n371 ^ 1'b0 ;
  assign n37814 = n26484 ^ n1991 ^ 1'b0 ;
  assign n37815 = n28745 | n33835 ;
  assign n37816 = n14130 ^ n1999 ^ n1688 ;
  assign n37817 = ~n20292 & n37816 ;
  assign n37818 = n12112 ^ n2529 ^ 1'b0 ;
  assign n37819 = ~n13544 & n37818 ;
  assign n37820 = n12665 & n36522 ;
  assign n37821 = n2787 | n4789 ;
  assign n37822 = n12299 | n37821 ;
  assign n37823 = n23225 ^ n17336 ^ 1'b0 ;
  assign n37824 = n37822 & n37823 ;
  assign n37825 = n3706 & n13770 ;
  assign n37826 = ~n13770 & n37825 ;
  assign n37827 = n4184 | n9865 ;
  assign n37828 = n37826 & ~n37827 ;
  assign n37829 = ( n10709 & n20700 ) | ( n10709 & ~n37828 ) | ( n20700 & ~n37828 ) ;
  assign n37830 = ( n3383 & n37420 ) | ( n3383 & ~n37829 ) | ( n37420 & ~n37829 ) ;
  assign n37831 = ( ~n6425 & n17625 ) | ( ~n6425 & n37830 ) | ( n17625 & n37830 ) ;
  assign n37832 = n29296 ^ n13609 ^ 1'b0 ;
  assign n37833 = n10026 & n17948 ;
  assign n37834 = n37833 ^ n36072 ^ 1'b0 ;
  assign n37835 = n10582 & ~n37834 ;
  assign n37836 = n26989 ^ n21709 ^ 1'b0 ;
  assign n37837 = n907 & n37836 ;
  assign n37838 = n33348 & ~n37837 ;
  assign n37839 = n30071 ^ n4579 ^ 1'b0 ;
  assign n37840 = n34579 & n37839 ;
  assign n37841 = n5445 | n6389 ;
  assign n37842 = n8976 | n9862 ;
  assign n37843 = n2057 & n15437 ;
  assign n37844 = ( n21338 & n37842 ) | ( n21338 & ~n37843 ) | ( n37842 & ~n37843 ) ;
  assign n37845 = ( n13837 & n37841 ) | ( n13837 & n37844 ) | ( n37841 & n37844 ) ;
  assign n37846 = n16144 & n28299 ;
  assign n37847 = n37845 & n37846 ;
  assign n37848 = n17942 ^ n14747 ^ n14114 ;
  assign n37849 = n14613 ^ n2191 ^ 1'b0 ;
  assign n37850 = ( n12841 & n37848 ) | ( n12841 & ~n37849 ) | ( n37848 & ~n37849 ) ;
  assign n37851 = n37850 ^ n32745 ^ n4440 ;
  assign n37852 = n35961 ^ n34347 ^ n2929 ;
  assign n37853 = n28576 ^ n12778 ^ n747 ;
  assign n37855 = n4742 | n21275 ;
  assign n37856 = n6420 & ~n37855 ;
  assign n37854 = n5636 & ~n26322 ;
  assign n37857 = n37856 ^ n37854 ^ 1'b0 ;
  assign n37858 = ~n22478 & n25250 ;
  assign n37859 = n37858 ^ n22415 ^ 1'b0 ;
  assign n37860 = ~n3362 & n19232 ;
  assign n37861 = n37860 ^ n6338 ^ 1'b0 ;
  assign n37862 = ~n3048 & n10178 ;
  assign n37863 = n37862 ^ n28077 ^ 1'b0 ;
  assign n37864 = n23595 ^ n18207 ^ n11109 ;
  assign n37865 = ( ~n30513 & n37863 ) | ( ~n30513 & n37864 ) | ( n37863 & n37864 ) ;
  assign n37866 = ( n2428 & n14612 ) | ( n2428 & ~n28484 ) | ( n14612 & ~n28484 ) ;
  assign n37867 = n17694 ^ n3642 ^ 1'b0 ;
  assign n37868 = n4331 & ~n37867 ;
  assign n37869 = n3198 ^ n706 ^ 1'b0 ;
  assign n37870 = n22443 ^ n12189 ^ 1'b0 ;
  assign n37871 = n3473 & n37870 ;
  assign n37872 = n11266 & n37871 ;
  assign n37873 = n37872 ^ n7604 ^ 1'b0 ;
  assign n37874 = n6450 & n21210 ;
  assign n37875 = ~n37873 & n37874 ;
  assign n37876 = n18202 & ~n37875 ;
  assign n37877 = n15964 ^ n10585 ^ 1'b0 ;
  assign n37878 = n2553 ^ n1340 ^ 1'b0 ;
  assign n37879 = n11657 | n37878 ;
  assign n37880 = ( ~n10493 & n27136 ) | ( ~n10493 & n37879 ) | ( n27136 & n37879 ) ;
  assign n37881 = ~n302 & n4165 ;
  assign n37882 = n37881 ^ n34801 ^ 1'b0 ;
  assign n37883 = n37882 ^ n10501 ^ 1'b0 ;
  assign n37884 = n29935 ^ n10660 ^ 1'b0 ;
  assign n37885 = x196 & ~n37884 ;
  assign n37886 = n2907 & ~n26351 ;
  assign n37887 = n37886 ^ n23915 ^ 1'b0 ;
  assign n37888 = n28747 & n37887 ;
  assign n37889 = ( n12229 & n17418 ) | ( n12229 & ~n34673 ) | ( n17418 & ~n34673 ) ;
  assign n37893 = n5031 | n12899 ;
  assign n37890 = n10634 | n21812 ;
  assign n37891 = n17570 & ~n37890 ;
  assign n37892 = n37891 ^ n10305 ^ 1'b0 ;
  assign n37894 = n37893 ^ n37892 ^ n12082 ;
  assign n37895 = n17523 & ~n31480 ;
  assign n37896 = n4830 & n6348 ;
  assign n37897 = n34466 ^ n11169 ^ 1'b0 ;
  assign n37898 = n1808 | n37897 ;
  assign n37899 = n37898 ^ n24000 ^ 1'b0 ;
  assign n37900 = n11063 | n25609 ;
  assign n37901 = n37900 ^ n9018 ^ 1'b0 ;
  assign n37902 = ( n734 & n10961 ) | ( n734 & n37901 ) | ( n10961 & n37901 ) ;
  assign n37903 = n5207 ^ n4927 ^ 1'b0 ;
  assign n37904 = ~n3205 & n25634 ;
  assign n37905 = n37904 ^ n27598 ^ 1'b0 ;
  assign n37906 = ~n6381 & n11000 ;
  assign n37907 = n9429 & ~n37906 ;
  assign n37908 = n37907 ^ n23894 ^ 1'b0 ;
  assign n37909 = n22568 & ~n37908 ;
  assign n37910 = n37777 & n37909 ;
  assign n37911 = n4615 | n18303 ;
  assign n37912 = n22408 ^ n856 ^ 1'b0 ;
  assign n37913 = n25935 ^ n10689 ^ 1'b0 ;
  assign n37914 = n1046 | n37913 ;
  assign n37915 = n13930 & ~n37914 ;
  assign n37916 = n6724 ^ n4630 ^ 1'b0 ;
  assign n37917 = n37916 ^ n1024 ^ 1'b0 ;
  assign n37918 = ~n13603 & n37917 ;
  assign n37919 = n21358 ^ n13793 ^ 1'b0 ;
  assign n37920 = n6177 | n11161 ;
  assign n37921 = n13967 & ~n37920 ;
  assign n37922 = n16129 | n16307 ;
  assign n37923 = ~n23656 & n26046 ;
  assign n37924 = n37923 ^ n28021 ^ 1'b0 ;
  assign n37925 = n37922 | n37924 ;
  assign n37926 = n11792 ^ n11168 ^ 1'b0 ;
  assign n37931 = ~n7897 & n8594 ;
  assign n37932 = n2355 & ~n37931 ;
  assign n37927 = n3975 | n31027 ;
  assign n37928 = n20847 | n37927 ;
  assign n37929 = ~n20268 & n37928 ;
  assign n37930 = n37929 ^ n16343 ^ 1'b0 ;
  assign n37933 = n37932 ^ n37930 ^ x65 ;
  assign n37934 = n10464 ^ n5319 ^ 1'b0 ;
  assign n37935 = n37934 ^ n28265 ^ n3499 ;
  assign n37936 = n9314 | n20721 ;
  assign n37937 = n15933 ^ n4137 ^ 1'b0 ;
  assign n37938 = n37937 ^ n18265 ^ 1'b0 ;
  assign n37939 = ~n5095 & n37938 ;
  assign n37940 = ~n5496 & n21078 ;
  assign n37941 = n15258 ^ n12080 ^ 1'b0 ;
  assign n37942 = n5790 | n37941 ;
  assign n37943 = n37942 ^ n3530 ^ 1'b0 ;
  assign n37944 = n10095 ^ n4775 ^ 1'b0 ;
  assign n37945 = n13057 & ~n37944 ;
  assign n37946 = ~n37943 & n37945 ;
  assign n37947 = ( n16604 & n29497 ) | ( n16604 & n37946 ) | ( n29497 & n37946 ) ;
  assign n37948 = n4969 & ~n21937 ;
  assign n37949 = n5720 & n37948 ;
  assign n37950 = n23456 | n37949 ;
  assign n37951 = n37950 ^ n12760 ^ 1'b0 ;
  assign n37952 = ~n756 & n33248 ;
  assign n37953 = ~n37951 & n37952 ;
  assign n37954 = n36579 ^ n16489 ^ 1'b0 ;
  assign n37955 = n35921 & n37954 ;
  assign n37956 = n17859 & ~n20678 ;
  assign n37957 = n34122 & n37956 ;
  assign n37958 = n24914 ^ n8262 ^ 1'b0 ;
  assign n37959 = n2915 | n8399 ;
  assign n37960 = n37958 & ~n37959 ;
  assign n37962 = n556 | n29160 ;
  assign n37963 = n12121 | n37962 ;
  assign n37961 = n28829 ^ n8899 ^ n4984 ;
  assign n37964 = n37963 ^ n37961 ^ 1'b0 ;
  assign n37965 = n10233 & n14746 ;
  assign n37966 = ( ~n15654 & n18665 ) | ( ~n15654 & n37965 ) | ( n18665 & n37965 ) ;
  assign n37967 = n16820 | n26906 ;
  assign n37968 = ~n9280 & n35429 ;
  assign n37969 = n3133 & n37968 ;
  assign n37970 = n2553 | n37969 ;
  assign n37971 = n2218 & ~n10155 ;
  assign n37972 = n1851 & n37971 ;
  assign n37973 = n27976 | n29169 ;
  assign n37974 = n37972 | n37973 ;
  assign n37975 = n24576 & ~n37974 ;
  assign n37976 = n37970 | n37975 ;
  assign n37977 = n19161 ^ n10902 ^ 1'b0 ;
  assign n37978 = ~n1858 & n18857 ;
  assign n37979 = n7360 & n37978 ;
  assign n37980 = n1096 | n19029 ;
  assign n37981 = ~n21064 & n26512 ;
  assign n37982 = n8296 | n26137 ;
  assign n37983 = n3056 | n11923 ;
  assign n37984 = n13674 ^ n4758 ^ 1'b0 ;
  assign n37985 = n27496 ^ n4895 ^ 1'b0 ;
  assign n37986 = n11231 ^ n9413 ^ 1'b0 ;
  assign n37987 = n14278 & n37986 ;
  assign n37988 = n23949 & n37987 ;
  assign n37989 = ~n8537 & n24390 ;
  assign n37990 = n10532 | n12691 ;
  assign n37991 = n1550 & ~n13632 ;
  assign n37992 = ~n32624 & n37991 ;
  assign n37996 = n33924 ^ n25340 ^ n2726 ;
  assign n37997 = ( n21064 & n29370 ) | ( n21064 & ~n37996 ) | ( n29370 & ~n37996 ) ;
  assign n37993 = ~n10400 & n19940 ;
  assign n37994 = n29619 ^ n1483 ^ 1'b0 ;
  assign n37995 = ~n37993 & n37994 ;
  assign n37998 = n37997 ^ n37995 ^ n18789 ;
  assign n37999 = n32586 ^ n22302 ^ 1'b0 ;
  assign n38001 = n28443 ^ n3362 ^ 1'b0 ;
  assign n38000 = n8585 | n24273 ;
  assign n38002 = n38001 ^ n38000 ^ 1'b0 ;
  assign n38003 = n2829 & n29159 ;
  assign n38004 = ~n34332 & n38003 ;
  assign n38005 = n1618 & n16668 ;
  assign n38006 = ~n25422 & n38005 ;
  assign n38007 = n909 & n38006 ;
  assign n38008 = n16879 ^ n1376 ^ 1'b0 ;
  assign n38009 = ( n6057 & n32482 ) | ( n6057 & n38008 ) | ( n32482 & n38008 ) ;
  assign n38010 = n9544 & ~n25953 ;
  assign n38011 = n2592 & n38010 ;
  assign n38012 = n642 & ~n24937 ;
  assign n38013 = n33866 ^ n6372 ^ 1'b0 ;
  assign n38014 = n6035 | n14092 ;
  assign n38015 = ( n4378 & ~n8898 ) | ( n4378 & n38014 ) | ( ~n8898 & n38014 ) ;
  assign n38016 = n27386 & n38015 ;
  assign n38017 = n38016 ^ n17178 ^ 1'b0 ;
  assign n38018 = n30871 ^ n10050 ^ 1'b0 ;
  assign n38019 = ~n3288 & n6609 ;
  assign n38020 = ~n17398 & n38019 ;
  assign n38021 = ( n25461 & ~n27296 ) | ( n25461 & n38020 ) | ( ~n27296 & n38020 ) ;
  assign n38022 = n11973 & ~n13744 ;
  assign n38023 = n38022 ^ n18867 ^ 1'b0 ;
  assign n38024 = n4537 & n35866 ;
  assign n38025 = ~n277 & n38024 ;
  assign n38026 = n5775 | n13353 ;
  assign n38027 = n38026 ^ n16407 ^ 1'b0 ;
  assign n38028 = n11758 | n33680 ;
  assign n38029 = ~n286 & n18089 ;
  assign n38030 = ~n11317 & n38029 ;
  assign n38031 = n20196 ^ n3362 ^ 1'b0 ;
  assign n38032 = ~n4903 & n38031 ;
  assign n38033 = n6610 ^ n1406 ^ 1'b0 ;
  assign n38034 = n2103 & n38033 ;
  assign n38035 = n38034 ^ n23151 ^ n13856 ;
  assign n38036 = n32292 | n37573 ;
  assign n38037 = x250 & ~n4397 ;
  assign n38038 = n38037 ^ n19510 ^ 1'b0 ;
  assign n38039 = n5672 ^ n3942 ^ 1'b0 ;
  assign n38040 = n38038 | n38039 ;
  assign n38041 = n5895 & n6615 ;
  assign n38042 = n31052 & n38041 ;
  assign n38043 = n3453 & ~n5151 ;
  assign n38044 = n38043 ^ n14949 ^ 1'b0 ;
  assign n38045 = n38042 | n38044 ;
  assign n38046 = n19245 ^ n11638 ^ 1'b0 ;
  assign n38047 = ~n11394 & n38046 ;
  assign n38048 = n6372 | n37284 ;
  assign n38049 = ( n7012 & n8372 ) | ( n7012 & n34654 ) | ( n8372 & n34654 ) ;
  assign n38050 = n38049 ^ n3333 ^ 1'b0 ;
  assign n38051 = n29971 ^ n16126 ^ 1'b0 ;
  assign n38052 = n25512 ^ n20425 ^ 1'b0 ;
  assign n38053 = n7826 | n9611 ;
  assign n38054 = n9113 ^ n6200 ^ 1'b0 ;
  assign n38055 = n4759 | n38054 ;
  assign n38056 = n38055 ^ n1524 ^ 1'b0 ;
  assign n38057 = n38053 | n38056 ;
  assign n38058 = ~n10486 & n21739 ;
  assign n38059 = n38058 ^ n27064 ^ 1'b0 ;
  assign n38060 = n12961 ^ n6910 ^ 1'b0 ;
  assign n38061 = ~n10917 & n38060 ;
  assign n38062 = ( ~n311 & n6863 ) | ( ~n311 & n9429 ) | ( n6863 & n9429 ) ;
  assign n38063 = n38062 ^ n9447 ^ 1'b0 ;
  assign n38064 = n38061 & n38063 ;
  assign n38065 = ~n13404 & n38064 ;
  assign n38066 = n38065 ^ n1729 ^ 1'b0 ;
  assign n38067 = ~n6096 & n22987 ;
  assign n38068 = ( n20747 & n28320 ) | ( n20747 & ~n38067 ) | ( n28320 & ~n38067 ) ;
  assign n38069 = n25091 ^ n3685 ^ 1'b0 ;
  assign n38070 = n38068 & ~n38069 ;
  assign n38071 = n34166 ^ x0 ^ 1'b0 ;
  assign n38072 = n38071 ^ n2411 ^ 1'b0 ;
  assign n38073 = ~n768 & n38072 ;
  assign n38074 = n6972 & ~n9772 ;
  assign n38075 = ~n38073 & n38074 ;
  assign n38076 = n38075 ^ n10835 ^ n5594 ;
  assign n38077 = n37374 ^ n2732 ^ 1'b0 ;
  assign n38078 = ~n30746 & n34527 ;
  assign n38079 = n20832 & n38078 ;
  assign n38080 = n20755 ^ n10598 ^ 1'b0 ;
  assign n38081 = n1965 | n38080 ;
  assign n38082 = n1486 & ~n23964 ;
  assign n38083 = n38081 & n38082 ;
  assign n38085 = ~n19765 & n36617 ;
  assign n38084 = n18449 | n22759 ;
  assign n38086 = n38085 ^ n38084 ^ 1'b0 ;
  assign n38087 = n19034 ^ n9451 ^ 1'b0 ;
  assign n38088 = n11458 & ~n38087 ;
  assign n38089 = n3926 ^ n283 ^ 1'b0 ;
  assign n38090 = n38088 & n38089 ;
  assign n38091 = n8451 ^ n4260 ^ 1'b0 ;
  assign n38092 = n8216 & ~n38091 ;
  assign n38093 = n31950 ^ n30760 ^ n1603 ;
  assign n38094 = n38093 ^ n18867 ^ n480 ;
  assign n38095 = n694 | n7306 ;
  assign n38096 = n2814 & ~n38095 ;
  assign n38097 = n5639 | n38096 ;
  assign n38098 = n7475 | n38097 ;
  assign n38099 = ~n17391 & n38098 ;
  assign n38100 = n20850 & n22449 ;
  assign n38101 = n3469 & ~n13004 ;
  assign n38102 = n38101 ^ n16127 ^ 1'b0 ;
  assign n38103 = ( n9012 & n31397 ) | ( n9012 & n38102 ) | ( n31397 & n38102 ) ;
  assign n38104 = n31717 & ~n38103 ;
  assign n38105 = n38104 ^ n5953 ^ 1'b0 ;
  assign n38106 = n20464 ^ n10079 ^ n7708 ;
  assign n38107 = n13706 ^ n1720 ^ 1'b0 ;
  assign n38108 = n38107 ^ n13181 ^ n423 ;
  assign n38110 = ~n3032 & n16563 ;
  assign n38109 = n2738 & ~n12942 ;
  assign n38111 = n38110 ^ n38109 ^ 1'b0 ;
  assign n38112 = n38111 ^ n13921 ^ n7842 ;
  assign n38113 = n15460 | n28488 ;
  assign n38114 = n38112 & n38113 ;
  assign n38115 = n4806 ^ x10 ^ 1'b0 ;
  assign n38116 = n7997 | n13167 ;
  assign n38117 = n29982 ^ n1557 ^ 1'b0 ;
  assign n38118 = n38116 | n38117 ;
  assign n38119 = n4298 | n8018 ;
  assign n38120 = ~n5441 & n26390 ;
  assign n38121 = n6912 ^ n5410 ^ 1'b0 ;
  assign n38122 = n38121 ^ n20427 ^ 1'b0 ;
  assign n38123 = ( n5538 & ~n9786 ) | ( n5538 & n10923 ) | ( ~n9786 & n10923 ) ;
  assign n38124 = n12486 ^ n1572 ^ 1'b0 ;
  assign n38125 = n16022 & n35429 ;
  assign n38126 = n15542 ^ n2642 ^ n1343 ;
  assign n38127 = n37312 ^ n15803 ^ 1'b0 ;
  assign n38128 = ~n2296 & n4749 ;
  assign n38129 = n15183 ^ n10609 ^ 1'b0 ;
  assign n38130 = n38128 | n38129 ;
  assign n38131 = n23408 ^ n22859 ^ 1'b0 ;
  assign n38132 = n12562 | n38131 ;
  assign n38133 = ~n6617 & n38132 ;
  assign n38134 = ~n9249 & n23776 ;
  assign n38135 = n38134 ^ n10434 ^ 1'b0 ;
  assign n38136 = n38135 ^ n5019 ^ 1'b0 ;
  assign n38137 = n22510 ^ n5248 ^ 1'b0 ;
  assign n38138 = n38136 & n38137 ;
  assign n38139 = n35328 ^ n7313 ^ 1'b0 ;
  assign n38140 = n2322 & ~n19658 ;
  assign n38141 = ( n4879 & n8178 ) | ( n4879 & n31782 ) | ( n8178 & n31782 ) ;
  assign n38142 = n38140 | n38141 ;
  assign n38143 = n21921 ^ n18119 ^ 1'b0 ;
  assign n38144 = ( ~n24548 & n25656 ) | ( ~n24548 & n38143 ) | ( n25656 & n38143 ) ;
  assign n38145 = n6453 & n26501 ;
  assign n38146 = n38145 ^ n24079 ^ 1'b0 ;
  assign n38147 = n38146 ^ n7095 ^ n3097 ;
  assign n38148 = n23688 ^ n11863 ^ 1'b0 ;
  assign n38149 = n4628 & n20544 ;
  assign n38150 = n462 & n4342 ;
  assign n38151 = n8215 | n38150 ;
  assign n38153 = ( n16413 & ~n19367 ) | ( n16413 & n35295 ) | ( ~n19367 & n35295 ) ;
  assign n38152 = n22579 & ~n35826 ;
  assign n38154 = n38153 ^ n38152 ^ 1'b0 ;
  assign n38155 = n29413 ^ n2847 ^ 1'b0 ;
  assign n38156 = ( ~n7613 & n14325 ) | ( ~n7613 & n33781 ) | ( n14325 & n33781 ) ;
  assign n38157 = n9379 & n18812 ;
  assign n38158 = n38157 ^ n11912 ^ 1'b0 ;
  assign n38159 = n38158 ^ n11359 ^ n10840 ;
  assign n38160 = n13637 | n38159 ;
  assign n38161 = n32452 & ~n34930 ;
  assign n38162 = n12177 | n15836 ;
  assign n38163 = n24625 ^ n9482 ^ 1'b0 ;
  assign n38164 = ~n38162 & n38163 ;
  assign n38167 = ~n288 & n13284 ;
  assign n38165 = n6369 | n23865 ;
  assign n38166 = n12357 & ~n38165 ;
  assign n38168 = n38167 ^ n38166 ^ 1'b0 ;
  assign n38169 = ~n4286 & n8672 ;
  assign n38170 = n15887 & n38169 ;
  assign n38171 = n38170 ^ n24328 ^ 1'b0 ;
  assign n38172 = ( n27501 & n29477 ) | ( n27501 & n38171 ) | ( n29477 & n38171 ) ;
  assign n38173 = n20036 ^ n634 ^ 1'b0 ;
  assign n38174 = n13708 | n38173 ;
  assign n38175 = n2107 & ~n38174 ;
  assign n38176 = n22408 | n26098 ;
  assign n38177 = n1722 & ~n7700 ;
  assign n38178 = n38177 ^ n30679 ^ 1'b0 ;
  assign n38179 = n24537 & n30169 ;
  assign n38180 = n29438 & n38179 ;
  assign n38181 = n12937 | n29275 ;
  assign n38182 = n38181 ^ n478 ^ 1'b0 ;
  assign n38183 = n16118 & ~n38182 ;
  assign n38184 = n38183 ^ n32432 ^ 1'b0 ;
  assign n38185 = ~n29193 & n38184 ;
  assign n38186 = n15983 & n38185 ;
  assign n38187 = n5020 & n6443 ;
  assign n38188 = n38187 ^ n8554 ^ 1'b0 ;
  assign n38189 = n38188 ^ n22907 ^ n3773 ;
  assign n38190 = n1010 & ~n11228 ;
  assign n38191 = n6997 & n38190 ;
  assign n38192 = ( ~n9316 & n36994 ) | ( ~n9316 & n38191 ) | ( n36994 & n38191 ) ;
  assign n38193 = n12921 & n38192 ;
  assign n38194 = n4070 | n23698 ;
  assign n38195 = n38194 ^ n31638 ^ 1'b0 ;
  assign n38196 = ( n12774 & n14732 ) | ( n12774 & ~n22067 ) | ( n14732 & ~n22067 ) ;
  assign n38197 = n38196 ^ n16676 ^ n11434 ;
  assign n38198 = n38197 ^ n11259 ^ 1'b0 ;
  assign n38199 = n1543 & n13070 ;
  assign n38200 = n5176 & n38199 ;
  assign n38201 = ~n10227 & n38200 ;
  assign n38202 = ~n10228 & n17369 ;
  assign n38203 = n16261 & n38202 ;
  assign n38204 = n38203 ^ n5243 ^ 1'b0 ;
  assign n38205 = n13581 ^ n8245 ^ 1'b0 ;
  assign n38206 = n31739 ^ n26855 ^ n1270 ;
  assign n38207 = n1401 | n8956 ;
  assign n38208 = n29663 | n34760 ;
  assign n38209 = ( n2006 & ~n2748 ) | ( n2006 & n8694 ) | ( ~n2748 & n8694 ) ;
  assign n38210 = n10539 | n11249 ;
  assign n38211 = n21278 | n38210 ;
  assign n38212 = n38211 ^ n17489 ^ 1'b0 ;
  assign n38213 = n38209 & n38212 ;
  assign n38216 = n18516 ^ n3775 ^ 1'b0 ;
  assign n38217 = n15876 | n38216 ;
  assign n38214 = n2052 | n6947 ;
  assign n38215 = ( ~n2810 & n13380 ) | ( ~n2810 & n38214 ) | ( n13380 & n38214 ) ;
  assign n38218 = n38217 ^ n38215 ^ 1'b0 ;
  assign n38219 = n14846 & ~n15408 ;
  assign n38220 = n9011 & n38219 ;
  assign n38221 = n10573 & ~n24449 ;
  assign n38222 = n38221 ^ n5818 ^ 1'b0 ;
  assign n38223 = ~n38220 & n38222 ;
  assign n38224 = ~n12566 & n38223 ;
  assign n38225 = n8914 ^ n6035 ^ 1'b0 ;
  assign n38226 = n11954 ^ n2486 ^ 1'b0 ;
  assign n38227 = n1736 & n38226 ;
  assign n38228 = ( n5039 & n37622 ) | ( n5039 & n38227 ) | ( n37622 & n38227 ) ;
  assign n38229 = n13733 ^ n5804 ^ x83 ;
  assign n38230 = n38229 ^ n19778 ^ 1'b0 ;
  assign n38231 = n38230 ^ n18610 ^ n3725 ;
  assign n38232 = n284 & n22343 ;
  assign n38233 = n38232 ^ n33109 ^ n9401 ;
  assign n38234 = n16607 & ~n27449 ;
  assign n38235 = n9097 & n38234 ;
  assign n38236 = n23441 ^ n19033 ^ 1'b0 ;
  assign n38237 = ~n5288 & n38236 ;
  assign n38238 = x222 & ~n34970 ;
  assign n38239 = n38238 ^ n26276 ^ 1'b0 ;
  assign n38240 = ( n5051 & n11807 ) | ( n5051 & n16335 ) | ( n11807 & n16335 ) ;
  assign n38241 = n15140 & ~n19438 ;
  assign n38242 = n7752 & n38241 ;
  assign n38243 = n17225 | n33913 ;
  assign n38244 = n500 & ~n38243 ;
  assign n38245 = ( ~n35108 & n37059 ) | ( ~n35108 & n38244 ) | ( n37059 & n38244 ) ;
  assign n38246 = n29545 ^ n307 ^ 1'b0 ;
  assign n38247 = n17243 ^ n15705 ^ 1'b0 ;
  assign n38248 = n12718 ^ n10709 ^ 1'b0 ;
  assign n38250 = n1049 | n3104 ;
  assign n38251 = n3814 & ~n38250 ;
  assign n38252 = ( n4302 & n4641 ) | ( n4302 & n38251 ) | ( n4641 & n38251 ) ;
  assign n38249 = ~n1120 & n5817 ;
  assign n38253 = n38252 ^ n38249 ^ 1'b0 ;
  assign n38254 = n38253 ^ n12344 ^ 1'b0 ;
  assign n38255 = ~n835 & n38254 ;
  assign n38256 = n2816 & ~n25045 ;
  assign n38257 = ( n19551 & ~n29122 ) | ( n19551 & n38256 ) | ( ~n29122 & n38256 ) ;
  assign n38258 = n11934 & ~n38257 ;
  assign n38259 = ~n38255 & n38258 ;
  assign n38260 = n608 & ~n9995 ;
  assign n38261 = n38260 ^ n28257 ^ 1'b0 ;
  assign n38262 = n1377 & ~n24815 ;
  assign n38263 = ~n25493 & n38262 ;
  assign n38264 = n7787 & ~n34968 ;
  assign n38265 = n23353 ^ n15462 ^ 1'b0 ;
  assign n38266 = n29128 & n33597 ;
  assign n38267 = ~n5350 & n32630 ;
  assign n38268 = n38267 ^ n21515 ^ 1'b0 ;
  assign n38269 = n38266 | n38268 ;
  assign n38270 = n4343 & ~n25892 ;
  assign n38271 = n30462 ^ n27693 ^ n11305 ;
  assign n38272 = n8066 ^ n4240 ^ 1'b0 ;
  assign n38273 = n3803 ^ n2735 ^ 1'b0 ;
  assign n38274 = n38273 ^ n2664 ^ 1'b0 ;
  assign n38275 = x5 & n11519 ;
  assign n38276 = n32432 ^ n5710 ^ 1'b0 ;
  assign n38277 = n22559 & n38276 ;
  assign n38279 = n19026 ^ n12212 ^ n5586 ;
  assign n38278 = n5986 & ~n21293 ;
  assign n38280 = n38279 ^ n38278 ^ 1'b0 ;
  assign n38281 = n5213 | n23432 ;
  assign n38282 = ~n4031 & n38281 ;
  assign n38283 = n12261 & n22172 ;
  assign n38284 = ~n14445 & n38283 ;
  assign n38285 = n8653 & ~n38284 ;
  assign n38286 = n38285 ^ n16001 ^ 1'b0 ;
  assign n38287 = n26715 ^ n11073 ^ n9702 ;
  assign n38289 = n2174 ^ n1369 ^ 1'b0 ;
  assign n38288 = n26339 ^ n18498 ^ 1'b0 ;
  assign n38290 = n38289 ^ n38288 ^ n3236 ;
  assign n38291 = n9639 & n24535 ;
  assign n38292 = ~n4136 & n38291 ;
  assign n38293 = n38292 ^ n24900 ^ 1'b0 ;
  assign n38294 = n11341 | n18768 ;
  assign n38295 = n10348 ^ n7534 ^ 1'b0 ;
  assign n38296 = n19757 & ~n38295 ;
  assign n38297 = n3023 & ~n8294 ;
  assign n38298 = n3662 & n38297 ;
  assign n38299 = n10632 | n18279 ;
  assign n38300 = ( n3499 & n9215 ) | ( n3499 & n10081 ) | ( n9215 & n10081 ) ;
  assign n38301 = ( n6997 & n19317 ) | ( n6997 & n38300 ) | ( n19317 & n38300 ) ;
  assign n38302 = n38301 ^ n7398 ^ 1'b0 ;
  assign n38303 = ~n38299 & n38302 ;
  assign n38304 = ~n35424 & n38303 ;
  assign n38305 = n8101 ^ x41 ^ 1'b0 ;
  assign n38306 = n10363 ^ n5907 ^ n2495 ;
  assign n38307 = n7930 & n38306 ;
  assign n38308 = n5865 & n38307 ;
  assign n38309 = n1574 & ~n38308 ;
  assign n38310 = n12500 ^ n5327 ^ 1'b0 ;
  assign n38311 = n38310 ^ n37304 ^ n4765 ;
  assign n38312 = n12503 & n26244 ;
  assign n38314 = ~n3675 & n17375 ;
  assign n38313 = n20349 ^ n16821 ^ n7031 ;
  assign n38315 = n38314 ^ n38313 ^ n32441 ;
  assign n38316 = ~n4729 & n6936 ;
  assign n38317 = n31704 ^ n9338 ^ 1'b0 ;
  assign n38318 = ~n38316 & n38317 ;
  assign n38319 = n29212 & n37602 ;
  assign n38320 = n38319 ^ n2347 ^ 1'b0 ;
  assign n38321 = ~n28311 & n34224 ;
  assign n38322 = n38321 ^ n3683 ^ 1'b0 ;
  assign n38323 = n9790 | n12039 ;
  assign n38324 = n7575 | n38323 ;
  assign n38325 = n30407 & n38324 ;
  assign n38326 = n15159 | n35258 ;
  assign n38328 = ( n9945 & n13844 ) | ( n9945 & n15087 ) | ( n13844 & n15087 ) ;
  assign n38329 = n10560 & ~n38328 ;
  assign n38330 = n17023 & n38329 ;
  assign n38331 = n13492 & ~n38330 ;
  assign n38327 = ~n10586 & n16735 ;
  assign n38332 = n38331 ^ n38327 ^ 1'b0 ;
  assign n38333 = ( n24392 & n25480 ) | ( n24392 & ~n38332 ) | ( n25480 & ~n38332 ) ;
  assign n38334 = ~n13589 & n18424 ;
  assign n38335 = n38334 ^ n1553 ^ 1'b0 ;
  assign n38336 = ~n6319 & n38335 ;
  assign n38337 = n4868 & ~n25218 ;
  assign n38338 = ~n19191 & n38337 ;
  assign n38339 = n5791 & n6607 ;
  assign n38340 = n38339 ^ n26258 ^ n3079 ;
  assign n38341 = n11509 ^ n2930 ^ 1'b0 ;
  assign n38342 = n25682 & ~n38341 ;
  assign n38343 = n38340 & n38342 ;
  assign n38344 = ~n10555 & n17266 ;
  assign n38345 = n1155 | n4694 ;
  assign n38346 = ~n38344 & n38345 ;
  assign n38347 = n3659 & n38346 ;
  assign n38348 = n5102 & n37324 ;
  assign n38349 = n11344 | n38348 ;
  assign n38350 = n6696 & ~n18465 ;
  assign n38351 = n38350 ^ n25167 ^ n15080 ;
  assign n38352 = n12080 ^ n9788 ^ 1'b0 ;
  assign n38353 = n34588 & ~n38352 ;
  assign n38354 = n37182 ^ n2739 ^ 1'b0 ;
  assign n38355 = n26280 & n29207 ;
  assign n38356 = n36828 & n38355 ;
  assign n38357 = ~n6057 & n13483 ;
  assign n38364 = n1884 | n7724 ;
  assign n38365 = x160 & ~n38364 ;
  assign n38362 = n30548 ^ n5893 ^ x76 ;
  assign n38358 = ~n9911 & n19054 ;
  assign n38359 = n38358 ^ n35183 ^ 1'b0 ;
  assign n38360 = n20269 ^ n8288 ^ 1'b0 ;
  assign n38361 = n38359 & ~n38360 ;
  assign n38363 = n38362 ^ n38361 ^ n13733 ;
  assign n38366 = n38365 ^ n38363 ^ n1347 ;
  assign n38367 = n22139 ^ n4969 ^ n4582 ;
  assign n38368 = n22769 ^ n16284 ^ 1'b0 ;
  assign n38369 = ~x110 & n5386 ;
  assign n38370 = n35760 & ~n38369 ;
  assign n38371 = n38370 ^ n22394 ^ 1'b0 ;
  assign n38372 = ( n4732 & n21673 ) | ( n4732 & n24872 ) | ( n21673 & n24872 ) ;
  assign n38373 = n38372 ^ n25320 ^ 1'b0 ;
  assign n38374 = n30225 | n33837 ;
  assign n38375 = n5920 & n29879 ;
  assign n38376 = ~n16764 & n38375 ;
  assign n38377 = n29220 & ~n38376 ;
  assign n38378 = x118 & ~n896 ;
  assign n38379 = ~n21644 & n38378 ;
  assign n38380 = ~n9747 & n25221 ;
  assign n38381 = n38380 ^ n15197 ^ 1'b0 ;
  assign n38382 = n14909 ^ n1281 ^ 1'b0 ;
  assign n38383 = x192 & n38382 ;
  assign n38384 = n38383 ^ n8030 ^ 1'b0 ;
  assign n38385 = n20841 & n35552 ;
  assign n38386 = ~n32746 & n38385 ;
  assign n38387 = n6833 | n33566 ;
  assign n38388 = n14955 & ~n33431 ;
  assign n38389 = n27714 & n38388 ;
  assign n38391 = ~n4896 & n18690 ;
  assign n38390 = n2499 & n22566 ;
  assign n38392 = n38391 ^ n38390 ^ n21851 ;
  assign n38393 = ( n3193 & n4819 ) | ( n3193 & n8891 ) | ( n4819 & n8891 ) ;
  assign n38394 = n4124 & ~n6725 ;
  assign n38395 = n38393 & n38394 ;
  assign n38396 = n38395 ^ n12209 ^ n7146 ;
  assign n38397 = n12204 & ~n26781 ;
  assign n38398 = ~n18348 & n34078 ;
  assign n38399 = n38398 ^ n17846 ^ 1'b0 ;
  assign n38400 = ~n2966 & n38199 ;
  assign n38401 = n38400 ^ n21245 ^ n16883 ;
  assign n38402 = n27940 ^ n8067 ^ 1'b0 ;
  assign n38403 = n18003 & ~n38402 ;
  assign n38404 = ~n26323 & n35673 ;
  assign n38405 = n38335 & n38404 ;
  assign n38406 = n16739 ^ n8471 ^ 1'b0 ;
  assign n38408 = n24355 ^ n8768 ^ 1'b0 ;
  assign n38407 = ( n3403 & n5415 ) | ( n3403 & ~n33360 ) | ( n5415 & ~n33360 ) ;
  assign n38409 = n38408 ^ n38407 ^ 1'b0 ;
  assign n38410 = n16217 & n38409 ;
  assign n38411 = n16914 & n38410 ;
  assign n38412 = n6646 & n11838 ;
  assign n38413 = ~n2658 & n38412 ;
  assign n38414 = n20675 ^ n7968 ^ 1'b0 ;
  assign n38415 = ~n15520 & n38414 ;
  assign n38416 = n2727 | n38415 ;
  assign n38417 = n18254 & ~n38416 ;
  assign n38418 = n38417 ^ n6520 ^ 1'b0 ;
  assign n38419 = n27587 | n38418 ;
  assign n38420 = n38419 ^ n4508 ^ 1'b0 ;
  assign n38421 = ( n4347 & ~n6964 ) | ( n4347 & n8022 ) | ( ~n6964 & n8022 ) ;
  assign n38422 = n38421 ^ n24707 ^ n3474 ;
  assign n38423 = n9680 | n38422 ;
  assign n38424 = ~n12733 & n38423 ;
  assign n38426 = n4884 | n5826 ;
  assign n38427 = ~n3884 & n4674 ;
  assign n38428 = n38426 & n38427 ;
  assign n38425 = n1782 & n5145 ;
  assign n38429 = n38428 ^ n38425 ^ 1'b0 ;
  assign n38430 = n23866 | n33307 ;
  assign n38431 = n20826 ^ n751 ^ 1'b0 ;
  assign n38432 = n38354 ^ n24275 ^ 1'b0 ;
  assign n38433 = n1831 & ~n5673 ;
  assign n38434 = n38433 ^ n29578 ^ 1'b0 ;
  assign n38435 = n25250 & n38434 ;
  assign n38436 = n26668 ^ n21374 ^ n18320 ;
  assign n38437 = ( ~n6624 & n21736 ) | ( ~n6624 & n38436 ) | ( n21736 & n38436 ) ;
  assign n38438 = ( n732 & ~n1432 ) | ( n732 & n2202 ) | ( ~n1432 & n2202 ) ;
  assign n38443 = n4458 & n4656 ;
  assign n38444 = n21951 & n38443 ;
  assign n38445 = n38444 ^ n28325 ^ n12283 ;
  assign n38446 = n17125 & ~n38445 ;
  assign n38439 = n26492 ^ n15649 ^ n4021 ;
  assign n38440 = n38439 ^ n13172 ^ 1'b0 ;
  assign n38441 = n29326 | n38440 ;
  assign n38442 = n1310 & ~n38441 ;
  assign n38447 = n38446 ^ n38442 ^ 1'b0 ;
  assign n38448 = n38438 | n38447 ;
  assign n38449 = n28573 ^ n14537 ^ 1'b0 ;
  assign n38450 = n31611 & n38449 ;
  assign n38451 = n26876 | n37704 ;
  assign n38452 = n38451 ^ n6122 ^ 1'b0 ;
  assign n38453 = ~n19808 & n22901 ;
  assign n38454 = n38453 ^ n3104 ^ 1'b0 ;
  assign n38455 = n21036 & n38454 ;
  assign n38456 = ~n7233 & n38455 ;
  assign n38457 = ~n22219 & n38456 ;
  assign n38458 = n18595 ^ n11290 ^ 1'b0 ;
  assign n38459 = n10321 & ~n38458 ;
  assign n38460 = ~n12704 & n38459 ;
  assign n38461 = ~n1900 & n4294 ;
  assign n38462 = n22996 & n38461 ;
  assign n38463 = n30702 ^ n3434 ^ 1'b0 ;
  assign n38464 = n38462 & n38463 ;
  assign n38465 = n8683 ^ n1648 ^ 1'b0 ;
  assign n38466 = n27568 ^ n3686 ^ 1'b0 ;
  assign n38467 = n11379 & n18205 ;
  assign n38468 = n1462 & ~n9640 ;
  assign n38469 = ( n32039 & n36355 ) | ( n32039 & ~n38468 ) | ( n36355 & ~n38468 ) ;
  assign n38470 = n24969 ^ n20976 ^ n13612 ;
  assign n38471 = ( n15326 & ~n23244 ) | ( n15326 & n24306 ) | ( ~n23244 & n24306 ) ;
  assign n38472 = n38471 ^ n32487 ^ 1'b0 ;
  assign n38473 = ( ~n5166 & n32718 ) | ( ~n5166 & n33183 ) | ( n32718 & n33183 ) ;
  assign n38474 = n38473 ^ n1406 ^ 1'b0 ;
  assign n38475 = n1091 & n38474 ;
  assign n38476 = n38472 & n38475 ;
  assign n38477 = n11656 & ~n26513 ;
  assign n38478 = n30551 ^ n28614 ^ 1'b0 ;
  assign n38479 = n7836 & n38478 ;
  assign n38480 = ~n2406 & n38479 ;
  assign n38481 = n38480 ^ n27506 ^ 1'b0 ;
  assign n38482 = n10529 | n20706 ;
  assign n38483 = n10095 & ~n38482 ;
  assign n38484 = ( n970 & n12002 ) | ( n970 & ~n38483 ) | ( n12002 & ~n38483 ) ;
  assign n38485 = n38484 ^ n10996 ^ n3572 ;
  assign n38486 = n38485 ^ n21150 ^ 1'b0 ;
  assign n38487 = n31236 ^ n15569 ^ n6388 ;
  assign n38488 = n22715 ^ n11963 ^ 1'b0 ;
  assign n38489 = n27033 | n38488 ;
  assign n38490 = n2744 & ~n38489 ;
  assign n38491 = n34266 ^ n27034 ^ 1'b0 ;
  assign n38492 = n38490 & ~n38491 ;
  assign n38493 = n38487 & n38492 ;
  assign n38494 = n33435 ^ n16859 ^ n8813 ;
  assign n38495 = n14914 | n33953 ;
  assign n38496 = n8209 ^ n4799 ^ n3315 ;
  assign n38497 = ~n2354 & n18171 ;
  assign n38498 = ~n33272 & n38497 ;
  assign n38499 = n15119 & ~n38393 ;
  assign n38500 = ~n21799 & n38499 ;
  assign n38501 = n38500 ^ n27482 ^ 1'b0 ;
  assign n38506 = ( n3169 & ~n10032 ) | ( n3169 & n27527 ) | ( ~n10032 & n27527 ) ;
  assign n38507 = ~n19191 & n38506 ;
  assign n38502 = ~n6424 & n10453 ;
  assign n38503 = ~n6624 & n38502 ;
  assign n38504 = n7841 | n27032 ;
  assign n38505 = n38503 & ~n38504 ;
  assign n38508 = n38507 ^ n38505 ^ 1'b0 ;
  assign n38509 = n13426 ^ n7664 ^ 1'b0 ;
  assign n38510 = n21593 | n38509 ;
  assign n38511 = n6513 | n24845 ;
  assign n38512 = n15992 ^ n1191 ^ 1'b0 ;
  assign n38513 = ~n5400 & n11718 ;
  assign n38514 = n32462 ^ n13024 ^ n304 ;
  assign n38515 = n6100 & n17430 ;
  assign n38516 = n13992 ^ n4911 ^ 1'b0 ;
  assign n38517 = n37574 & ~n38408 ;
  assign n38518 = n6565 | n26099 ;
  assign n38519 = n14957 & n28586 ;
  assign n38520 = ( ~n4458 & n30172 ) | ( ~n4458 & n38519 ) | ( n30172 & n38519 ) ;
  assign n38521 = n2953 | n19276 ;
  assign n38522 = n731 | n9324 ;
  assign n38523 = n38521 & ~n38522 ;
  assign n38524 = n32292 ^ n9971 ^ 1'b0 ;
  assign n38525 = n7599 & ~n38227 ;
  assign n38526 = ~x70 & n38525 ;
  assign n38527 = ~n8487 & n19134 ;
  assign n38528 = n38527 ^ n9506 ^ 1'b0 ;
  assign n38529 = n531 | n14957 ;
  assign n38530 = ~n19186 & n23677 ;
  assign n38531 = n38530 ^ n8748 ^ 1'b0 ;
  assign n38532 = n28552 | n38531 ;
  assign n38533 = n38532 ^ n25298 ^ 1'b0 ;
  assign n38534 = n38533 ^ n1779 ^ 1'b0 ;
  assign n38535 = n38534 ^ n23316 ^ n14668 ;
  assign n38536 = n16836 ^ n9912 ^ x200 ;
  assign n38537 = n38536 ^ n32398 ^ 1'b0 ;
  assign n38538 = n31643 ^ n25358 ^ n10713 ;
  assign n38539 = n4287 & ~n38538 ;
  assign n38540 = ~n1370 & n4359 ;
  assign n38541 = n38540 ^ n30866 ^ 1'b0 ;
  assign n38542 = n11937 | n23949 ;
  assign n38543 = n2380 | n6647 ;
  assign n38544 = n38543 ^ n25327 ^ 1'b0 ;
  assign n38545 = n1234 & ~n37481 ;
  assign n38546 = n24937 ^ n6795 ^ 1'b0 ;
  assign n38547 = ~n11597 & n38546 ;
  assign n38548 = n38547 ^ n35168 ^ 1'b0 ;
  assign n38549 = n21290 & ~n36115 ;
  assign n38550 = ~n21036 & n38549 ;
  assign n38551 = ~n9610 & n34670 ;
  assign n38553 = ~n7254 & n10455 ;
  assign n38552 = n19514 | n34618 ;
  assign n38554 = n38553 ^ n38552 ^ 1'b0 ;
  assign n38555 = n17170 ^ n8961 ^ 1'b0 ;
  assign n38556 = n681 & ~n8866 ;
  assign n38558 = ~n2262 & n4806 ;
  assign n38559 = n38558 ^ n9964 ^ 1'b0 ;
  assign n38557 = n677 | n17994 ;
  assign n38560 = n38559 ^ n38557 ^ 1'b0 ;
  assign n38561 = n20101 & n36703 ;
  assign n38562 = ~n28249 & n31528 ;
  assign n38563 = n38562 ^ n4721 ^ 1'b0 ;
  assign n38564 = n5051 & ~n19722 ;
  assign n38565 = n38564 ^ n10154 ^ 1'b0 ;
  assign n38566 = n4374 & ~n5680 ;
  assign n38567 = n12310 ^ n10303 ^ 1'b0 ;
  assign n38568 = ( ~n38565 & n38566 ) | ( ~n38565 & n38567 ) | ( n38566 & n38567 ) ;
  assign n38569 = n2067 | n12302 ;
  assign n38570 = n38569 ^ n23902 ^ 1'b0 ;
  assign n38571 = ( n15357 & n16939 ) | ( n15357 & n38570 ) | ( n16939 & n38570 ) ;
  assign n38572 = n7739 ^ n5558 ^ n4823 ;
  assign n38573 = n24058 & n38572 ;
  assign n38574 = n28431 & n31934 ;
  assign n38575 = n38574 ^ n23161 ^ 1'b0 ;
  assign n38576 = ( n1459 & ~n7015 ) | ( n1459 & n14615 ) | ( ~n7015 & n14615 ) ;
  assign n38577 = n10036 & n38576 ;
  assign n38578 = n1044 & n4468 ;
  assign n38579 = n38578 ^ n14106 ^ 1'b0 ;
  assign n38580 = n19893 & n38579 ;
  assign n38581 = ~n5350 & n13740 ;
  assign n38582 = n38581 ^ n27144 ^ 1'b0 ;
  assign n38583 = ( n7917 & n30257 ) | ( n7917 & n38582 ) | ( n30257 & n38582 ) ;
  assign n38584 = n15383 ^ n9807 ^ 1'b0 ;
  assign n38585 = ( n25473 & ~n28982 ) | ( n25473 & n38584 ) | ( ~n28982 & n38584 ) ;
  assign n38586 = n19664 ^ n18096 ^ n6730 ;
  assign n38587 = ~n1192 & n29413 ;
  assign n38588 = n15542 | n17263 ;
  assign n38589 = n27388 ^ n21593 ^ 1'b0 ;
  assign n38590 = n27253 | n38589 ;
  assign n38591 = n11631 ^ n593 ^ 1'b0 ;
  assign n38592 = ~n4752 & n38591 ;
  assign n38593 = n38592 ^ n28678 ^ n17568 ;
  assign n38594 = n9212 & ~n38593 ;
  assign n38595 = n12008 & n30538 ;
  assign n38596 = n3061 & ~n16181 ;
  assign n38597 = n1797 & n38596 ;
  assign n38598 = n22696 ^ n20870 ^ 1'b0 ;
  assign n38599 = n6704 & ~n19778 ;
  assign n38600 = ( n15281 & n38598 ) | ( n15281 & ~n38599 ) | ( n38598 & ~n38599 ) ;
  assign n38601 = ~n5531 & n23946 ;
  assign n38602 = n38423 ^ n22595 ^ 1'b0 ;
  assign n38603 = ~n29042 & n38602 ;
  assign n38604 = n24006 ^ n4984 ^ 1'b0 ;
  assign n38607 = n2359 & ~n18296 ;
  assign n38605 = n13985 & n25908 ;
  assign n38606 = n38605 ^ n24114 ^ 1'b0 ;
  assign n38608 = n38607 ^ n38606 ^ n24931 ;
  assign n38609 = n1297 ^ x49 ^ 1'b0 ;
  assign n38610 = n24436 | n38609 ;
  assign n38611 = n36469 ^ n3460 ^ 1'b0 ;
  assign n38613 = n3568 & ~n12546 ;
  assign n38614 = n10867 & ~n38613 ;
  assign n38615 = n38614 ^ n6401 ^ 1'b0 ;
  assign n38612 = n24263 | n37330 ;
  assign n38616 = n38615 ^ n38612 ^ n33988 ;
  assign n38617 = n14510 | n34527 ;
  assign n38618 = ( n1188 & n27144 ) | ( n1188 & ~n38617 ) | ( n27144 & ~n38617 ) ;
  assign n38619 = n29330 ^ n3927 ^ 1'b0 ;
  assign n38620 = n28311 & n29159 ;
  assign n38621 = n38620 ^ n12057 ^ 1'b0 ;
  assign n38622 = n33623 ^ n17267 ^ 1'b0 ;
  assign n38623 = n35968 ^ n25260 ^ 1'b0 ;
  assign n38624 = n30755 | n38623 ;
  assign n38625 = n4242 & ~n10036 ;
  assign n38626 = n38625 ^ n19722 ^ 1'b0 ;
  assign n38627 = n10292 & ~n14639 ;
  assign n38628 = n38627 ^ n19506 ^ n9793 ;
  assign n38629 = n38626 & ~n38628 ;
  assign n38630 = ~n5277 & n8336 ;
  assign n38631 = ~n38629 & n38630 ;
  assign n38632 = n17373 & n30253 ;
  assign n38633 = n9093 & n38632 ;
  assign n38634 = ~n18670 & n22042 ;
  assign n38635 = n12302 & n38634 ;
  assign n38636 = n29522 | n38635 ;
  assign n38637 = n38636 ^ n6998 ^ 1'b0 ;
  assign n38638 = n20563 & n29812 ;
  assign n38639 = n24793 ^ n18851 ^ 1'b0 ;
  assign n38640 = n24352 ^ n4481 ^ 1'b0 ;
  assign n38641 = ~n4959 & n38640 ;
  assign n38642 = n7645 & n35652 ;
  assign n38643 = n7273 ^ n4556 ^ 1'b0 ;
  assign n38644 = n25748 & ~n38643 ;
  assign n38645 = n27874 & n38644 ;
  assign n38646 = ~n29202 & n38645 ;
  assign n38647 = n17192 & ~n27423 ;
  assign n38648 = n15290 & n38647 ;
  assign n38649 = n9287 | n15464 ;
  assign n38650 = n3540 | n38649 ;
  assign n38651 = n38650 ^ n22009 ^ n6303 ;
  assign n38653 = ~n11838 & n38383 ;
  assign n38654 = n38653 ^ n6681 ^ 1'b0 ;
  assign n38652 = n14010 ^ n10088 ^ 1'b0 ;
  assign n38655 = n38654 ^ n38652 ^ n4470 ;
  assign n38656 = n19821 ^ n4474 ^ 1'b0 ;
  assign n38657 = ~n29689 & n38656 ;
  assign n38658 = ( ~n6128 & n29914 ) | ( ~n6128 & n38657 ) | ( n29914 & n38657 ) ;
  assign n38659 = n8899 ^ n3068 ^ 1'b0 ;
  assign n38660 = n16560 ^ n8850 ^ 1'b0 ;
  assign n38661 = ~n16958 & n38660 ;
  assign n38662 = ( n27970 & n38659 ) | ( n27970 & ~n38661 ) | ( n38659 & ~n38661 ) ;
  assign n38663 = n38662 ^ n28741 ^ 1'b0 ;
  assign n38664 = n19992 & ~n35410 ;
  assign n38665 = ~n13955 & n14644 ;
  assign n38666 = n38665 ^ n16948 ^ 1'b0 ;
  assign n38667 = n6936 & ~n18933 ;
  assign n38668 = n38667 ^ n4468 ^ 1'b0 ;
  assign n38674 = n16098 ^ n13925 ^ n5624 ;
  assign n38671 = n821 & n1550 ;
  assign n38672 = ~n18409 & n38671 ;
  assign n38673 = n38672 ^ n17694 ^ 1'b0 ;
  assign n38669 = n33307 ^ n21087 ^ 1'b0 ;
  assign n38670 = n21082 & n38669 ;
  assign n38675 = n38674 ^ n38673 ^ n38670 ;
  assign n38676 = n13570 ^ n9961 ^ 1'b0 ;
  assign n38677 = n17143 ^ n14320 ^ 1'b0 ;
  assign n38678 = n1767 & n11503 ;
  assign n38679 = n11153 & ~n38678 ;
  assign n38680 = n38679 ^ n4535 ^ 1'b0 ;
  assign n38681 = ~n5048 & n18529 ;
  assign n38682 = n26377 ^ n456 ^ 1'b0 ;
  assign n38683 = n11930 ^ n1929 ^ 1'b0 ;
  assign n38684 = n14766 | n38683 ;
  assign n38685 = n38684 ^ n37704 ^ n18387 ;
  assign n38686 = ~n13048 & n38685 ;
  assign n38687 = n8562 & n38686 ;
  assign n38688 = n11344 ^ n4390 ^ 1'b0 ;
  assign n38689 = n10873 | n17784 ;
  assign n38690 = n27111 | n38689 ;
  assign n38691 = ~n9099 & n20941 ;
  assign n38692 = n5244 ^ n471 ^ 1'b0 ;
  assign n38693 = n23513 & ~n38692 ;
  assign n38694 = n38693 ^ n6332 ^ 1'b0 ;
  assign n38695 = n12611 & ~n37404 ;
  assign n38696 = n2715 & n29428 ;
  assign n38697 = n1332 | n38696 ;
  assign n38698 = n38697 ^ n14481 ^ 1'b0 ;
  assign n38699 = ~n38695 & n38698 ;
  assign n38700 = n2843 & n29604 ;
  assign n38701 = n12724 & n18967 ;
  assign n38702 = ( n15415 & ~n38700 ) | ( n15415 & n38701 ) | ( ~n38700 & n38701 ) ;
  assign n38703 = n2144 | n19244 ;
  assign n38704 = n31370 & ~n38703 ;
  assign n38705 = n4491 & ~n38704 ;
  assign n38706 = ~n3132 & n33287 ;
  assign n38707 = n4487 ^ n2108 ^ 1'b0 ;
  assign n38708 = n33886 | n38707 ;
  assign n38709 = n5122 ^ n1626 ^ 1'b0 ;
  assign n38710 = n38708 | n38709 ;
  assign n38711 = n24531 ^ n20736 ^ 1'b0 ;
  assign n38712 = ~n20952 & n38711 ;
  assign n38713 = n38710 | n38712 ;
  assign n38714 = n20809 | n24500 ;
  assign n38715 = ~n22444 & n28788 ;
  assign n38716 = n22754 ^ n9025 ^ 1'b0 ;
  assign n38717 = n8933 ^ n5518 ^ 1'b0 ;
  assign n38718 = n3032 & ~n4954 ;
  assign n38719 = n5014 | n6122 ;
  assign n38720 = n8018 & ~n17218 ;
  assign n38721 = n29720 ^ n28257 ^ 1'b0 ;
  assign n38722 = n38721 ^ n10146 ^ 1'b0 ;
  assign n38723 = n30703 & n38722 ;
  assign n38724 = n6975 ^ n3617 ^ 1'b0 ;
  assign n38725 = n18874 & ~n20529 ;
  assign n38726 = n4089 & n38725 ;
  assign n38727 = n38726 ^ n27253 ^ 1'b0 ;
  assign n38728 = n1969 & n38727 ;
  assign n38729 = ( ~n18622 & n38724 ) | ( ~n18622 & n38728 ) | ( n38724 & n38728 ) ;
  assign n38730 = n25069 ^ n4925 ^ 1'b0 ;
  assign n38731 = n28838 ^ n11193 ^ 1'b0 ;
  assign n38732 = n16330 & ~n29649 ;
  assign n38733 = n16521 & ~n29344 ;
  assign n38734 = ~n17178 & n25071 ;
  assign n38735 = ~n29153 & n38734 ;
  assign n38736 = ~n1038 & n11067 ;
  assign n38737 = n30663 & n38736 ;
  assign n38738 = n2489 & ~n38737 ;
  assign n38739 = ~n3126 & n38738 ;
  assign n38740 = n5837 & ~n10636 ;
  assign n38741 = n38740 ^ n3059 ^ 1'b0 ;
  assign n38742 = ~n5433 & n38741 ;
  assign n38743 = ~n29577 & n38742 ;
  assign n38744 = n9023 & ~n38743 ;
  assign n38745 = n38744 ^ n1803 ^ 1'b0 ;
  assign n38746 = n11285 & n22800 ;
  assign n38747 = n28854 ^ n13733 ^ 1'b0 ;
  assign n38748 = n37173 & ~n38747 ;
  assign n38749 = ( n1630 & n13756 ) | ( n1630 & ~n14139 ) | ( n13756 & ~n14139 ) ;
  assign n38750 = ( n5805 & n20553 ) | ( n5805 & ~n38749 ) | ( n20553 & ~n38749 ) ;
  assign n38751 = n13004 | n21354 ;
  assign n38752 = n20314 & ~n38751 ;
  assign n38753 = ( n11932 & ~n23337 ) | ( n11932 & n38752 ) | ( ~n23337 & n38752 ) ;
  assign n38754 = n37876 ^ x40 ^ 1'b0 ;
  assign n38755 = ~n6605 & n34881 ;
  assign n38756 = ~n9309 & n38755 ;
  assign n38757 = n21055 ^ n7317 ^ 1'b0 ;
  assign n38758 = n7017 | n19285 ;
  assign n38759 = n38758 ^ n22499 ^ 1'b0 ;
  assign n38760 = ~n23511 & n38759 ;
  assign n38761 = n23471 & n38760 ;
  assign n38762 = n38761 ^ n2692 ^ 1'b0 ;
  assign n38763 = n24919 ^ n18213 ^ 1'b0 ;
  assign n38764 = n14978 | n38763 ;
  assign n38765 = n38764 ^ n22696 ^ n22465 ;
  assign n38766 = ( n1475 & ~n6656 ) | ( n1475 & n10237 ) | ( ~n6656 & n10237 ) ;
  assign n38767 = n12474 ^ n8330 ^ 1'b0 ;
  assign n38768 = ~n2005 & n38767 ;
  assign n38769 = ~n15418 & n38768 ;
  assign n38770 = n3369 ^ n1164 ^ 1'b0 ;
  assign n38771 = ~n22064 & n38770 ;
  assign n38772 = n25143 ^ n9231 ^ 1'b0 ;
  assign n38773 = ~n8938 & n26140 ;
  assign n38774 = n6001 & n10366 ;
  assign n38775 = ~n7466 & n38774 ;
  assign n38776 = n12433 & n38775 ;
  assign n38777 = n11377 | n38776 ;
  assign n38778 = n4518 | n18508 ;
  assign n38779 = n3883 | n38778 ;
  assign n38780 = n1314 & n4047 ;
  assign n38781 = n38780 ^ n16534 ^ 1'b0 ;
  assign n38782 = n2537 & ~n16484 ;
  assign n38783 = n38782 ^ n24158 ^ n519 ;
  assign n38784 = n21105 & ~n21132 ;
  assign n38785 = n38784 ^ n14833 ^ 1'b0 ;
  assign n38786 = n7723 & ~n29041 ;
  assign n38787 = n38785 & n38786 ;
  assign n38788 = n38783 & n38787 ;
  assign n38789 = n24833 & n33698 ;
  assign n38790 = n38789 ^ n29135 ^ 1'b0 ;
  assign n38791 = n11067 ^ n8022 ^ 1'b0 ;
  assign n38792 = n38790 & n38791 ;
  assign n38793 = n17548 | n30531 ;
  assign n38794 = n20345 ^ n9652 ^ n5223 ;
  assign n38795 = ~n13197 & n38794 ;
  assign n38796 = ~n38793 & n38795 ;
  assign n38797 = n19050 ^ n9088 ^ 1'b0 ;
  assign n38800 = ( n6597 & n9453 ) | ( n6597 & ~n18876 ) | ( n9453 & ~n18876 ) ;
  assign n38798 = n7316 ^ n5006 ^ 1'b0 ;
  assign n38799 = ~n4267 & n38798 ;
  assign n38801 = n38800 ^ n38799 ^ n19239 ;
  assign n38802 = n822 | n2106 ;
  assign n38803 = n36090 | n38802 ;
  assign n38804 = n27948 ^ n24271 ^ 1'b0 ;
  assign n38805 = n17369 & ~n38804 ;
  assign n38806 = ~n4762 & n5824 ;
  assign n38807 = ( n20166 & n28296 ) | ( n20166 & n38806 ) | ( n28296 & n38806 ) ;
  assign n38808 = n31432 ^ n2686 ^ 1'b0 ;
  assign n38809 = n14930 & ~n18367 ;
  assign n38810 = n18313 ^ n14991 ^ 1'b0 ;
  assign n38811 = n38810 ^ n31336 ^ 1'b0 ;
  assign n38812 = ~n9342 & n34374 ;
  assign n38813 = n38812 ^ n29698 ^ 1'b0 ;
  assign n38814 = n7138 & ~n8093 ;
  assign n38815 = n2689 & ~n33223 ;
  assign n38816 = n38815 ^ n33574 ^ 1'b0 ;
  assign n38817 = ~n13932 & n38816 ;
  assign n38818 = n460 & n38817 ;
  assign n38819 = n10939 & ~n37229 ;
  assign n38820 = n29616 ^ n8001 ^ n1702 ;
  assign n38821 = n38820 ^ n18415 ^ 1'b0 ;
  assign n38822 = n24479 ^ n7756 ^ 1'b0 ;
  assign n38823 = n8066 ^ n3481 ^ 1'b0 ;
  assign n38824 = ( n22567 & ~n38822 ) | ( n22567 & n38823 ) | ( ~n38822 & n38823 ) ;
  assign n38825 = n873 | n2307 ;
  assign n38826 = n13990 | n38825 ;
  assign n38827 = n35707 | n37124 ;
  assign n38828 = n24457 ^ n3362 ^ n3328 ;
  assign n38829 = n38828 ^ n10117 ^ 1'b0 ;
  assign n38830 = n24765 | n38829 ;
  assign n38831 = n11281 & ~n37312 ;
  assign n38832 = n38831 ^ n9440 ^ 1'b0 ;
  assign n38833 = n38832 ^ n16416 ^ x45 ;
  assign n38834 = n890 & n38833 ;
  assign n38835 = ~n18121 & n19181 ;
  assign n38836 = n38834 & n38835 ;
  assign n38837 = n8531 ^ n2363 ^ 1'b0 ;
  assign n38838 = n38837 ^ n2819 ^ 1'b0 ;
  assign n38839 = n12877 & ~n30798 ;
  assign n38840 = n13386 | n15130 ;
  assign n38841 = n30026 | n38840 ;
  assign n38843 = n27575 ^ n26593 ^ n23814 ;
  assign n38844 = n2232 | n14151 ;
  assign n38845 = n38843 | n38844 ;
  assign n38842 = ~n1339 & n28529 ;
  assign n38846 = n38845 ^ n38842 ^ 1'b0 ;
  assign n38847 = n2739 | n8449 ;
  assign n38848 = n38847 ^ n10176 ^ 1'b0 ;
  assign n38849 = ( n18805 & ~n22610 ) | ( n18805 & n38848 ) | ( ~n22610 & n38848 ) ;
  assign n38850 = n33493 | n38849 ;
  assign n38851 = n38846 | n38850 ;
  assign n38852 = n32010 ^ n1665 ^ 1'b0 ;
  assign n38853 = n21949 | n38852 ;
  assign n38854 = n6747 | n38853 ;
  assign n38855 = n11718 & ~n38854 ;
  assign n38856 = n35139 & n38855 ;
  assign n38857 = n10881 | n10907 ;
  assign n38858 = n2847 | n19470 ;
  assign n38859 = ( ~n14994 & n26937 ) | ( ~n14994 & n38858 ) | ( n26937 & n38858 ) ;
  assign n38860 = ~n6801 & n25082 ;
  assign n38861 = n38860 ^ n31559 ^ 1'b0 ;
  assign n38862 = n34721 ^ n34037 ^ n3149 ;
  assign n38863 = n38862 ^ n13215 ^ 1'b0 ;
  assign n38864 = ( n5731 & n18725 ) | ( n5731 & n27485 ) | ( n18725 & n27485 ) ;
  assign n38865 = n38864 ^ n18015 ^ 1'b0 ;
  assign n38866 = n24144 & n38865 ;
  assign n38871 = n2887 | n10186 ;
  assign n38867 = n11703 ^ n513 ^ 1'b0 ;
  assign n38868 = ( n5315 & n20137 ) | ( n5315 & ~n38867 ) | ( n20137 & ~n38867 ) ;
  assign n38869 = n13264 & n38868 ;
  assign n38870 = n8855 & n38869 ;
  assign n38872 = n38871 ^ n38870 ^ 1'b0 ;
  assign n38873 = n16718 & n24176 ;
  assign n38874 = ( n3588 & n10600 ) | ( n3588 & ~n38873 ) | ( n10600 & ~n38873 ) ;
  assign n38875 = n22605 ^ n3318 ^ x206 ;
  assign n38876 = n38875 ^ n24329 ^ n288 ;
  assign n38877 = ~x203 & n19260 ;
  assign n38878 = ~n21424 & n38877 ;
  assign n38879 = n38878 ^ n6755 ^ 1'b0 ;
  assign n38880 = n38879 ^ n5791 ^ 1'b0 ;
  assign n38881 = ~n13469 & n14816 ;
  assign n38882 = n10459 & n38881 ;
  assign n38883 = n38882 ^ n20755 ^ 1'b0 ;
  assign n38886 = n31855 ^ n13281 ^ 1'b0 ;
  assign n38884 = n13609 ^ n4895 ^ 1'b0 ;
  assign n38885 = n27051 & ~n38884 ;
  assign n38887 = n38886 ^ n38885 ^ 1'b0 ;
  assign n38888 = n5780 | n13900 ;
  assign n38889 = n12885 & ~n38888 ;
  assign n38890 = n23822 | n27639 ;
  assign n38891 = n33430 ^ n21540 ^ n10657 ;
  assign n38892 = n7585 & n29741 ;
  assign n38893 = n38892 ^ n26961 ^ n8742 ;
  assign n38894 = n38893 ^ n11956 ^ 1'b0 ;
  assign n38895 = ~n22068 & n38894 ;
  assign n38896 = n8691 | n11088 ;
  assign n38897 = n15383 | n26293 ;
  assign n38898 = n7839 | n12394 ;
  assign n38899 = ( n38896 & n38897 ) | ( n38896 & ~n38898 ) | ( n38897 & ~n38898 ) ;
  assign n38900 = ( n24329 & n38895 ) | ( n24329 & ~n38899 ) | ( n38895 & ~n38899 ) ;
  assign n38902 = n2179 | n27970 ;
  assign n38903 = ~n3884 & n18194 ;
  assign n38904 = ~n38902 & n38903 ;
  assign n38901 = n4398 & n31936 ;
  assign n38905 = n38904 ^ n38901 ^ 1'b0 ;
  assign n38906 = n4534 ^ n2437 ^ 1'b0 ;
  assign n38907 = n27207 | n38906 ;
  assign n38908 = n579 & n28165 ;
  assign n38909 = ~n26197 & n38908 ;
  assign n38910 = n11656 | n17486 ;
  assign n38913 = n14746 ^ n3029 ^ 1'b0 ;
  assign n38912 = n5461 | n27384 ;
  assign n38914 = n38913 ^ n38912 ^ 1'b0 ;
  assign n38911 = n10338 ^ n9526 ^ n6656 ;
  assign n38915 = n38914 ^ n38911 ^ n11069 ;
  assign n38916 = x144 | n451 ;
  assign n38917 = n38916 ^ n15028 ^ n8171 ;
  assign n38918 = ( ~n9895 & n13566 ) | ( ~n9895 & n26245 ) | ( n13566 & n26245 ) ;
  assign n38919 = n38917 & ~n38918 ;
  assign n38920 = n38915 & n38919 ;
  assign n38921 = ~n557 & n38917 ;
  assign n38922 = ( n1930 & ~n3554 ) | ( n1930 & n3617 ) | ( ~n3554 & n3617 ) ;
  assign n38923 = n38922 ^ n15465 ^ 1'b0 ;
  assign n38924 = ~n8664 & n38923 ;
  assign n38925 = n704 | n1323 ;
  assign n38926 = n38925 ^ n12025 ^ 1'b0 ;
  assign n38927 = n33055 | n38926 ;
  assign n38928 = n38927 ^ n21313 ^ 1'b0 ;
  assign n38929 = n12241 ^ n8044 ^ 1'b0 ;
  assign n38930 = ~n16004 & n21483 ;
  assign n38931 = n21687 ^ n14403 ^ n1421 ;
  assign n38932 = ~n1396 & n38931 ;
  assign n38933 = n38930 & n38932 ;
  assign n38934 = n6331 ^ n629 ^ 1'b0 ;
  assign n38935 = n38934 ^ n11372 ^ 1'b0 ;
  assign n38936 = n12959 & ~n38935 ;
  assign n38937 = n38936 ^ n30245 ^ 1'b0 ;
  assign n38938 = n15104 & ~n38937 ;
  assign n38940 = n3545 & n20455 ;
  assign n38941 = n38940 ^ n14693 ^ 1'b0 ;
  assign n38942 = ~n38461 & n38941 ;
  assign n38939 = ~n2134 & n37288 ;
  assign n38943 = n38942 ^ n38939 ^ 1'b0 ;
  assign n38944 = n11726 & ~n32981 ;
  assign n38945 = n27282 ^ n16261 ^ n15908 ;
  assign n38946 = n1377 ^ n790 ^ 1'b0 ;
  assign n38947 = ~n1715 & n16684 ;
  assign n38948 = n3027 & n38947 ;
  assign n38949 = n38946 | n38948 ;
  assign n38950 = ~n8911 & n19050 ;
  assign n38951 = n38950 ^ n8815 ^ 1'b0 ;
  assign n38952 = n17013 & n24942 ;
  assign n38953 = x162 & n1182 ;
  assign n38954 = ~x162 & n38953 ;
  assign n38955 = n790 & ~n38954 ;
  assign n38956 = n38955 ^ n3272 ^ 1'b0 ;
  assign n38957 = ~n16539 & n38956 ;
  assign n38958 = n11361 & n38957 ;
  assign n38959 = n38958 ^ n16075 ^ 1'b0 ;
  assign n38960 = n10043 & ~n13606 ;
  assign n38961 = ~n38959 & n38960 ;
  assign n38962 = n16838 | n38897 ;
  assign n38963 = n38961 & ~n38962 ;
  assign n38964 = ~n3082 & n6290 ;
  assign n38966 = n7693 | n13198 ;
  assign n38967 = n38966 ^ n16902 ^ 1'b0 ;
  assign n38965 = n11628 & n33807 ;
  assign n38968 = n38967 ^ n38965 ^ 1'b0 ;
  assign n38969 = ~n38964 & n38968 ;
  assign n38970 = n38969 ^ n27684 ^ n13563 ;
  assign n38971 = n17052 ^ n10267 ^ 1'b0 ;
  assign n38972 = ( n3702 & n18528 ) | ( n3702 & n36283 ) | ( n18528 & n36283 ) ;
  assign n38973 = n9356 | n13328 ;
  assign n38974 = n26252 | n38973 ;
  assign n38975 = n13447 & ~n27661 ;
  assign n38976 = n1506 & ~n27943 ;
  assign n38977 = n38976 ^ n5306 ^ 1'b0 ;
  assign n38978 = n38977 ^ n10715 ^ 1'b0 ;
  assign n38981 = n3414 & n3776 ;
  assign n38982 = n31361 & n38981 ;
  assign n38979 = n30258 ^ n2564 ^ 1'b0 ;
  assign n38980 = n25203 | n38979 ;
  assign n38983 = n38982 ^ n38980 ^ 1'b0 ;
  assign n38984 = x15 | n10182 ;
  assign n38985 = n11960 | n38984 ;
  assign n38986 = ~n13391 & n38985 ;
  assign n38987 = ~n20233 & n27846 ;
  assign n38988 = ~n4124 & n38987 ;
  assign n38989 = n2548 ^ n570 ^ 1'b0 ;
  assign n38990 = n5311 | n38989 ;
  assign n38991 = n29038 & ~n38990 ;
  assign n38992 = n9110 & n38991 ;
  assign n38993 = n388 & ~n1806 ;
  assign n38994 = n38993 ^ n16181 ^ 1'b0 ;
  assign n38995 = n2754 & ~n38994 ;
  assign n38996 = ( ~n9849 & n11357 ) | ( ~n9849 & n38995 ) | ( n11357 & n38995 ) ;
  assign n38997 = n36012 ^ n32849 ^ n2958 ;
  assign n38998 = n22671 ^ n2821 ^ 1'b0 ;
  assign n38999 = n5464 & n38998 ;
  assign n39000 = ~n4907 & n31840 ;
  assign n39001 = n38999 & n39000 ;
  assign n39002 = n39001 ^ n30084 ^ 1'b0 ;
  assign n39003 = n2824 & n14795 ;
  assign n39004 = n7106 ^ n3829 ^ 1'b0 ;
  assign n39005 = n15227 & n39004 ;
  assign n39006 = n27684 ^ n19746 ^ 1'b0 ;
  assign n39007 = n15186 & ~n18188 ;
  assign n39008 = ~n13885 & n38170 ;
  assign n39009 = ( n1029 & n15583 ) | ( n1029 & ~n24904 ) | ( n15583 & ~n24904 ) ;
  assign n39010 = n39009 ^ n38085 ^ n35995 ;
  assign n39011 = n9793 & ~n22894 ;
  assign n39012 = n39011 ^ n18848 ^ 1'b0 ;
  assign n39015 = n17129 ^ n14177 ^ 1'b0 ;
  assign n39016 = n22861 & ~n39015 ;
  assign n39013 = n20161 & n22611 ;
  assign n39014 = n19021 | n39013 ;
  assign n39017 = n39016 ^ n39014 ^ 1'b0 ;
  assign n39018 = n24460 ^ n4900 ^ 1'b0 ;
  assign n39019 = ~n12353 & n39018 ;
  assign n39020 = n12937 | n13211 ;
  assign n39021 = n39020 ^ n301 ^ 1'b0 ;
  assign n39022 = n39019 | n39021 ;
  assign n39023 = n39022 ^ n14417 ^ 1'b0 ;
  assign n39024 = n6540 | n39023 ;
  assign n39025 = ~n6980 & n14120 ;
  assign n39026 = n27494 ^ n21664 ^ 1'b0 ;
  assign n39027 = n11443 | n39026 ;
  assign n39028 = n39025 & n39027 ;
  assign n39029 = n34901 ^ n12923 ^ n4249 ;
  assign n39030 = ( n836 & n2002 ) | ( n836 & n6363 ) | ( n2002 & n6363 ) ;
  assign n39031 = n15229 | n39030 ;
  assign n39032 = n28169 & n39031 ;
  assign n39033 = ( n8851 & n23133 ) | ( n8851 & ~n39032 ) | ( n23133 & ~n39032 ) ;
  assign n39034 = ~n16587 & n26770 ;
  assign n39035 = n28562 ^ n24001 ^ 1'b0 ;
  assign n39036 = n10746 & n39035 ;
  assign n39037 = n39036 ^ n9002 ^ 1'b0 ;
  assign n39038 = n31312 | n39037 ;
  assign n39039 = n32900 | n36943 ;
  assign n39040 = ( ~n1843 & n6285 ) | ( ~n1843 & n31120 ) | ( n6285 & n31120 ) ;
  assign n39041 = n37433 ^ n11425 ^ 1'b0 ;
  assign n39042 = n39040 | n39041 ;
  assign n39043 = n5534 | n13563 ;
  assign n39044 = n14401 ^ n8740 ^ 1'b0 ;
  assign n39045 = ~n32197 & n39044 ;
  assign n39046 = n32527 ^ n11646 ^ 1'b0 ;
  assign n39047 = n36652 ^ n34664 ^ 1'b0 ;
  assign n39048 = n13119 ^ n10464 ^ 1'b0 ;
  assign n39049 = ~n8148 & n12906 ;
  assign n39050 = n39049 ^ n16754 ^ 1'b0 ;
  assign n39051 = ~n16857 & n39050 ;
  assign n39052 = ( n6715 & ~n7897 ) | ( n6715 & n36709 ) | ( ~n7897 & n36709 ) ;
  assign n39053 = ( ~n10194 & n31097 ) | ( ~n10194 & n39052 ) | ( n31097 & n39052 ) ;
  assign n39054 = n17352 ^ n6223 ^ n4293 ;
  assign n39055 = ~n15051 & n39054 ;
  assign n39056 = ~n39053 & n39055 ;
  assign n39057 = n27649 & ~n39056 ;
  assign n39058 = ~n30474 & n39057 ;
  assign n39059 = n5304 & n23209 ;
  assign n39060 = n8255 & ~n39059 ;
  assign n39061 = n8113 & n29928 ;
  assign n39062 = x209 & ~n4614 ;
  assign n39063 = n39062 ^ n28076 ^ n4628 ;
  assign n39064 = n39063 ^ n32314 ^ n29692 ;
  assign n39065 = n13536 & ~n24858 ;
  assign n39066 = ~n6704 & n39065 ;
  assign n39067 = n22542 ^ n7135 ^ 1'b0 ;
  assign n39068 = ~n2648 & n39067 ;
  assign n39069 = n39068 ^ n18455 ^ 1'b0 ;
  assign n39070 = n32112 & ~n39069 ;
  assign n39071 = n39066 & n39070 ;
  assign n39072 = ~n22046 & n27581 ;
  assign n39073 = ~n18776 & n39072 ;
  assign n39074 = n10298 | n39073 ;
  assign n39075 = n36398 & ~n39074 ;
  assign n39076 = n491 | n7237 ;
  assign n39077 = ~n20548 & n39076 ;
  assign n39078 = ( n2207 & ~n10186 ) | ( n2207 & n17949 ) | ( ~n10186 & n17949 ) ;
  assign n39079 = n9056 ^ n7603 ^ 1'b0 ;
  assign n39080 = n4555 ^ n2670 ^ n1953 ;
  assign n39081 = n38721 ^ n6284 ^ 1'b0 ;
  assign n39082 = ~n22978 & n39081 ;
  assign n39083 = n39082 ^ n30267 ^ 1'b0 ;
  assign n39084 = n31290 ^ n26207 ^ n14119 ;
  assign n39085 = n4303 & n39084 ;
  assign n39086 = n836 & ~n4529 ;
  assign n39087 = n39086 ^ n13735 ^ 1'b0 ;
  assign n39088 = n8902 | n16311 ;
  assign n39089 = n39088 ^ n30282 ^ 1'b0 ;
  assign n39090 = n7559 ^ n770 ^ n671 ;
  assign n39091 = n18451 ^ n3773 ^ 1'b0 ;
  assign n39092 = ( n4514 & ~n11665 ) | ( n4514 & n39091 ) | ( ~n11665 & n39091 ) ;
  assign n39093 = n27032 | n39092 ;
  assign n39094 = n39093 ^ n33032 ^ 1'b0 ;
  assign n39095 = n35345 ^ n27738 ^ 1'b0 ;
  assign n39096 = n20845 & ~n33440 ;
  assign n39097 = ~n33822 & n39096 ;
  assign n39098 = ~n5758 & n39097 ;
  assign n39099 = n4189 | n26320 ;
  assign n39100 = n39099 ^ n8780 ^ 1'b0 ;
  assign n39101 = n36915 & n39100 ;
  assign n39102 = ( n8858 & n13232 ) | ( n8858 & n28067 ) | ( n13232 & n28067 ) ;
  assign n39103 = n19157 ^ n7507 ^ 1'b0 ;
  assign n39104 = n8661 & n17968 ;
  assign n39105 = ~n39103 & n39104 ;
  assign n39106 = n3626 | n24305 ;
  assign n39107 = n39106 ^ n13715 ^ 1'b0 ;
  assign n39108 = n35076 ^ n16712 ^ n3296 ;
  assign n39109 = n5159 & ~n39108 ;
  assign n39110 = n30487 ^ n1636 ^ 1'b0 ;
  assign n39111 = n10222 & ~n39110 ;
  assign n39112 = n24169 & n24726 ;
  assign n39113 = n30221 ^ n19504 ^ 1'b0 ;
  assign n39114 = n9461 | n10112 ;
  assign n39115 = n39114 ^ n30772 ^ 1'b0 ;
  assign n39116 = n11608 | n35301 ;
  assign n39117 = n17522 & ~n36568 ;
  assign n39118 = n39116 & n39117 ;
  assign n39119 = n4137 & n18095 ;
  assign n39120 = n21705 ^ n18409 ^ 1'b0 ;
  assign n39121 = n11488 & n20684 ;
  assign n39122 = n39121 ^ x105 ^ 1'b0 ;
  assign n39123 = n23004 | n29557 ;
  assign n39124 = n556 | n3675 ;
  assign n39125 = n39124 ^ n11064 ^ 1'b0 ;
  assign n39126 = n39125 ^ n14419 ^ 1'b0 ;
  assign n39127 = n32872 & n39126 ;
  assign n39128 = ( n19677 & n27666 ) | ( n19677 & ~n39127 ) | ( n27666 & ~n39127 ) ;
  assign n39129 = n23230 ^ n5145 ^ 1'b0 ;
  assign n39130 = n5051 & ~n39129 ;
  assign n39131 = n39130 ^ n26529 ^ n15772 ;
  assign n39132 = n4544 & n16228 ;
  assign n39133 = n39132 ^ n23647 ^ 1'b0 ;
  assign n39134 = n1489 & n30563 ;
  assign n39135 = n39134 ^ n14421 ^ 1'b0 ;
  assign n39136 = n7046 & n39135 ;
  assign n39137 = n39136 ^ n5264 ^ 1'b0 ;
  assign n39138 = n37450 & n39137 ;
  assign n39139 = n28378 & n39138 ;
  assign n39140 = n39139 ^ n31161 ^ 1'b0 ;
  assign n39141 = n33379 ^ n1312 ^ 1'b0 ;
  assign n39142 = n21675 & n39141 ;
  assign n39143 = n5361 & n39142 ;
  assign n39144 = n12193 & n22814 ;
  assign n39145 = n39144 ^ n21590 ^ 1'b0 ;
  assign n39146 = ~n39143 & n39145 ;
  assign n39147 = n3073 & n14286 ;
  assign n39149 = n14250 ^ n10011 ^ 1'b0 ;
  assign n39148 = n27597 & ~n32922 ;
  assign n39150 = n39149 ^ n39148 ^ 1'b0 ;
  assign n39151 = ( ~n2685 & n3175 ) | ( ~n2685 & n39150 ) | ( n3175 & n39150 ) ;
  assign n39152 = n1284 | n10939 ;
  assign n39153 = n39152 ^ n5225 ^ n5031 ;
  assign n39154 = n39153 ^ n9960 ^ 1'b0 ;
  assign n39155 = ( ~n5543 & n16812 ) | ( ~n5543 & n39154 ) | ( n16812 & n39154 ) ;
  assign n39156 = n7700 | n9589 ;
  assign n39157 = n39156 ^ x187 ^ 1'b0 ;
  assign n39158 = n39157 ^ n5544 ^ 1'b0 ;
  assign n39159 = n21959 ^ n9008 ^ 1'b0 ;
  assign n39160 = n18115 | n39159 ;
  assign n39161 = ( n3078 & ~n5141 ) | ( n3078 & n13780 ) | ( ~n5141 & n13780 ) ;
  assign n39162 = n8137 & ~n24159 ;
  assign n39163 = n39162 ^ n20851 ^ n4759 ;
  assign n39164 = ( ~n10292 & n10513 ) | ( ~n10292 & n18069 ) | ( n10513 & n18069 ) ;
  assign n39165 = n39164 ^ n18881 ^ n18440 ;
  assign n39166 = ~n2955 & n11518 ;
  assign n39167 = n39166 ^ n27163 ^ 1'b0 ;
  assign n39168 = n7960 | n29922 ;
  assign n39169 = n11265 & ~n39168 ;
  assign n39170 = n32214 ^ n19895 ^ 1'b0 ;
  assign n39171 = ~n38159 & n39170 ;
  assign n39176 = n10844 | n11512 ;
  assign n39177 = n19554 & ~n39176 ;
  assign n39178 = n39177 ^ n14421 ^ n10776 ;
  assign n39174 = n4419 & ~n7305 ;
  assign n39172 = ~x241 & n2692 ;
  assign n39173 = n39172 ^ n2769 ^ 1'b0 ;
  assign n39175 = n39174 ^ n39173 ^ n31910 ;
  assign n39179 = n39178 ^ n39175 ^ 1'b0 ;
  assign n39180 = n14036 & ~n39179 ;
  assign n39181 = n39180 ^ n6607 ^ 1'b0 ;
  assign n39182 = n22068 ^ n780 ^ 1'b0 ;
  assign n39183 = n24340 & ~n39182 ;
  assign n39184 = n11050 & n39183 ;
  assign n39188 = n19579 ^ n12059 ^ 1'b0 ;
  assign n39185 = n10028 & ~n10770 ;
  assign n39186 = n4412 & n39185 ;
  assign n39187 = ~n10679 & n39186 ;
  assign n39189 = n39188 ^ n39187 ^ n19922 ;
  assign n39190 = ( ~n15919 & n33911 ) | ( ~n15919 & n39189 ) | ( n33911 & n39189 ) ;
  assign n39191 = n7581 & ~n12915 ;
  assign n39192 = ~n2847 & n39191 ;
  assign n39193 = n39192 ^ n39080 ^ 1'b0 ;
  assign n39194 = n33331 ^ n5164 ^ 1'b0 ;
  assign n39195 = n11127 ^ n698 ^ 1'b0 ;
  assign n39196 = n27324 & ~n39195 ;
  assign n39197 = n8507 | n13848 ;
  assign n39198 = n15282 | n39197 ;
  assign n39199 = n39198 ^ n35371 ^ 1'b0 ;
  assign n39201 = n6085 & n11913 ;
  assign n39202 = n39201 ^ n13517 ^ 1'b0 ;
  assign n39203 = n39202 ^ n7426 ^ 1'b0 ;
  assign n39200 = n29971 | n30072 ;
  assign n39204 = n39203 ^ n39200 ^ 1'b0 ;
  assign n39205 = n12427 ^ n11153 ^ n10512 ;
  assign n39206 = n12253 ^ n4247 ^ 1'b0 ;
  assign n39207 = n39206 ^ n1430 ^ 1'b0 ;
  assign n39208 = n13048 & n32428 ;
  assign n39209 = n13597 & n39208 ;
  assign n39210 = n24086 | n33417 ;
  assign n39211 = ( n5537 & n17849 ) | ( n5537 & ~n21198 ) | ( n17849 & ~n21198 ) ;
  assign n39212 = n21937 | n39211 ;
  assign n39213 = n39212 ^ n18492 ^ 1'b0 ;
  assign n39214 = n984 & ~n14429 ;
  assign n39215 = ~n10935 & n39214 ;
  assign n39216 = ~n3708 & n6601 ;
  assign n39217 = n39216 ^ n6856 ^ n2543 ;
  assign n39218 = n19884 ^ n9307 ^ 1'b0 ;
  assign n39219 = ~n29608 & n39218 ;
  assign n39220 = ~x144 & n39219 ;
  assign n39221 = ( n20944 & n39217 ) | ( n20944 & ~n39220 ) | ( n39217 & ~n39220 ) ;
  assign n39222 = n19138 & n39221 ;
  assign n39223 = n36494 ^ n20798 ^ 1'b0 ;
  assign n39224 = n6730 & ~n24699 ;
  assign n39225 = n17435 & ~n29232 ;
  assign n39226 = ~n10054 & n39225 ;
  assign n39227 = n5731 | n8352 ;
  assign n39228 = n39226 & ~n39227 ;
  assign n39229 = n5843 | n9946 ;
  assign n39230 = n39229 ^ n783 ^ 1'b0 ;
  assign n39231 = n1145 & ~n39230 ;
  assign n39232 = n37729 ^ n22163 ^ 1'b0 ;
  assign n39233 = n39231 & n39232 ;
  assign n39234 = ( n1880 & n15912 ) | ( n1880 & n35168 ) | ( n15912 & n35168 ) ;
  assign n39235 = n39234 ^ n16330 ^ n5010 ;
  assign n39236 = n12489 ^ n4253 ^ 1'b0 ;
  assign n39237 = n9729 & ~n39236 ;
  assign n39238 = ~n9074 & n23203 ;
  assign n39239 = n39238 ^ n9720 ^ 1'b0 ;
  assign n39240 = ( ~n20481 & n34957 ) | ( ~n20481 & n36043 ) | ( n34957 & n36043 ) ;
  assign n39241 = n9133 & ~n39240 ;
  assign n39242 = n11278 ^ n10717 ^ 1'b0 ;
  assign n39243 = n20347 ^ n6528 ^ 1'b0 ;
  assign n39244 = n33575 & n39243 ;
  assign n39245 = ~n6451 & n39244 ;
  assign n39246 = n28870 & n37739 ;
  assign n39247 = ~n2690 & n39246 ;
  assign n39248 = n30493 & ~n39247 ;
  assign n39249 = n29103 ^ n26985 ^ 1'b0 ;
  assign n39250 = ~n20797 & n39249 ;
  assign n39251 = n12514 | n27634 ;
  assign n39252 = n39251 ^ n18731 ^ 1'b0 ;
  assign n39253 = n1959 & ~n39252 ;
  assign n39254 = n11350 ^ n9367 ^ 1'b0 ;
  assign n39255 = ~n4454 & n14244 ;
  assign n39256 = n39255 ^ n19281 ^ n10525 ;
  assign n39257 = n5398 ^ n5227 ^ 1'b0 ;
  assign n39258 = n39257 ^ n20845 ^ 1'b0 ;
  assign n39259 = n11290 & ~n39258 ;
  assign n39260 = n23617 ^ n1719 ^ 1'b0 ;
  assign n39261 = n39260 ^ n3985 ^ 1'b0 ;
  assign n39262 = n20957 & n30444 ;
  assign n39263 = n37916 ^ n23145 ^ 1'b0 ;
  assign n39264 = ~n1797 & n39263 ;
  assign n39265 = ( n6929 & n27172 ) | ( n6929 & n39264 ) | ( n27172 & n39264 ) ;
  assign n39266 = n3134 ^ n3055 ^ n400 ;
  assign n39267 = n24928 ^ n19234 ^ 1'b0 ;
  assign n39268 = ~n4915 & n39267 ;
  assign n39269 = ~n39266 & n39268 ;
  assign n39270 = n39269 ^ n2732 ^ 1'b0 ;
  assign n39271 = n13441 | n29522 ;
  assign n39272 = n13712 | n35707 ;
  assign n39273 = n2337 & n24708 ;
  assign n39274 = n25621 | n28564 ;
  assign n39275 = n6665 | n39274 ;
  assign n39276 = n32034 & n39275 ;
  assign n39277 = ~n17296 & n23110 ;
  assign n39278 = n39277 ^ n9856 ^ 1'b0 ;
  assign n39279 = ( n4907 & n33506 ) | ( n4907 & ~n39278 ) | ( n33506 & ~n39278 ) ;
  assign n39280 = n1913 | n9608 ;
  assign n39281 = n1920 | n39280 ;
  assign n39282 = n39281 ^ n10925 ^ 1'b0 ;
  assign n39283 = n39282 ^ n4168 ^ n439 ;
  assign n39284 = n25688 | n33274 ;
  assign n39285 = n7508 & n39284 ;
  assign n39286 = n12888 ^ n5711 ^ 1'b0 ;
  assign n39287 = n16981 ^ n3283 ^ n3193 ;
  assign n39288 = n39287 ^ n21383 ^ 1'b0 ;
  assign n39289 = n3254 ^ n1227 ^ 1'b0 ;
  assign n39290 = n553 | n39289 ;
  assign n39291 = n10573 & ~n39290 ;
  assign n39292 = n35191 ^ n11646 ^ n1571 ;
  assign n39293 = n2349 ^ n1651 ^ 1'b0 ;
  assign n39294 = n39293 ^ n9640 ^ 1'b0 ;
  assign n39295 = ~n4550 & n12359 ;
  assign n39296 = n15182 | n24955 ;
  assign n39297 = n283 | n18868 ;
  assign n39298 = n24544 & n39297 ;
  assign n39299 = ~n3391 & n20039 ;
  assign n39300 = ~n14903 & n39299 ;
  assign n39301 = n2621 & ~n39300 ;
  assign n39302 = ~n3272 & n39301 ;
  assign n39303 = n8791 ^ n880 ^ 1'b0 ;
  assign n39304 = n39302 | n39303 ;
  assign n39305 = n39304 ^ n34695 ^ n30383 ;
  assign n39306 = ( ~n3688 & n14677 ) | ( ~n3688 & n25534 ) | ( n14677 & n25534 ) ;
  assign n39307 = n1600 | n5887 ;
  assign n39308 = n24403 ^ n7060 ^ n2050 ;
  assign n39309 = n15509 ^ n15227 ^ 1'b0 ;
  assign n39310 = n39308 | n39309 ;
  assign n39311 = ( n11419 & n39307 ) | ( n11419 & ~n39310 ) | ( n39307 & ~n39310 ) ;
  assign n39312 = ( ~n10935 & n39306 ) | ( ~n10935 & n39311 ) | ( n39306 & n39311 ) ;
  assign n39313 = ( n5864 & n10230 ) | ( n5864 & n28067 ) | ( n10230 & n28067 ) ;
  assign n39314 = n13343 & ~n35136 ;
  assign n39315 = n11091 ^ n2855 ^ 1'b0 ;
  assign n39316 = ~n11887 & n39315 ;
  assign n39317 = n5532 & ~n33627 ;
  assign n39318 = n39317 ^ n26593 ^ n25471 ;
  assign n39319 = n37546 ^ n16608 ^ n7253 ;
  assign n39324 = n3943 & n8019 ;
  assign n39325 = n7826 & n39324 ;
  assign n39323 = n14687 | n37566 ;
  assign n39326 = n39325 ^ n39323 ^ 1'b0 ;
  assign n39320 = n20694 & ~n31383 ;
  assign n39321 = n39320 ^ n23944 ^ 1'b0 ;
  assign n39322 = n26295 & ~n39321 ;
  assign n39327 = n39326 ^ n39322 ^ 1'b0 ;
  assign n39328 = n39327 ^ n12440 ^ 1'b0 ;
  assign n39329 = n36485 ^ n30978 ^ 1'b0 ;
  assign n39330 = n15741 & n19237 ;
  assign n39331 = n39330 ^ n11974 ^ 1'b0 ;
  assign n39332 = n16925 ^ n13508 ^ 1'b0 ;
  assign n39333 = n9790 & n39332 ;
  assign n39334 = n26267 ^ n22186 ^ 1'b0 ;
  assign n39335 = n39266 | n39334 ;
  assign n39336 = ( ~n9181 & n24725 ) | ( ~n9181 & n26664 ) | ( n24725 & n26664 ) ;
  assign n39337 = n4981 ^ n1330 ^ 1'b0 ;
  assign n39338 = n3706 & n7495 ;
  assign n39339 = n39338 ^ n22177 ^ 1'b0 ;
  assign n39340 = n27290 ^ n17137 ^ 1'b0 ;
  assign n39341 = n39339 & n39340 ;
  assign n39342 = n17198 ^ n8734 ^ 1'b0 ;
  assign n39343 = n33189 ^ n15413 ^ n1312 ;
  assign n39346 = ( n581 & ~n12144 ) | ( n581 & n14909 ) | ( ~n12144 & n14909 ) ;
  assign n39344 = n31576 ^ n8474 ^ 1'b0 ;
  assign n39345 = n39344 ^ n10414 ^ 1'b0 ;
  assign n39347 = n39346 ^ n39345 ^ n38849 ;
  assign n39348 = n20103 | n21461 ;
  assign n39349 = n39348 ^ n19166 ^ 1'b0 ;
  assign n39350 = n20009 | n20684 ;
  assign n39351 = n32072 ^ n19142 ^ n18645 ;
  assign n39352 = n39350 | n39351 ;
  assign n39353 = n39349 | n39352 ;
  assign n39354 = n22433 ^ n10243 ^ 1'b0 ;
  assign n39355 = n2909 & n39354 ;
  assign n39356 = n11246 | n12592 ;
  assign n39357 = n10125 | n33200 ;
  assign n39358 = n10022 | n39357 ;
  assign n39359 = n39358 ^ n26650 ^ 1'b0 ;
  assign n39360 = n36359 ^ n16602 ^ 1'b0 ;
  assign n39366 = n9259 ^ n7937 ^ 1'b0 ;
  assign n39361 = ~n2661 & n5905 ;
  assign n39362 = n357 & n39361 ;
  assign n39363 = n11692 | n39362 ;
  assign n39364 = n39363 ^ n18869 ^ 1'b0 ;
  assign n39365 = n24196 & ~n39364 ;
  assign n39367 = n39366 ^ n39365 ^ 1'b0 ;
  assign n39368 = n2501 ^ n2497 ^ 1'b0 ;
  assign n39369 = n6382 | n39368 ;
  assign n39370 = n39369 ^ n806 ^ 1'b0 ;
  assign n39371 = n25381 ^ n9709 ^ 1'b0 ;
  assign n39372 = ~n36139 & n39371 ;
  assign n39373 = ~n4775 & n10848 ;
  assign n39374 = n39373 ^ n34763 ^ 1'b0 ;
  assign n39375 = n19948 ^ n15240 ^ 1'b0 ;
  assign n39376 = ( n1160 & ~n5746 ) | ( n1160 & n17192 ) | ( ~n5746 & n17192 ) ;
  assign n39377 = n25996 | n39376 ;
  assign n39378 = n30304 ^ n5722 ^ 1'b0 ;
  assign n39379 = ~n26604 & n39378 ;
  assign n39380 = n2623 | n23562 ;
  assign n39381 = n39380 ^ n32135 ^ 1'b0 ;
  assign n39382 = n1421 & n18371 ;
  assign n39383 = n39382 ^ n2644 ^ 1'b0 ;
  assign n39384 = n39381 | n39383 ;
  assign n39385 = n27496 ^ n10262 ^ 1'b0 ;
  assign n39386 = n39384 | n39385 ;
  assign n39387 = n11394 & ~n35060 ;
  assign n39388 = n39387 ^ n5852 ^ 1'b0 ;
  assign n39389 = n16093 ^ n5040 ^ 1'b0 ;
  assign n39390 = n6622 | n39389 ;
  assign n39391 = ( n1164 & n2661 ) | ( n1164 & ~n39390 ) | ( n2661 & ~n39390 ) ;
  assign n39392 = n15102 & ~n23362 ;
  assign n39393 = ~n2307 & n35554 ;
  assign n39394 = n39393 ^ n7839 ^ 1'b0 ;
  assign n39395 = n30776 & ~n39394 ;
  assign n39396 = ~n20847 & n39395 ;
  assign n39397 = n2888 & ~n27450 ;
  assign n39398 = ~n6353 & n7743 ;
  assign n39399 = n29970 ^ n14379 ^ 1'b0 ;
  assign n39400 = n39398 & ~n39399 ;
  assign n39401 = n28884 ^ n5081 ^ 1'b0 ;
  assign n39402 = n12209 & ~n39401 ;
  assign n39403 = n39402 ^ n13889 ^ n2875 ;
  assign n39404 = n39400 & ~n39403 ;
  assign n39405 = n10994 ^ n7776 ^ 1'b0 ;
  assign n39406 = n13621 & n28530 ;
  assign n39407 = ~n39405 & n39406 ;
  assign n39408 = n39307 & n39407 ;
  assign n39409 = ~n9725 & n27403 ;
  assign n39410 = n39408 & n39409 ;
  assign n39412 = n7593 | n31289 ;
  assign n39413 = n39412 ^ n12710 ^ 1'b0 ;
  assign n39414 = n39413 ^ n28087 ^ n7468 ;
  assign n39411 = ~n5230 & n30924 ;
  assign n39415 = n39414 ^ n39411 ^ 1'b0 ;
  assign n39416 = ~n511 & n39080 ;
  assign n39417 = n1671 & n39416 ;
  assign n39418 = ( ~n407 & n11239 ) | ( ~n407 & n39417 ) | ( n11239 & n39417 ) ;
  assign n39419 = n24471 ^ n11844 ^ n7917 ;
  assign n39420 = ( ~x13 & n19852 ) | ( ~x13 & n39419 ) | ( n19852 & n39419 ) ;
  assign n39421 = n2173 & n30809 ;
  assign n39422 = n39421 ^ n5721 ^ 1'b0 ;
  assign n39423 = ( ~n3751 & n4832 ) | ( ~n3751 & n39422 ) | ( n4832 & n39422 ) ;
  assign n39424 = n4406 & n10563 ;
  assign n39425 = n28327 ^ n1866 ^ 1'b0 ;
  assign n39426 = ~n9572 & n39425 ;
  assign n39427 = ~n39424 & n39426 ;
  assign n39428 = n39423 | n39427 ;
  assign n39429 = n36188 ^ n28342 ^ n9667 ;
  assign n39430 = ~n4876 & n39429 ;
  assign n39431 = n34766 ^ n12579 ^ 1'b0 ;
  assign n39432 = n11938 | n39431 ;
  assign n39433 = n2966 & n11345 ;
  assign n39434 = n39433 ^ n5285 ^ 1'b0 ;
  assign n39435 = ~n2246 & n8296 ;
  assign n39436 = n39435 ^ n22853 ^ 1'b0 ;
  assign n39437 = n13135 & ~n21286 ;
  assign n39438 = n27267 ^ n1551 ^ 1'b0 ;
  assign n39439 = ~n39437 & n39438 ;
  assign n39440 = n26489 & n39439 ;
  assign n39441 = ~n4236 & n39440 ;
  assign n39442 = n5762 & n15847 ;
  assign n39443 = n23518 ^ n17170 ^ 1'b0 ;
  assign n39444 = n8432 & n28979 ;
  assign n39445 = ~n6561 & n39444 ;
  assign n39446 = n39445 ^ n12957 ^ 1'b0 ;
  assign n39447 = n39446 ^ n16186 ^ 1'b0 ;
  assign n39448 = ( n39442 & n39443 ) | ( n39442 & n39447 ) | ( n39443 & n39447 ) ;
  assign n39449 = n23659 & ~n26457 ;
  assign n39450 = n21773 ^ n16140 ^ 1'b0 ;
  assign n39451 = n541 & n27629 ;
  assign n39452 = n11530 ^ n7661 ^ 1'b0 ;
  assign n39453 = n35312 & ~n39452 ;
  assign n39454 = n2061 & n39453 ;
  assign n39455 = n959 & n39454 ;
  assign n39456 = n39455 ^ n2866 ^ 1'b0 ;
  assign n39457 = n7062 & n27128 ;
  assign n39458 = n39457 ^ n26951 ^ 1'b0 ;
  assign n39459 = n18083 & ~n37855 ;
  assign n39460 = n39459 ^ n8848 ^ 1'b0 ;
  assign n39461 = n20828 & n39460 ;
  assign n39462 = n712 | n5731 ;
  assign n39463 = n5432 & ~n39462 ;
  assign n39464 = n21117 ^ n16218 ^ 1'b0 ;
  assign n39465 = n39463 | n39464 ;
  assign n39466 = n39465 ^ n27598 ^ 1'b0 ;
  assign n39467 = ~n28457 & n36394 ;
  assign n39468 = n30727 ^ n17694 ^ 1'b0 ;
  assign n39469 = n3095 & n39468 ;
  assign n39470 = ~n35002 & n39469 ;
  assign n39471 = n24681 ^ n10313 ^ 1'b0 ;
  assign n39472 = ~n10088 & n39471 ;
  assign n39473 = ~n4216 & n5051 ;
  assign n39474 = n11740 & n39473 ;
  assign n39475 = n27932 ^ n21931 ^ x221 ;
  assign n39476 = n39475 ^ n29643 ^ 1'b0 ;
  assign n39477 = n7573 & ~n12297 ;
  assign n39478 = n13757 & n27947 ;
  assign n39479 = ~n39477 & n39478 ;
  assign n39480 = n33742 ^ n14302 ^ 1'b0 ;
  assign n39481 = n38359 & n39480 ;
  assign n39482 = n10582 & ~n11580 ;
  assign n39483 = n39482 ^ n17853 ^ 1'b0 ;
  assign n39485 = n1582 & ~n3707 ;
  assign n39484 = n5869 & ~n23242 ;
  assign n39486 = n39485 ^ n39484 ^ 1'b0 ;
  assign n39487 = n32901 ^ n29277 ^ 1'b0 ;
  assign n39488 = n14917 & n39487 ;
  assign n39489 = ~n16800 & n29879 ;
  assign n39490 = n39489 ^ n16625 ^ 1'b0 ;
  assign n39491 = x197 & ~n9613 ;
  assign n39492 = ~n6355 & n39491 ;
  assign n39493 = n11853 | n39492 ;
  assign n39494 = n7017 | n39493 ;
  assign n39495 = n39494 ^ n29795 ^ 1'b0 ;
  assign n39496 = n2651 & n13757 ;
  assign n39497 = n39496 ^ n6240 ^ 1'b0 ;
  assign n39498 = n5221 & n16920 ;
  assign n39499 = ~n39497 & n39498 ;
  assign n39500 = ~n18629 & n39499 ;
  assign n39501 = ~n14830 & n18283 ;
  assign n39502 = n39501 ^ n15656 ^ 1'b0 ;
  assign n39503 = n39502 ^ n1875 ^ 1'b0 ;
  assign n39504 = n8756 | n39503 ;
  assign n39505 = n38489 ^ n36729 ^ 1'b0 ;
  assign n39506 = n7466 ^ n5841 ^ 1'b0 ;
  assign n39507 = n32745 ^ n16205 ^ n10221 ;
  assign n39508 = n5988 | n11083 ;
  assign n39509 = n39507 & ~n39508 ;
  assign n39510 = n9127 & n30100 ;
  assign n39511 = n8435 | n39510 ;
  assign n39512 = n8270 | n39511 ;
  assign n39513 = ~n10102 & n39068 ;
  assign n39514 = ~n31656 & n39513 ;
  assign n39515 = n39514 ^ n10408 ^ 1'b0 ;
  assign n39517 = n7469 ^ n589 ^ 1'b0 ;
  assign n39518 = n23983 | n39517 ;
  assign n39516 = ~n4507 & n14449 ;
  assign n39519 = n39518 ^ n39516 ^ n31640 ;
  assign n39520 = n31003 ^ n6007 ^ 1'b0 ;
  assign n39521 = n21186 | n25627 ;
  assign n39522 = n13589 & ~n39521 ;
  assign n39523 = n27499 & ~n29032 ;
  assign n39524 = n8485 & ~n12377 ;
  assign n39525 = ~n5338 & n39524 ;
  assign n39526 = ~n1805 & n39525 ;
  assign n39527 = n13068 ^ n5929 ^ 1'b0 ;
  assign n39528 = ( n6597 & n33404 ) | ( n6597 & ~n39527 ) | ( n33404 & ~n39527 ) ;
  assign n39529 = n39528 ^ n31234 ^ n3681 ;
  assign n39530 = n4335 & n39529 ;
  assign n39531 = n39526 | n39530 ;
  assign n39532 = n9260 | n29656 ;
  assign n39533 = n3895 & ~n39532 ;
  assign n39534 = n20166 | n27194 ;
  assign n39535 = ~n8654 & n19998 ;
  assign n39536 = ~n16827 & n39535 ;
  assign n39537 = n39536 ^ n8243 ^ 1'b0 ;
  assign n39538 = n4218 & ~n39537 ;
  assign n39539 = n39538 ^ n18544 ^ n3850 ;
  assign n39540 = n39539 ^ n1976 ^ 1'b0 ;
  assign n39541 = n15550 ^ n11983 ^ 1'b0 ;
  assign n39542 = n9979 ^ n8066 ^ 1'b0 ;
  assign n39543 = ~n39541 & n39542 ;
  assign n39544 = n2843 & n39543 ;
  assign n39545 = n18164 ^ n2547 ^ 1'b0 ;
  assign n39546 = n16665 ^ n4353 ^ x20 ;
  assign n39547 = n10142 & ~n37946 ;
  assign n39548 = n39547 ^ n28319 ^ 1'b0 ;
  assign n39549 = ( ~n19247 & n20968 ) | ( ~n19247 & n28129 ) | ( n20968 & n28129 ) ;
  assign n39550 = n16865 & ~n39549 ;
  assign n39551 = n39252 ^ n9528 ^ 1'b0 ;
  assign n39552 = n4824 | n39551 ;
  assign n39553 = ~n30388 & n37243 ;
  assign n39554 = n39552 & n39553 ;
  assign n39555 = n17344 & ~n20539 ;
  assign n39556 = n12011 & n39555 ;
  assign n39559 = n16174 & n19220 ;
  assign n39557 = ( ~n5974 & n13744 ) | ( ~n5974 & n15717 ) | ( n13744 & n15717 ) ;
  assign n39558 = n1041 & ~n39557 ;
  assign n39560 = n39559 ^ n39558 ^ n8751 ;
  assign n39561 = n2603 ^ n2176 ^ 1'b0 ;
  assign n39562 = n6849 & ~n39561 ;
  assign n39563 = n30380 & n34561 ;
  assign n39564 = n39563 ^ n19746 ^ 1'b0 ;
  assign n39565 = ( n3011 & ~n5138 ) | ( n3011 & n8493 ) | ( ~n5138 & n8493 ) ;
  assign n39566 = n34812 ^ n2202 ^ 1'b0 ;
  assign n39567 = ~n39565 & n39566 ;
  assign n39568 = ( ~n39562 & n39564 ) | ( ~n39562 & n39567 ) | ( n39564 & n39567 ) ;
  assign n39569 = n13704 ^ n4795 ^ 1'b0 ;
  assign n39570 = n9299 & n39569 ;
  assign n39571 = n15388 ^ n10767 ^ 1'b0 ;
  assign n39572 = n39570 & ~n39571 ;
  assign n39573 = ~n34871 & n39572 ;
  assign n39578 = n37204 ^ n24803 ^ 1'b0 ;
  assign n39574 = n4338 & ~n15124 ;
  assign n39575 = n27570 & n31093 ;
  assign n39576 = n39575 ^ n35677 ^ 1'b0 ;
  assign n39577 = n39574 & ~n39576 ;
  assign n39579 = n39578 ^ n39577 ^ 1'b0 ;
  assign n39580 = n10991 | n39579 ;
  assign n39581 = n3427 & n21041 ;
  assign n39582 = n8075 & n39581 ;
  assign n39583 = x3 | n22622 ;
  assign n39584 = n29046 | n39583 ;
  assign n39585 = n5167 & n7881 ;
  assign n39586 = ~n39584 & n39585 ;
  assign n39587 = n25213 ^ n2719 ^ 1'b0 ;
  assign n39588 = n13017 ^ n12361 ^ n10444 ;
  assign n39589 = n5226 & ~n14204 ;
  assign n39590 = n39589 ^ n32594 ^ n20946 ;
  assign n39591 = n818 & ~n29469 ;
  assign n39592 = ~n1744 & n26141 ;
  assign n39593 = n39592 ^ n18889 ^ 1'b0 ;
  assign n39594 = n15682 ^ n6644 ^ 1'b0 ;
  assign n39595 = n29461 ^ n5496 ^ n376 ;
  assign n39596 = ( n2561 & n9866 ) | ( n2561 & ~n37029 ) | ( n9866 & ~n37029 ) ;
  assign n39597 = n31205 ^ n18609 ^ 1'b0 ;
  assign n39598 = n20622 | n39597 ;
  assign n39599 = n2609 | n16805 ;
  assign n39600 = n18835 ^ n2949 ^ 1'b0 ;
  assign n39601 = n19917 | n22831 ;
  assign n39603 = n612 | n5597 ;
  assign n39604 = n39603 ^ n17625 ^ 1'b0 ;
  assign n39602 = ~n8654 & n9810 ;
  assign n39605 = n39604 ^ n39602 ^ 1'b0 ;
  assign n39606 = n38731 | n39605 ;
  assign n39607 = n10071 & ~n39606 ;
  assign n39608 = n22422 ^ n10771 ^ n455 ;
  assign n39609 = n24556 ^ n1835 ^ 1'b0 ;
  assign n39610 = n20586 | n39609 ;
  assign n39611 = n30608 ^ n15975 ^ n993 ;
  assign n39612 = n12112 ^ n11143 ^ 1'b0 ;
  assign n39615 = n34472 ^ n22139 ^ n13555 ;
  assign n39613 = n33820 ^ n11348 ^ 1'b0 ;
  assign n39614 = n38299 | n39613 ;
  assign n39616 = n39615 ^ n39614 ^ 1'b0 ;
  assign n39617 = n3927 & n4719 ;
  assign n39618 = n1473 | n1975 ;
  assign n39619 = n39618 ^ n8430 ^ 1'b0 ;
  assign n39620 = n39619 ^ n14644 ^ 1'b0 ;
  assign n39621 = n18457 | n20662 ;
  assign n39622 = n13941 ^ n6798 ^ 1'b0 ;
  assign n39623 = ~n17046 & n39622 ;
  assign n39624 = n39623 ^ n10872 ^ 1'b0 ;
  assign n39625 = n33947 ^ n21991 ^ 1'b0 ;
  assign n39626 = n16090 ^ n10879 ^ 1'b0 ;
  assign n39627 = n16045 | n39626 ;
  assign n39628 = n39627 ^ n31028 ^ n11791 ;
  assign n39629 = n19264 | n39405 ;
  assign n39630 = n39629 ^ n7710 ^ 1'b0 ;
  assign n39631 = n29402 ^ n8785 ^ 1'b0 ;
  assign n39632 = n1266 & ~n39631 ;
  assign n39633 = ( n673 & n6451 ) | ( n673 & n7420 ) | ( n6451 & n7420 ) ;
  assign n39634 = n39633 ^ n9804 ^ 1'b0 ;
  assign n39635 = n39632 & ~n39634 ;
  assign n39636 = n8478 ^ n2436 ^ 1'b0 ;
  assign n39637 = n9009 ^ n6590 ^ 1'b0 ;
  assign n39638 = n13031 | n39637 ;
  assign n39639 = n32075 | n39638 ;
  assign n39640 = n39639 ^ n20868 ^ 1'b0 ;
  assign n39641 = ( ~n8058 & n24292 ) | ( ~n8058 & n29424 ) | ( n24292 & n29424 ) ;
  assign n39642 = n2799 & ~n5988 ;
  assign n39643 = n39642 ^ n23239 ^ n11699 ;
  assign n39644 = n3244 & n39643 ;
  assign n39645 = ( x239 & n30948 ) | ( x239 & n39644 ) | ( n30948 & n39644 ) ;
  assign n39646 = n22658 ^ n5760 ^ 1'b0 ;
  assign n39647 = ~n30512 & n39646 ;
  assign n39648 = n11332 ^ n3294 ^ 1'b0 ;
  assign n39649 = x114 & n39648 ;
  assign n39650 = ~n5594 & n39649 ;
  assign n39651 = n1286 & n28322 ;
  assign n39652 = n39650 & n39651 ;
  assign n39653 = n5298 & ~n17062 ;
  assign n39654 = n39653 ^ n5987 ^ 1'b0 ;
  assign n39655 = n22737 & ~n39654 ;
  assign n39656 = n27731 & n39655 ;
  assign n39657 = n824 & ~n39656 ;
  assign n39658 = n6877 & n39657 ;
  assign n39659 = n6515 | n22089 ;
  assign n39660 = n7433 & ~n22863 ;
  assign n39666 = n20233 & ~n29165 ;
  assign n39661 = n2360 ^ n697 ^ 1'b0 ;
  assign n39662 = n7171 ^ n2096 ^ 1'b0 ;
  assign n39663 = ~n8535 & n39662 ;
  assign n39664 = n15080 & n39663 ;
  assign n39665 = n39661 & n39664 ;
  assign n39667 = n39666 ^ n39665 ^ n16711 ;
  assign n39668 = ( ~n2142 & n6539 ) | ( ~n2142 & n21952 ) | ( n6539 & n21952 ) ;
  assign n39669 = n8428 & ~n22980 ;
  assign n39670 = ~n39668 & n39669 ;
  assign n39671 = x210 & ~n39670 ;
  assign n39682 = ~n1124 & n3182 ;
  assign n39683 = ~n3182 & n39682 ;
  assign n39684 = n1760 & ~n39683 ;
  assign n39685 = n39683 & n39684 ;
  assign n39686 = n1742 & ~n39685 ;
  assign n39687 = n39685 & n39686 ;
  assign n39688 = n1469 & ~n2124 ;
  assign n39689 = n39687 & n39688 ;
  assign n39690 = n2402 | n3919 ;
  assign n39691 = n39689 & ~n39690 ;
  assign n39692 = n8227 & ~n39691 ;
  assign n39693 = n39691 & n39692 ;
  assign n39672 = x11 & n736 ;
  assign n39673 = ~n736 & n39672 ;
  assign n39674 = x82 & ~n1210 ;
  assign n39675 = n1210 & n39674 ;
  assign n39676 = n39675 ^ n829 ^ 1'b0 ;
  assign n39677 = x238 & n39676 ;
  assign n39678 = n39673 & n39677 ;
  assign n39679 = n13763 & ~n39678 ;
  assign n39680 = n39678 & n39679 ;
  assign n39681 = n21526 & ~n39680 ;
  assign n39694 = n39693 ^ n39681 ^ 1'b0 ;
  assign n39695 = n12213 & n39183 ;
  assign n39696 = n948 & n39695 ;
  assign n39697 = n4136 & ~n39696 ;
  assign n39698 = n39697 ^ n21020 ^ 1'b0 ;
  assign n39699 = n14589 & n18728 ;
  assign n39700 = ~n332 & n11153 ;
  assign n39701 = n2073 & n39700 ;
  assign n39702 = n1281 & n12121 ;
  assign n39703 = n39702 ^ n3081 ^ 1'b0 ;
  assign n39704 = n29525 | n39703 ;
  assign n39705 = n39704 ^ n9316 ^ 1'b0 ;
  assign n39706 = n10808 & ~n33062 ;
  assign n39707 = n39705 & n39706 ;
  assign n39708 = n1596 | n2029 ;
  assign n39709 = n15902 & ~n19564 ;
  assign n39710 = ~n20923 & n39709 ;
  assign n39711 = n19948 ^ n9180 ^ n3747 ;
  assign n39712 = n28683 ^ n14102 ^ n791 ;
  assign n39713 = ~n35513 & n39712 ;
  assign n39714 = n39711 & n39713 ;
  assign n39715 = n23462 ^ n5674 ^ 1'b0 ;
  assign n39716 = n7369 & ~n39715 ;
  assign n39717 = n39716 ^ n8620 ^ 1'b0 ;
  assign n39718 = n3686 & n29136 ;
  assign n39719 = n39718 ^ n6536 ^ 1'b0 ;
  assign n39720 = n15391 & n39719 ;
  assign n39721 = n39720 ^ n3278 ^ 1'b0 ;
  assign n39722 = n5415 & ~n28233 ;
  assign n39723 = n39722 ^ n11833 ^ 1'b0 ;
  assign n39724 = n17185 ^ n535 ^ 1'b0 ;
  assign n39725 = n39723 | n39724 ;
  assign n39726 = n29194 ^ n3228 ^ 1'b0 ;
  assign n39727 = ~n28891 & n39726 ;
  assign n39728 = n8992 | n11724 ;
  assign n39729 = ~n15612 & n39728 ;
  assign n39730 = n15058 & ~n20204 ;
  assign n39731 = ~n19757 & n39730 ;
  assign n39732 = n3220 | n7156 ;
  assign n39733 = n8226 & ~n12011 ;
  assign n39734 = n39733 ^ n20700 ^ 1'b0 ;
  assign n39735 = n20395 | n39734 ;
  assign n39736 = n39735 ^ n30922 ^ 1'b0 ;
  assign n39737 = x41 & ~n1378 ;
  assign n39738 = n39737 ^ n6613 ^ 1'b0 ;
  assign n39739 = ~n15621 & n38935 ;
  assign n39740 = n6563 | n29502 ;
  assign n39741 = n39740 ^ n7861 ^ 1'b0 ;
  assign n39743 = n11745 & ~n29879 ;
  assign n39742 = ~n6613 & n11842 ;
  assign n39744 = n39743 ^ n39742 ^ 1'b0 ;
  assign n39745 = n9451 ^ n4095 ^ n860 ;
  assign n39746 = ~n706 & n39745 ;
  assign n39747 = n18161 & ~n39746 ;
  assign n39749 = n740 & n2991 ;
  assign n39750 = ~n4768 & n39749 ;
  assign n39748 = ~n4654 & n5932 ;
  assign n39751 = n39750 ^ n39748 ^ 1'b0 ;
  assign n39752 = n39751 ^ n25466 ^ n8539 ;
  assign n39753 = n39752 ^ n26168 ^ 1'b0 ;
  assign n39754 = ~n16516 & n23302 ;
  assign n39755 = n39754 ^ n21661 ^ 1'b0 ;
  assign n39756 = n26817 ^ n16867 ^ 1'b0 ;
  assign n39757 = n14698 & n39756 ;
  assign n39758 = n26810 ^ x251 ^ 1'b0 ;
  assign n39759 = n716 & ~n39758 ;
  assign n39760 = n5092 ^ n2416 ^ 1'b0 ;
  assign n39761 = ~n4780 & n39760 ;
  assign n39762 = n39761 ^ n38824 ^ 1'b0 ;
  assign n39763 = n39759 & n39762 ;
  assign n39764 = n5869 & ~n21268 ;
  assign n39765 = n39764 ^ n8381 ^ 1'b0 ;
  assign n39766 = n22015 & n27866 ;
  assign n39767 = ~n9757 & n38530 ;
  assign n39768 = n2606 & n11469 ;
  assign n39769 = ~n17884 & n39768 ;
  assign n39770 = ( n4852 & n30209 ) | ( n4852 & ~n39769 ) | ( n30209 & ~n39769 ) ;
  assign n39771 = n18697 ^ n12788 ^ 1'b0 ;
  assign n39772 = n26099 & ~n29591 ;
  assign n39773 = ~n39771 & n39772 ;
  assign n39774 = n26320 ^ n13201 ^ 1'b0 ;
  assign n39775 = n15427 | n21075 ;
  assign n39776 = ( n3654 & n11967 ) | ( n3654 & ~n13757 ) | ( n11967 & ~n13757 ) ;
  assign n39777 = n11123 | n39776 ;
  assign n39778 = n24381 & ~n33817 ;
  assign n39779 = ~n39777 & n39778 ;
  assign n39780 = n17809 & ~n23843 ;
  assign n39781 = n39780 ^ n2096 ^ 1'b0 ;
  assign n39782 = n32208 ^ n3633 ^ 1'b0 ;
  assign n39783 = n29598 ^ n16324 ^ 1'b0 ;
  assign n39784 = n13447 ^ n5328 ^ 1'b0 ;
  assign n39785 = n30885 | n39784 ;
  assign n39786 = n21056 ^ n3326 ^ 1'b0 ;
  assign n39787 = n39786 ^ n36990 ^ n4597 ;
  assign n39788 = ~n2961 & n39787 ;
  assign n39789 = n39788 ^ n16585 ^ 1'b0 ;
  assign n39790 = ( n5114 & n12597 ) | ( n5114 & n30826 ) | ( n12597 & n30826 ) ;
  assign n39791 = ~n6101 & n12449 ;
  assign n39792 = n39791 ^ n7152 ^ 1'b0 ;
  assign n39793 = x30 & ~n10655 ;
  assign n39794 = ~n31732 & n39793 ;
  assign n39795 = n3099 & n39794 ;
  assign n39796 = n39795 ^ n31470 ^ 1'b0 ;
  assign n39797 = ~n11461 & n39796 ;
  assign n39798 = n20424 & ~n22647 ;
  assign n39799 = n39798 ^ n17247 ^ 1'b0 ;
  assign n39800 = n21460 ^ n8261 ^ 1'b0 ;
  assign n39801 = n21424 & ~n39800 ;
  assign n39802 = ~n4842 & n13780 ;
  assign n39803 = n23004 ^ n13342 ^ 1'b0 ;
  assign n39804 = n20908 | n39803 ;
  assign n39805 = n15920 | n28650 ;
  assign n39806 = n39805 ^ n22588 ^ n17504 ;
  assign n39807 = n25461 ^ n10333 ^ n9595 ;
  assign n39808 = n21359 & n39807 ;
  assign n39809 = n39808 ^ n9451 ^ 1'b0 ;
  assign n39811 = n3767 & ~n10600 ;
  assign n39812 = ~n20193 & n39811 ;
  assign n39813 = n8800 ^ n6592 ^ 1'b0 ;
  assign n39814 = n39812 | n39813 ;
  assign n39810 = x66 & ~n18301 ;
  assign n39815 = n39814 ^ n39810 ^ 1'b0 ;
  assign n39816 = n12251 | n33610 ;
  assign n39817 = n26743 ^ n15151 ^ n10092 ;
  assign n39818 = n39817 ^ n9469 ^ 1'b0 ;
  assign n39819 = n18338 ^ n5294 ^ 1'b0 ;
  assign n39820 = n9986 & n39819 ;
  assign n39821 = n39820 ^ n14884 ^ 1'b0 ;
  assign n39822 = ( ~n6361 & n29217 ) | ( ~n6361 & n35854 ) | ( n29217 & n35854 ) ;
  assign n39823 = n7489 | n39822 ;
  assign n39824 = n26745 & ~n36742 ;
  assign n39825 = n10787 & n17075 ;
  assign n39826 = n18575 & n39825 ;
  assign n39827 = ( n1603 & n26666 ) | ( n1603 & n32518 ) | ( n26666 & n32518 ) ;
  assign n39828 = n18379 | n39776 ;
  assign n39829 = n39828 ^ n17500 ^ x121 ;
  assign n39830 = n12755 & n14656 ;
  assign n39831 = n39830 ^ n3716 ^ 1'b0 ;
  assign n39832 = n15534 | n39831 ;
  assign n39833 = n18881 ^ n4636 ^ 1'b0 ;
  assign n39834 = n8340 & ~n39833 ;
  assign n39835 = n5542 | n6108 ;
  assign n39836 = n39835 ^ n36745 ^ 1'b0 ;
  assign n39837 = n39836 ^ n5508 ^ 1'b0 ;
  assign n39838 = n39834 & n39837 ;
  assign n39839 = n17358 & n32285 ;
  assign n39840 = ~n5924 & n35185 ;
  assign n39843 = ~x76 & n7058 ;
  assign n39844 = n14359 & ~n24270 ;
  assign n39845 = ~n39843 & n39844 ;
  assign n39841 = n10746 & ~n27630 ;
  assign n39842 = ~n12282 & n39841 ;
  assign n39846 = n39845 ^ n39842 ^ 1'b0 ;
  assign n39849 = ~n16566 & n30587 ;
  assign n39850 = ~n10025 & n39849 ;
  assign n39847 = n1024 & ~n30549 ;
  assign n39848 = ~n842 & n39847 ;
  assign n39851 = n39850 ^ n39848 ^ 1'b0 ;
  assign n39852 = ( n5177 & n25289 ) | ( n5177 & ~n30398 ) | ( n25289 & ~n30398 ) ;
  assign n39853 = n18784 ^ n8154 ^ 1'b0 ;
  assign n39854 = n11866 & n39853 ;
  assign n39855 = n39854 ^ n38504 ^ n16883 ;
  assign n39856 = n2757 | n4446 ;
  assign n39857 = ( ~n14926 & n34736 ) | ( ~n14926 & n39856 ) | ( n34736 & n39856 ) ;
  assign n39858 = n1691 | n36037 ;
  assign n39859 = n22421 & ~n39858 ;
  assign n39860 = n8332 ^ n2423 ^ n407 ;
  assign n39861 = n32358 & ~n39860 ;
  assign n39862 = n27547 & n39861 ;
  assign n39863 = n18818 | n19692 ;
  assign n39864 = n39562 ^ n12221 ^ n11236 ;
  assign n39865 = n37659 ^ n18901 ^ 1'b0 ;
  assign n39866 = ~n21951 & n39865 ;
  assign n39867 = n39866 ^ n9204 ^ 1'b0 ;
  assign n39868 = n36584 & ~n39867 ;
  assign n39869 = n39864 & n39868 ;
  assign n39870 = n39869 ^ n1593 ^ 1'b0 ;
  assign n39871 = ~n1453 & n15204 ;
  assign n39872 = n39871 ^ n17180 ^ 1'b0 ;
  assign n39873 = n14314 | n28049 ;
  assign n39874 = n39873 ^ n18465 ^ 1'b0 ;
  assign n39875 = n21087 ^ n18183 ^ n1136 ;
  assign n39876 = n39875 ^ n17820 ^ 1'b0 ;
  assign n39877 = n19850 & ~n20761 ;
  assign n39879 = n9779 | n21305 ;
  assign n39880 = n17775 | n39879 ;
  assign n39881 = n39880 ^ n3269 ^ 1'b0 ;
  assign n39882 = n7877 & ~n39881 ;
  assign n39878 = ( n1809 & n3357 ) | ( n1809 & n6375 ) | ( n3357 & n6375 ) ;
  assign n39883 = n39882 ^ n39878 ^ 1'b0 ;
  assign n39884 = n33491 ^ n6898 ^ 1'b0 ;
  assign n39885 = ( n759 & n9471 ) | ( n759 & ~n16171 ) | ( n9471 & ~n16171 ) ;
  assign n39886 = n39885 ^ n28063 ^ 1'b0 ;
  assign n39887 = n39886 ^ n11723 ^ 1'b0 ;
  assign n39888 = ~n27055 & n39887 ;
  assign n39889 = n30460 ^ n20700 ^ 1'b0 ;
  assign n39890 = n39888 & ~n39889 ;
  assign n39891 = n37477 ^ n26626 ^ n11651 ;
  assign n39892 = ~n3650 & n39297 ;
  assign n39893 = n8636 & n25640 ;
  assign n39894 = n39893 ^ x44 ^ 1'b0 ;
  assign n39895 = n16217 & n22733 ;
  assign n39896 = n18720 & n24258 ;
  assign n39897 = n39896 ^ n30100 ^ 1'b0 ;
  assign n39898 = n30468 ^ n4833 ^ n2349 ;
  assign n39899 = n404 & ~n2246 ;
  assign n39900 = n5892 | n39899 ;
  assign n39901 = n10164 | n39900 ;
  assign n39902 = n30341 ^ n22452 ^ 1'b0 ;
  assign n39903 = n39902 ^ n24921 ^ n4430 ;
  assign n39904 = n31414 | n39903 ;
  assign n39905 = n6544 | n6949 ;
  assign n39906 = n6561 & ~n39905 ;
  assign n39907 = n6881 ^ n5354 ^ 1'b0 ;
  assign n39908 = n32451 ^ n6736 ^ 1'b0 ;
  assign n39909 = n1930 & n10995 ;
  assign n39910 = n38531 & n39909 ;
  assign n39911 = n39910 ^ n17759 ^ n14802 ;
  assign n39912 = n39911 ^ n36232 ^ n18058 ;
  assign n39913 = ( n24208 & n28426 ) | ( n24208 & ~n38150 ) | ( n28426 & ~n38150 ) ;
  assign n39914 = ~n6577 & n8312 ;
  assign n39915 = n39914 ^ n1365 ^ 1'b0 ;
  assign n39916 = n17672 & ~n39915 ;
  assign n39917 = n17887 | n39916 ;
  assign n39918 = n9309 & ~n29404 ;
  assign n39919 = n17343 & n39918 ;
  assign n39920 = ~n9925 & n39741 ;
  assign n39921 = n33604 & n39920 ;
  assign n39923 = ( n4759 & n5586 ) | ( n4759 & ~n5793 ) | ( n5586 & ~n5793 ) ;
  assign n39922 = n21138 & ~n31554 ;
  assign n39924 = n39923 ^ n39922 ^ 1'b0 ;
  assign n39925 = n9267 & ~n11024 ;
  assign n39926 = n39925 ^ n6249 ^ 1'b0 ;
  assign n39927 = n39924 & ~n39926 ;
  assign n39928 = n27747 ^ n21446 ^ 1'b0 ;
  assign n39929 = ( ~n16284 & n21767 ) | ( ~n16284 & n39928 ) | ( n21767 & n39928 ) ;
  assign n39930 = n33013 ^ n11959 ^ 1'b0 ;
  assign n39931 = n3797 | n39930 ;
  assign n39932 = n34236 ^ n8029 ^ 1'b0 ;
  assign n39933 = ~n12167 & n13846 ;
  assign n39934 = n39933 ^ n32756 ^ 1'b0 ;
  assign n39935 = n34104 ^ n4832 ^ 1'b0 ;
  assign n39936 = n28463 ^ n2350 ^ n622 ;
  assign n39937 = n39936 ^ n14051 ^ 1'b0 ;
  assign n39938 = ~n19868 & n39937 ;
  assign n39940 = n27331 ^ n12625 ^ 1'b0 ;
  assign n39941 = ~n33732 & n39940 ;
  assign n39939 = n898 | n11580 ;
  assign n39942 = n39941 ^ n39939 ^ n10273 ;
  assign n39943 = n39942 ^ n23490 ^ 1'b0 ;
  assign n39944 = n5979 & n39925 ;
  assign n39945 = n21592 | n39776 ;
  assign n39946 = ( n4089 & ~n33563 ) | ( n4089 & n33575 ) | ( ~n33563 & n33575 ) ;
  assign n39947 = n7569 & n10172 ;
  assign n39948 = n1362 & n1975 ;
  assign n39949 = n39948 ^ n15479 ^ n5246 ;
  assign n39950 = n39949 ^ n29473 ^ 1'b0 ;
  assign n39951 = ~n39947 & n39950 ;
  assign n39952 = ( n1500 & n14974 ) | ( n1500 & ~n21965 ) | ( n14974 & ~n21965 ) ;
  assign n39953 = n19367 & ~n39952 ;
  assign n39954 = n39953 ^ n39622 ^ 1'b0 ;
  assign n39955 = n14502 & n21635 ;
  assign n39956 = n39955 ^ n2682 ^ 1'b0 ;
  assign n39957 = n21716 ^ n18731 ^ n15168 ;
  assign n39958 = n39957 ^ n17461 ^ n1382 ;
  assign n39959 = n28206 ^ n12836 ^ n7954 ;
  assign n39960 = n39959 ^ n26997 ^ 1'b0 ;
  assign n39961 = n7072 & n9848 ;
  assign n39962 = n6645 ^ n1189 ^ 1'b0 ;
  assign n39963 = n39961 & ~n39962 ;
  assign n39964 = n38608 | n39963 ;
  assign n39965 = n8264 & ~n10775 ;
  assign n39966 = ~n20082 & n32448 ;
  assign n39967 = ~n24489 & n39966 ;
  assign n39970 = n5804 & ~n7310 ;
  assign n39968 = n5134 & ~n13357 ;
  assign n39969 = ~n21759 & n39968 ;
  assign n39971 = n39970 ^ n39969 ^ 1'b0 ;
  assign n39972 = n39971 ^ n7113 ^ 1'b0 ;
  assign n39973 = n2162 | n37399 ;
  assign n39974 = n8417 & ~n39973 ;
  assign n39975 = n6084 & n26544 ;
  assign n39976 = n39975 ^ x147 ^ 1'b0 ;
  assign n39977 = ( n1091 & ~n3195 ) | ( n1091 & n4179 ) | ( ~n3195 & n4179 ) ;
  assign n39978 = ~n30916 & n39977 ;
  assign n39979 = ~n18716 & n39978 ;
  assign n39980 = n39979 ^ n30365 ^ 1'b0 ;
  assign n39981 = n39980 ^ n35907 ^ 1'b0 ;
  assign n39982 = ~n13046 & n39981 ;
  assign n39983 = n1742 & n6156 ;
  assign n39984 = n34738 ^ n22019 ^ n4932 ;
  assign n39985 = n2085 ^ n1869 ^ 1'b0 ;
  assign n39986 = ( n39983 & n39984 ) | ( n39983 & ~n39985 ) | ( n39984 & ~n39985 ) ;
  assign n39987 = ~n6969 & n9656 ;
  assign n39988 = n39987 ^ n15246 ^ 1'b0 ;
  assign n39989 = ~n20429 & n26280 ;
  assign n39990 = n39989 ^ n39108 ^ 1'b0 ;
  assign n39991 = n7487 ^ n1297 ^ 1'b0 ;
  assign n39992 = n30353 & ~n35177 ;
  assign n39993 = ~n1946 & n39992 ;
  assign n39994 = ~n39991 & n39993 ;
  assign n39995 = n5635 & ~n21381 ;
  assign n39996 = n27546 ^ n7014 ^ n6781 ;
  assign n39997 = n2921 | n39996 ;
  assign n39998 = ~n7464 & n14625 ;
  assign n39999 = n7027 & n39998 ;
  assign n40000 = ( n8707 & ~n36199 ) | ( n8707 & n39999 ) | ( ~n36199 & n39999 ) ;
  assign n40001 = ~n20137 & n20225 ;
  assign n40002 = n8039 & n40001 ;
  assign n40003 = n1296 & n12018 ;
  assign n40004 = n40002 & n40003 ;
  assign n40005 = n5858 & n11949 ;
  assign n40006 = n13041 & n40005 ;
  assign n40007 = n526 & n1547 ;
  assign n40008 = n40007 ^ n32838 ^ 1'b0 ;
  assign n40009 = ~n30456 & n40008 ;
  assign n40010 = n38093 ^ n5009 ^ 1'b0 ;
  assign n40011 = n38527 & ~n40010 ;
  assign n40012 = n1151 & n1993 ;
  assign n40013 = n31517 ^ n5667 ^ 1'b0 ;
  assign n40014 = n40012 & ~n40013 ;
  assign n40015 = n39630 | n40014 ;
  assign n40016 = n33667 ^ n6242 ^ 1'b0 ;
  assign n40017 = n4471 & n5850 ;
  assign n40018 = n18937 & ~n28363 ;
  assign n40019 = ~n40017 & n40018 ;
  assign n40020 = ( n5766 & n35264 ) | ( n5766 & n40019 ) | ( n35264 & n40019 ) ;
  assign n40021 = n1536 & n6888 ;
  assign n40022 = n40021 ^ n25847 ^ n7918 ;
  assign n40023 = n40022 ^ n2804 ^ 1'b0 ;
  assign n40024 = n2080 & ~n40023 ;
  assign n40025 = ( ~n9977 & n13937 ) | ( ~n9977 & n40024 ) | ( n13937 & n40024 ) ;
  assign n40026 = ~n19568 & n26005 ;
  assign n40027 = n40026 ^ n7781 ^ 1'b0 ;
  assign n40028 = n40027 ^ n27580 ^ 1'b0 ;
  assign n40029 = n22647 ^ n16665 ^ n7769 ;
  assign n40030 = n17771 ^ n8038 ^ 1'b0 ;
  assign n40031 = n40029 | n40030 ;
  assign n40032 = n33342 ^ n29038 ^ 1'b0 ;
  assign n40033 = n12238 | n21508 ;
  assign n40034 = n23739 & ~n40033 ;
  assign n40035 = n6361 & ~n40034 ;
  assign n40036 = n40035 ^ n4145 ^ 1'b0 ;
  assign n40037 = n3557 & ~n10598 ;
  assign n40038 = n3241 & n40037 ;
  assign n40039 = n40038 ^ n15141 ^ n7475 ;
  assign n40040 = n14507 ^ n4990 ^ 1'b0 ;
  assign n40041 = n39769 ^ n33101 ^ n3723 ;
  assign n40042 = n7026 ^ n1655 ^ 1'b0 ;
  assign n40043 = n5668 & n37634 ;
  assign n40044 = ~n683 & n10352 ;
  assign n40045 = ~n24510 & n36590 ;
  assign n40046 = n40044 & n40045 ;
  assign n40047 = n3590 | n7881 ;
  assign n40048 = n14454 ^ n2274 ^ n646 ;
  assign n40049 = n40048 ^ n29136 ^ n9172 ;
  assign n40052 = n32438 ^ n2402 ^ 1'b0 ;
  assign n40050 = n6268 ^ n804 ^ 1'b0 ;
  assign n40051 = ( n10655 & ~n37961 ) | ( n10655 & n40050 ) | ( ~n37961 & n40050 ) ;
  assign n40053 = n40052 ^ n40051 ^ n21531 ;
  assign n40054 = n36349 ^ n9501 ^ n4077 ;
  assign n40058 = n13729 ^ n5994 ^ 1'b0 ;
  assign n40059 = n28259 & n40058 ;
  assign n40055 = n4231 | n30274 ;
  assign n40056 = n2592 & ~n8393 ;
  assign n40057 = n40055 & n40056 ;
  assign n40060 = n40059 ^ n40057 ^ 1'b0 ;
  assign n40061 = ( x220 & ~n6528 ) | ( x220 & n10354 ) | ( ~n6528 & n10354 ) ;
  assign n40062 = n37284 | n40061 ;
  assign n40063 = n25029 & ~n40062 ;
  assign n40064 = n21271 ^ n4010 ^ 1'b0 ;
  assign n40065 = n5298 & ~n18339 ;
  assign n40066 = n34871 ^ n7303 ^ 1'b0 ;
  assign n40067 = ~n4167 & n40066 ;
  assign n40068 = n1783 & n17006 ;
  assign n40069 = n26477 | n38544 ;
  assign n40070 = n40069 ^ n17903 ^ 1'b0 ;
  assign n40071 = n19322 ^ n17654 ^ n2345 ;
  assign n40072 = n31061 & n40071 ;
  assign n40073 = n40072 ^ n19056 ^ 1'b0 ;
  assign n40074 = ~n19687 & n25274 ;
  assign n40075 = n40074 ^ n19261 ^ 1'b0 ;
  assign n40076 = n40075 ^ n20527 ^ n12059 ;
  assign n40077 = ( n18193 & ~n40073 ) | ( n18193 & n40076 ) | ( ~n40073 & n40076 ) ;
  assign n40078 = n12698 ^ n2471 ^ 1'b0 ;
  assign n40079 = n15378 | n40078 ;
  assign n40080 = n40079 ^ n9531 ^ 1'b0 ;
  assign n40081 = n37617 ^ n7244 ^ n751 ;
  assign n40082 = n5836 & n16919 ;
  assign n40083 = n11734 ^ n4129 ^ 1'b0 ;
  assign n40084 = n4077 & n40083 ;
  assign n40085 = ~n14873 & n40084 ;
  assign n40086 = n21487 ^ n9117 ^ 1'b0 ;
  assign n40087 = n4661 | n29481 ;
  assign n40088 = n40087 ^ n28473 ^ 1'b0 ;
  assign n40089 = n18948 | n30247 ;
  assign n40090 = ( ~n9856 & n14894 ) | ( ~n9856 & n33942 ) | ( n14894 & n33942 ) ;
  assign n40091 = n40090 ^ n19773 ^ 1'b0 ;
  assign n40092 = n40091 ^ n20011 ^ 1'b0 ;
  assign n40093 = n4073 & n40092 ;
  assign n40094 = n8946 | n12685 ;
  assign n40095 = n40094 ^ n4422 ^ n634 ;
  assign n40096 = n16502 ^ n7731 ^ 1'b0 ;
  assign n40097 = ( n2552 & n20362 ) | ( n2552 & ~n40096 ) | ( n20362 & ~n40096 ) ;
  assign n40098 = n17678 ^ n8125 ^ n6804 ;
  assign n40099 = n33374 ^ n24156 ^ n22434 ;
  assign n40100 = n37157 & ~n40099 ;
  assign n40101 = n14059 ^ n9561 ^ 1'b0 ;
  assign n40102 = n15360 & ~n40101 ;
  assign n40103 = ~n13733 & n30072 ;
  assign n40104 = n15188 & n40103 ;
  assign n40105 = n19047 | n40104 ;
  assign n40106 = n34098 & ~n40105 ;
  assign n40109 = n19659 ^ n3731 ^ 1'b0 ;
  assign n40110 = ( n8316 & n22780 ) | ( n8316 & n40109 ) | ( n22780 & n40109 ) ;
  assign n40107 = n3874 & n8587 ;
  assign n40108 = n40107 ^ n5927 ^ 1'b0 ;
  assign n40111 = n40110 ^ n40108 ^ n28585 ;
  assign n40112 = n16159 ^ x247 ^ 1'b0 ;
  assign n40113 = n17958 & n24584 ;
  assign n40114 = n27952 & ~n40113 ;
  assign n40115 = n11587 ^ n11317 ^ 1'b0 ;
  assign n40116 = n23110 & n40115 ;
  assign n40117 = n40116 ^ n33007 ^ 1'b0 ;
  assign n40118 = n292 | n21096 ;
  assign n40119 = n32202 | n40118 ;
  assign n40120 = n19849 ^ n1727 ^ 1'b0 ;
  assign n40121 = n40120 ^ n6917 ^ 1'b0 ;
  assign n40122 = n34204 & n36727 ;
  assign n40123 = n40121 & n40122 ;
  assign n40124 = n1840 | n2127 ;
  assign n40125 = n14660 ^ n1574 ^ 1'b0 ;
  assign n40126 = n40115 & n40125 ;
  assign n40127 = n40126 ^ n17558 ^ n10992 ;
  assign n40128 = n26504 ^ n21515 ^ 1'b0 ;
  assign n40129 = ~n3979 & n7415 ;
  assign n40130 = n40129 ^ n2829 ^ 1'b0 ;
  assign n40131 = n12693 | n40130 ;
  assign n40132 = n31926 | n40131 ;
  assign n40133 = n4943 & n24380 ;
  assign n40134 = n40133 ^ n1433 ^ 1'b0 ;
  assign n40135 = ( n944 & n17296 ) | ( n944 & ~n30156 ) | ( n17296 & ~n30156 ) ;
  assign n40136 = n40135 ^ n11932 ^ 1'b0 ;
  assign n40137 = n40134 & n40136 ;
  assign n40138 = n8839 & ~n21733 ;
  assign n40139 = n40138 ^ n18081 ^ 1'b0 ;
  assign n40140 = ~n11402 & n28739 ;
  assign n40141 = n40140 ^ n24967 ^ 1'b0 ;
  assign n40142 = n917 & ~n8915 ;
  assign n40143 = n40142 ^ n17270 ^ 1'b0 ;
  assign n40144 = n40141 | n40143 ;
  assign n40145 = x110 & ~n9594 ;
  assign n40146 = n8370 & n40145 ;
  assign n40147 = n12850 ^ n2078 ^ 1'b0 ;
  assign n40148 = ~n40146 & n40147 ;
  assign n40149 = n15696 & ~n40148 ;
  assign n40150 = n40149 ^ n26328 ^ n22781 ;
  assign n40151 = n21455 ^ n4205 ^ 1'b0 ;
  assign n40152 = n40151 ^ n25203 ^ 1'b0 ;
  assign n40153 = ~n6074 & n21128 ;
  assign n40154 = n24081 ^ n17572 ^ 1'b0 ;
  assign n40155 = ( n27684 & n40153 ) | ( n27684 & n40154 ) | ( n40153 & n40154 ) ;
  assign n40156 = n40155 ^ n36813 ^ 1'b0 ;
  assign n40157 = ~n35623 & n36945 ;
  assign n40158 = ~n14003 & n40157 ;
  assign n40159 = n17699 ^ n9693 ^ n8942 ;
  assign n40160 = n30072 & n40159 ;
  assign n40161 = n9435 | n40160 ;
  assign n40162 = n30865 ^ n22698 ^ 1'b0 ;
  assign n40163 = n40161 | n40162 ;
  assign n40164 = ~n1865 & n11426 ;
  assign n40165 = n29557 & n40164 ;
  assign n40166 = n12265 & n19706 ;
  assign n40167 = n40166 ^ n840 ^ 1'b0 ;
  assign n40168 = ~n9051 & n13416 ;
  assign n40169 = n35997 ^ n1957 ^ 1'b0 ;
  assign n40170 = n34310 & n40169 ;
  assign n40171 = n24468 | n40170 ;
  assign n40172 = ( n13889 & ~n22733 ) | ( n13889 & n35823 ) | ( ~n22733 & n35823 ) ;
  assign n40173 = n6968 & ~n18926 ;
  assign n40174 = ~n10257 & n40173 ;
  assign n40175 = n40174 ^ n35612 ^ 1'b0 ;
  assign n40176 = n33736 ^ n3174 ^ 1'b0 ;
  assign n40177 = n10917 ^ n1313 ^ 1'b0 ;
  assign n40178 = n40177 ^ n10973 ^ 1'b0 ;
  assign n40179 = n30587 ^ n14780 ^ 1'b0 ;
  assign n40180 = n9151 & ~n40179 ;
  assign n40181 = n40180 ^ n1920 ^ 1'b0 ;
  assign n40182 = n17309 ^ n10614 ^ 1'b0 ;
  assign n40183 = ( ~x35 & n4180 ) | ( ~x35 & n15119 ) | ( n4180 & n15119 ) ;
  assign n40184 = ~n30267 & n40183 ;
  assign n40185 = ~n40182 & n40184 ;
  assign n40187 = n27653 ^ n9636 ^ 1'b0 ;
  assign n40186 = n5689 & ~n33296 ;
  assign n40188 = n40187 ^ n40186 ^ 1'b0 ;
  assign n40189 = n11963 | n13464 ;
  assign n40190 = n5991 & ~n35217 ;
  assign n40191 = n16124 & n22175 ;
  assign n40192 = ( ~n1571 & n10532 ) | ( ~n1571 & n40191 ) | ( n10532 & n40191 ) ;
  assign n40193 = ( n7473 & n11686 ) | ( n7473 & n17856 ) | ( n11686 & n17856 ) ;
  assign n40194 = n15962 & ~n40193 ;
  assign n40195 = ~n29923 & n34871 ;
  assign n40196 = ( n5610 & n7364 ) | ( n5610 & ~n10855 ) | ( n7364 & ~n10855 ) ;
  assign n40197 = n6998 ^ n2250 ^ x3 ;
  assign n40198 = ( n17045 & n24685 ) | ( n17045 & n33415 ) | ( n24685 & n33415 ) ;
  assign n40199 = n40198 ^ n18832 ^ 1'b0 ;
  assign n40200 = ~n3107 & n40199 ;
  assign n40201 = n35677 ^ n15608 ^ 1'b0 ;
  assign n40202 = ( n40197 & n40200 ) | ( n40197 & ~n40201 ) | ( n40200 & ~n40201 ) ;
  assign n40203 = n28124 ^ n10562 ^ 1'b0 ;
  assign n40204 = ~n20185 & n40203 ;
  assign n40205 = n9217 & ~n36238 ;
  assign n40206 = ~n12075 & n14815 ;
  assign n40207 = n40206 ^ n6727 ^ 1'b0 ;
  assign n40208 = n40207 ^ n2715 ^ 1'b0 ;
  assign n40209 = n13279 ^ n4789 ^ 1'b0 ;
  assign n40210 = n16879 & ~n18313 ;
  assign n40211 = n27222 & n40210 ;
  assign n40212 = n40211 ^ n1551 ^ 1'b0 ;
  assign n40213 = n2722 | n3330 ;
  assign n40214 = n15970 & ~n40213 ;
  assign n40215 = n40214 ^ n5175 ^ 1'b0 ;
  assign n40216 = n2684 | n40215 ;
  assign n40217 = ( n1472 & ~n5051 ) | ( n1472 & n40216 ) | ( ~n5051 & n40216 ) ;
  assign n40218 = n18315 | n40217 ;
  assign n40219 = n15829 & n40218 ;
  assign n40220 = ~n12647 & n32100 ;
  assign n40221 = n9707 & ~n35508 ;
  assign n40222 = n40220 & ~n40221 ;
  assign n40223 = n8301 ^ n5446 ^ 1'b0 ;
  assign n40224 = n6167 | n40223 ;
  assign n40225 = ~n6724 & n21291 ;
  assign n40226 = n40224 & n40225 ;
  assign n40227 = n23377 | n40226 ;
  assign n40228 = ~n345 & n5973 ;
  assign n40229 = n7426 & n8892 ;
  assign n40230 = ~n27413 & n40229 ;
  assign n40231 = n13117 | n40230 ;
  assign n40232 = n4245 | n40231 ;
  assign n40233 = ~n25269 & n29237 ;
  assign n40234 = n23161 & n40233 ;
  assign n40235 = n40234 ^ n26911 ^ 1'b0 ;
  assign n40236 = n12638 & ~n40235 ;
  assign n40237 = ( n7261 & n13397 ) | ( n7261 & ~n34019 ) | ( n13397 & ~n34019 ) ;
  assign n40238 = ( n23912 & ~n26867 ) | ( n23912 & n35212 ) | ( ~n26867 & n35212 ) ;
  assign n40239 = n592 | n5588 ;
  assign n40240 = n24271 & ~n40239 ;
  assign n40241 = ( n8715 & n15635 ) | ( n8715 & ~n18955 ) | ( n15635 & ~n18955 ) ;
  assign n40242 = n25360 & ~n40241 ;
  assign n40243 = ~n6291 & n32525 ;
  assign n40244 = n40243 ^ n40142 ^ 1'b0 ;
  assign n40245 = n9132 ^ x90 ^ 1'b0 ;
  assign n40246 = n27702 | n40245 ;
  assign n40247 = n13419 & n30015 ;
  assign n40252 = ( ~n15986 & n18411 ) | ( ~n15986 & n34849 ) | ( n18411 & n34849 ) ;
  assign n40248 = n7523 & n15569 ;
  assign n40249 = n40248 ^ n6829 ^ 1'b0 ;
  assign n40250 = ( n8634 & ~n17495 ) | ( n8634 & n40249 ) | ( ~n17495 & n40249 ) ;
  assign n40251 = n8564 | n40250 ;
  assign n40253 = n40252 ^ n40251 ^ 1'b0 ;
  assign n40254 = n40253 ^ n33347 ^ n24267 ;
  assign n40255 = n22828 ^ n3064 ^ 1'b0 ;
  assign n40256 = ~n12957 & n21993 ;
  assign n40257 = n21959 ^ n6101 ^ 1'b0 ;
  assign n40258 = ~n17614 & n25937 ;
  assign n40259 = n16427 & n40258 ;
  assign n40260 = ~n2518 & n26238 ;
  assign n40261 = n8632 & n40260 ;
  assign n40262 = n19832 ^ n4754 ^ 1'b0 ;
  assign n40263 = n2756 & n40262 ;
  assign n40264 = n40263 ^ n14205 ^ 1'b0 ;
  assign n40265 = ~n721 & n9373 ;
  assign n40266 = ~n26903 & n40265 ;
  assign n40267 = ( n24699 & n40264 ) | ( n24699 & n40266 ) | ( n40264 & n40266 ) ;
  assign n40268 = n31136 ^ n13676 ^ 1'b0 ;
  assign n40269 = ~n3201 & n6468 ;
  assign n40270 = n40269 ^ n37473 ^ 1'b0 ;
  assign n40271 = n10464 | n20669 ;
  assign n40272 = n16753 & ~n40271 ;
  assign n40273 = n13268 | n26156 ;
  assign n40274 = n40273 ^ n19019 ^ 1'b0 ;
  assign n40275 = n12908 & ~n40274 ;
  assign n40276 = ~n33617 & n40275 ;
  assign n40277 = n647 | n15699 ;
  assign n40278 = n40277 ^ n17302 ^ 1'b0 ;
  assign n40279 = ( n4177 & n20307 ) | ( n4177 & n34999 ) | ( n20307 & n34999 ) ;
  assign n40280 = n11933 & ~n28591 ;
  assign n40281 = ( n25865 & n37545 ) | ( n25865 & n40280 ) | ( n37545 & n40280 ) ;
  assign n40282 = n33320 ^ n29252 ^ 1'b0 ;
  assign n40283 = n18449 ^ n5313 ^ 1'b0 ;
  assign n40284 = n12934 & n40283 ;
  assign n40285 = n982 & n40284 ;
  assign n40286 = n2627 ^ x70 ^ 1'b0 ;
  assign n40287 = ~n19275 & n40286 ;
  assign n40288 = n24428 | n40287 ;
  assign n40289 = n33118 ^ n22635 ^ 1'b0 ;
  assign n40290 = n11174 & n18832 ;
  assign n40291 = n11882 & ~n21390 ;
  assign n40292 = n39642 & n40291 ;
  assign n40293 = n19272 ^ x159 ^ 1'b0 ;
  assign n40294 = ( ~n4858 & n12793 ) | ( ~n4858 & n25390 ) | ( n12793 & n25390 ) ;
  assign n40295 = n40294 ^ n9322 ^ 1'b0 ;
  assign n40296 = ( ~n13610 & n21165 ) | ( ~n13610 & n25811 ) | ( n21165 & n25811 ) ;
  assign n40297 = n5210 | n8512 ;
  assign n40298 = n1579 & n38001 ;
  assign n40299 = n14338 & ~n17921 ;
  assign n40300 = ~n40298 & n40299 ;
  assign n40301 = n12048 ^ n1232 ^ 1'b0 ;
  assign n40302 = n27098 ^ n23773 ^ 1'b0 ;
  assign n40303 = n13568 | n14663 ;
  assign n40304 = n40303 ^ n15696 ^ 1'b0 ;
  assign n40305 = ( n25434 & n27085 ) | ( n25434 & ~n35002 ) | ( n27085 & ~n35002 ) ;
  assign n40306 = ( n374 & ~n4573 ) | ( n374 & n29879 ) | ( ~n4573 & n29879 ) ;
  assign n40308 = n22083 ^ n5071 ^ 1'b0 ;
  assign n40309 = n5229 & n40308 ;
  assign n40307 = n32200 & n40056 ;
  assign n40310 = n40309 ^ n40307 ^ 1'b0 ;
  assign n40311 = n4948 & ~n8423 ;
  assign n40312 = ~n4542 & n40311 ;
  assign n40313 = n39137 ^ n27529 ^ 1'b0 ;
  assign n40314 = n34835 | n40313 ;
  assign n40315 = n2024 & ~n18420 ;
  assign n40316 = n40315 ^ n20199 ^ 1'b0 ;
  assign n40317 = n13517 ^ n1801 ^ 1'b0 ;
  assign n40318 = n1590 & n40317 ;
  assign n40319 = n40318 ^ n36111 ^ 1'b0 ;
  assign n40320 = ~n5866 & n16170 ;
  assign n40321 = ~n15463 & n40320 ;
  assign n40322 = n17442 ^ n7482 ^ 1'b0 ;
  assign n40323 = ~n40321 & n40322 ;
  assign n40324 = n2208 | n40323 ;
  assign n40325 = n3316 | n40324 ;
  assign n40326 = n27859 ^ n18425 ^ 1'b0 ;
  assign n40327 = ~n11722 & n40326 ;
  assign n40328 = n6945 | n17614 ;
  assign n40329 = n7497 ^ n4135 ^ 1'b0 ;
  assign n40330 = n4451 & n15226 ;
  assign n40331 = ~n6348 & n25197 ;
  assign n40332 = ( n444 & n31834 ) | ( n444 & ~n40331 ) | ( n31834 & ~n40331 ) ;
  assign n40333 = ~n5591 & n11149 ;
  assign n40334 = n13577 ^ n1010 ^ 1'b0 ;
  assign n40335 = n6641 & ~n40334 ;
  assign n40336 = n10779 | n40335 ;
  assign n40337 = n35866 ^ n27481 ^ 1'b0 ;
  assign n40338 = n7527 | n15833 ;
  assign n40339 = n16290 | n40338 ;
  assign n40340 = n2712 ^ n1440 ^ 1'b0 ;
  assign n40341 = n15350 | n40340 ;
  assign n40342 = n40341 ^ n2053 ^ 1'b0 ;
  assign n40343 = n40339 & ~n40342 ;
  assign n40344 = n12004 | n29947 ;
  assign n40345 = n28776 ^ n24258 ^ n15749 ;
  assign n40346 = n7118 ^ n2114 ^ 1'b0 ;
  assign n40347 = n12882 ^ n12797 ^ n791 ;
  assign n40348 = n40347 ^ n11443 ^ 1'b0 ;
  assign n40349 = n8215 & ~n40348 ;
  assign n40350 = n3445 & n40349 ;
  assign n40351 = n40350 ^ n12574 ^ 1'b0 ;
  assign n40352 = n5738 | n12648 ;
  assign n40353 = ~n26396 & n40352 ;
  assign n40354 = n27222 & n40353 ;
  assign n40355 = n40354 ^ n18776 ^ 1'b0 ;
  assign n40356 = n12105 | n32543 ;
  assign n40357 = n13419 & ~n16943 ;
  assign n40358 = n40357 ^ n12856 ^ 1'b0 ;
  assign n40359 = n10940 | n40358 ;
  assign n40360 = n40359 ^ n7124 ^ 1'b0 ;
  assign n40361 = ~n5857 & n6009 ;
  assign n40362 = ~n39589 & n40361 ;
  assign n40363 = n10537 ^ n9993 ^ n9708 ;
  assign n40364 = ( n5051 & n10919 ) | ( n5051 & n40363 ) | ( n10919 & n40363 ) ;
  assign n40365 = n28231 & n40364 ;
  assign n40366 = n376 | n13363 ;
  assign n40367 = n40366 ^ n28893 ^ n21016 ;
  assign n40368 = n5303 & n14742 ;
  assign n40369 = n40368 ^ n16168 ^ n387 ;
  assign n40370 = ~n6114 & n23479 ;
  assign n40371 = n32878 | n40370 ;
  assign n40372 = ~n9750 & n10143 ;
  assign n40373 = ~n39114 & n40372 ;
  assign n40374 = n15717 & n40373 ;
  assign n40375 = ~n1475 & n3747 ;
  assign n40376 = ~n12906 & n40375 ;
  assign n40377 = n5491 & n38151 ;
  assign n40378 = n40376 & n40377 ;
  assign n40379 = ( ~x36 & n13760 ) | ( ~x36 & n19612 ) | ( n13760 & n19612 ) ;
  assign n40380 = n39424 ^ n17573 ^ n12226 ;
  assign n40381 = n23698 | n30097 ;
  assign n40382 = n4613 & ~n40381 ;
  assign n40383 = n3712 | n40382 ;
  assign n40385 = n10750 & ~n16798 ;
  assign n40386 = n30562 & n40385 ;
  assign n40384 = n3118 & ~n11141 ;
  assign n40387 = n40386 ^ n40384 ^ 1'b0 ;
  assign n40391 = ~n572 & n20004 ;
  assign n40389 = n4182 & ~n39247 ;
  assign n40390 = n40389 ^ n12522 ^ 1'b0 ;
  assign n40388 = n2380 & ~n21569 ;
  assign n40392 = n40391 ^ n40390 ^ n40388 ;
  assign n40393 = n20563 ^ n6388 ^ 1'b0 ;
  assign n40394 = n40393 ^ n13641 ^ n10166 ;
  assign n40395 = n20909 ^ n14429 ^ n11394 ;
  assign n40396 = n40395 ^ n1358 ^ 1'b0 ;
  assign n40397 = n40396 ^ n22503 ^ n7756 ;
  assign n40398 = n27242 & n40397 ;
  assign n40399 = n17154 & n40398 ;
  assign n40400 = n10234 & n13000 ;
  assign n40401 = n2444 ^ n275 ^ 1'b0 ;
  assign n40402 = ~n23632 & n40401 ;
  assign n40403 = n34037 ^ n22933 ^ n14598 ;
  assign n40404 = n14569 & ~n40403 ;
  assign n40405 = n40404 ^ n19285 ^ 1'b0 ;
  assign n40407 = n12808 ^ n11227 ^ 1'b0 ;
  assign n40406 = n12059 & n13573 ;
  assign n40408 = n40407 ^ n40406 ^ 1'b0 ;
  assign n40409 = n9874 & n22756 ;
  assign n40410 = n40409 ^ n20042 ^ 1'b0 ;
  assign n40411 = ( n9469 & n10870 ) | ( n9469 & ~n40410 ) | ( n10870 & ~n40410 ) ;
  assign n40412 = n1731 & n21095 ;
  assign n40413 = ~n13164 & n30709 ;
  assign n40414 = n1651 & ~n21508 ;
  assign n40415 = n14020 & n40414 ;
  assign n40416 = n14619 | n21098 ;
  assign n40417 = n15234 | n40416 ;
  assign n40418 = n33446 ^ n8329 ^ 1'b0 ;
  assign n40419 = n3504 & n5538 ;
  assign n40420 = n38695 & n40419 ;
  assign n40421 = n40420 ^ n33822 ^ n27451 ;
  assign n40422 = ( n23612 & ~n36187 ) | ( n23612 & n40421 ) | ( ~n36187 & n40421 ) ;
  assign n40423 = n36780 ^ n1403 ^ 1'b0 ;
  assign n40424 = n5650 & ~n40423 ;
  assign n40425 = n40424 ^ n32183 ^ n13495 ;
  assign n40426 = n19623 & ~n36748 ;
  assign n40427 = n38798 ^ n4375 ^ 1'b0 ;
  assign n40428 = n10818 & n40427 ;
  assign n40429 = n40428 ^ n6467 ^ 1'b0 ;
  assign n40432 = n22692 ^ n374 ^ 1'b0 ;
  assign n40430 = n6063 & n13281 ;
  assign n40431 = n4995 & ~n40430 ;
  assign n40433 = n40432 ^ n40431 ^ 1'b0 ;
  assign n40434 = ( n4052 & ~n15551 ) | ( n4052 & n37393 ) | ( ~n15551 & n37393 ) ;
  assign n40435 = x34 & ~n7130 ;
  assign n40436 = n8231 & ~n35292 ;
  assign n40437 = ( n16925 & n40435 ) | ( n16925 & ~n40436 ) | ( n40435 & ~n40436 ) ;
  assign n40438 = n27495 & ~n36511 ;
  assign n40439 = n40438 ^ n6360 ^ 1'b0 ;
  assign n40440 = ( ~n11661 & n18005 ) | ( ~n11661 & n32674 ) | ( n18005 & n32674 ) ;
  assign n40441 = n492 | n15618 ;
  assign n40442 = n2376 & ~n40441 ;
  assign n40443 = n40442 ^ n5099 ^ 1'b0 ;
  assign n40444 = n40440 | n40443 ;
  assign n40445 = n7145 & ~n33382 ;
  assign n40446 = ~n6964 & n40445 ;
  assign n40447 = n16517 ^ n12950 ^ 1'b0 ;
  assign n40448 = ( ~n8148 & n18121 ) | ( ~n8148 & n33370 ) | ( n18121 & n33370 ) ;
  assign n40449 = n10387 & ~n21743 ;
  assign n40450 = n9355 & n40449 ;
  assign n40451 = n3627 ^ n3230 ^ 1'b0 ;
  assign n40452 = n4002 & ~n40451 ;
  assign n40453 = n40452 ^ n6912 ^ 1'b0 ;
  assign n40454 = ~n729 & n12338 ;
  assign n40455 = n40454 ^ n8719 ^ 1'b0 ;
  assign n40456 = ~n13048 & n15365 ;
  assign n40457 = n22989 & n40456 ;
  assign n40458 = n20516 ^ n19526 ^ n8984 ;
  assign n40459 = n31790 ^ n19554 ^ 1'b0 ;
  assign n40460 = n40458 & n40459 ;
  assign n40461 = n8924 | n24355 ;
  assign n40462 = n12625 ^ n12479 ^ 1'b0 ;
  assign n40463 = n24738 ^ n20533 ^ 1'b0 ;
  assign n40464 = n40462 | n40463 ;
  assign n40465 = n40464 ^ n30727 ^ n8194 ;
  assign n40466 = x21 & ~n31414 ;
  assign n40467 = n3951 | n10451 ;
  assign n40468 = n18555 & n20455 ;
  assign n40469 = n40468 ^ n677 ^ 1'b0 ;
  assign n40470 = n5644 ^ n1203 ^ 1'b0 ;
  assign n40471 = n40469 | n40470 ;
  assign n40472 = n25486 ^ n23436 ^ 1'b0 ;
  assign n40473 = n21873 | n40472 ;
  assign n40474 = n40473 ^ n15646 ^ 1'b0 ;
  assign n40475 = ( ~n7267 & n8893 ) | ( ~n7267 & n21343 ) | ( n8893 & n21343 ) ;
  assign n40476 = n40475 ^ n32499 ^ 1'b0 ;
  assign n40477 = n15276 & n40476 ;
  assign n40478 = ~n40474 & n40477 ;
  assign n40479 = n5264 | n9055 ;
  assign n40481 = ~n15179 & n19470 ;
  assign n40482 = n40481 ^ n6268 ^ 1'b0 ;
  assign n40483 = n983 | n40482 ;
  assign n40484 = n6193 | n40483 ;
  assign n40485 = n40484 ^ n21932 ^ 1'b0 ;
  assign n40480 = n17013 | n20637 ;
  assign n40486 = n40485 ^ n40480 ^ 1'b0 ;
  assign n40487 = n14390 & ~n27051 ;
  assign n40488 = n2573 ^ n2124 ^ 1'b0 ;
  assign n40489 = n35045 | n40488 ;
  assign n40490 = n40487 | n40489 ;
  assign n40491 = n7306 & ~n8756 ;
  assign n40492 = ~n23255 & n40491 ;
  assign n40493 = n40492 ^ n30922 ^ 1'b0 ;
  assign n40494 = n37732 ^ n7277 ^ n3922 ;
  assign n40495 = n9411 ^ x115 ^ 1'b0 ;
  assign n40496 = n12415 & n14581 ;
  assign n40497 = n27421 ^ n22911 ^ 1'b0 ;
  assign n40498 = n40497 ^ n15557 ^ n4015 ;
  assign n40499 = ~n11879 & n40498 ;
  assign n40500 = n40499 ^ n21873 ^ 1'b0 ;
  assign n40501 = n7653 & n27827 ;
  assign n40502 = n40501 ^ n7974 ^ 1'b0 ;
  assign n40503 = n22096 ^ n18311 ^ 1'b0 ;
  assign n40504 = n3728 & n12689 ;
  assign n40505 = n40504 ^ n34419 ^ 1'b0 ;
  assign n40506 = n21796 ^ n14278 ^ n8029 ;
  assign n40507 = n28272 | n40506 ;
  assign n40508 = n2991 | n3246 ;
  assign n40509 = n3246 & ~n40508 ;
  assign n40510 = n40509 ^ n1546 ^ 1'b0 ;
  assign n40511 = n17245 & ~n40510 ;
  assign n40512 = n40511 ^ n27469 ^ 1'b0 ;
  assign n40513 = n27065 ^ n650 ^ 1'b0 ;
  assign n40514 = n33647 & n40513 ;
  assign n40515 = ~n311 & n7431 ;
  assign n40516 = n30562 ^ n14566 ^ x217 ;
  assign n40517 = n5522 & n15270 ;
  assign n40518 = n40517 ^ n19272 ^ 1'b0 ;
  assign n40519 = n10939 | n29970 ;
  assign n40520 = n40518 & ~n40519 ;
  assign n40521 = n4812 | n5303 ;
  assign n40522 = ~n10329 & n25783 ;
  assign n40523 = n34384 ^ n15865 ^ n6683 ;
  assign n40524 = n11827 ^ n5731 ^ 1'b0 ;
  assign n40525 = n40523 & n40524 ;
  assign n40526 = n14229 & ~n34464 ;
  assign n40527 = n39227 & n40526 ;
  assign n40528 = n30824 ^ n18648 ^ 1'b0 ;
  assign n40529 = n11556 & ~n40528 ;
  assign n40530 = n40529 ^ n28099 ^ 1'b0 ;
  assign n40531 = n6720 & n40530 ;
  assign n40532 = n9977 | n18715 ;
  assign n40533 = n4027 & ~n40532 ;
  assign n40534 = n40533 ^ n34031 ^ 1'b0 ;
  assign n40535 = n1518 & n4858 ;
  assign n40536 = n23885 | n27959 ;
  assign n40537 = ~n7259 & n10886 ;
  assign n40538 = ( n24500 & n26213 ) | ( n24500 & n40537 ) | ( n26213 & n40537 ) ;
  assign n40539 = n40538 ^ n26089 ^ 1'b0 ;
  assign n40540 = n40539 ^ n25187 ^ n12704 ;
  assign n40541 = n40540 ^ n3064 ^ 1'b0 ;
  assign n40543 = ~n1409 & n4850 ;
  assign n40542 = n5329 & ~n19848 ;
  assign n40544 = n40543 ^ n40542 ^ 1'b0 ;
  assign n40545 = n12774 ^ n2689 ^ 1'b0 ;
  assign n40546 = ~n1935 & n35185 ;
  assign n40547 = ~n12557 & n17192 ;
  assign n40548 = n40547 ^ n14465 ^ 1'b0 ;
  assign n40549 = ( n4245 & ~n31882 ) | ( n4245 & n40548 ) | ( ~n31882 & n40548 ) ;
  assign n40550 = n11201 & ~n21196 ;
  assign n40551 = n1181 & ~n9057 ;
  assign n40552 = ~n28692 & n40551 ;
  assign n40553 = n1350 & ~n40552 ;
  assign n40554 = ~n16992 & n40553 ;
  assign n40555 = n3405 & ~n4207 ;
  assign n40556 = n8134 & n40555 ;
  assign n40557 = n11236 ^ n704 ^ 1'b0 ;
  assign n40558 = ( n3291 & n40556 ) | ( n3291 & n40557 ) | ( n40556 & n40557 ) ;
  assign n40559 = n5748 & ~n40558 ;
  assign n40560 = n8734 & n40559 ;
  assign n40561 = n11580 | n30622 ;
  assign n40562 = n5321 & ~n40561 ;
  assign n40563 = n17622 & n40562 ;
  assign n40564 = ( n1013 & n6910 ) | ( n1013 & n36520 ) | ( n6910 & n36520 ) ;
  assign n40565 = n13212 ^ n3348 ^ 1'b0 ;
  assign n40566 = n9502 & ~n40565 ;
  assign n40567 = n2132 & n32641 ;
  assign n40568 = n38828 ^ n2808 ^ 1'b0 ;
  assign n40569 = n37625 & ~n38021 ;
  assign n40570 = ~n33360 & n40569 ;
  assign n40571 = n20634 & ~n32626 ;
  assign n40572 = n28949 ^ n20022 ^ 1'b0 ;
  assign n40578 = n13780 & n23362 ;
  assign n40576 = ( ~n2970 & n8785 ) | ( ~n2970 & n37283 ) | ( n8785 & n37283 ) ;
  assign n40573 = n14928 & n26694 ;
  assign n40574 = ~n11125 & n40573 ;
  assign n40575 = n10946 & ~n40574 ;
  assign n40577 = n40576 ^ n40575 ^ 1'b0 ;
  assign n40579 = n40578 ^ n40577 ^ 1'b0 ;
  assign n40580 = n3648 & ~n10525 ;
  assign n40581 = n40580 ^ n21436 ^ 1'b0 ;
  assign n40582 = n7774 & ~n26001 ;
  assign n40583 = ~n19899 & n40582 ;
  assign n40584 = n40583 ^ n5741 ^ 1'b0 ;
  assign n40585 = n13742 | n40584 ;
  assign n40586 = n9134 | n40585 ;
  assign n40587 = n16767 & ~n40586 ;
  assign n40588 = n29859 ^ n5850 ^ 1'b0 ;
  assign n40589 = ~n40587 & n40588 ;
  assign n40590 = ( n2720 & ~n4526 ) | ( n2720 & n23368 ) | ( ~n4526 & n23368 ) ;
  assign n40591 = n20654 & ~n40590 ;
  assign n40592 = n40591 ^ n27951 ^ 1'b0 ;
  assign n40593 = ( n2522 & ~n10324 ) | ( n2522 & n14618 ) | ( ~n10324 & n14618 ) ;
  assign n40594 = n9546 & n40593 ;
  assign n40595 = n40592 & n40594 ;
  assign n40596 = ( ~n3917 & n10879 ) | ( ~n3917 & n32257 ) | ( n10879 & n32257 ) ;
  assign n40597 = ( n9545 & ~n12228 ) | ( n9545 & n27309 ) | ( ~n12228 & n27309 ) ;
  assign n40598 = n6589 | n19803 ;
  assign n40599 = n38855 & ~n40598 ;
  assign n40600 = n40599 ^ n7785 ^ 1'b0 ;
  assign n40601 = n26541 | n40600 ;
  assign n40602 = n25944 & ~n29471 ;
  assign n40603 = n40602 ^ n33331 ^ 1'b0 ;
  assign n40604 = n1508 & n24183 ;
  assign n40605 = n40604 ^ n11620 ^ 1'b0 ;
  assign n40606 = n2810 | n40605 ;
  assign n40607 = n40603 & ~n40606 ;
  assign n40608 = n11231 & n16096 ;
  assign n40609 = n40608 ^ n10906 ^ 1'b0 ;
  assign n40610 = n14870 & n40609 ;
  assign n40611 = n18324 & ~n19486 ;
  assign n40612 = ~n18645 & n40611 ;
  assign n40613 = n9366 & n9644 ;
  assign n40614 = n40613 ^ n17011 ^ 1'b0 ;
  assign n40615 = n2135 ^ x254 ^ 1'b0 ;
  assign n40616 = ( n930 & n2291 ) | ( n930 & ~n6968 ) | ( n2291 & ~n6968 ) ;
  assign n40617 = n40616 ^ n36023 ^ n840 ;
  assign n40618 = n40533 ^ n14814 ^ 1'b0 ;
  assign n40619 = n1147 ^ n959 ^ 1'b0 ;
  assign n40621 = n1228 | n2789 ;
  assign n40620 = n1239 & n25517 ;
  assign n40622 = n40621 ^ n40620 ^ 1'b0 ;
  assign n40623 = n40622 ^ n16983 ^ 1'b0 ;
  assign n40624 = n39705 | n40623 ;
  assign n40625 = n6414 | n40624 ;
  assign n40626 = n7923 & n21880 ;
  assign n40627 = n20424 ^ n16427 ^ n7372 ;
  assign n40628 = ( n16733 & n26703 ) | ( n16733 & ~n40627 ) | ( n26703 & ~n40627 ) ;
  assign n40629 = n20289 ^ n18095 ^ 1'b0 ;
  assign n40630 = n40629 ^ n37279 ^ n19673 ;
  assign n40631 = n21888 ^ n10636 ^ 1'b0 ;
  assign n40632 = n6159 | n25768 ;
  assign n40633 = n40632 ^ n5453 ^ 1'b0 ;
  assign n40634 = ~n417 & n27591 ;
  assign n40635 = n40634 ^ n16452 ^ 1'b0 ;
  assign n40636 = n10862 ^ n6309 ^ 1'b0 ;
  assign n40637 = n40636 ^ n12415 ^ n2774 ;
  assign n40638 = n28555 & n40637 ;
  assign n40640 = n3251 & ~n4815 ;
  assign n40639 = n40318 ^ n22126 ^ 1'b0 ;
  assign n40641 = n40640 ^ n40639 ^ n31773 ;
  assign n40642 = n15462 ^ n12350 ^ 1'b0 ;
  assign n40643 = n29046 ^ n26800 ^ n22901 ;
  assign n40644 = n14505 | n22046 ;
  assign n40645 = n38877 | n40644 ;
  assign n40646 = n1152 | n24268 ;
  assign n40647 = n40645 | n40646 ;
  assign n40648 = n6111 | n6745 ;
  assign n40649 = n40648 ^ n36085 ^ 1'b0 ;
  assign n40650 = n735 | n1587 ;
  assign n40651 = ~n10138 & n40650 ;
  assign n40652 = ~n40649 & n40651 ;
  assign n40657 = ( n2728 & ~n9913 ) | ( n2728 & n27219 ) | ( ~n9913 & n27219 ) ;
  assign n40653 = n3449 | n6873 ;
  assign n40654 = n40653 ^ n8231 ^ 1'b0 ;
  assign n40655 = ( ~n1443 & n6520 ) | ( ~n1443 & n6877 ) | ( n6520 & n6877 ) ;
  assign n40656 = n40654 & ~n40655 ;
  assign n40658 = n40657 ^ n40656 ^ 1'b0 ;
  assign n40659 = ~n12579 & n16766 ;
  assign n40660 = n40659 ^ n10626 ^ 1'b0 ;
  assign n40661 = n13826 ^ n8318 ^ n7632 ;
  assign n40662 = n24489 | n40661 ;
  assign n40663 = n5042 ^ n1882 ^ 1'b0 ;
  assign n40664 = n6085 & n8309 ;
  assign n40665 = ~n8309 & n40664 ;
  assign n40666 = n11242 | n40665 ;
  assign n40667 = n40666 ^ n18587 ^ 1'b0 ;
  assign n40668 = n14246 ^ n10940 ^ 1'b0 ;
  assign n40669 = ~n18697 & n40668 ;
  assign n40670 = n14161 & n40669 ;
  assign n40671 = n40670 ^ n16715 ^ 1'b0 ;
  assign n40672 = ~n14133 & n25459 ;
  assign n40673 = n40672 ^ n12758 ^ 1'b0 ;
  assign n40674 = n2226 & ~n40673 ;
  assign n40675 = ~n15869 & n40674 ;
  assign n40676 = n9810 ^ n4462 ^ 1'b0 ;
  assign n40677 = n19756 & n40676 ;
  assign n40678 = n16612 & n40677 ;
  assign n40679 = n40678 ^ n40154 ^ 1'b0 ;
  assign n40682 = n11724 & n23866 ;
  assign n40683 = n21240 ^ n14254 ^ 1'b0 ;
  assign n40684 = n40682 & ~n40683 ;
  assign n40680 = n5281 | n19298 ;
  assign n40681 = n15987 & n40680 ;
  assign n40685 = n40684 ^ n40681 ^ 1'b0 ;
  assign n40686 = ~n4627 & n10164 ;
  assign n40687 = n8556 & n39295 ;
  assign n40688 = ~n40686 & n40687 ;
  assign n40689 = ~n3404 & n20695 ;
  assign n40690 = n40689 ^ n10560 ^ 1'b0 ;
  assign n40691 = n25778 & n40690 ;
  assign n40692 = ( n9600 & n24441 ) | ( n9600 & ~n38559 ) | ( n24441 & ~n38559 ) ;
  assign n40693 = n22630 ^ n13262 ^ n6725 ;
  assign n40694 = n13598 | n16451 ;
  assign n40695 = n40694 ^ n12480 ^ 1'b0 ;
  assign n40696 = n5363 & ~n34126 ;
  assign n40697 = n34080 & n40696 ;
  assign n40698 = ~x162 & n3506 ;
  assign n40699 = n5064 & n34377 ;
  assign n40700 = ~n31528 & n40699 ;
  assign n40701 = n3283 ^ n320 ^ 1'b0 ;
  assign n40702 = ( n24124 & n28025 ) | ( n24124 & n38941 ) | ( n28025 & n38941 ) ;
  assign n40703 = ~n11756 & n34086 ;
  assign n40704 = n40703 ^ n14134 ^ 1'b0 ;
  assign n40705 = n3848 ^ n2512 ^ 1'b0 ;
  assign n40706 = n6874 | n22092 ;
  assign n40707 = n40706 ^ n6700 ^ 1'b0 ;
  assign n40708 = n40705 & ~n40707 ;
  assign n40709 = ~n5127 & n8124 ;
  assign n40710 = n3273 & ~n5077 ;
  assign n40711 = n40710 ^ n2986 ^ 1'b0 ;
  assign n40712 = n40711 ^ n31342 ^ 1'b0 ;
  assign n40713 = n33831 | n40712 ;
  assign n40714 = n19645 ^ n19621 ^ 1'b0 ;
  assign n40715 = n11041 & ~n40714 ;
  assign n40716 = n40715 ^ n36867 ^ n4724 ;
  assign n40717 = x66 | n40716 ;
  assign n40718 = n28784 ^ n14690 ^ n8245 ;
  assign n40719 = n11724 & n32147 ;
  assign n40720 = n905 & n15880 ;
  assign n40721 = n40720 ^ n23276 ^ 1'b0 ;
  assign n40722 = n10334 | n18547 ;
  assign n40723 = n40722 ^ n13371 ^ 1'b0 ;
  assign n40724 = n6205 ^ n3664 ^ 1'b0 ;
  assign n40725 = n1913 & n40724 ;
  assign n40726 = n15500 & n40725 ;
  assign n40729 = n11332 ^ n10052 ^ 1'b0 ;
  assign n40730 = ~n31007 & n40729 ;
  assign n40727 = n5550 & n15657 ;
  assign n40728 = ~n23937 & n40727 ;
  assign n40731 = n40730 ^ n40728 ^ 1'b0 ;
  assign n40732 = x55 | n30803 ;
  assign n40733 = n40731 & ~n40732 ;
  assign n40734 = n20594 ^ n19992 ^ n19099 ;
  assign n40735 = n34654 ^ n4072 ^ 1'b0 ;
  assign n40736 = n28162 | n40735 ;
  assign n40737 = n40736 ^ n2797 ^ 1'b0 ;
  assign n40738 = n3551 | n13328 ;
  assign n40739 = n21107 ^ n2873 ^ 1'b0 ;
  assign n40740 = n18520 & n40739 ;
  assign n40741 = n21086 ^ n12574 ^ 1'b0 ;
  assign n40742 = n7955 & n40741 ;
  assign n40743 = ~n19398 & n40742 ;
  assign n40744 = n1199 | n17458 ;
  assign n40745 = n30092 | n40744 ;
  assign n40746 = n32185 ^ n4242 ^ 1'b0 ;
  assign n40747 = n34428 & ~n40746 ;
  assign n40748 = ~n13921 & n40747 ;
  assign n40749 = n40748 ^ n26593 ^ 1'b0 ;
  assign n40750 = n37011 ^ n3754 ^ x84 ;
  assign n40751 = n18458 & n24217 ;
  assign n40752 = x241 & n40751 ;
  assign n40755 = n1575 & ~n30898 ;
  assign n40756 = ~n358 & n40755 ;
  assign n40753 = n5068 | n7445 ;
  assign n40754 = n5583 | n40753 ;
  assign n40757 = n40756 ^ n40754 ^ 1'b0 ;
  assign n40758 = n31478 & n35235 ;
  assign n40759 = n1827 & n17873 ;
  assign n40760 = n31066 & ~n40759 ;
  assign n40761 = ~n5514 & n40760 ;
  assign n40762 = n13689 & ~n28422 ;
  assign n40763 = n6937 & n7824 ;
  assign n40764 = n40763 ^ n5601 ^ 1'b0 ;
  assign n40765 = n40764 ^ n8441 ^ 1'b0 ;
  assign n40766 = ( n2672 & n7012 ) | ( n2672 & ~n18623 ) | ( n7012 & ~n18623 ) ;
  assign n40767 = n40766 ^ n4397 ^ 1'b0 ;
  assign n40768 = n5263 & n33313 ;
  assign n40769 = n40768 ^ n28857 ^ 1'b0 ;
  assign n40770 = ( ~n7849 & n21862 ) | ( ~n7849 & n29651 ) | ( n21862 & n29651 ) ;
  assign n40771 = n25835 ^ n5063 ^ 1'b0 ;
  assign n40772 = ~n21225 & n40771 ;
  assign n40773 = n10684 ^ n9814 ^ 1'b0 ;
  assign n40774 = ( n301 & ~n16617 ) | ( n301 & n28737 ) | ( ~n16617 & n28737 ) ;
  assign n40775 = n2442 & ~n40774 ;
  assign n40776 = n40775 ^ n27418 ^ 1'b0 ;
  assign n40777 = n16967 & ~n19986 ;
  assign n40778 = n20747 ^ n2389 ^ 1'b0 ;
  assign n40779 = n26144 ^ n24150 ^ n9851 ;
  assign n40780 = ( ~n5875 & n5987 ) | ( ~n5875 & n9077 ) | ( n5987 & n9077 ) ;
  assign n40781 = n16187 ^ n6331 ^ 1'b0 ;
  assign n40782 = n13320 & ~n40781 ;
  assign n40783 = ~n40780 & n40782 ;
  assign n40784 = n39831 ^ n5006 ^ 1'b0 ;
  assign n40785 = ~n3156 & n40784 ;
  assign n40786 = ( ~n7405 & n9012 ) | ( ~n7405 & n18200 ) | ( n9012 & n18200 ) ;
  assign n40787 = n33800 & ~n40786 ;
  assign n40788 = ~n9103 & n17384 ;
  assign n40789 = n40788 ^ n22671 ^ 1'b0 ;
  assign n40790 = n30323 | n30869 ;
  assign n40791 = ( n12034 & n16564 ) | ( n12034 & ~n33349 ) | ( n16564 & ~n33349 ) ;
  assign n40792 = n40791 ^ n17369 ^ 1'b0 ;
  assign n40793 = n32845 ^ n2513 ^ 1'b0 ;
  assign n40794 = n10078 & ~n11489 ;
  assign n40795 = n34980 ^ n16879 ^ 1'b0 ;
  assign n40796 = n2497 | n40795 ;
  assign n40797 = ~n19275 & n40796 ;
  assign n40798 = n21379 ^ n14507 ^ 1'b0 ;
  assign n40799 = n20555 & n40798 ;
  assign n40800 = n11831 | n16523 ;
  assign n40801 = n766 & ~n40800 ;
  assign n40802 = n22822 & n23465 ;
  assign n40803 = ~n1499 & n15780 ;
  assign n40804 = n2243 & ~n40803 ;
  assign n40805 = n40804 ^ n18945 ^ 1'b0 ;
  assign n40806 = n40802 & ~n40805 ;
  assign n40807 = n37177 ^ n2877 ^ 1'b0 ;
  assign n40808 = n40807 ^ n17907 ^ n12901 ;
  assign n40809 = n12888 ^ n11761 ^ n11591 ;
  assign n40810 = n5388 | n26475 ;
  assign n40811 = n5596 & ~n8619 ;
  assign n40812 = n24007 ^ n13284 ^ n7213 ;
  assign n40813 = n40811 & ~n40812 ;
  assign n40814 = ~n24969 & n38462 ;
  assign n40815 = n40814 ^ n10146 ^ 1'b0 ;
  assign n40816 = ( n9480 & n23072 ) | ( n9480 & n28130 ) | ( n23072 & n28130 ) ;
  assign n40817 = ~n8235 & n12470 ;
  assign n40818 = n37557 & n40817 ;
  assign n40819 = n7012 | n24854 ;
  assign n40820 = n29209 ^ n16925 ^ 1'b0 ;
  assign n40821 = n17749 & n18368 ;
  assign n40822 = n40820 & n40821 ;
  assign n40823 = n8048 ^ n2294 ^ 1'b0 ;
  assign n40824 = n40823 ^ n30193 ^ 1'b0 ;
  assign n40825 = n40822 | n40824 ;
  assign n40826 = n40819 & ~n40825 ;
  assign n40828 = n668 | n4746 ;
  assign n40827 = n5495 & ~n9327 ;
  assign n40829 = n40828 ^ n40827 ^ 1'b0 ;
  assign n40830 = n8889 | n16470 ;
  assign n40831 = n40830 ^ n9494 ^ 1'b0 ;
  assign n40832 = ~n29151 & n40831 ;
  assign n40833 = n40832 ^ n35062 ^ n4456 ;
  assign n40837 = ~n15426 & n15689 ;
  assign n40838 = n2632 & n40837 ;
  assign n40834 = ~n3168 & n39527 ;
  assign n40835 = n9653 ^ n5632 ^ 1'b0 ;
  assign n40836 = n40834 & ~n40835 ;
  assign n40839 = n40838 ^ n40836 ^ n19380 ;
  assign n40840 = n1594 & ~n2040 ;
  assign n40841 = ~n7063 & n17155 ;
  assign n40842 = ~n6784 & n40841 ;
  assign n40843 = ( n3336 & ~n10969 ) | ( n3336 & n16024 ) | ( ~n10969 & n16024 ) ;
  assign n40844 = n13161 & n24906 ;
  assign n40845 = n18004 ^ n6408 ^ 1'b0 ;
  assign n40846 = n40364 ^ n25945 ^ n14272 ;
  assign n40847 = n20418 & ~n21838 ;
  assign n40848 = n40847 ^ n33409 ^ 1'b0 ;
  assign n40849 = ( ~n5817 & n22538 ) | ( ~n5817 & n40848 ) | ( n22538 & n40848 ) ;
  assign n40850 = n13746 ^ n4425 ^ 1'b0 ;
  assign n40851 = n36575 ^ n35185 ^ 1'b0 ;
  assign n40852 = n34660 ^ n30169 ^ n20300 ;
  assign n40853 = n32953 ^ n16605 ^ n3778 ;
  assign n40854 = n3738 & ~n40853 ;
  assign n40855 = n3923 & ~n5511 ;
  assign n40856 = n5133 | n18228 ;
  assign n40857 = n15532 & ~n40856 ;
  assign n40858 = n20657 ^ n9541 ^ n1633 ;
  assign n40859 = n11252 & ~n28504 ;
  assign n40860 = n40859 ^ n23316 ^ 1'b0 ;
  assign n40861 = n33719 ^ n16133 ^ 1'b0 ;
  assign n40862 = ( ~n5986 & n25205 ) | ( ~n5986 & n37604 ) | ( n25205 & n37604 ) ;
  assign n40863 = n12971 & ~n17424 ;
  assign n40864 = n21390 ^ n15422 ^ 1'b0 ;
  assign n40865 = n40863 | n40864 ;
  assign n40866 = n40865 ^ n10357 ^ 1'b0 ;
  assign n40867 = n40866 ^ n21341 ^ n6141 ;
  assign n40868 = n14498 & ~n19748 ;
  assign n40869 = ( n6929 & n40867 ) | ( n6929 & ~n40868 ) | ( n40867 & ~n40868 ) ;
  assign n40870 = n27894 ^ n3723 ^ 1'b0 ;
  assign n40871 = n27790 & ~n38613 ;
  assign n40872 = ~n1006 & n40871 ;
  assign n40873 = n13232 & ~n14236 ;
  assign n40874 = n40873 ^ n7890 ^ 1'b0 ;
  assign n40875 = n3683 | n40874 ;
  assign n40876 = n39040 & ~n40875 ;
  assign n40877 = n29260 ^ n14154 ^ 1'b0 ;
  assign n40878 = n7863 & ~n40877 ;
  assign n40879 = x133 & n9733 ;
  assign n40880 = n40879 ^ n5338 ^ 1'b0 ;
  assign n40881 = n1237 & ~n7457 ;
  assign n40882 = n30916 & n40881 ;
  assign n40883 = n5343 & ~n6019 ;
  assign n40884 = n15364 & n40883 ;
  assign n40885 = n18091 | n40884 ;
  assign n40886 = n12638 & ~n40885 ;
  assign n40887 = n40050 ^ n30538 ^ n397 ;
  assign n40888 = n37126 ^ n9198 ^ 1'b0 ;
  assign n40889 = ( n6463 & n6919 ) | ( n6463 & n40505 ) | ( n6919 & n40505 ) ;
  assign n40890 = ~n4493 & n40889 ;
  assign n40891 = n21031 & ~n33055 ;
  assign n40892 = ~n24537 & n40891 ;
  assign n40893 = n25973 ^ n3924 ^ 1'b0 ;
  assign n40894 = n29049 & n36412 ;
  assign n40895 = n21064 & n40894 ;
  assign n40896 = n10856 ^ n2335 ^ x146 ;
  assign n40897 = n20684 & ~n29928 ;
  assign n40898 = ~n4777 & n9559 ;
  assign n40899 = n40898 ^ n23766 ^ 1'b0 ;
  assign n40900 = n3174 & n36458 ;
  assign n40901 = n2234 & n40900 ;
  assign n40902 = ~x155 & n1594 ;
  assign n40903 = n39059 ^ n12332 ^ 1'b0 ;
  assign n40904 = n21539 & n29661 ;
  assign n40905 = ~n11469 & n40904 ;
  assign n40906 = n2548 | n40815 ;
  assign n40907 = n40905 & ~n40906 ;
  assign n40908 = n15664 ^ n7994 ^ 1'b0 ;
  assign n40909 = ( ~n13357 & n29888 ) | ( ~n13357 & n40908 ) | ( n29888 & n40908 ) ;
  assign n40910 = n33435 ^ n3763 ^ 1'b0 ;
  assign n40911 = n1558 | n2711 ;
  assign n40912 = n40911 ^ n1716 ^ 1'b0 ;
  assign n40913 = ~n38252 & n40912 ;
  assign n40914 = ~n1038 & n9559 ;
  assign n40915 = n40914 ^ n16767 ^ 1'b0 ;
  assign n40916 = n1440 & n33503 ;
  assign n40917 = ( n9790 & n11483 ) | ( n9790 & ~n37086 ) | ( n11483 & ~n37086 ) ;
  assign n40918 = n8218 & n25892 ;
  assign n40919 = n36194 & n40918 ;
  assign n40920 = n40919 ^ n35126 ^ 1'b0 ;
  assign n40921 = ~n5636 & n36106 ;
  assign n40922 = n7578 & n40921 ;
  assign n40923 = n30338 ^ n23426 ^ 1'b0 ;
  assign n40924 = ~n14974 & n40923 ;
  assign n40925 = n40924 ^ n11633 ^ 1'b0 ;
  assign n40926 = n9842 | n40925 ;
  assign n40927 = n12922 ^ n11393 ^ 1'b0 ;
  assign n40928 = n38923 & ~n40927 ;
  assign n40929 = n18741 & n34128 ;
  assign n40930 = ~n29851 & n40929 ;
  assign n40931 = n14246 & ~n40930 ;
  assign n40932 = n11810 | n13575 ;
  assign n40933 = n4315 & ~n40932 ;
  assign n40934 = n32405 ^ n12608 ^ 1'b0 ;
  assign n40935 = n40933 | n40934 ;
  assign n40936 = ( n11386 & n33579 ) | ( n11386 & ~n38816 ) | ( n33579 & ~n38816 ) ;
  assign n40937 = ~n5022 & n40936 ;
  assign n40938 = n40937 ^ n7755 ^ 1'b0 ;
  assign n40939 = x215 & ~n40938 ;
  assign n40940 = n1869 & ~n2437 ;
  assign n40941 = n40940 ^ n21446 ^ 1'b0 ;
  assign n40942 = n18495 ^ n9638 ^ n7172 ;
  assign n40943 = n5903 & n13069 ;
  assign n40944 = ~n36627 & n40943 ;
  assign n40945 = n13359 & n19258 ;
  assign n40946 = n34818 ^ n16441 ^ n1876 ;
  assign n40947 = ~n9952 & n40946 ;
  assign n40948 = n39220 ^ n14584 ^ 1'b0 ;
  assign n40949 = ~n10068 & n19602 ;
  assign n40955 = n25420 ^ n16688 ^ 1'b0 ;
  assign n40950 = n18509 ^ n18267 ^ n1692 ;
  assign n40951 = n6979 | n38764 ;
  assign n40952 = n10246 | n40951 ;
  assign n40953 = n40952 ^ n28813 ^ 1'b0 ;
  assign n40954 = n40950 & n40953 ;
  assign n40956 = n40955 ^ n40954 ^ 1'b0 ;
  assign n40957 = n25077 & ~n31419 ;
  assign n40958 = n11824 | n40880 ;
  assign n40959 = x55 & ~n21690 ;
  assign n40960 = n40959 ^ n16164 ^ 1'b0 ;
  assign n40961 = ( ~n13900 & n21773 ) | ( ~n13900 & n40960 ) | ( n21773 & n40960 ) ;
  assign n40962 = n36254 ^ n25931 ^ n16352 ;
  assign n40963 = n35114 ^ n16123 ^ n1605 ;
  assign n40964 = n40963 ^ n8098 ^ x251 ;
  assign n40965 = n33348 ^ n5669 ^ 1'b0 ;
  assign n40966 = ~n12167 & n40965 ;
  assign n40967 = n40964 & n40966 ;
  assign n40968 = n6031 & n14326 ;
  assign n40969 = n38800 & n40968 ;
  assign n40970 = n12275 | n22828 ;
  assign n40971 = n40970 ^ n37426 ^ 1'b0 ;
  assign n40972 = n28731 ^ n3193 ^ 1'b0 ;
  assign n40973 = n19245 & n40972 ;
  assign n40974 = n27414 ^ n6778 ^ 1'b0 ;
  assign n40975 = n40973 & ~n40974 ;
  assign n40976 = ( n17769 & n26603 ) | ( n17769 & ~n31226 ) | ( n26603 & ~n31226 ) ;
  assign n40977 = n39108 ^ n10236 ^ 1'b0 ;
  assign n40978 = ~n15337 & n38712 ;
  assign n40979 = n40978 ^ n3776 ^ 1'b0 ;
  assign n40980 = n8578 | n21559 ;
  assign n40981 = ~n29037 & n40980 ;
  assign n40982 = ( ~n11831 & n28015 ) | ( ~n11831 & n37729 ) | ( n28015 & n37729 ) ;
  assign n40983 = n40982 ^ n40650 ^ n31931 ;
  assign n40984 = n2910 ^ n1166 ^ 1'b0 ;
  assign n40985 = n7047 & ~n20802 ;
  assign n40986 = n5976 | n27796 ;
  assign n40987 = n28307 ^ n26252 ^ 1'b0 ;
  assign n40989 = n8775 & ~n33735 ;
  assign n40988 = n22152 & n29578 ;
  assign n40990 = n40989 ^ n40988 ^ 1'b0 ;
  assign n40991 = ( n18690 & ~n24817 ) | ( n18690 & n38696 ) | ( ~n24817 & n38696 ) ;
  assign n40992 = n7844 ^ n5588 ^ 1'b0 ;
  assign n40994 = n15597 & n29385 ;
  assign n40993 = ( n2085 & n10168 ) | ( n2085 & n33379 ) | ( n10168 & n33379 ) ;
  assign n40995 = n40994 ^ n40993 ^ n18574 ;
  assign n40996 = n5685 & ~n13749 ;
  assign n40997 = n40996 ^ n18045 ^ 1'b0 ;
  assign n40998 = n40997 ^ n29151 ^ n3898 ;
  assign n40999 = n11912 & ~n40998 ;
  assign n41000 = n15025 ^ n5068 ^ 1'b0 ;
  assign n41001 = ~n19414 & n41000 ;
  assign n41002 = ( n26194 & n40153 ) | ( n26194 & ~n41001 ) | ( n40153 & ~n41001 ) ;
  assign n41003 = n33517 ^ n27499 ^ x67 ;
  assign n41004 = ~n41002 & n41003 ;
  assign n41005 = n21787 ^ n16839 ^ n3954 ;
  assign n41007 = n693 | n913 ;
  assign n41006 = x83 & ~n1056 ;
  assign n41008 = n41007 ^ n41006 ^ 1'b0 ;
  assign n41009 = n41008 ^ n34093 ^ n749 ;
  assign n41010 = n5988 & n22228 ;
  assign n41011 = n41010 ^ n8682 ^ 1'b0 ;
  assign n41012 = ( n6520 & n18050 ) | ( n6520 & n23131 ) | ( n18050 & n23131 ) ;
  assign n41013 = n41012 ^ n28583 ^ 1'b0 ;
  assign n41014 = n18938 ^ n5164 ^ 1'b0 ;
  assign n41015 = ~n11109 & n16925 ;
  assign n41016 = ~n2586 & n41015 ;
  assign n41018 = n37916 ^ n15002 ^ 1'b0 ;
  assign n41017 = ( n12478 & n20651 ) | ( n12478 & ~n33602 ) | ( n20651 & ~n33602 ) ;
  assign n41019 = n41018 ^ n41017 ^ n38471 ;
  assign n41020 = n41019 ^ n2585 ^ 1'b0 ;
  assign n41021 = n12932 & n39218 ;
  assign n41022 = n41020 & n41021 ;
  assign n41023 = n3126 & ~n4627 ;
  assign n41024 = n19138 ^ n6851 ^ 1'b0 ;
  assign n41025 = n41023 & n41024 ;
  assign n41026 = n2082 & n5610 ;
  assign n41027 = n41026 ^ n5345 ^ 1'b0 ;
  assign n41028 = n41027 ^ n37536 ^ 1'b0 ;
  assign n41029 = n40716 ^ n12068 ^ 1'b0 ;
  assign n41030 = n25048 ^ n6461 ^ 1'b0 ;
  assign n41031 = n10825 | n25115 ;
  assign n41032 = ( n17302 & ~n30727 ) | ( n17302 & n32108 ) | ( ~n30727 & n32108 ) ;
  assign n41033 = n41032 ^ n20797 ^ 1'b0 ;
  assign n41034 = ~n11723 & n41033 ;
  assign n41035 = ~n1106 & n26861 ;
  assign n41036 = ~n41034 & n41035 ;
  assign n41037 = ~n12925 & n25607 ;
  assign n41038 = n21207 ^ n11903 ^ 1'b0 ;
  assign n41039 = n18587 & ~n41038 ;
  assign n41040 = n14677 & ~n19438 ;
  assign n41041 = ~n41039 & n41040 ;
  assign n41042 = n11286 ^ n6953 ^ 1'b0 ;
  assign n41043 = n41042 ^ n12552 ^ 1'b0 ;
  assign n41044 = n26133 & ~n41043 ;
  assign n41045 = n8513 ^ n4242 ^ 1'b0 ;
  assign n41046 = n37923 & n41045 ;
  assign n41047 = n17716 | n20235 ;
  assign n41048 = n41047 ^ n28424 ^ 1'b0 ;
  assign n41049 = n8298 | n24531 ;
  assign n41050 = n18601 & ~n41049 ;
  assign n41052 = n344 & n7250 ;
  assign n41053 = n41052 ^ n8772 ^ 1'b0 ;
  assign n41054 = n41053 ^ n36939 ^ n34157 ;
  assign n41051 = n5084 & ~n19856 ;
  assign n41055 = n41054 ^ n41051 ^ 1'b0 ;
  assign n41056 = n2337 & n32680 ;
  assign n41057 = n1015 & n41056 ;
  assign n41058 = n1055 | n33482 ;
  assign n41059 = n17646 & n18758 ;
  assign n41060 = ~n15140 & n41059 ;
  assign n41061 = n33480 & ~n41060 ;
  assign n41062 = n28510 & n30036 ;
  assign n41063 = n2218 & n15983 ;
  assign n41064 = n7721 ^ n1665 ^ 1'b0 ;
  assign n41065 = n16409 | n41064 ;
  assign n41066 = n5522 & ~n16142 ;
  assign n41067 = n34032 & n41066 ;
  assign n41068 = n15555 & ~n41067 ;
  assign n41069 = ~n20721 & n41068 ;
  assign n41070 = n30385 ^ n26630 ^ 1'b0 ;
  assign n41071 = ~n41069 & n41070 ;
  assign n41072 = n16352 ^ n10343 ^ 1'b0 ;
  assign n41073 = n5423 & n41072 ;
  assign n41074 = n4394 | n41073 ;
  assign n41076 = n2648 & n3103 ;
  assign n41075 = n19097 & ~n24711 ;
  assign n41077 = n41076 ^ n41075 ^ n16427 ;
  assign n41078 = n32322 ^ n15835 ^ 1'b0 ;
  assign n41079 = ~n32922 & n38481 ;
  assign n41080 = n41079 ^ n7306 ^ 1'b0 ;
  assign n41081 = n15080 & ~n31901 ;
  assign n41082 = n7554 & n41081 ;
  assign n41083 = n2250 & ~n13725 ;
  assign n41084 = n36463 & n41083 ;
  assign n41085 = ~n365 & n7126 ;
  assign n41086 = n15793 & n41085 ;
  assign n41087 = ~n13266 & n41086 ;
  assign n41088 = n5135 & n39949 ;
  assign n41089 = n2957 & n21591 ;
  assign n41090 = n16964 & n41089 ;
  assign n41091 = n9187 | n21462 ;
  assign n41092 = n41091 ^ n9594 ^ 1'b0 ;
  assign n41093 = n14922 ^ n1304 ^ 1'b0 ;
  assign n41094 = n2924 & ~n41093 ;
  assign n41095 = ~n5926 & n41094 ;
  assign n41096 = n30083 & n41095 ;
  assign n41097 = n15847 & ~n29471 ;
  assign n41098 = ~n35870 & n41097 ;
  assign n41099 = n13740 ^ n8352 ^ 1'b0 ;
  assign n41100 = n9838 | n20212 ;
  assign n41101 = n3275 | n41100 ;
  assign n41102 = ( n9177 & n17076 ) | ( n9177 & n41101 ) | ( n17076 & n41101 ) ;
  assign n41103 = n15418 ^ n3405 ^ 1'b0 ;
  assign n41104 = ~n24847 & n41103 ;
  assign n41105 = n8678 & n18978 ;
  assign n41106 = ~n20824 & n41105 ;
  assign n41107 = n31496 ^ n7426 ^ 1'b0 ;
  assign n41108 = n9273 | n17068 ;
  assign n41109 = ( n8659 & ~n41107 ) | ( n8659 & n41108 ) | ( ~n41107 & n41108 ) ;
  assign n41110 = ~n13932 & n41109 ;
  assign n41111 = n38471 & n41110 ;
  assign n41112 = n22293 & ~n33574 ;
  assign n41113 = ~x244 & n29758 ;
  assign n41114 = n41113 ^ n37510 ^ 1'b0 ;
  assign n41115 = n11833 & n17241 ;
  assign n41116 = ( n1486 & n23698 ) | ( n1486 & n24928 ) | ( n23698 & n24928 ) ;
  assign n41117 = n12908 & ~n41116 ;
  assign n41118 = n41117 ^ n27496 ^ 1'b0 ;
  assign n41119 = n13450 & n41118 ;
  assign n41120 = n34311 & n41119 ;
  assign n41121 = n10627 ^ n9353 ^ 1'b0 ;
  assign n41122 = n17192 & ~n41121 ;
  assign n41123 = n9693 ^ n6398 ^ 1'b0 ;
  assign n41124 = n474 & n18025 ;
  assign n41125 = n41124 ^ n5885 ^ 1'b0 ;
  assign n41126 = n11988 & n40682 ;
  assign n41127 = ~n41125 & n41126 ;
  assign n41128 = n10408 & ~n25390 ;
  assign n41129 = n41127 & n41128 ;
  assign n41130 = n29711 ^ n15620 ^ 1'b0 ;
  assign n41131 = ( n2777 & n4343 ) | ( n2777 & n6842 ) | ( n4343 & n6842 ) ;
  assign n41132 = ~n2621 & n41131 ;
  assign n41133 = n41132 ^ n40749 ^ n32034 ;
  assign n41134 = n14979 & n29249 ;
  assign n41135 = n41134 ^ n8239 ^ 1'b0 ;
  assign n41136 = ~x149 & n6129 ;
  assign n41137 = n8318 ^ n5773 ^ 1'b0 ;
  assign n41138 = ~n2782 & n13460 ;
  assign n41139 = n41138 ^ n16691 ^ 1'b0 ;
  assign n41140 = n41139 ^ n26929 ^ 1'b0 ;
  assign n41141 = n4705 & n11581 ;
  assign n41142 = n41141 ^ n35469 ^ 1'b0 ;
  assign n41143 = n13171 & n29542 ;
  assign n41144 = n40008 ^ n34398 ^ 1'b0 ;
  assign n41145 = n20056 ^ n10422 ^ 1'b0 ;
  assign n41146 = n41145 ^ n5131 ^ n704 ;
  assign n41147 = ( ~n5586 & n8541 ) | ( ~n5586 & n12612 ) | ( n8541 & n12612 ) ;
  assign n41148 = n3894 & ~n16338 ;
  assign n41149 = ~n2614 & n3638 ;
  assign n41150 = n5042 & n41149 ;
  assign n41151 = n7793 ^ n663 ^ 1'b0 ;
  assign n41152 = n41150 | n41151 ;
  assign n41153 = n8027 & ~n11397 ;
  assign n41154 = n41153 ^ n31919 ^ 1'b0 ;
  assign n41155 = ( ~n1444 & n1458 ) | ( ~n1444 & n30871 ) | ( n1458 & n30871 ) ;
  assign n41156 = n11196 & ~n27029 ;
  assign n41157 = n29495 ^ n2081 ^ 1'b0 ;
  assign n41158 = n41156 | n41157 ;
  assign n41159 = n6329 & ~n13000 ;
  assign n41160 = n35739 ^ n8413 ^ 1'b0 ;
  assign n41161 = ~n41159 & n41160 ;
  assign n41162 = n41161 ^ n19606 ^ n18020 ;
  assign n41163 = ( n19998 & n41158 ) | ( n19998 & ~n41162 ) | ( n41158 & ~n41162 ) ;
  assign n41164 = n20850 & n32254 ;
  assign n41165 = ~x120 & n41164 ;
  assign n41166 = ~n4699 & n13202 ;
  assign n41167 = n41166 ^ n11616 ^ 1'b0 ;
  assign n41168 = n30210 ^ n5244 ^ 1'b0 ;
  assign n41169 = n41167 & n41168 ;
  assign n41170 = ~n1202 & n3721 ;
  assign n41171 = n41170 ^ n29037 ^ 1'b0 ;
  assign n41172 = n41169 & n41171 ;
  assign n41173 = n37875 ^ n34395 ^ 1'b0 ;
  assign n41174 = n10940 & ~n23035 ;
  assign n41175 = ~n9952 & n41174 ;
  assign n41176 = ~n581 & n6967 ;
  assign n41177 = n19538 | n24145 ;
  assign n41178 = n30260 ^ n2378 ^ 1'b0 ;
  assign n41179 = n9496 & n13467 ;
  assign n41180 = n41179 ^ n17961 ^ n6045 ;
  assign n41181 = ~n7700 & n10004 ;
  assign n41182 = ~n24482 & n41181 ;
  assign n41183 = n41182 ^ n12253 ^ 1'b0 ;
  assign n41184 = n41183 ^ n11072 ^ n6053 ;
  assign n41185 = n41184 ^ n18891 ^ n8484 ;
  assign n41186 = n12802 & n33498 ;
  assign n41187 = n41186 ^ n28132 ^ 1'b0 ;
  assign n41188 = n32777 ^ n8594 ^ n622 ;
  assign n41189 = n2993 & n21385 ;
  assign n41190 = n41188 & n41189 ;
  assign n41191 = n1947 | n18994 ;
  assign n41192 = n6103 | n41191 ;
  assign n41193 = n41190 & ~n41192 ;
  assign n41194 = n15390 ^ n10469 ^ 1'b0 ;
  assign n41195 = n40019 | n41194 ;
  assign n41196 = n4050 & ~n4152 ;
  assign n41197 = n41196 ^ n8900 ^ 1'b0 ;
  assign n41198 = n4167 | n5352 ;
  assign n41199 = n41197 | n41198 ;
  assign n41200 = n10777 & n30995 ;
  assign n41202 = n24086 ^ n8037 ^ n7342 ;
  assign n41203 = n19625 & ~n41202 ;
  assign n41201 = ~n13492 & n18394 ;
  assign n41204 = n41203 ^ n41201 ^ 1'b0 ;
  assign n41205 = n6296 & n13843 ;
  assign n41206 = ~n8856 & n27889 ;
  assign n41207 = n37485 ^ n23001 ^ 1'b0 ;
  assign n41208 = n17748 ^ n8226 ^ 1'b0 ;
  assign n41209 = ~n5949 & n41208 ;
  assign n41210 = n41209 ^ n37092 ^ 1'b0 ;
  assign n41213 = n3256 | n5996 ;
  assign n41214 = n41213 ^ n2133 ^ 1'b0 ;
  assign n41211 = n27038 ^ n3874 ^ 1'b0 ;
  assign n41212 = n41211 ^ n36828 ^ n1339 ;
  assign n41215 = n41214 ^ n41212 ^ n39888 ;
  assign n41216 = n20868 ^ n2819 ^ 1'b0 ;
  assign n41217 = n17938 ^ n11649 ^ 1'b0 ;
  assign n41218 = n10759 | n15608 ;
  assign n41219 = n15608 & ~n41218 ;
  assign n41220 = ~x242 & n21569 ;
  assign n41221 = n37944 ^ n20301 ^ 1'b0 ;
  assign n41222 = n11575 & n41221 ;
  assign n41223 = n6833 & ~n8842 ;
  assign n41224 = ~n14138 & n41223 ;
  assign n41225 = n20561 ^ n1036 ^ 1'b0 ;
  assign n41226 = ( n5463 & n41224 ) | ( n5463 & n41225 ) | ( n41224 & n41225 ) ;
  assign n41227 = ~n35012 & n38631 ;
  assign n41228 = n11587 ^ n6995 ^ 1'b0 ;
  assign n41229 = ~n38251 & n41228 ;
  assign n41230 = n41229 ^ n19856 ^ n10382 ;
  assign n41231 = n41230 ^ n34935 ^ n21362 ;
  assign n41232 = n41231 ^ x36 ^ 1'b0 ;
  assign n41233 = n32740 ^ n7939 ^ 1'b0 ;
  assign n41234 = n17483 ^ n12505 ^ 1'b0 ;
  assign n41235 = ~n28032 & n41234 ;
  assign n41236 = n41235 ^ n33987 ^ 1'b0 ;
  assign n41237 = n17124 ^ n2279 ^ 1'b0 ;
  assign n41238 = n6719 & ~n41237 ;
  assign n41239 = n12355 ^ n9352 ^ 1'b0 ;
  assign n41240 = ~n4931 & n41239 ;
  assign n41241 = n4545 & ~n6800 ;
  assign n41242 = ( n9782 & n10288 ) | ( n9782 & ~n41241 ) | ( n10288 & ~n41241 ) ;
  assign n41243 = n38033 ^ n4750 ^ 1'b0 ;
  assign n41244 = ~n13948 & n28007 ;
  assign n41245 = ~n3335 & n35219 ;
  assign n41246 = n2650 | n14738 ;
  assign n41247 = n41246 ^ n16684 ^ 1'b0 ;
  assign n41248 = n18124 ^ n13920 ^ 1'b0 ;
  assign n41249 = n3695 & ~n41248 ;
  assign n41250 = n33416 ^ n15353 ^ 1'b0 ;
  assign n41251 = n13806 ^ n7598 ^ 1'b0 ;
  assign n41252 = n41251 ^ n25253 ^ n10771 ;
  assign n41254 = n8403 & n31042 ;
  assign n41253 = n2360 | n5043 ;
  assign n41255 = n41254 ^ n41253 ^ x86 ;
  assign n41256 = n14918 & ~n24614 ;
  assign n41257 = ~n17934 & n41256 ;
  assign n41258 = n41257 ^ n27942 ^ n11070 ;
  assign n41259 = n23890 ^ n13581 ^ 1'b0 ;
  assign n41260 = ~n11951 & n30293 ;
  assign n41261 = n41260 ^ n6906 ^ 1'b0 ;
  assign n41262 = n29010 | n29959 ;
  assign n41263 = ~n22327 & n41262 ;
  assign n41264 = n1521 & n22414 ;
  assign n41265 = ~n14102 & n17038 ;
  assign n41266 = n8433 | n41265 ;
  assign n41267 = ~n23583 & n33381 ;
  assign n41268 = n41267 ^ n23318 ^ 1'b0 ;
  assign n41269 = n4315 & ~n9123 ;
  assign n41270 = n41269 ^ n1460 ^ 1'b0 ;
  assign n41271 = n41268 | n41270 ;
  assign n41272 = ~n1518 & n23698 ;
  assign n41273 = n31209 ^ n6784 ^ 1'b0 ;
  assign n41274 = ( n959 & ~n1991 ) | ( n959 & n2506 ) | ( ~n1991 & n2506 ) ;
  assign n41275 = n1421 & n41274 ;
  assign n41276 = n20546 & n41275 ;
  assign n41277 = n10332 & n41276 ;
  assign n41278 = ( n14405 & n25181 ) | ( n14405 & n41277 ) | ( n25181 & n41277 ) ;
  assign n41279 = n6866 & n12554 ;
  assign n41280 = n41279 ^ n7572 ^ 1'b0 ;
  assign n41281 = ~n6253 & n21264 ;
  assign n41282 = n41281 ^ n10900 ^ 1'b0 ;
  assign n41283 = n28449 & ~n41282 ;
  assign n41284 = n41280 & n41283 ;
  assign n41285 = n4948 | n41284 ;
  assign n41286 = n6225 & n9529 ;
  assign n41287 = n41286 ^ n11505 ^ 1'b0 ;
  assign n41288 = n41287 ^ n9345 ^ 1'b0 ;
  assign n41289 = ~n3690 & n33226 ;
  assign n41290 = n18808 ^ n4777 ^ 1'b0 ;
  assign n41291 = n3757 | n41290 ;
  assign n41292 = n34367 ^ n18697 ^ 1'b0 ;
  assign n41293 = n9919 | n27488 ;
  assign n41294 = n41293 ^ n21121 ^ n14028 ;
  assign n41295 = ~n26426 & n41294 ;
  assign n41296 = n9877 ^ n6751 ^ 1'b0 ;
  assign n41297 = n21899 ^ n7732 ^ n4826 ;
  assign n41298 = n41297 ^ n20469 ^ 1'b0 ;
  assign n41299 = n11819 & ~n41298 ;
  assign n41300 = n8432 | n19085 ;
  assign n41301 = n37463 | n41300 ;
  assign n41302 = n10315 & n41301 ;
  assign n41303 = ~n31136 & n41302 ;
  assign n41304 = ~n2266 & n40946 ;
  assign n41305 = n1462 & ~n23108 ;
  assign n41306 = n20777 & n41305 ;
  assign n41307 = n7658 ^ n3604 ^ 1'b0 ;
  assign n41310 = n9355 ^ n6756 ^ 1'b0 ;
  assign n41308 = n7074 & ~n21089 ;
  assign n41309 = n41308 ^ n20979 ^ 1'b0 ;
  assign n41311 = n41310 ^ n41309 ^ n21481 ;
  assign n41312 = n39578 ^ n23005 ^ 1'b0 ;
  assign n41313 = n11815 & n23533 ;
  assign n41314 = n11897 & n41313 ;
  assign n41315 = n18539 ^ n16781 ^ 1'b0 ;
  assign n41316 = n7170 & n41315 ;
  assign n41317 = n38790 ^ n34342 ^ n6321 ;
  assign n41318 = n35304 ^ n11653 ^ n5895 ;
  assign n41319 = n18942 ^ n4790 ^ 1'b0 ;
  assign n41320 = n41319 ^ n7899 ^ n3985 ;
  assign n41321 = n41320 ^ n29179 ^ 1'b0 ;
  assign n41322 = n41321 ^ n12411 ^ 1'b0 ;
  assign n41323 = n4977 & n41322 ;
  assign n41325 = n3998 & n24721 ;
  assign n41324 = n17672 & n20470 ;
  assign n41326 = n41325 ^ n41324 ^ 1'b0 ;
  assign n41327 = ~n7393 & n41326 ;
  assign n41328 = n30286 ^ n15846 ^ 1'b0 ;
  assign n41329 = n1295 & n4480 ;
  assign n41332 = ~n18775 & n22122 ;
  assign n41333 = n8080 & n41332 ;
  assign n41330 = n835 & n18189 ;
  assign n41331 = n41330 ^ n35103 ^ 1'b0 ;
  assign n41334 = n41333 ^ n41331 ^ n1991 ;
  assign n41339 = n34526 ^ n20508 ^ 1'b0 ;
  assign n41340 = n15988 | n41339 ;
  assign n41341 = n33427 & ~n41340 ;
  assign n41337 = n11070 ^ n7668 ^ 1'b0 ;
  assign n41335 = n10169 ^ n6569 ^ 1'b0 ;
  assign n41336 = n15341 & ~n41335 ;
  assign n41338 = n41337 ^ n41336 ^ 1'b0 ;
  assign n41342 = n41341 ^ n41338 ^ n5725 ;
  assign n41343 = n28826 ^ n14421 ^ n9259 ;
  assign n41345 = n18520 ^ n12346 ^ n4366 ;
  assign n41344 = n608 & n23689 ;
  assign n41346 = n41345 ^ n41344 ^ 1'b0 ;
  assign n41347 = n16003 & ~n23511 ;
  assign n41348 = n27578 ^ n26636 ^ 1'b0 ;
  assign n41349 = ~n30117 & n41348 ;
  assign n41350 = n28784 ^ n19830 ^ 1'b0 ;
  assign n41351 = n1478 & n8762 ;
  assign n41352 = ~n38794 & n41351 ;
  assign n41353 = n11620 | n40831 ;
  assign n41354 = ~n15624 & n39846 ;
  assign n41355 = n41354 ^ n5675 ^ 1'b0 ;
  assign n41356 = n12123 | n29198 ;
  assign n41357 = n28132 & n41356 ;
  assign n41358 = n33321 ^ n23786 ^ 1'b0 ;
  assign n41359 = n4284 & n24302 ;
  assign n41360 = n2418 & n14502 ;
  assign n41361 = ~n631 & n41360 ;
  assign n41362 = n27411 ^ n11559 ^ 1'b0 ;
  assign n41363 = ~n1582 & n41362 ;
  assign n41364 = n29922 & n41363 ;
  assign n41365 = n557 & n38314 ;
  assign n41366 = n11145 | n12766 ;
  assign n41367 = n4864 ^ n931 ^ 1'b0 ;
  assign n41368 = n18260 ^ n1304 ^ 1'b0 ;
  assign n41369 = ~n23760 & n41358 ;
  assign n41370 = n41369 ^ n41157 ^ 1'b0 ;
  assign n41371 = n10120 & ~n24759 ;
  assign n41372 = n35758 ^ n8597 ^ 1'b0 ;
  assign n41373 = n26787 | n34031 ;
  assign n41374 = ~n25446 & n41373 ;
  assign n41375 = ~n13188 & n41374 ;
  assign n41376 = n41375 ^ n25263 ^ n14762 ;
  assign n41377 = n28695 ^ n24706 ^ 1'b0 ;
  assign n41378 = n41376 & ~n41377 ;
  assign n41379 = ( n12382 & n41372 ) | ( n12382 & n41378 ) | ( n41372 & n41378 ) ;
  assign n41380 = n16715 & n41379 ;
  assign n41381 = ~n41371 & n41380 ;
  assign n41382 = ( n4170 & n4211 ) | ( n4170 & ~n34568 ) | ( n4211 & ~n34568 ) ;
  assign n41387 = n15302 ^ n761 ^ 1'b0 ;
  assign n41388 = ~n5260 & n41387 ;
  assign n41383 = ( n10248 & ~n10966 ) | ( n10248 & n18427 ) | ( ~n10966 & n18427 ) ;
  assign n41384 = n41383 ^ n34870 ^ 1'b0 ;
  assign n41385 = ~n28488 & n41384 ;
  assign n41386 = ( ~n22167 & n32805 ) | ( ~n22167 & n41385 ) | ( n32805 & n41385 ) ;
  assign n41389 = n41388 ^ n41386 ^ 1'b0 ;
  assign n41390 = n24780 ^ n12669 ^ n4042 ;
  assign n41391 = n13140 ^ n2598 ^ 1'b0 ;
  assign n41392 = x76 & ~n21593 ;
  assign n41393 = n41392 ^ n3365 ^ 1'b0 ;
  assign n41394 = n8785 ^ n5133 ^ n3201 ;
  assign n41395 = n6728 | n26832 ;
  assign n41396 = n1653 & ~n24263 ;
  assign n41397 = n15442 | n32035 ;
  assign n41398 = n30520 & ~n41397 ;
  assign n41399 = n36971 & n41398 ;
  assign n41400 = n22475 ^ n15580 ^ 1'b0 ;
  assign n41401 = n41400 ^ n6541 ^ 1'b0 ;
  assign n41402 = n11642 | n41401 ;
  assign n41403 = n4473 & n7854 ;
  assign n41404 = ~n4259 & n19706 ;
  assign n41405 = n41404 ^ n17527 ^ 1'b0 ;
  assign n41406 = ~n41403 & n41405 ;
  assign n41408 = ( ~n17000 & n27519 ) | ( ~n17000 & n30001 ) | ( n27519 & n30001 ) ;
  assign n41409 = ( n16990 & ~n17124 ) | ( n16990 & n41408 ) | ( ~n17124 & n41408 ) ;
  assign n41407 = n2173 & ~n30280 ;
  assign n41410 = n41409 ^ n41407 ^ 1'b0 ;
  assign n41411 = n5129 & ~n31963 ;
  assign n41412 = n41411 ^ n12923 ^ 1'b0 ;
  assign n41413 = n40804 & ~n41412 ;
  assign n41414 = n18724 ^ n4767 ^ 1'b0 ;
  assign n41415 = n4828 | n41414 ;
  assign n41416 = n13505 ^ n2587 ^ 1'b0 ;
  assign n41417 = ~n1969 & n10764 ;
  assign n41418 = n26725 ^ n1059 ^ 1'b0 ;
  assign n41419 = ( n41416 & n41417 ) | ( n41416 & ~n41418 ) | ( n41417 & ~n41418 ) ;
  assign n41420 = n20349 ^ n7000 ^ 1'b0 ;
  assign n41421 = n15326 ^ n7185 ^ 1'b0 ;
  assign n41422 = n19681 | n41421 ;
  assign n41423 = n41422 ^ n5391 ^ 1'b0 ;
  assign n41424 = n31823 & ~n41423 ;
  assign n41425 = ~n2900 & n21898 ;
  assign n41426 = n41425 ^ n19748 ^ 1'b0 ;
  assign n41427 = n41426 ^ n29823 ^ 1'b0 ;
  assign n41428 = n40021 ^ n16194 ^ n4033 ;
  assign n41429 = n34062 ^ n31117 ^ n9396 ;
  assign n41430 = ~n20375 & n25647 ;
  assign n41431 = ~n18503 & n41430 ;
  assign n41432 = ~n32270 & n38792 ;
  assign n41433 = n41432 ^ n26922 ^ 1'b0 ;
  assign n41434 = n14790 ^ n4418 ^ 1'b0 ;
  assign n41435 = n500 & ~n17518 ;
  assign n41436 = n41434 & n41435 ;
  assign n41437 = n19561 & ~n35172 ;
  assign n41438 = ( n7109 & n29019 ) | ( n7109 & ~n35826 ) | ( n29019 & ~n35826 ) ;
  assign n41440 = n16396 | n19140 ;
  assign n41441 = n26112 | n41440 ;
  assign n41442 = n3972 | n41441 ;
  assign n41443 = n41442 ^ n15971 ^ n5313 ;
  assign n41439 = n32804 ^ n8386 ^ 1'b0 ;
  assign n41444 = n41443 ^ n41439 ^ n23518 ;
  assign n41445 = ( n12524 & n27096 ) | ( n12524 & ~n37699 ) | ( n27096 & ~n37699 ) ;
  assign n41446 = n14289 & ~n22588 ;
  assign n41447 = n41446 ^ n34141 ^ 1'b0 ;
  assign n41448 = n3367 & ~n24838 ;
  assign n41449 = n15277 & n41448 ;
  assign n41450 = n15322 ^ n2469 ^ 1'b0 ;
  assign n41451 = n4977 & ~n41450 ;
  assign n41452 = n22494 ^ n13318 ^ 1'b0 ;
  assign n41453 = ~n35300 & n41452 ;
  assign n41454 = ( n9232 & ~n16628 ) | ( n9232 & n41453 ) | ( ~n16628 & n41453 ) ;
  assign n41455 = n41454 ^ n20828 ^ 1'b0 ;
  assign n41456 = n41451 & ~n41455 ;
  assign n41457 = n10600 | n19465 ;
  assign n41458 = n36548 & ~n41457 ;
  assign n41459 = n19052 & n32348 ;
  assign n41460 = n3650 ^ n1153 ^ 1'b0 ;
  assign n41461 = n41460 ^ n1984 ^ 1'b0 ;
  assign n41462 = n34129 | n41461 ;
  assign n41465 = n28057 ^ n987 ^ 1'b0 ;
  assign n41466 = n23041 | n41465 ;
  assign n41463 = n29431 ^ n3712 ^ 1'b0 ;
  assign n41464 = n28878 | n41463 ;
  assign n41467 = n41466 ^ n41464 ^ 1'b0 ;
  assign n41468 = n5918 | n41467 ;
  assign n41469 = n41462 & n41468 ;
  assign n41470 = n41469 ^ n21004 ^ 1'b0 ;
  assign n41474 = ~n1396 & n23670 ;
  assign n41475 = n41474 ^ n22787 ^ 1'b0 ;
  assign n41471 = n26656 ^ n15168 ^ n5161 ;
  assign n41472 = n41471 ^ n40955 ^ 1'b0 ;
  assign n41473 = n41472 ^ n33531 ^ 1'b0 ;
  assign n41476 = n41475 ^ n41473 ^ n34992 ;
  assign n41481 = n5420 & n12420 ;
  assign n41482 = n41481 ^ n40230 ^ 1'b0 ;
  assign n41477 = n5028 & ~n14038 ;
  assign n41478 = n41477 ^ n36877 ^ 1'b0 ;
  assign n41479 = ( n721 & n15723 ) | ( n721 & ~n41478 ) | ( n15723 & ~n41478 ) ;
  assign n41480 = n10088 | n41479 ;
  assign n41483 = n41482 ^ n41480 ^ 1'b0 ;
  assign n41484 = ~n8833 & n24482 ;
  assign n41485 = n41484 ^ n29133 ^ 1'b0 ;
  assign n41486 = ~n19694 & n41485 ;
  assign n41487 = ~n2118 & n41486 ;
  assign n41488 = n26979 ^ n20156 ^ 1'b0 ;
  assign n41489 = n11070 & n41488 ;
  assign n41490 = ~n32204 & n41489 ;
  assign n41491 = n41487 & n41490 ;
  assign n41492 = n31021 | n36194 ;
  assign n41493 = n5732 & ~n41492 ;
  assign n41494 = ~n1685 & n16410 ;
  assign n41495 = ( n790 & n36450 ) | ( n790 & n41494 ) | ( n36450 & n41494 ) ;
  assign n41496 = n24329 ^ n1519 ^ 1'b0 ;
  assign n41497 = n2299 & ~n41496 ;
  assign n41498 = n1546 | n19737 ;
  assign n41499 = n13192 & n29914 ;
  assign n41500 = n1673 & n26704 ;
  assign n41501 = n20976 | n29902 ;
  assign n41502 = n41501 ^ n2299 ^ 1'b0 ;
  assign n41503 = n31330 ^ n14764 ^ 1'b0 ;
  assign n41504 = n41502 & ~n41503 ;
  assign n41505 = n4256 | n7794 ;
  assign n41506 = n41505 ^ n36716 ^ 1'b0 ;
  assign n41507 = n19404 | n22062 ;
  assign n41508 = n6372 & ~n7663 ;
  assign n41509 = n29093 & n41508 ;
  assign n41510 = n23205 & n23903 ;
  assign n41511 = n41510 ^ n5546 ^ 1'b0 ;
  assign n41512 = n915 & ~n12360 ;
  assign n41514 = n9341 ^ n2124 ^ x157 ;
  assign n41513 = n4800 | n7148 ;
  assign n41515 = n41514 ^ n41513 ^ 1'b0 ;
  assign n41516 = n13494 & ~n41515 ;
  assign n41517 = n13446 & n34718 ;
  assign n41518 = ~n17022 & n41517 ;
  assign n41519 = n41518 ^ n11030 ^ 1'b0 ;
  assign n41520 = n41519 ^ n32316 ^ n20932 ;
  assign n41521 = n10498 ^ n10447 ^ 1'b0 ;
  assign n41522 = n41521 ^ n4135 ^ 1'b0 ;
  assign n41523 = n2956 & ~n41522 ;
  assign n41524 = ~n17748 & n41523 ;
  assign n41525 = n1559 & ~n12974 ;
  assign n41526 = ~n15398 & n25245 ;
  assign n41527 = ( n1027 & n13717 ) | ( n1027 & ~n19099 ) | ( n13717 & ~n19099 ) ;
  assign n41528 = ~n6149 & n21504 ;
  assign n41529 = n41527 & n41528 ;
  assign n41530 = ( ~n2250 & n13621 ) | ( ~n2250 & n31518 ) | ( n13621 & n31518 ) ;
  assign n41531 = n41530 ^ n1313 ^ 1'b0 ;
  assign n41532 = n22552 & ~n41531 ;
  assign n41533 = n19503 & n30828 ;
  assign n41534 = n14917 & n24585 ;
  assign n41535 = ~n37916 & n41534 ;
  assign n41536 = n17435 & n35666 ;
  assign n41537 = ( n4913 & n13140 ) | ( n4913 & n41536 ) | ( n13140 & n41536 ) ;
  assign n41538 = ~n3156 & n26273 ;
  assign n41539 = n33937 & n41538 ;
  assign n41540 = n15158 & ~n34424 ;
  assign n41541 = ~n29597 & n41540 ;
  assign n41542 = n19702 | n19738 ;
  assign n41543 = n35637 & n36926 ;
  assign n41544 = ~n2577 & n36565 ;
  assign n41545 = ~n21457 & n41544 ;
  assign n41546 = n4977 & ~n32534 ;
  assign n41548 = n20777 ^ n19438 ^ 1'b0 ;
  assign n41549 = n41383 & ~n41548 ;
  assign n41547 = ~n5008 & n13458 ;
  assign n41550 = n41549 ^ n41547 ^ 1'b0 ;
  assign n41551 = n23380 ^ n854 ^ 1'b0 ;
  assign n41552 = x208 & ~n2795 ;
  assign n41553 = ~n41551 & n41552 ;
  assign n41554 = n41553 ^ n16972 ^ 1'b0 ;
  assign n41555 = n5217 & n33469 ;
  assign n41556 = n41555 ^ n24606 ^ 1'b0 ;
  assign n41557 = ~n23915 & n35004 ;
  assign n41558 = n41557 ^ n33278 ^ 1'b0 ;
  assign n41559 = n2635 & ~n11251 ;
  assign n41560 = ( n10125 & n32092 ) | ( n10125 & ~n32519 ) | ( n32092 & ~n32519 ) ;
  assign n41564 = n1489 | n15314 ;
  assign n41561 = n12713 & ~n19469 ;
  assign n41562 = n34133 ^ n1847 ^ 1'b0 ;
  assign n41563 = n41561 & ~n41562 ;
  assign n41565 = n41564 ^ n41563 ^ n16427 ;
  assign n41566 = ( n4353 & ~n13077 ) | ( n4353 & n26204 ) | ( ~n13077 & n26204 ) ;
  assign n41567 = n10252 | n25781 ;
  assign n41568 = n40207 | n41567 ;
  assign n41569 = n17568 & n30922 ;
  assign n41570 = ~n4241 & n20694 ;
  assign n41571 = n13668 & ~n41570 ;
  assign n41572 = n41571 ^ n30572 ^ 1'b0 ;
  assign n41573 = n673 | n2376 ;
  assign n41574 = n41573 ^ n342 ^ 1'b0 ;
  assign n41575 = n6903 & n26933 ;
  assign n41576 = ~n11285 & n41575 ;
  assign n41578 = n20738 ^ n16735 ^ n3912 ;
  assign n41577 = n12417 | n38444 ;
  assign n41579 = n41578 ^ n41577 ^ 1'b0 ;
  assign n41580 = n6188 ^ n1145 ^ 1'b0 ;
  assign n41581 = ~n5857 & n26049 ;
  assign n41582 = n41581 ^ n21350 ^ 1'b0 ;
  assign n41583 = ~n9394 & n30836 ;
  assign n41584 = ~n22159 & n41583 ;
  assign n41585 = n41584 ^ n19893 ^ 1'b0 ;
  assign n41586 = n6493 ^ n2623 ^ 1'b0 ;
  assign n41587 = n17578 ^ n2181 ^ 1'b0 ;
  assign n41588 = n19640 | n41587 ;
  assign n41589 = ~n41586 & n41588 ;
  assign n41590 = n1518 & ~n11039 ;
  assign n41591 = ~n15936 & n41590 ;
  assign n41592 = n41591 ^ n33345 ^ n23226 ;
  assign n41593 = n4996 & ~n25320 ;
  assign n41594 = n16959 & ~n41593 ;
  assign n41595 = n1147 & ~n25724 ;
  assign n41596 = n41595 ^ n1689 ^ 1'b0 ;
  assign n41597 = n25800 ^ n10217 ^ 1'b0 ;
  assign n41599 = ~n5391 & n21264 ;
  assign n41598 = n5129 & n32641 ;
  assign n41600 = n41599 ^ n41598 ^ 1'b0 ;
  assign n41601 = ( ~n547 & n32012 ) | ( ~n547 & n37909 ) | ( n32012 & n37909 ) ;
  assign n41602 = n3382 | n16651 ;
  assign n41603 = n32707 & n41602 ;
  assign n41604 = n31092 ^ n8551 ^ 1'b0 ;
  assign n41605 = n9169 ^ n7925 ^ 1'b0 ;
  assign n41606 = n9456 ^ n2759 ^ 1'b0 ;
  assign n41607 = ( ~n6455 & n12126 ) | ( ~n6455 & n41606 ) | ( n12126 & n41606 ) ;
  assign n41608 = n919 | n41607 ;
  assign n41609 = ( n12265 & ~n14270 ) | ( n12265 & n27735 ) | ( ~n14270 & n27735 ) ;
  assign n41610 = n41609 ^ n10311 ^ 1'b0 ;
  assign n41611 = n38359 & ~n41610 ;
  assign n41613 = n7481 | n11658 ;
  assign n41612 = n6514 & n37158 ;
  assign n41614 = n41613 ^ n41612 ^ 1'b0 ;
  assign n41615 = n41614 ^ n780 ^ 1'b0 ;
  assign n41616 = ~n11640 & n41615 ;
  assign n41622 = n2801 & ~n17388 ;
  assign n41623 = n41622 ^ n30722 ^ 1'b0 ;
  assign n41617 = n16703 ^ n7622 ^ 1'b0 ;
  assign n41618 = n10371 & ~n41617 ;
  assign n41619 = ~n9767 & n41618 ;
  assign n41620 = ~n27411 & n41619 ;
  assign n41621 = n2757 & ~n41620 ;
  assign n41624 = n41623 ^ n41621 ^ 1'b0 ;
  assign n41625 = n399 & ~n33866 ;
  assign n41626 = n33903 & n41625 ;
  assign n41627 = ~x0 & n23102 ;
  assign n41628 = n15715 ^ n14538 ^ 1'b0 ;
  assign n41629 = ~n3304 & n27644 ;
  assign n41630 = n41629 ^ n7810 ^ 1'b0 ;
  assign n41631 = n7314 | n37734 ;
  assign n41632 = n8565 | n41631 ;
  assign n41633 = n39961 & ~n40595 ;
  assign n41634 = n41633 ^ n8141 ^ 1'b0 ;
  assign n41635 = n5658 & ~n5864 ;
  assign n41636 = n17815 & ~n29573 ;
  assign n41637 = ( ~n16454 & n23981 ) | ( ~n16454 & n29209 ) | ( n23981 & n29209 ) ;
  assign n41638 = n13216 ^ n967 ^ 1'b0 ;
  assign n41639 = n25360 ^ n1596 ^ 1'b0 ;
  assign n41640 = ~n428 & n41639 ;
  assign n41641 = ( n4340 & n11631 ) | ( n4340 & n41640 ) | ( n11631 & n41640 ) ;
  assign n41642 = ~n17124 & n41641 ;
  assign n41643 = n41638 & n41642 ;
  assign n41644 = n17714 & n26150 ;
  assign n41645 = ~n16912 & n30192 ;
  assign n41646 = n41645 ^ n6371 ^ 1'b0 ;
  assign n41647 = n37955 & ~n41646 ;
  assign n41648 = n16170 ^ n8585 ^ 1'b0 ;
  assign n41650 = ~n9073 & n11239 ;
  assign n41649 = n32903 | n36425 ;
  assign n41651 = n41650 ^ n41649 ^ 1'b0 ;
  assign n41652 = n41651 ^ n36001 ^ 1'b0 ;
  assign n41653 = n12256 & ~n41652 ;
  assign n41654 = n41416 ^ n3059 ^ 1'b0 ;
  assign n41655 = n28303 ^ n23225 ^ n18565 ;
  assign n41656 = ( n3229 & n38362 ) | ( n3229 & ~n41655 ) | ( n38362 & ~n41655 ) ;
  assign n41657 = n12908 & n32900 ;
  assign n41658 = ( n1961 & n18018 ) | ( n1961 & n28516 ) | ( n18018 & n28516 ) ;
  assign n41659 = n36825 ^ n18375 ^ 1'b0 ;
  assign n41660 = n15025 | n41659 ;
  assign n41661 = n41658 | n41660 ;
  assign n41662 = n35823 ^ n6196 ^ 1'b0 ;
  assign n41663 = n9891 & ~n19102 ;
  assign n41664 = n41663 ^ n5146 ^ 1'b0 ;
  assign n41665 = n41664 ^ n26922 ^ n20611 ;
  assign n41666 = n19237 & ~n41665 ;
  assign n41667 = n39977 ^ n9973 ^ n6857 ;
  assign n41668 = ~n8014 & n41667 ;
  assign n41669 = n21276 ^ n19982 ^ 1'b0 ;
  assign n41670 = ~n34591 & n41669 ;
  assign n41671 = ~n13144 & n41670 ;
  assign n41672 = ~n16126 & n41671 ;
  assign n41673 = n7508 ^ n6257 ^ 1'b0 ;
  assign n41674 = n40372 ^ n29458 ^ 1'b0 ;
  assign n41675 = ( n14558 & n18623 ) | ( n14558 & n20196 ) | ( n18623 & n20196 ) ;
  assign n41676 = n19455 ^ x227 ^ 1'b0 ;
  assign n41677 = n8932 & ~n13795 ;
  assign n41678 = n12594 & ~n41677 ;
  assign n41679 = ~n22172 & n41678 ;
  assign n41680 = n3560 & ~n41679 ;
  assign n41681 = ~n25663 & n35329 ;
  assign n41682 = n38655 ^ n8539 ^ 1'b0 ;
  assign n41683 = n11080 & ~n18723 ;
  assign n41684 = ~n3126 & n41683 ;
  assign n41685 = n3411 & n8772 ;
  assign n41686 = n41685 ^ n21494 ^ 1'b0 ;
  assign n41687 = n25531 ^ n21377 ^ 1'b0 ;
  assign n41688 = ~n7282 & n41687 ;
  assign n41689 = n6352 & n33452 ;
  assign n41690 = ( n24060 & n29833 ) | ( n24060 & n41689 ) | ( n29833 & n41689 ) ;
  assign n41691 = n11333 ^ n7687 ^ n1823 ;
  assign n41693 = n886 | n4049 ;
  assign n41694 = n5610 & ~n41693 ;
  assign n41692 = ~n14677 & n15990 ;
  assign n41695 = n41694 ^ n41692 ^ n22755 ;
  assign n41696 = ~n2272 & n22976 ;
  assign n41697 = n24482 | n25728 ;
  assign n41698 = n27211 & n28680 ;
  assign n41699 = n41698 ^ n6388 ^ 1'b0 ;
  assign n41700 = n12074 | n23388 ;
  assign n41701 = n7788 & ~n41700 ;
  assign n41702 = n4880 | n12460 ;
  assign n41703 = n41701 & ~n41702 ;
  assign n41704 = n3624 | n41703 ;
  assign n41705 = n41704 ^ n23365 ^ 1'b0 ;
  assign n41706 = n13957 | n13988 ;
  assign n41707 = n2440 & ~n41706 ;
  assign n41708 = n11435 ^ n4208 ^ 1'b0 ;
  assign n41709 = n1913 & n41708 ;
  assign n41710 = n10374 | n41709 ;
  assign n41711 = n19204 & ~n28477 ;
  assign n41712 = ~n41710 & n41711 ;
  assign n41713 = ( n24017 & n41707 ) | ( n24017 & n41712 ) | ( n41707 & n41712 ) ;
  assign n41714 = n21075 ^ n8187 ^ n6185 ;
  assign n41715 = ( n2054 & n19278 ) | ( n2054 & ~n41714 ) | ( n19278 & ~n41714 ) ;
  assign n41716 = n14239 ^ n1337 ^ 1'b0 ;
  assign n41717 = ( ~n6517 & n17256 ) | ( ~n6517 & n41716 ) | ( n17256 & n41716 ) ;
  assign n41718 = n41717 ^ n29965 ^ n21093 ;
  assign n41719 = n7876 | n16296 ;
  assign n41720 = n33907 & ~n41719 ;
  assign n41721 = n1263 | n24337 ;
  assign n41722 = ~n18534 & n41721 ;
  assign n41723 = ~n17164 & n41722 ;
  assign n41724 = n30316 ^ n29002 ^ 1'b0 ;
  assign n41725 = n674 & n2253 ;
  assign n41726 = n673 ^ x74 ^ 1'b0 ;
  assign n41727 = ~n4947 & n41726 ;
  assign n41728 = n3343 | n41727 ;
  assign n41729 = n35517 ^ n7210 ^ 1'b0 ;
  assign n41734 = n1733 & n13157 ;
  assign n41735 = n41734 ^ n33480 ^ 1'b0 ;
  assign n41736 = n8899 | n41735 ;
  assign n41730 = n32634 | n36359 ;
  assign n41731 = n41730 ^ n27324 ^ 1'b0 ;
  assign n41732 = ~n13291 & n41731 ;
  assign n41733 = n41732 ^ n12171 ^ 1'b0 ;
  assign n41737 = n41736 ^ n41733 ^ n11540 ;
  assign n41738 = n36720 ^ n18006 ^ 1'b0 ;
  assign n41739 = n3692 | n9925 ;
  assign n41740 = n39578 & ~n41739 ;
  assign n41741 = n37566 ^ n7190 ^ n1323 ;
  assign n41742 = ~n8972 & n35477 ;
  assign n41743 = ~n31655 & n41742 ;
  assign n41744 = n41743 ^ n36072 ^ 1'b0 ;
  assign n41745 = n41741 & ~n41744 ;
  assign n41746 = n15196 | n41745 ;
  assign n41747 = n21793 ^ n5372 ^ 1'b0 ;
  assign n41748 = n38455 & ~n41485 ;
  assign n41749 = n26215 & ~n39073 ;
  assign n41750 = ~n7214 & n41749 ;
  assign n41752 = n22992 ^ n610 ^ 1'b0 ;
  assign n41751 = ~n4256 & n26192 ;
  assign n41753 = n41752 ^ n41751 ^ 1'b0 ;
  assign n41754 = n17397 ^ n12766 ^ 1'b0 ;
  assign n41755 = ~n20515 & n41754 ;
  assign n41756 = n9708 ^ n3271 ^ 1'b0 ;
  assign n41757 = n9544 & n41756 ;
  assign n41758 = ~n9561 & n41757 ;
  assign n41761 = n1453 ^ n1270 ^ 1'b0 ;
  assign n41762 = n12707 & n41761 ;
  assign n41763 = ~n41761 & n41762 ;
  assign n41759 = n40198 ^ n20117 ^ n5255 ;
  assign n41760 = n7123 & n41759 ;
  assign n41764 = n41763 ^ n41760 ^ 1'b0 ;
  assign n41765 = ~n14479 & n16398 ;
  assign n41766 = n14750 & n41765 ;
  assign n41767 = n36486 ^ n20700 ^ 1'b0 ;
  assign n41768 = n41766 | n41767 ;
  assign n41769 = n31704 ^ n14828 ^ 1'b0 ;
  assign n41770 = n37052 ^ n14713 ^ n10932 ;
  assign n41771 = ( n2483 & ~n4626 ) | ( n2483 & n40780 ) | ( ~n4626 & n40780 ) ;
  assign n41772 = n22370 ^ n3633 ^ 1'b0 ;
  assign n41773 = n15430 ^ n4561 ^ 1'b0 ;
  assign n41774 = ~n8201 & n41773 ;
  assign n41775 = ~n34568 & n41774 ;
  assign n41776 = ~n15467 & n41373 ;
  assign n41777 = n41776 ^ n9916 ^ 1'b0 ;
  assign n41778 = n9686 | n41777 ;
  assign n41779 = ( ~n5829 & n10964 ) | ( ~n5829 & n20747 ) | ( n10964 & n20747 ) ;
  assign n41780 = n7318 | n35191 ;
  assign n41781 = n41779 | n41780 ;
  assign n41782 = ~n1763 & n34825 ;
  assign n41783 = n27258 & n41782 ;
  assign n41784 = n5037 ^ n908 ^ 1'b0 ;
  assign n41785 = n41784 ^ n19822 ^ n11864 ;
  assign n41786 = n9155 & ~n32022 ;
  assign n41787 = n2829 | n30020 ;
  assign n41788 = n4626 & ~n41787 ;
  assign n41789 = n41788 ^ n14133 ^ n4777 ;
  assign n41790 = n41789 ^ n29915 ^ n1217 ;
  assign n41791 = n25509 ^ n21390 ^ n17230 ;
  assign n41792 = n28739 ^ n8711 ^ n610 ;
  assign n41793 = n32790 ^ n11888 ^ 1'b0 ;
  assign n41794 = n9172 | n41793 ;
  assign n41795 = n41794 ^ n8125 ^ 1'b0 ;
  assign n41799 = n9726 | n11196 ;
  assign n41796 = n15241 | n24148 ;
  assign n41797 = n21060 & ~n41796 ;
  assign n41798 = n4929 & ~n41797 ;
  assign n41800 = n41799 ^ n41798 ^ 1'b0 ;
  assign n41801 = n3889 ^ n1646 ^ n441 ;
  assign n41802 = n20783 & ~n41801 ;
  assign n41803 = ( n15737 & n18628 ) | ( n15737 & ~n26405 ) | ( n18628 & ~n26405 ) ;
  assign n41804 = n41803 ^ n10273 ^ 1'b0 ;
  assign n41805 = n13907 | n41804 ;
  assign n41806 = n23218 & ~n41805 ;
  assign n41807 = ~n15002 & n41806 ;
  assign n41808 = ~n18818 & n32482 ;
  assign n41809 = ~n1527 & n41808 ;
  assign n41810 = n18350 ^ n8790 ^ 1'b0 ;
  assign n41811 = n10855 & n41810 ;
  assign n41812 = n11852 | n14258 ;
  assign n41813 = n41812 ^ n20185 ^ n13887 ;
  assign n41814 = ( n35223 & n41811 ) | ( n35223 & n41813 ) | ( n41811 & n41813 ) ;
  assign n41818 = n14683 ^ x100 ^ 1'b0 ;
  assign n41815 = n4694 | n28819 ;
  assign n41816 = n29484 ^ n9734 ^ 1'b0 ;
  assign n41817 = n41815 | n41816 ;
  assign n41819 = n41818 ^ n41817 ^ n5748 ;
  assign n41820 = ~n15389 & n26488 ;
  assign n41821 = n41820 ^ n13854 ^ 1'b0 ;
  assign n41822 = n3747 & n41821 ;
  assign n41824 = ~n4936 & n7546 ;
  assign n41823 = ( n1110 & ~n1590 ) | ( n1110 & n7678 ) | ( ~n1590 & n7678 ) ;
  assign n41825 = n41824 ^ n41823 ^ n5785 ;
  assign n41826 = n19462 ^ n5770 ^ 1'b0 ;
  assign n41827 = n12293 | n41826 ;
  assign n41828 = n39801 | n41827 ;
  assign n41829 = n41825 & ~n41828 ;
  assign n41830 = n39576 ^ n23427 ^ 1'b0 ;
  assign n41831 = n31634 & ~n41830 ;
  assign n41835 = n24277 ^ n3210 ^ 1'b0 ;
  assign n41836 = n41835 ^ n41422 ^ 1'b0 ;
  assign n41832 = n17817 & ~n31420 ;
  assign n41833 = n41832 ^ n6029 ^ 1'b0 ;
  assign n41834 = n28559 & n41833 ;
  assign n41837 = n41836 ^ n41834 ^ 1'b0 ;
  assign n41838 = n41837 ^ n6481 ^ 1'b0 ;
  assign n41839 = n3085 | n18987 ;
  assign n41840 = n41839 ^ n20269 ^ 1'b0 ;
  assign n41841 = n9782 | n41840 ;
  assign n41842 = n15168 ^ n1102 ^ 1'b0 ;
  assign n41843 = ~n1350 & n32365 ;
  assign n41844 = ( ~n29720 & n38696 ) | ( ~n29720 & n41843 ) | ( n38696 & n41843 ) ;
  assign n41845 = n12697 & ~n16820 ;
  assign n41847 = n20420 ^ n18253 ^ 1'b0 ;
  assign n41846 = n27958 & n40220 ;
  assign n41848 = n41847 ^ n41846 ^ 1'b0 ;
  assign n41849 = n22486 ^ n6779 ^ 1'b0 ;
  assign n41850 = n23752 & n41849 ;
  assign n41851 = n6821 & n41850 ;
  assign n41852 = n434 | n25471 ;
  assign n41853 = n33336 & ~n41852 ;
  assign n41854 = n20302 ^ n7549 ^ 1'b0 ;
  assign n41855 = n25431 | n41854 ;
  assign n41856 = ~n7112 & n11007 ;
  assign n41857 = n29236 ^ n2698 ^ 1'b0 ;
  assign n41858 = ~n41856 & n41857 ;
  assign n41859 = ~n28216 & n38609 ;
  assign n41860 = n13812 ^ n671 ^ 1'b0 ;
  assign n41861 = n17161 ^ n12148 ^ 1'b0 ;
  assign n41862 = n8105 | n9490 ;
  assign n41863 = n32672 ^ n5063 ^ 1'b0 ;
  assign n41864 = x64 & n5569 ;
  assign n41865 = ~n8277 & n41864 ;
  assign n41867 = n21504 ^ n14030 ^ n2116 ;
  assign n41868 = n41867 ^ n38864 ^ n8748 ;
  assign n41866 = ~n20335 & n33389 ;
  assign n41869 = n41868 ^ n41866 ^ 1'b0 ;
  assign n41870 = n19180 ^ n10088 ^ 1'b0 ;
  assign n41871 = n28096 | n41870 ;
  assign n41872 = n7984 | n19670 ;
  assign n41873 = n755 & ~n36876 ;
  assign n41874 = ~n41872 & n41873 ;
  assign n41875 = n18686 & ~n41874 ;
  assign n41876 = n2627 & n41875 ;
  assign n41877 = n41871 & n41876 ;
  assign n41878 = n40407 ^ n33757 ^ 1'b0 ;
  assign n41879 = n24506 ^ n15281 ^ n8989 ;
  assign n41880 = n10515 ^ n7054 ^ 1'b0 ;
  assign n41881 = n6264 | n6452 ;
  assign n41882 = n4776 & ~n30543 ;
  assign n41883 = ( n41880 & n41881 ) | ( n41880 & n41882 ) | ( n41881 & n41882 ) ;
  assign n41884 = n26127 | n36572 ;
  assign n41885 = n41884 ^ n908 ^ 1'b0 ;
  assign n41886 = n18420 & ~n21681 ;
  assign n41887 = ~n7360 & n9820 ;
  assign n41888 = n41887 ^ n4792 ^ 1'b0 ;
  assign n41889 = n1004 | n41284 ;
  assign n41890 = n41889 ^ n11449 ^ 1'b0 ;
  assign n41891 = n7546 ^ n1343 ^ 1'b0 ;
  assign n41892 = n41891 ^ n34965 ^ 1'b0 ;
  assign n41893 = n9068 ^ n6688 ^ 1'b0 ;
  assign n41894 = ~n10688 & n41893 ;
  assign n41895 = ( ~n1166 & n6891 ) | ( ~n1166 & n41894 ) | ( n6891 & n41894 ) ;
  assign n41896 = n14479 & n15096 ;
  assign n41897 = n41896 ^ n33054 ^ n13056 ;
  assign n41898 = n2902 & ~n10947 ;
  assign n41899 = ( ~n24963 & n36393 ) | ( ~n24963 & n41898 ) | ( n36393 & n41898 ) ;
  assign n41900 = n22812 & n35858 ;
  assign n41901 = n32147 & ~n32626 ;
  assign n41903 = n2140 & n4160 ;
  assign n41904 = n41903 ^ n2586 ^ 1'b0 ;
  assign n41905 = n2384 | n41904 ;
  assign n41906 = n2882 | n41905 ;
  assign n41907 = ~n22806 & n41906 ;
  assign n41902 = n14773 | n35836 ;
  assign n41908 = n41907 ^ n41902 ^ 1'b0 ;
  assign n41909 = n10246 | n14016 ;
  assign n41910 = n28868 & ~n41909 ;
  assign n41911 = n41910 ^ n1110 ^ 1'b0 ;
  assign n41912 = n35845 & ~n40386 ;
  assign n41913 = n41912 ^ n27295 ^ 1'b0 ;
  assign n41914 = n17713 & n27548 ;
  assign n41915 = n1239 & ~n3501 ;
  assign n41916 = n26504 & ~n41915 ;
  assign n41917 = ~n3600 & n41916 ;
  assign n41918 = n407 | n707 ;
  assign n41919 = n26539 & n41918 ;
  assign n41920 = ~n5075 & n6459 ;
  assign n41921 = ( n29475 & n31588 ) | ( n29475 & n41920 ) | ( n31588 & n41920 ) ;
  assign n41922 = ( ~n5931 & n26245 ) | ( ~n5931 & n35004 ) | ( n26245 & n35004 ) ;
  assign n41923 = n21912 ^ n18775 ^ 1'b0 ;
  assign n41924 = n27295 & n41923 ;
  assign n41925 = n41924 ^ n22116 ^ 1'b0 ;
  assign n41926 = n10992 & n41925 ;
  assign n41927 = n20572 ^ n11583 ^ 1'b0 ;
  assign n41928 = n16700 ^ n1304 ^ 1'b0 ;
  assign n41929 = n529 | n41928 ;
  assign n41930 = n3445 | n41929 ;
  assign n41933 = n12900 & n17316 ;
  assign n41934 = ~n6880 & n41933 ;
  assign n41931 = n14470 ^ n5404 ^ 1'b0 ;
  assign n41932 = n19464 & ~n41931 ;
  assign n41935 = n41934 ^ n41932 ^ 1'b0 ;
  assign n41936 = ( n6435 & n37059 ) | ( n6435 & n41935 ) | ( n37059 & n41935 ) ;
  assign n41937 = n26787 ^ n3922 ^ 1'b0 ;
  assign n41938 = n18778 ^ n11591 ^ n7067 ;
  assign n41939 = ~n3716 & n38014 ;
  assign n41940 = n33732 ^ n12183 ^ 1'b0 ;
  assign n41941 = n23992 ^ n6312 ^ 1'b0 ;
  assign n41942 = ~n22924 & n41941 ;
  assign n41943 = ~n4060 & n24174 ;
  assign n41944 = n41943 ^ n13418 ^ 1'b0 ;
  assign n41945 = ~n11183 & n17417 ;
  assign n41946 = ~n41944 & n41945 ;
  assign n41947 = n15155 | n27780 ;
  assign n41948 = n41947 ^ n20319 ^ 1'b0 ;
  assign n41949 = n41948 ^ n18668 ^ 1'b0 ;
  assign n41950 = ( n3316 & n18013 ) | ( n3316 & ~n31354 ) | ( n18013 & ~n31354 ) ;
  assign n41951 = n11226 & n20372 ;
  assign n41952 = n41951 ^ n9079 ^ 1'b0 ;
  assign n41953 = n41952 ^ n34382 ^ 1'b0 ;
  assign n41954 = n41953 ^ n18930 ^ n12347 ;
  assign n41955 = n19202 | n36136 ;
  assign n41957 = n5804 | n10012 ;
  assign n41958 = n20245 & ~n41957 ;
  assign n41956 = n7439 & n12169 ;
  assign n41959 = n41958 ^ n41956 ^ 1'b0 ;
  assign n41960 = n6895 ^ n5798 ^ 1'b0 ;
  assign n41961 = n30945 | n41960 ;
  assign n41962 = ~n41959 & n41961 ;
  assign n41963 = n25935 ^ n18418 ^ 1'b0 ;
  assign n41964 = n275 & n8391 ;
  assign n41965 = n41964 ^ n9352 ^ 1'b0 ;
  assign n41966 = n33149 ^ n13766 ^ 1'b0 ;
  assign n41967 = n4872 & n31157 ;
  assign n41968 = n41966 & n41967 ;
  assign n41969 = n4150 | n10200 ;
  assign n41970 = n10962 & ~n41969 ;
  assign n41971 = ~n3742 & n41970 ;
  assign n41972 = n23985 & n30063 ;
  assign n41973 = n41972 ^ n5313 ^ 1'b0 ;
  assign n41974 = n6088 | n8369 ;
  assign n41975 = n1129 & n9651 ;
  assign n41976 = ( n4434 & n18636 ) | ( n4434 & ~n41975 ) | ( n18636 & ~n41975 ) ;
  assign n41977 = ( ~n6295 & n28291 ) | ( ~n6295 & n41976 ) | ( n28291 & n41976 ) ;
  assign n41978 = n41977 ^ n8708 ^ 1'b0 ;
  assign n41979 = n2337 & n41978 ;
  assign n41980 = n13766 & n31953 ;
  assign n41981 = n604 & n41980 ;
  assign n41982 = n26422 ^ n7850 ^ 1'b0 ;
  assign n41983 = n17629 & ~n31603 ;
  assign n41984 = n41983 ^ n8245 ^ 1'b0 ;
  assign n41985 = ( n2151 & n9401 ) | ( n2151 & n41984 ) | ( n9401 & n41984 ) ;
  assign n41986 = ( n8925 & n8978 ) | ( n8925 & n41985 ) | ( n8978 & n41985 ) ;
  assign n41990 = ~n4584 & n7843 ;
  assign n41991 = n2492 & n41990 ;
  assign n41987 = n23532 ^ n11692 ^ 1'b0 ;
  assign n41988 = n27545 | n41987 ;
  assign n41989 = n3292 & ~n41988 ;
  assign n41992 = n41991 ^ n41989 ^ n41966 ;
  assign n41993 = n441 & ~n3534 ;
  assign n41994 = n41993 ^ n2785 ^ 1'b0 ;
  assign n41995 = ( n21017 & ~n29788 ) | ( n21017 & n41994 ) | ( ~n29788 & n41994 ) ;
  assign n41997 = n5087 & ~n8145 ;
  assign n41996 = n4905 & n10093 ;
  assign n41998 = n41997 ^ n41996 ^ 1'b0 ;
  assign n41999 = n38810 ^ n15672 ^ 1'b0 ;
  assign n42000 = n30147 | n41999 ;
  assign n42001 = n8081 | n20712 ;
  assign n42002 = n42001 ^ n4339 ^ 1'b0 ;
  assign n42003 = n2076 | n13937 ;
  assign n42004 = n42002 | n42003 ;
  assign n42005 = n4150 ^ x220 ^ 1'b0 ;
  assign n42006 = n7339 & ~n42005 ;
  assign n42007 = n42006 ^ n27132 ^ 1'b0 ;
  assign n42008 = n10742 & ~n42007 ;
  assign n42009 = ~n3543 & n33978 ;
  assign n42010 = n42009 ^ n5517 ^ 1'b0 ;
  assign n42011 = n31629 ^ n24424 ^ n15369 ;
  assign n42012 = n42011 ^ n36411 ^ 1'b0 ;
  assign n42013 = n42012 ^ n37115 ^ n8274 ;
  assign n42014 = n24272 ^ n14110 ^ 1'b0 ;
  assign n42015 = n20908 & ~n35441 ;
  assign n42016 = n17011 & n31972 ;
  assign n42017 = n24215 ^ n606 ^ 1'b0 ;
  assign n42018 = n296 & n42017 ;
  assign n42019 = n4241 & n42018 ;
  assign n42020 = n24034 & n32611 ;
  assign n42021 = n25479 & n42020 ;
  assign n42022 = n18387 ^ x187 ^ 1'b0 ;
  assign n42023 = n12674 & n29473 ;
  assign n42027 = n19002 | n31638 ;
  assign n42028 = ~n21600 & n42027 ;
  assign n42024 = n2483 & ~n9483 ;
  assign n42025 = ~n34801 & n42024 ;
  assign n42026 = n42025 ^ n473 ^ 1'b0 ;
  assign n42029 = n42028 ^ n42026 ^ n24046 ;
  assign n42030 = n42029 ^ n27401 ^ n17627 ;
  assign n42031 = ( n29931 & ~n30857 ) | ( n29931 & n33651 ) | ( ~n30857 & n33651 ) ;
  assign n42032 = n41573 ^ n33984 ^ n14057 ;
  assign n42036 = n6341 & n8756 ;
  assign n42033 = n17473 ^ n8932 ^ 1'b0 ;
  assign n42034 = n42033 ^ n25039 ^ n13256 ;
  assign n42035 = ( n1943 & n41097 ) | ( n1943 & n42034 ) | ( n41097 & n42034 ) ;
  assign n42037 = n42036 ^ n42035 ^ 1'b0 ;
  assign n42038 = n27343 & n42037 ;
  assign n42039 = n29731 ^ n3827 ^ 1'b0 ;
  assign n42040 = n10888 & ~n42039 ;
  assign n42041 = n13750 & n29201 ;
  assign n42042 = n23645 ^ n2995 ^ 1'b0 ;
  assign n42043 = n18334 | n42042 ;
  assign n42044 = n14636 ^ n4614 ^ 1'b0 ;
  assign n42045 = ~n42043 & n42044 ;
  assign n42046 = ~n9672 & n25296 ;
  assign n42047 = n42046 ^ n39311 ^ n2718 ;
  assign n42048 = n36176 ^ n31171 ^ n10015 ;
  assign n42049 = ( n5965 & ~n6571 ) | ( n5965 & n11865 ) | ( ~n6571 & n11865 ) ;
  assign n42050 = ~n30281 & n42049 ;
  assign n42051 = n42050 ^ n16262 ^ 1'b0 ;
  assign n42052 = n14110 ^ n5711 ^ 1'b0 ;
  assign n42053 = n13955 | n42052 ;
  assign n42054 = n23253 | n42053 ;
  assign n42055 = n42054 ^ n36789 ^ 1'b0 ;
  assign n42056 = n4797 & n16251 ;
  assign n42057 = ~n10926 & n20359 ;
  assign n42058 = n23280 ^ n6281 ^ 1'b0 ;
  assign n42059 = n19398 | n20761 ;
  assign n42060 = n12799 & ~n42059 ;
  assign n42061 = n17807 & ~n29344 ;
  assign n42062 = n8704 & n42061 ;
  assign n42063 = ( n3727 & n42060 ) | ( n3727 & ~n42062 ) | ( n42060 & ~n42062 ) ;
  assign n42064 = n25887 ^ n22985 ^ n6371 ;
  assign n42065 = n13390 | n17124 ;
  assign n42066 = n16257 & ~n42065 ;
  assign n42067 = n6535 & n21530 ;
  assign n42068 = n2201 & n42067 ;
  assign n42069 = n13000 & n42068 ;
  assign n42070 = n4931 & ~n18642 ;
  assign n42071 = n42070 ^ n11849 ^ 1'b0 ;
  assign n42072 = ~n5396 & n42071 ;
  assign n42073 = n17373 ^ n6703 ^ n279 ;
  assign n42074 = n11137 | n42073 ;
  assign n42075 = n1792 & n4200 ;
  assign n42076 = n42075 ^ n5687 ^ 1'b0 ;
  assign n42077 = n42076 ^ n8198 ^ 1'b0 ;
  assign n42078 = n37173 | n42077 ;
  assign n42079 = ( n3545 & ~n3862 ) | ( n3545 & n5725 ) | ( ~n3862 & n5725 ) ;
  assign n42080 = n13780 & n18296 ;
  assign n42081 = ~n4638 & n42080 ;
  assign n42082 = n42081 ^ n25920 ^ n2384 ;
  assign n42083 = n17060 ^ n13324 ^ 1'b0 ;
  assign n42084 = ( n27852 & n35995 ) | ( n27852 & n42083 ) | ( n35995 & n42083 ) ;
  assign n42085 = n18629 ^ x142 ^ 1'b0 ;
  assign n42086 = n736 & ~n42085 ;
  assign n42087 = n29453 & n42086 ;
  assign n42088 = ~n2701 & n42087 ;
  assign n42089 = ~n14490 & n21856 ;
  assign n42090 = n4932 & n13446 ;
  assign n42091 = n42090 ^ n9660 ^ 1'b0 ;
  assign n42092 = ~n8119 & n41147 ;
  assign n42093 = n42092 ^ n8438 ^ 1'b0 ;
  assign n42094 = n5543 & ~n9161 ;
  assign n42095 = n579 & n42094 ;
  assign n42096 = n42095 ^ n1269 ^ 1'b0 ;
  assign n42097 = n768 & n8330 ;
  assign n42098 = ~n10702 & n42097 ;
  assign n42099 = n18392 & n20557 ;
  assign n42100 = n42099 ^ n41097 ^ n3490 ;
  assign n42101 = n1228 & n18292 ;
  assign n42102 = n42101 ^ n19962 ^ 1'b0 ;
  assign n42103 = x81 & n2471 ;
  assign n42104 = n5610 & n42103 ;
  assign n42108 = n13237 ^ n2569 ^ 1'b0 ;
  assign n42105 = n10011 ^ n2521 ^ 1'b0 ;
  assign n42106 = n26664 & n42105 ;
  assign n42107 = n3106 & n42106 ;
  assign n42109 = n42108 ^ n42107 ^ 1'b0 ;
  assign n42110 = n4213 & n16001 ;
  assign n42111 = n42110 ^ n1872 ^ 1'b0 ;
  assign n42112 = ~n30805 & n38088 ;
  assign n42113 = ~n4222 & n42112 ;
  assign n42114 = n31219 & n32079 ;
  assign n42115 = ~n11452 & n42114 ;
  assign n42116 = n1484 & ~n42115 ;
  assign n42117 = n3504 | n21593 ;
  assign n42118 = n2675 | n42117 ;
  assign n42119 = n42118 ^ n15455 ^ 1'b0 ;
  assign n42120 = n42116 & ~n42119 ;
  assign n42121 = n37630 | n40144 ;
  assign n42122 = n42121 ^ n4812 ^ 1'b0 ;
  assign n42123 = n10298 & n29458 ;
  assign n42124 = n42123 ^ n11111 ^ 1'b0 ;
  assign n42125 = n15351 | n42124 ;
  assign n42126 = n42125 ^ n22473 ^ n9638 ;
  assign n42127 = n15446 | n34818 ;
  assign n42128 = n7798 & n16415 ;
  assign n42129 = ~n6731 & n42128 ;
  assign n42130 = n20531 ^ n8695 ^ 1'b0 ;
  assign n42131 = n42129 | n42130 ;
  assign n42132 = ( n38093 & n42127 ) | ( n38093 & ~n42131 ) | ( n42127 & ~n42131 ) ;
  assign n42133 = ~n21627 & n27128 ;
  assign n42134 = n6124 & n42133 ;
  assign n42135 = ~n8637 & n13462 ;
  assign n42136 = n37044 & n42135 ;
  assign n42137 = n42136 ^ n10975 ^ 1'b0 ;
  assign n42138 = ( n8294 & n25294 ) | ( n8294 & ~n42137 ) | ( n25294 & ~n42137 ) ;
  assign n42139 = n42138 ^ n13609 ^ 1'b0 ;
  assign n42140 = n17782 ^ n17700 ^ 1'b0 ;
  assign n42141 = n42139 | n42140 ;
  assign n42142 = ~n2142 & n20285 ;
  assign n42143 = n19635 & n22691 ;
  assign n42144 = ~n29157 & n42143 ;
  assign n42145 = n42144 ^ n19322 ^ n12897 ;
  assign n42146 = n14669 ^ n2967 ^ 1'b0 ;
  assign n42147 = ~n4540 & n8977 ;
  assign n42148 = n42147 ^ n26178 ^ 1'b0 ;
  assign n42149 = n14477 & n42148 ;
  assign n42150 = n42149 ^ n3113 ^ 1'b0 ;
  assign n42151 = n2979 ^ x75 ^ 1'b0 ;
  assign n42152 = n1809 & n42151 ;
  assign n42154 = n9044 & ~n21853 ;
  assign n42155 = n21853 & n42154 ;
  assign n42153 = n37569 | n40823 ;
  assign n42156 = n42155 ^ n42153 ^ 1'b0 ;
  assign n42157 = n16402 & n39188 ;
  assign n42158 = n42157 ^ n4257 ^ 1'b0 ;
  assign n42159 = ~n20798 & n25694 ;
  assign n42160 = n1033 & n25947 ;
  assign n42161 = n42160 ^ n2006 ^ 1'b0 ;
  assign n42162 = n1015 & n29475 ;
  assign n42163 = n42162 ^ n17350 ^ n10472 ;
  assign n42164 = n22564 ^ n13915 ^ n4924 ;
  assign n42165 = n9783 ^ n8589 ^ 1'b0 ;
  assign n42166 = n18085 & ~n42165 ;
  assign n42167 = n11324 | n28681 ;
  assign n42168 = n30335 & ~n42167 ;
  assign n42169 = n29604 ^ n28140 ^ 1'b0 ;
  assign n42170 = n42169 ^ n9220 ^ n1496 ;
  assign n42171 = n24361 ^ n7578 ^ 1'b0 ;
  assign n42172 = n42170 & n42171 ;
  assign n42173 = ~n2789 & n3550 ;
  assign n42174 = ~n13056 & n42173 ;
  assign n42175 = n42174 ^ n18194 ^ 1'b0 ;
  assign n42176 = n14909 | n22338 ;
  assign n42177 = n42176 ^ n6483 ^ 1'b0 ;
  assign n42178 = ~n34819 & n40077 ;
  assign n42179 = n42178 ^ n27284 ^ 1'b0 ;
  assign n42180 = n39712 ^ n18925 ^ 1'b0 ;
  assign n42181 = n30036 ^ n320 ^ 1'b0 ;
  assign n42182 = n42181 ^ n9298 ^ n7326 ;
  assign n42183 = n42182 ^ n9884 ^ 1'b0 ;
  assign n42184 = n20688 & ~n42183 ;
  assign n42185 = n42184 ^ n1055 ^ x15 ;
  assign n42186 = n17226 ^ n10339 ^ n7325 ;
  assign n42187 = n1875 & n38284 ;
  assign n42188 = ( n608 & n25244 ) | ( n608 & n31490 ) | ( n25244 & n31490 ) ;
  assign n42189 = n14115 ^ x25 ^ 1'b0 ;
  assign n42190 = ~n42188 & n42189 ;
  assign n42191 = n42190 ^ n4561 ^ n3202 ;
  assign n42192 = n42191 ^ n23303 ^ 1'b0 ;
  assign n42193 = n39166 ^ n27232 ^ 1'b0 ;
  assign n42194 = n6859 | n42193 ;
  assign n42195 = n42194 ^ n37746 ^ 1'b0 ;
  assign n42196 = n3005 & n17483 ;
  assign n42197 = n2817 ^ n1858 ^ 1'b0 ;
  assign n42198 = ~n41549 & n42197 ;
  assign n42199 = ~n1409 & n1486 ;
  assign n42200 = n42199 ^ n20524 ^ 1'b0 ;
  assign n42201 = n27178 & ~n42200 ;
  assign n42202 = n42201 ^ n6717 ^ 1'b0 ;
  assign n42203 = n21185 | n42202 ;
  assign n42204 = n7559 | n42203 ;
  assign n42205 = n15960 ^ n2544 ^ x203 ;
  assign n42206 = n38116 ^ n28828 ^ 1'b0 ;
  assign n42207 = n14851 ^ n13832 ^ 1'b0 ;
  assign n42208 = ~n7573 & n13584 ;
  assign n42209 = n14439 | n42208 ;
  assign n42210 = n23472 ^ n6926 ^ 1'b0 ;
  assign n42211 = n42209 & ~n42210 ;
  assign n42212 = ~n3430 & n30643 ;
  assign n42213 = ~n27003 & n42212 ;
  assign n42214 = ~n2165 & n14662 ;
  assign n42215 = n31003 & n42214 ;
  assign n42216 = n14138 ^ n7830 ^ 1'b0 ;
  assign n42217 = n18831 ^ n13475 ^ n3359 ;
  assign n42218 = n8735 | n42217 ;
  assign n42219 = n24151 | n35076 ;
  assign n42220 = ~n31029 & n42219 ;
  assign n42221 = n1001 & ~n18736 ;
  assign n42222 = n2968 & n42221 ;
  assign n42223 = ( ~n6819 & n17053 ) | ( ~n6819 & n32718 ) | ( n17053 & n32718 ) ;
  assign n42224 = n42223 ^ n30884 ^ x7 ;
  assign n42225 = n11735 ^ n2024 ^ 1'b0 ;
  assign n42226 = n42224 & n42225 ;
  assign n42227 = ~n6389 & n14867 ;
  assign n42228 = n2588 | n10723 ;
  assign n42229 = n9902 | n42228 ;
  assign n42230 = ~n2521 & n5802 ;
  assign n42231 = n8833 | n42230 ;
  assign n42232 = n23402 | n28883 ;
  assign n42233 = n4976 | n42232 ;
  assign n42234 = n42233 ^ n3782 ^ 1'b0 ;
  assign n42235 = ~n42231 & n42234 ;
  assign n42239 = n1439 | n13218 ;
  assign n42236 = n22534 ^ n9645 ^ 1'b0 ;
  assign n42237 = n9331 & ~n42236 ;
  assign n42238 = ~n3814 & n42237 ;
  assign n42240 = n42239 ^ n42238 ^ 1'b0 ;
  assign n42241 = n9997 | n24120 ;
  assign n42242 = n15529 | n32620 ;
  assign n42243 = n42242 ^ n8860 ^ n7593 ;
  assign n42244 = n2982 & ~n9470 ;
  assign n42245 = n42244 ^ n26218 ^ 1'b0 ;
  assign n42246 = n42245 ^ n23815 ^ n17958 ;
  assign n42247 = n3124 & n35920 ;
  assign n42248 = n42247 ^ n27156 ^ n20382 ;
  assign n42252 = n33547 | n40756 ;
  assign n42253 = n42252 ^ n12547 ^ 1'b0 ;
  assign n42249 = ~n10405 & n15541 ;
  assign n42250 = n34226 ^ n18301 ^ 1'b0 ;
  assign n42251 = ~n42249 & n42250 ;
  assign n42254 = n42253 ^ n42251 ^ 1'b0 ;
  assign n42255 = n35663 ^ n24267 ^ 1'b0 ;
  assign n42257 = n7199 ^ n681 ^ 1'b0 ;
  assign n42258 = n35744 | n42257 ;
  assign n42259 = n2173 & ~n7690 ;
  assign n42260 = ~n2173 & n42259 ;
  assign n42261 = n345 & ~n1766 ;
  assign n42262 = ~n345 & n42261 ;
  assign n42263 = x229 & ~n42262 ;
  assign n42264 = ~x229 & n42263 ;
  assign n42265 = n42264 ^ n10472 ^ 1'b0 ;
  assign n42266 = n42260 | n42265 ;
  assign n42267 = n42260 & ~n42266 ;
  assign n42268 = n1917 | n5512 ;
  assign n42269 = ( n42258 & n42267 ) | ( n42258 & ~n42268 ) | ( n42267 & ~n42268 ) ;
  assign n42256 = n28012 & n31729 ;
  assign n42270 = n42269 ^ n42256 ^ 1'b0 ;
  assign n42271 = n13880 ^ n10174 ^ 1'b0 ;
  assign n42272 = n32445 ^ n10169 ^ 1'b0 ;
  assign n42273 = n27998 | n42272 ;
  assign n42274 = n6373 | n20541 ;
  assign n42275 = n42273 & ~n42274 ;
  assign n42276 = ( n14581 & n23780 ) | ( n14581 & n31069 ) | ( n23780 & n31069 ) ;
  assign n42277 = ( ~n29464 & n33564 ) | ( ~n29464 & n42276 ) | ( n33564 & n42276 ) ;
  assign n42278 = ( n2259 & n38774 ) | ( n2259 & ~n42277 ) | ( n38774 & ~n42277 ) ;
  assign n42279 = n42278 ^ n12600 ^ n5370 ;
  assign n42280 = n29324 & n38884 ;
  assign n42281 = n6888 ^ n3256 ^ 1'b0 ;
  assign n42282 = n4153 & ~n42281 ;
  assign n42283 = ( n12862 & ~n32821 ) | ( n12862 & n42282 ) | ( ~n32821 & n42282 ) ;
  assign n42284 = ~n942 & n42283 ;
  assign n42285 = ~n12981 & n38855 ;
  assign n42286 = n25296 | n39746 ;
  assign n42287 = n39788 | n42286 ;
  assign n42290 = n14933 | n24216 ;
  assign n42288 = n1442 | n3308 ;
  assign n42289 = n3881 & ~n42288 ;
  assign n42291 = n42290 ^ n42289 ^ n32253 ;
  assign n42297 = ~n3227 & n10253 ;
  assign n42292 = n6042 & n36882 ;
  assign n42293 = n8589 & n42292 ;
  assign n42294 = n42293 ^ n12125 ^ 1'b0 ;
  assign n42295 = n42294 ^ n14961 ^ 1'b0 ;
  assign n42296 = n35467 & ~n42295 ;
  assign n42298 = n42297 ^ n42296 ^ 1'b0 ;
  assign n42299 = n21661 & n38344 ;
  assign n42300 = n24144 & n24482 ;
  assign n42301 = ~n42299 & n42300 ;
  assign n42303 = ~n455 & n16513 ;
  assign n42304 = n25290 & n42303 ;
  assign n42302 = n10534 & n16532 ;
  assign n42305 = n42304 ^ n42302 ^ 1'b0 ;
  assign n42306 = n19285 | n21680 ;
  assign n42307 = n42306 ^ n22533 ^ 1'b0 ;
  assign n42308 = n28082 & n42307 ;
  assign n42309 = n42308 ^ n3543 ^ 1'b0 ;
  assign n42310 = n2197 | n42309 ;
  assign n42311 = ~n6512 & n26949 ;
  assign n42312 = ~n21775 & n42311 ;
  assign n42314 = ~n1046 & n20440 ;
  assign n42315 = n42314 ^ n35174 ^ 1'b0 ;
  assign n42313 = n29159 & n36040 ;
  assign n42316 = n42315 ^ n42313 ^ 1'b0 ;
  assign n42317 = n18911 | n18981 ;
  assign n42318 = n42317 ^ n4144 ^ 1'b0 ;
  assign n42319 = n3692 | n42318 ;
  assign n42321 = n10311 ^ n10255 ^ n7556 ;
  assign n42322 = ~n29240 & n42321 ;
  assign n42323 = n25728 | n42322 ;
  assign n42324 = n4409 & ~n42323 ;
  assign n42325 = ( n2118 & n10457 ) | ( n2118 & ~n42324 ) | ( n10457 & ~n42324 ) ;
  assign n42320 = n20523 ^ n527 ^ 1'b0 ;
  assign n42326 = n42325 ^ n42320 ^ n7675 ;
  assign n42327 = n1401 & ~n13577 ;
  assign n42328 = n22527 ^ n3040 ^ 1'b0 ;
  assign n42329 = n20130 | n42328 ;
  assign n42330 = n2345 & ~n42329 ;
  assign n42331 = ~n15951 & n21257 ;
  assign n42332 = n42331 ^ n36728 ^ 1'b0 ;
  assign n42333 = n13048 & ~n42332 ;
  assign n42334 = n42333 ^ n38887 ^ 1'b0 ;
  assign n42335 = n3773 | n5142 ;
  assign n42336 = n42335 ^ n2006 ^ 1'b0 ;
  assign n42337 = n5725 | n25798 ;
  assign n42338 = n37082 ^ n998 ^ 1'b0 ;
  assign n42339 = n42337 & ~n42338 ;
  assign n42340 = ~n8929 & n23834 ;
  assign n42341 = n42340 ^ n32774 ^ 1'b0 ;
  assign n42342 = ~n733 & n35626 ;
  assign n42343 = n39384 & n42342 ;
  assign n42344 = n26502 ^ n2681 ^ n1413 ;
  assign n42345 = n24587 ^ n3995 ^ 1'b0 ;
  assign n42346 = n42345 ^ n40766 ^ n15902 ;
  assign n42347 = ( n3960 & n8319 ) | ( n3960 & ~n10902 ) | ( n8319 & ~n10902 ) ;
  assign n42348 = n10111 ^ n5927 ^ 1'b0 ;
  assign n42349 = n42347 | n42348 ;
  assign n42350 = n40887 ^ n33498 ^ 1'b0 ;
  assign n42351 = ~n7180 & n42350 ;
  assign n42352 = n9472 | n10457 ;
  assign n42353 = n3929 & ~n42352 ;
  assign n42354 = ( n5230 & ~n14736 ) | ( n5230 & n18387 ) | ( ~n14736 & n18387 ) ;
  assign n42355 = ~n36095 & n42354 ;
  assign n42356 = n36189 & n42355 ;
  assign n42357 = ~n11136 & n42356 ;
  assign n42358 = n42357 ^ n7777 ^ 1'b0 ;
  assign n42359 = n17298 ^ n1961 ^ 1'b0 ;
  assign n42361 = n5718 & ~n12728 ;
  assign n42362 = n42361 ^ n562 ^ 1'b0 ;
  assign n42363 = n42362 ^ n11688 ^ n2409 ;
  assign n42360 = n36159 ^ n19575 ^ n10534 ;
  assign n42364 = n42363 ^ n42360 ^ n7303 ;
  assign n42365 = n38936 ^ n36178 ^ 1'b0 ;
  assign n42366 = n12273 ^ n8578 ^ 1'b0 ;
  assign n42367 = n11993 & n42366 ;
  assign n42368 = ~n7081 & n21787 ;
  assign n42369 = ~n42367 & n42368 ;
  assign n42370 = n3430 & n14379 ;
  assign n42371 = ~n8103 & n42370 ;
  assign n42372 = n15196 ^ n10753 ^ 1'b0 ;
  assign n42373 = ~n2681 & n42372 ;
  assign n42374 = n1166 & n2836 ;
  assign n42375 = n9790 & n42374 ;
  assign n42376 = n42375 ^ n14541 ^ 1'b0 ;
  assign n42377 = ~n5809 & n42376 ;
  assign n42378 = n21003 | n42377 ;
  assign n42379 = n27064 ^ n12514 ^ 1'b0 ;
  assign n42380 = n3445 & ~n42379 ;
  assign n42381 = n16091 ^ n13752 ^ 1'b0 ;
  assign n42382 = n21816 | n42381 ;
  assign n42383 = n19408 ^ n10766 ^ 1'b0 ;
  assign n42384 = ( n1767 & ~n31290 ) | ( n1767 & n35782 ) | ( ~n31290 & n35782 ) ;
  assign n42385 = ~n27925 & n42384 ;
  assign n42386 = n1377 & ~n1822 ;
  assign n42387 = n42386 ^ n28090 ^ n3993 ;
  assign n42388 = n25425 ^ n6985 ^ 1'b0 ;
  assign n42389 = n9442 | n9561 ;
  assign n42390 = ( n8980 & n25505 ) | ( n8980 & ~n37090 ) | ( n25505 & ~n37090 ) ;
  assign n42391 = n42390 ^ n32271 ^ 1'b0 ;
  assign n42392 = n20010 | n42391 ;
  assign n42393 = n9105 | n37748 ;
  assign n42394 = n4774 | n27246 ;
  assign n42395 = n39703 ^ n6234 ^ 1'b0 ;
  assign n42396 = n42394 | n42395 ;
  assign n42397 = n42396 ^ n12965 ^ 1'b0 ;
  assign n42398 = n42397 ^ n10713 ^ x58 ;
  assign n42399 = n30557 ^ n22487 ^ 1'b0 ;
  assign n42400 = n18551 ^ n7937 ^ n2020 ;
  assign n42401 = n32289 | n35987 ;
  assign n42402 = n20270 & ~n42401 ;
  assign n42403 = ~n10397 & n36113 ;
  assign n42404 = ~n5230 & n20197 ;
  assign n42405 = ~n42403 & n42404 ;
  assign n42406 = n29002 & ~n29689 ;
  assign n42407 = n15966 ^ n1256 ^ 1'b0 ;
  assign n42408 = ~n42406 & n42407 ;
  assign n42409 = ~n11191 & n41797 ;
  assign n42410 = n24985 & ~n34543 ;
  assign n42411 = ( n4287 & n18544 ) | ( n4287 & n18675 ) | ( n18544 & n18675 ) ;
  assign n42412 = n24551 ^ n7038 ^ 1'b0 ;
  assign n42413 = n4338 & n11171 ;
  assign n42414 = ~n42412 & n42413 ;
  assign n42415 = n5482 & n23151 ;
  assign n42416 = n15137 ^ n4163 ^ 1'b0 ;
  assign n42418 = n34538 ^ n16684 ^ n1113 ;
  assign n42417 = ~n4585 & n10560 ;
  assign n42419 = n42418 ^ n42417 ^ 1'b0 ;
  assign n42420 = n11339 & n28006 ;
  assign n42421 = n42420 ^ n13861 ^ 1'b0 ;
  assign n42422 = ( ~n9222 & n23966 ) | ( ~n9222 & n42421 ) | ( n23966 & n42421 ) ;
  assign n42423 = ~n3992 & n7004 ;
  assign n42424 = n6151 & n42423 ;
  assign n42425 = n38111 ^ n11033 ^ 1'b0 ;
  assign n42426 = n9088 & n42425 ;
  assign n42427 = n42426 ^ n24095 ^ n6435 ;
  assign n42428 = n4775 & n37267 ;
  assign n42429 = n42428 ^ n16452 ^ 1'b0 ;
  assign n42430 = n28449 ^ n23122 ^ 1'b0 ;
  assign n42431 = n5399 & n42430 ;
  assign n42432 = x22 & n30034 ;
  assign n42433 = ~n30034 & n42432 ;
  assign n42434 = n42433 ^ n1836 ^ 1'b0 ;
  assign n42435 = ~n5164 & n25238 ;
  assign n42436 = n19874 & n42435 ;
  assign n42437 = n9361 ^ n833 ^ 1'b0 ;
  assign n42438 = ( n9851 & n24208 ) | ( n9851 & n42437 ) | ( n24208 & n42437 ) ;
  assign n42439 = ( n4560 & n10955 ) | ( n4560 & n18367 ) | ( n10955 & n18367 ) ;
  assign n42440 = n30680 & ~n42439 ;
  assign n42441 = n3106 & ~n31387 ;
  assign n42442 = n42441 ^ n8797 ^ 1'b0 ;
  assign n42443 = n4395 & n18313 ;
  assign n42444 = n29403 ^ n2963 ^ 1'b0 ;
  assign n42445 = ~n26783 & n31699 ;
  assign n42446 = n36972 ^ n14747 ^ n11585 ;
  assign n42447 = ~n6370 & n10257 ;
  assign n42448 = n10850 & n42447 ;
  assign n42449 = n42448 ^ n18115 ^ n10097 ;
  assign n42450 = ~n9512 & n37732 ;
  assign n42451 = ~n42449 & n42450 ;
  assign n42452 = n42451 ^ n21888 ^ n21749 ;
  assign n42453 = n33338 ^ n1527 ^ 1'b0 ;
  assign n42454 = n33583 | n42453 ;
  assign n42455 = n13284 & n23076 ;
  assign n42458 = n7544 | n15511 ;
  assign n42459 = n42458 ^ n4415 ^ 1'b0 ;
  assign n42456 = n11876 ^ n725 ^ 1'b0 ;
  assign n42457 = n42456 ^ n28929 ^ 1'b0 ;
  assign n42460 = n42459 ^ n42457 ^ 1'b0 ;
  assign n42461 = n17716 ^ n13705 ^ 1'b0 ;
  assign n42462 = ~n4903 & n37596 ;
  assign n42463 = ~n42461 & n42462 ;
  assign n42475 = n40430 ^ n1242 ^ 1'b0 ;
  assign n42464 = n570 & ~n3256 ;
  assign n42465 = n3256 & n42464 ;
  assign n42466 = n42465 ^ n33995 ^ 1'b0 ;
  assign n42467 = ( n3089 & ~n10339 ) | ( n3089 & n42466 ) | ( ~n10339 & n42466 ) ;
  assign n42468 = ~n258 & n4892 ;
  assign n42469 = n11141 & n42468 ;
  assign n42470 = n13596 ^ n2924 ^ 1'b0 ;
  assign n42471 = ~n42469 & n42470 ;
  assign n42472 = ~n42467 & n42471 ;
  assign n42473 = n42472 ^ n41408 ^ 1'b0 ;
  assign n42474 = n26384 | n42473 ;
  assign n42476 = n42475 ^ n42474 ^ n31936 ;
  assign n42477 = n28903 | n30258 ;
  assign n42478 = n42477 ^ n20439 ^ 1'b0 ;
  assign n42479 = n42478 ^ n1611 ^ 1'b0 ;
  assign n42480 = n42479 ^ n25023 ^ 1'b0 ;
  assign n42481 = ~n5590 & n10625 ;
  assign n42482 = n11761 | n42481 ;
  assign n42483 = n5915 & n8308 ;
  assign n42484 = n42483 ^ n35368 ^ 1'b0 ;
  assign n42485 = n12881 & n14289 ;
  assign n42486 = n14680 & ~n24465 ;
  assign n42487 = n23264 ^ n5136 ^ 1'b0 ;
  assign n42488 = n3244 | n28562 ;
  assign n42489 = ~n39486 & n41209 ;
  assign n42490 = n42489 ^ n1991 ^ 1'b0 ;
  assign n42491 = n42488 & n42490 ;
  assign n42492 = n11781 & n31472 ;
  assign n42493 = ( ~n3555 & n5748 ) | ( ~n3555 & n42492 ) | ( n5748 & n42492 ) ;
  assign n42494 = n42493 ^ n36679 ^ n24060 ;
  assign n42495 = n12640 ^ n10677 ^ n5055 ;
  assign n42496 = n7986 & n10089 ;
  assign n42497 = n42496 ^ n27989 ^ 1'b0 ;
  assign n42498 = n22785 ^ n16907 ^ 1'b0 ;
  assign n42499 = n42497 & ~n42498 ;
  assign n42500 = n939 & ~n21170 ;
  assign n42501 = n6697 & n42500 ;
  assign n42502 = n32425 | n42501 ;
  assign n42503 = n10191 & ~n42502 ;
  assign n42504 = n4499 | n13384 ;
  assign n42505 = n1403 ^ n1215 ^ 1'b0 ;
  assign n42506 = n22779 ^ n13326 ^ n3632 ;
  assign n42507 = n7732 | n19214 ;
  assign n42508 = n42506 & ~n42507 ;
  assign n42509 = n4383 | n42508 ;
  assign n42510 = n42509 ^ n22354 ^ 1'b0 ;
  assign n42511 = n13817 & n21663 ;
  assign n42512 = ~n7318 & n42511 ;
  assign n42513 = n8659 & ~n42512 ;
  assign n42516 = ( n869 & n21136 ) | ( n869 & ~n33381 ) | ( n21136 & ~n33381 ) ;
  assign n42514 = ( n6068 & ~n7807 ) | ( n6068 & n31370 ) | ( ~n7807 & n31370 ) ;
  assign n42515 = ( n24705 & n34505 ) | ( n24705 & n42514 ) | ( n34505 & n42514 ) ;
  assign n42517 = n42516 ^ n42515 ^ n39860 ;
  assign n42518 = n32709 ^ n5591 ^ 1'b0 ;
  assign n42519 = n17143 ^ n13994 ^ 1'b0 ;
  assign n42520 = ~n550 & n4097 ;
  assign n42521 = n42520 ^ n14004 ^ 1'b0 ;
  assign n42522 = n42521 ^ n34395 ^ n10864 ;
  assign n42523 = ~n20355 & n42522 ;
  assign n42524 = n42523 ^ n7068 ^ 1'b0 ;
  assign n42525 = ~n1590 & n6513 ;
  assign n42528 = n12152 & ~n15465 ;
  assign n42526 = n33353 ^ n7035 ^ 1'b0 ;
  assign n42527 = n24175 & n42526 ;
  assign n42529 = n42528 ^ n42527 ^ 1'b0 ;
  assign n42530 = ( n740 & n35827 ) | ( n740 & n42529 ) | ( n35827 & n42529 ) ;
  assign n42531 = n42530 ^ x118 ^ 1'b0 ;
  assign n42532 = n42525 & n42531 ;
  assign n42533 = n2797 & n5986 ;
  assign n42534 = ~n6969 & n42533 ;
  assign n42535 = ~n16834 & n42534 ;
  assign n42536 = n17521 ^ n8689 ^ 1'b0 ;
  assign n42537 = n42536 ^ n19785 ^ n12118 ;
  assign n42538 = n41915 ^ n30567 ^ n19830 ;
  assign n42539 = n14487 & n22933 ;
  assign n42540 = n42539 ^ n4153 ^ 1'b0 ;
  assign n42541 = n19704 | n42540 ;
  assign n42542 = n42541 ^ n31752 ^ 1'b0 ;
  assign n42545 = n22999 ^ n22360 ^ 1'b0 ;
  assign n42546 = ( n15500 & n34511 ) | ( n15500 & ~n42545 ) | ( n34511 & ~n42545 ) ;
  assign n42543 = n3617 & ~n33964 ;
  assign n42544 = n42543 ^ n11599 ^ 1'b0 ;
  assign n42547 = n42546 ^ n42544 ^ 1'b0 ;
  assign n42548 = n26358 ^ n20272 ^ n11533 ;
  assign n42549 = n3878 & n42548 ;
  assign n42550 = n985 & n42549 ;
  assign n42551 = n18479 & n42550 ;
  assign n42552 = n12617 & n24275 ;
  assign n42553 = ~n39244 & n42552 ;
  assign n42554 = n27510 ^ n7749 ^ 1'b0 ;
  assign n42555 = n29488 | n42554 ;
  assign n42556 = n42553 & ~n42555 ;
  assign n42557 = n42556 ^ n31008 ^ 1'b0 ;
  assign n42558 = n35924 ^ n30468 ^ 1'b0 ;
  assign n42559 = n1081 & n10633 ;
  assign n42560 = n39257 | n42559 ;
  assign n42561 = n18329 ^ n12148 ^ 1'b0 ;
  assign n42562 = n24223 ^ n11591 ^ 1'b0 ;
  assign n42563 = ~n23940 & n42562 ;
  assign n42564 = n624 & ~n26126 ;
  assign n42565 = ( n18432 & n18781 ) | ( n18432 & ~n21044 ) | ( n18781 & ~n21044 ) ;
  assign n42566 = n42565 ^ n25870 ^ 1'b0 ;
  assign n42567 = ~n42564 & n42566 ;
  assign n42568 = n7203 & ~n14160 ;
  assign n42569 = n42568 ^ n22373 ^ 1'b0 ;
  assign n42570 = n42569 ^ n13454 ^ 1'b0 ;
  assign n42571 = ~n8960 & n42570 ;
  assign n42572 = ~n23738 & n42571 ;
  assign n42573 = n1400 & n42572 ;
  assign n42574 = n1281 & ~n6009 ;
  assign n42575 = n42574 ^ n8966 ^ 1'b0 ;
  assign n42576 = ~n5697 & n42575 ;
  assign n42577 = n15655 | n26081 ;
  assign n42578 = n42576 | n42577 ;
  assign n42579 = n21965 ^ n2556 ^ 1'b0 ;
  assign n42580 = n36584 ^ n29034 ^ 1'b0 ;
  assign n42581 = n6602 ^ n486 ^ 1'b0 ;
  assign n42582 = ~n1732 & n9260 ;
  assign n42583 = ~n4608 & n33936 ;
  assign n42584 = n14216 ^ x39 ^ 1'b0 ;
  assign n42585 = n29321 | n42584 ;
  assign n42586 = n37993 & ~n42585 ;
  assign n42587 = n36825 ^ n23406 ^ 1'b0 ;
  assign n42588 = n25463 ^ n11114 ^ 1'b0 ;
  assign n42589 = n14974 ^ n11747 ^ 1'b0 ;
  assign n42590 = n42589 ^ n38899 ^ n12134 ;
  assign n42591 = ~n20570 & n22959 ;
  assign n42592 = n17127 & n18503 ;
  assign n42593 = n2645 & n42592 ;
  assign n42594 = n39492 ^ n2893 ^ 1'b0 ;
  assign n42595 = n42593 | n42594 ;
  assign n42596 = n13271 | n23336 ;
  assign n42597 = n38267 | n42596 ;
  assign n42598 = n36784 ^ x167 ^ 1'b0 ;
  assign n42599 = n21462 | n42598 ;
  assign n42600 = n4531 | n39350 ;
  assign n42601 = n10203 & ~n42600 ;
  assign n42602 = n23007 ^ n1364 ^ 1'b0 ;
  assign n42603 = ( n2548 & ~n25753 ) | ( n2548 & n42602 ) | ( ~n25753 & n42602 ) ;
  assign n42604 = n24191 ^ n12773 ^ 1'b0 ;
  assign n42605 = n33561 | n42604 ;
  assign n42606 = n42605 ^ x200 ^ 1'b0 ;
  assign n42607 = ( n15088 & n21654 ) | ( n15088 & n25245 ) | ( n21654 & n25245 ) ;
  assign n42608 = n8190 & n10685 ;
  assign n42609 = n1246 & n42608 ;
  assign n42610 = n6134 & n26806 ;
  assign n42611 = n42610 ^ n9489 ^ 1'b0 ;
  assign n42612 = n7380 ^ n5067 ^ n1384 ;
  assign n42613 = n30402 ^ n6066 ^ 1'b0 ;
  assign n42614 = n42612 & ~n42613 ;
  assign n42615 = ( n18008 & n32878 ) | ( n18008 & n33971 ) | ( n32878 & n33971 ) ;
  assign n42616 = n42615 ^ n38559 ^ n6080 ;
  assign n42617 = n32455 ^ n12099 ^ x191 ;
  assign n42618 = n42617 ^ n28110 ^ n11258 ;
  assign n42619 = n2437 & ~n12679 ;
  assign n42620 = ~n5399 & n42619 ;
  assign n42621 = n5828 | n11593 ;
  assign n42622 = n10123 & ~n42621 ;
  assign n42623 = ~n34491 & n42622 ;
  assign n42624 = n1719 | n42623 ;
  assign n42625 = n42624 ^ n25637 ^ 1'b0 ;
  assign n42626 = n11219 ^ n6209 ^ 1'b0 ;
  assign n42630 = n2438 | n19295 ;
  assign n42631 = n42630 ^ n8278 ^ 1'b0 ;
  assign n42627 = ~n5736 & n12373 ;
  assign n42628 = n7417 & n42627 ;
  assign n42629 = n7518 & ~n42628 ;
  assign n42632 = n42631 ^ n42629 ^ 1'b0 ;
  assign n42633 = n42632 ^ n15260 ^ 1'b0 ;
  assign n42634 = n7102 ^ n2431 ^ 1'b0 ;
  assign n42635 = n32570 & ~n42634 ;
  assign n42636 = n23685 ^ n1453 ^ 1'b0 ;
  assign n42637 = n7522 ^ n4294 ^ 1'b0 ;
  assign n42638 = ( n6724 & n42636 ) | ( n6724 & ~n42637 ) | ( n42636 & ~n42637 ) ;
  assign n42639 = ( n15032 & n15582 ) | ( n15032 & ~n17326 ) | ( n15582 & ~n17326 ) ;
  assign n42640 = n42639 ^ n16468 ^ 1'b0 ;
  assign n42641 = n648 & ~n22438 ;
  assign n42642 = n42641 ^ n7680 ^ 1'b0 ;
  assign n42643 = n13495 & ~n42642 ;
  assign n42644 = n5167 & n32413 ;
  assign n42645 = ~n2743 & n42644 ;
  assign n42646 = n29105 ^ n20009 ^ 1'b0 ;
  assign n42647 = n6291 & n42646 ;
  assign n42648 = n22665 & ~n32384 ;
  assign n42649 = n42456 & n42648 ;
  assign n42650 = n42649 ^ n29587 ^ 1'b0 ;
  assign n42651 = ( n42645 & ~n42647 ) | ( n42645 & n42650 ) | ( ~n42647 & n42650 ) ;
  assign n42652 = n3335 & ~n23027 ;
  assign n42653 = n7441 & n12049 ;
  assign n42654 = n42653 ^ n25599 ^ 1'b0 ;
  assign n42655 = n23617 ^ n1757 ^ 1'b0 ;
  assign n42656 = n26605 & ~n42655 ;
  assign n42657 = n8391 & ~n13581 ;
  assign n42658 = n38688 & n42657 ;
  assign n42659 = n11319 & ~n39314 ;
  assign n42660 = n9978 ^ n7999 ^ x14 ;
  assign n42661 = n42660 ^ n4688 ^ 1'b0 ;
  assign n42662 = ( n18190 & ~n19670 ) | ( n18190 & n27324 ) | ( ~n19670 & n27324 ) ;
  assign n42663 = n42662 ^ n38361 ^ n13483 ;
  assign n42664 = n23933 ^ n7559 ^ n2970 ;
  assign n42666 = n33534 ^ n713 ^ 1'b0 ;
  assign n42667 = ~n11198 & n22031 ;
  assign n42668 = n42666 & n42667 ;
  assign n42665 = n8259 & n29380 ;
  assign n42669 = n42668 ^ n42665 ^ 1'b0 ;
  assign n42670 = n36399 ^ n15168 ^ 1'b0 ;
  assign n42671 = n3501 ^ n1466 ^ 1'b0 ;
  assign n42673 = n20783 ^ n20752 ^ 1'b0 ;
  assign n42672 = ~n11290 & n13989 ;
  assign n42674 = n42673 ^ n42672 ^ n2460 ;
  assign n42675 = n42674 ^ n25845 ^ 1'b0 ;
  assign n42676 = ~n10252 & n30424 ;
  assign n42677 = ~n5272 & n42676 ;
  assign n42678 = ( n20054 & n27184 ) | ( n20054 & ~n42677 ) | ( n27184 & ~n42677 ) ;
  assign n42682 = n604 | n19968 ;
  assign n42683 = n32382 | n42682 ;
  assign n42679 = ( n20586 & n26671 ) | ( n20586 & n30465 ) | ( n26671 & n30465 ) ;
  assign n42680 = n42679 ^ n18870 ^ 1'b0 ;
  assign n42681 = n3859 & n42680 ;
  assign n42684 = n42683 ^ n42681 ^ n8769 ;
  assign n42685 = n22818 & n39358 ;
  assign n42686 = n21015 | n30494 ;
  assign n42687 = x22 & ~n42686 ;
  assign n42688 = n1297 & ~n23857 ;
  assign n42689 = n4062 & ~n10576 ;
  assign n42690 = ~n36481 & n42689 ;
  assign n42691 = n20279 ^ n8645 ^ 1'b0 ;
  assign n42692 = ~n15970 & n42691 ;
  assign n42693 = n42692 ^ n23479 ^ 1'b0 ;
  assign n42694 = n42693 ^ n16673 ^ 1'b0 ;
  assign n42695 = n7323 & ~n21211 ;
  assign n42696 = ( ~n7260 & n42694 ) | ( ~n7260 & n42695 ) | ( n42694 & n42695 ) ;
  assign n42697 = n17687 ^ n6992 ^ 1'b0 ;
  assign n42698 = n8120 & n34600 ;
  assign n42699 = ( n23336 & n42697 ) | ( n23336 & ~n42698 ) | ( n42697 & ~n42698 ) ;
  assign n42700 = n3841 & ~n5905 ;
  assign n42701 = n16807 & n42700 ;
  assign n42702 = n42701 ^ n39900 ^ n27155 ;
  assign n42703 = n9872 ^ n6216 ^ 1'b0 ;
  assign n42704 = n40782 & ~n42703 ;
  assign n42705 = n22202 ^ n21265 ^ 1'b0 ;
  assign n42706 = n20524 & n42705 ;
  assign n42707 = n42706 ^ n10040 ^ 1'b0 ;
  assign n42709 = n19255 ^ n13440 ^ n8403 ;
  assign n42708 = n18869 & ~n24845 ;
  assign n42710 = n42709 ^ n42708 ^ n3300 ;
  assign n42711 = n8688 & ~n32102 ;
  assign n42712 = n42711 ^ n1850 ^ 1'b0 ;
  assign n42713 = n32263 ^ n30535 ^ n7559 ;
  assign n42714 = n26692 | n28685 ;
  assign n42715 = n8815 & n31291 ;
  assign n42716 = n39781 ^ n21726 ^ 1'b0 ;
  assign n42717 = ~n33156 & n41594 ;
  assign n42718 = ~n33090 & n37822 ;
  assign n42719 = n42718 ^ n12554 ^ n5457 ;
  assign n42720 = n42719 ^ n7311 ^ 1'b0 ;
  assign n42721 = n804 & ~n9422 ;
  assign n42722 = ~n19680 & n42721 ;
  assign n42723 = n42722 ^ n15258 ^ 1'b0 ;
  assign n42724 = n26119 | n42723 ;
  assign n42725 = n9350 & ~n9932 ;
  assign n42726 = n869 & n42725 ;
  assign n42727 = ~n42724 & n42726 ;
  assign n42728 = n24073 ^ n20844 ^ 1'b0 ;
  assign n42729 = ~n7906 & n42728 ;
  assign n42730 = n42729 ^ n22415 ^ 1'b0 ;
  assign n42731 = n29980 ^ n8276 ^ 1'b0 ;
  assign n42732 = n42730 & n42731 ;
  assign n42733 = n15096 ^ n14873 ^ 1'b0 ;
  assign n42734 = ~n12445 & n42733 ;
  assign n42735 = n41127 & n42734 ;
  assign n42736 = n13851 | n31771 ;
  assign n42737 = n3683 ^ n2783 ^ 1'b0 ;
  assign n42739 = n2777 & ~n8143 ;
  assign n42738 = n19375 & n21272 ;
  assign n42740 = n42739 ^ n42738 ^ 1'b0 ;
  assign n42741 = ~n23269 & n42740 ;
  assign n42742 = n2782 & ~n30963 ;
  assign n42743 = ( n3063 & n31421 ) | ( n3063 & n42742 ) | ( n31421 & n42742 ) ;
  assign n42744 = n8829 | n34818 ;
  assign n42745 = ( n20392 & ~n39805 ) | ( n20392 & n42744 ) | ( ~n39805 & n42744 ) ;
  assign n42746 = n23114 ^ n5996 ^ 1'b0 ;
  assign n42747 = n14701 | n42746 ;
  assign n42748 = n17179 | n30600 ;
  assign n42749 = n42748 ^ n13860 ^ 1'b0 ;
  assign n42750 = ( n39746 & n42747 ) | ( n39746 & n42749 ) | ( n42747 & n42749 ) ;
  assign n42751 = n7246 & n7748 ;
  assign n42752 = n12548 | n42751 ;
  assign n42753 = n42752 ^ n16047 ^ 1'b0 ;
  assign n42754 = ( n3659 & n5387 ) | ( n3659 & ~n16834 ) | ( n5387 & ~n16834 ) ;
  assign n42755 = n4840 | n19602 ;
  assign n42756 = n42754 & ~n42755 ;
  assign n42757 = n14181 & n35856 ;
  assign n42758 = ~n5731 & n6054 ;
  assign n42759 = n19934 & n42758 ;
  assign n42760 = ~n405 & n6192 ;
  assign n42761 = n2230 & n42760 ;
  assign n42762 = n822 & ~n42761 ;
  assign n42763 = n14918 | n42762 ;
  assign n42764 = n4602 & n40497 ;
  assign n42765 = n14992 & ~n24608 ;
  assign n42766 = ~n10535 & n18189 ;
  assign n42767 = n42766 ^ n22423 ^ 1'b0 ;
  assign n42768 = n19788 & ~n42767 ;
  assign n42769 = n42768 ^ n19462 ^ 1'b0 ;
  assign n42770 = n24042 ^ n2780 ^ 1'b0 ;
  assign n42771 = ~n13885 & n42770 ;
  assign n42772 = ~n3985 & n8725 ;
  assign n42773 = n42772 ^ n42694 ^ 1'b0 ;
  assign n42774 = n37194 ^ n30167 ^ 1'b0 ;
  assign n42775 = n28716 & ~n42774 ;
  assign n42776 = n13610 & ~n20592 ;
  assign n42777 = n24928 ^ n13442 ^ 1'b0 ;
  assign n42778 = ~n1023 & n42777 ;
  assign n42779 = ~n30617 & n42778 ;
  assign n42780 = n42779 ^ n15567 ^ 1'b0 ;
  assign n42781 = ( ~n14510 & n23672 ) | ( ~n14510 & n42780 ) | ( n23672 & n42780 ) ;
  assign n42782 = n18831 & ~n42781 ;
  assign n42783 = n17184 ^ n6930 ^ 1'b0 ;
  assign n42784 = n13742 ^ n7473 ^ 1'b0 ;
  assign n42785 = n2675 & n17364 ;
  assign n42786 = ~n42784 & n42785 ;
  assign n42787 = ~n4385 & n5637 ;
  assign n42788 = n698 & n42787 ;
  assign n42789 = n12930 ^ n9133 ^ n3905 ;
  assign n42790 = ( n1033 & n3088 ) | ( n1033 & n19195 ) | ( n3088 & n19195 ) ;
  assign n42791 = n8754 | n30158 ;
  assign n42792 = n10023 & ~n42791 ;
  assign n42793 = n42792 ^ n31404 ^ n14329 ;
  assign n42794 = n35493 ^ n19487 ^ 1'b0 ;
  assign n42795 = n17326 ^ n2142 ^ 1'b0 ;
  assign n42796 = n10095 | n13868 ;
  assign n42797 = n34830 & ~n42796 ;
  assign n42798 = n2571 | n20749 ;
  assign n42799 = n5326 & ~n42798 ;
  assign n42800 = n19760 ^ n10579 ^ 1'b0 ;
  assign n42801 = ~n42799 & n42800 ;
  assign n42802 = ~n20509 & n38267 ;
  assign n42803 = ~n42801 & n42802 ;
  assign n42804 = n10555 & ~n30628 ;
  assign n42805 = n42804 ^ n30726 ^ 1'b0 ;
  assign n42806 = n8549 & n17658 ;
  assign n42808 = n36548 ^ n24020 ^ 1'b0 ;
  assign n42809 = n20684 & ~n42808 ;
  assign n42807 = n31175 | n41724 ;
  assign n42810 = n42809 ^ n42807 ^ 1'b0 ;
  assign n42811 = n42810 ^ n13122 ^ n9874 ;
  assign n42812 = ( n4547 & n7974 ) | ( n4547 & ~n15168 ) | ( n7974 & ~n15168 ) ;
  assign n42813 = n2024 & n39982 ;
  assign n42814 = ~n10469 & n42813 ;
  assign n42815 = ( n3089 & n6421 ) | ( n3089 & ~n13996 ) | ( n6421 & ~n13996 ) ;
  assign n42816 = x241 | n1965 ;
  assign n42817 = n42815 & ~n42816 ;
  assign n42818 = n42817 ^ n18140 ^ 1'b0 ;
  assign n42819 = n11046 | n42818 ;
  assign n42820 = n42751 ^ n32989 ^ 1'b0 ;
  assign n42821 = n27438 & ~n42820 ;
  assign n42822 = n8125 ^ n5855 ^ 1'b0 ;
  assign n42823 = ( ~n1800 & n16810 ) | ( ~n1800 & n42115 ) | ( n16810 & n42115 ) ;
  assign n42824 = n21701 ^ n20914 ^ 1'b0 ;
  assign n42825 = x234 & n42824 ;
  assign n42826 = n11585 ^ n8785 ^ 1'b0 ;
  assign n42827 = n18894 ^ n1272 ^ 1'b0 ;
  assign n42828 = n28294 & ~n42827 ;
  assign n42829 = ~n16251 & n42828 ;
  assign n42830 = n42829 ^ n27036 ^ 1'b0 ;
  assign n42831 = n23376 ^ n2460 ^ 1'b0 ;
  assign n42832 = x253 & ~n3894 ;
  assign n42833 = n9865 & n42832 ;
  assign n42834 = n42833 ^ n489 ^ 1'b0 ;
  assign n42835 = ( n4686 & ~n7260 ) | ( n4686 & n42834 ) | ( ~n7260 & n42834 ) ;
  assign n42836 = n22148 ^ n3872 ^ 1'b0 ;
  assign n42837 = ~n42835 & n42836 ;
  assign n42838 = n6242 ^ n681 ^ 1'b0 ;
  assign n42839 = n4918 & ~n42838 ;
  assign n42841 = n3523 & n11316 ;
  assign n42840 = ~n11350 & n16651 ;
  assign n42842 = n42841 ^ n42840 ^ 1'b0 ;
  assign n42843 = n42842 ^ n20511 ^ 1'b0 ;
  assign n42844 = ( n17576 & ~n19129 ) | ( n17576 & n20693 ) | ( ~n19129 & n20693 ) ;
  assign n42845 = n14077 ^ n3422 ^ 1'b0 ;
  assign n42846 = n42845 ^ n38014 ^ n32498 ;
  assign n42847 = n2670 & n13441 ;
  assign n42848 = n42847 ^ n22261 ^ 1'b0 ;
  assign n42849 = n16804 & ~n28123 ;
  assign n42850 = ~n1247 & n42849 ;
  assign n42851 = n29270 & ~n37143 ;
  assign n42852 = n19399 ^ n12290 ^ 1'b0 ;
  assign n42853 = ~n13159 & n31648 ;
  assign n42854 = n30871 ^ n10801 ^ 1'b0 ;
  assign n42855 = n4293 & n42854 ;
  assign n42856 = n13063 | n27524 ;
  assign n42857 = n4762 & ~n42856 ;
  assign n42858 = n42857 ^ n12551 ^ 1'b0 ;
  assign n42859 = n12753 & n29856 ;
  assign n42860 = n20523 | n31230 ;
  assign n42861 = n42860 ^ n21649 ^ 1'b0 ;
  assign n42862 = n3953 & ~n14549 ;
  assign n42863 = n42862 ^ n2100 ^ 1'b0 ;
  assign n42864 = ~n39188 & n42863 ;
  assign n42865 = n32177 ^ n18691 ^ 1'b0 ;
  assign n42866 = n17374 & ~n31397 ;
  assign n42867 = ( ~n7843 & n8058 ) | ( ~n7843 & n42866 ) | ( n8058 & n42866 ) ;
  assign n42868 = n30434 ^ n6131 ^ 1'b0 ;
  assign n42869 = n31528 & ~n42868 ;
  assign n42870 = n15147 ^ n2440 ^ 1'b0 ;
  assign n42871 = n9373 & n42870 ;
  assign n42872 = n42871 ^ n40767 ^ 1'b0 ;
  assign n42873 = x58 & ~n42872 ;
  assign n42874 = n22186 ^ n10211 ^ 1'b0 ;
  assign n42875 = n18549 | n42874 ;
  assign n42876 = n15566 ^ n4370 ^ 1'b0 ;
  assign n42877 = ~n42875 & n42876 ;
  assign n42878 = ~n27451 & n35506 ;
  assign n42879 = ~n5157 & n8908 ;
  assign n42880 = n11317 & n18032 ;
  assign n42881 = n42880 ^ n15776 ^ 1'b0 ;
  assign n42882 = n24803 ^ n10920 ^ 1'b0 ;
  assign n42883 = n32549 & ~n42882 ;
  assign n42884 = ( n39382 & n42881 ) | ( n39382 & ~n42883 ) | ( n42881 & ~n42883 ) ;
  assign n42885 = n513 & ~n3957 ;
  assign n42886 = ~n11593 & n42885 ;
  assign n42887 = ( n3464 & n37972 ) | ( n3464 & n42886 ) | ( n37972 & n42886 ) ;
  assign n42888 = n2561 & ~n29983 ;
  assign n42889 = n14076 ^ n3228 ^ n917 ;
  assign n42890 = n42889 ^ n16207 ^ 1'b0 ;
  assign n42891 = ~n9965 & n16775 ;
  assign n42892 = n16516 | n27368 ;
  assign n42893 = n11420 | n42892 ;
  assign n42894 = n12357 ^ n11360 ^ 1'b0 ;
  assign n42895 = n39218 & n42894 ;
  assign n42897 = n4029 ^ n2592 ^ 1'b0 ;
  assign n42896 = ~n14665 & n24169 ;
  assign n42898 = n42897 ^ n42896 ^ 1'b0 ;
  assign n42899 = ~n3430 & n42898 ;
  assign n42900 = n10985 & ~n12199 ;
  assign n42901 = n8772 & n42900 ;
  assign n42902 = n42901 ^ n20594 ^ 1'b0 ;
  assign n42903 = n38220 ^ n4353 ^ n1779 ;
  assign n42904 = n11175 ^ n9476 ^ n4034 ;
  assign n42905 = n42904 ^ n22689 ^ 1'b0 ;
  assign n42906 = n14379 ^ n3711 ^ 1'b0 ;
  assign n42907 = n5788 ^ n4359 ^ 1'b0 ;
  assign n42908 = n42906 | n42907 ;
  assign n42909 = ( n3423 & n5308 ) | ( n3423 & ~n7897 ) | ( n5308 & ~n7897 ) ;
  assign n42910 = n27539 ^ n5915 ^ 1'b0 ;
  assign n42911 = ~n42909 & n42910 ;
  assign n42912 = n40564 ^ n20481 ^ 1'b0 ;
  assign n42913 = n42911 & n42912 ;
  assign n42914 = n22163 | n35134 ;
  assign n42915 = n42914 ^ n40576 ^ 1'b0 ;
  assign n42916 = n5864 | n21683 ;
  assign n42917 = n7017 & ~n40576 ;
  assign n42918 = n20260 & n42917 ;
  assign n42919 = ~n42916 & n42918 ;
  assign n42920 = n24847 ^ n14485 ^ 1'b0 ;
  assign n42921 = n16490 | n42920 ;
  assign n42922 = n5013 | n42921 ;
  assign n42923 = n17979 & ~n24835 ;
  assign n42924 = n26633 | n42923 ;
  assign n42925 = n42924 ^ n20666 ^ 1'b0 ;
  assign n42926 = n42925 ^ n11111 ^ n10019 ;
  assign n42927 = ~n4422 & n24776 ;
  assign n42928 = n32137 | n35022 ;
  assign n42929 = n38196 & ~n42928 ;
  assign n42930 = n10032 | n23470 ;
  assign n42931 = ~n26699 & n42930 ;
  assign n42932 = n42931 ^ n2296 ^ 1'b0 ;
  assign n42933 = ~n11674 & n13891 ;
  assign n42934 = ~n9942 & n42933 ;
  assign n42935 = n4247 & ~n20912 ;
  assign n42936 = n42935 ^ n14657 ^ 1'b0 ;
  assign n42937 = n7386 ^ n5449 ^ 1'b0 ;
  assign n42938 = n690 & ~n5782 ;
  assign n42939 = n840 & n42938 ;
  assign n42940 = n42939 ^ n17631 ^ n8778 ;
  assign n42941 = n11060 & ~n33627 ;
  assign n42942 = n15653 & n26447 ;
  assign n42943 = n5605 & n42942 ;
  assign n42944 = n17717 ^ n15516 ^ n7540 ;
  assign n42945 = ~n20223 & n42944 ;
  assign n42949 = n2066 & n3134 ;
  assign n42950 = ~n24403 & n42949 ;
  assign n42946 = n3737 ^ n878 ^ 1'b0 ;
  assign n42947 = n1651 & ~n42946 ;
  assign n42948 = ~n13523 & n42947 ;
  assign n42951 = n42950 ^ n42948 ^ 1'b0 ;
  assign n42952 = n42951 ^ n14218 ^ 1'b0 ;
  assign n42953 = n1991 & n41655 ;
  assign n42954 = n7656 | n9993 ;
  assign n42955 = n42954 ^ n9490 ^ 1'b0 ;
  assign n42956 = ~n6023 & n42955 ;
  assign n42957 = n42956 ^ n17320 ^ 1'b0 ;
  assign n42958 = n42035 ^ n30807 ^ n29854 ;
  assign n42959 = n25079 ^ n14027 ^ 1'b0 ;
  assign n42960 = n13920 ^ n3479 ^ 1'b0 ;
  assign n42961 = n427 & ~n26124 ;
  assign n42962 = ~n2098 & n42961 ;
  assign n42963 = n42962 ^ n8532 ^ n3129 ;
  assign n42964 = x149 & n27162 ;
  assign n42965 = n8709 & n24909 ;
  assign n42968 = n9838 ^ n8924 ^ n4684 ;
  assign n42966 = n21632 ^ n432 ^ 1'b0 ;
  assign n42967 = ~n20866 & n42966 ;
  assign n42969 = n42968 ^ n42967 ^ n24699 ;
  assign n42970 = n3770 & ~n29914 ;
  assign n42971 = n3528 | n8054 ;
  assign n42972 = n4719 | n42971 ;
  assign n42973 = n42972 ^ n23470 ^ n4446 ;
  assign n42974 = n2315 & n9170 ;
  assign n42975 = n681 & n42974 ;
  assign n42976 = n18639 & n38536 ;
  assign n42977 = n42976 ^ n13742 ^ 1'b0 ;
  assign n42978 = n8619 | n42977 ;
  assign n42979 = n26498 ^ n10460 ^ 1'b0 ;
  assign n42980 = n42979 ^ n23157 ^ 1'b0 ;
  assign n42981 = n42980 ^ n35352 ^ 1'b0 ;
  assign n42982 = ~n9075 & n42981 ;
  assign n42984 = n33926 | n35847 ;
  assign n42983 = n7810 & n33935 ;
  assign n42985 = n42984 ^ n42983 ^ 1'b0 ;
  assign n42986 = n23215 & ~n28233 ;
  assign n42987 = ~n29402 & n42986 ;
  assign n42988 = n14813 & n42917 ;
  assign n42989 = n42987 & n42988 ;
  assign n42990 = n1533 | n28484 ;
  assign n42991 = n15284 ^ n11935 ^ 1'b0 ;
  assign n42992 = n4309 & ~n42991 ;
  assign n42993 = ~n14693 & n42992 ;
  assign n42994 = n42993 ^ n39164 ^ n1957 ;
  assign n42995 = n28658 & n32320 ;
  assign n42996 = ~n6216 & n42995 ;
  assign n42997 = n12157 | n35048 ;
  assign n42998 = n10078 & ~n26377 ;
  assign n42999 = n38135 ^ n9843 ^ 1'b0 ;
  assign n43000 = ( n3733 & n5962 ) | ( n3733 & n18915 ) | ( n5962 & n18915 ) ;
  assign n43001 = ~n20523 & n23698 ;
  assign n43002 = ( n11165 & ~n11282 ) | ( n11165 & n43001 ) | ( ~n11282 & n43001 ) ;
  assign n43003 = n4549 & ~n36662 ;
  assign n43004 = n43003 ^ n39268 ^ 1'b0 ;
  assign n43005 = n12366 | n22078 ;
  assign n43006 = n43005 ^ n3313 ^ 1'b0 ;
  assign n43007 = n19056 | n43006 ;
  assign n43008 = n15795 ^ n5004 ^ 1'b0 ;
  assign n43009 = n17022 ^ n15639 ^ 1'b0 ;
  assign n43010 = n836 & n43009 ;
  assign n43011 = n43010 ^ n28018 ^ 1'b0 ;
  assign n43013 = n12776 ^ n12074 ^ 1'b0 ;
  assign n43014 = n6767 & ~n43013 ;
  assign n43012 = n1904 & ~n4846 ;
  assign n43015 = n43014 ^ n43012 ^ 1'b0 ;
  assign n43016 = n14659 & ~n19935 ;
  assign n43017 = n43016 ^ n10862 ^ 1'b0 ;
  assign n43018 = n15970 & ~n37889 ;
  assign n43019 = n43018 ^ n19564 ^ 1'b0 ;
  assign n43020 = n5667 | n13899 ;
  assign n43021 = n43020 ^ n8630 ^ 1'b0 ;
  assign n43022 = n1951 | n3515 ;
  assign n43023 = n43021 & ~n43022 ;
  assign n43024 = n9920 & ~n23396 ;
  assign n43025 = n13122 & n40095 ;
  assign n43026 = n43025 ^ n4996 ^ 1'b0 ;
  assign n43027 = n1332 | n5880 ;
  assign n43028 = n18942 | n43027 ;
  assign n43029 = n27998 ^ n5991 ^ 1'b0 ;
  assign n43030 = ( n17964 & n25621 ) | ( n17964 & n31469 ) | ( n25621 & n31469 ) ;
  assign n43031 = ( n1585 & n25221 ) | ( n1585 & ~n43030 ) | ( n25221 & ~n43030 ) ;
  assign n43033 = n2230 ^ x224 ^ 1'b0 ;
  assign n43032 = n13239 & ~n28630 ;
  assign n43034 = n43033 ^ n43032 ^ 1'b0 ;
  assign n43035 = n2675 & n6228 ;
  assign n43036 = n16922 & n43035 ;
  assign n43037 = n43036 ^ n26941 ^ 1'b0 ;
  assign n43038 = n13535 ^ n12323 ^ 1'b0 ;
  assign n43039 = n307 & ~n4505 ;
  assign n43040 = n30757 & n43039 ;
  assign n43041 = ( n12760 & n24565 ) | ( n12760 & n25807 ) | ( n24565 & n25807 ) ;
  assign n43042 = n42574 ^ n30656 ^ 1'b0 ;
  assign n43043 = ( n693 & n25601 ) | ( n693 & ~n31528 ) | ( n25601 & ~n31528 ) ;
  assign n43044 = n9121 & n28402 ;
  assign n43045 = n43044 ^ n5314 ^ 1'b0 ;
  assign n43046 = n43045 ^ n1777 ^ 1'b0 ;
  assign n43047 = n43043 | n43046 ;
  assign n43048 = ~n13201 & n43047 ;
  assign n43049 = n12035 | n35794 ;
  assign n43050 = n9299 | n43049 ;
  assign n43051 = n43050 ^ n38704 ^ n19552 ;
  assign n43052 = n43051 ^ n6286 ^ 1'b0 ;
  assign n43053 = n19734 ^ n8313 ^ 1'b0 ;
  assign n43054 = n43052 & n43053 ;
  assign n43055 = n4308 & n14711 ;
  assign n43056 = n4560 & n43055 ;
  assign n43057 = n43056 ^ n38519 ^ 1'b0 ;
  assign n43058 = n12763 ^ n3036 ^ 1'b0 ;
  assign n43059 = n10975 | n13757 ;
  assign n43060 = n43058 & ~n43059 ;
  assign n43061 = n43060 ^ n16205 ^ n8381 ;
  assign n43062 = n11784 ^ n6353 ^ n2281 ;
  assign n43063 = n21140 & n43062 ;
  assign n43064 = n11696 & n43063 ;
  assign n43065 = n5151 ^ n1404 ^ 1'b0 ;
  assign n43066 = n20633 | n43065 ;
  assign n43067 = n43064 & ~n43066 ;
  assign n43068 = ( n6458 & n28658 ) | ( n6458 & n43067 ) | ( n28658 & n43067 ) ;
  assign n43069 = n11011 & ~n26643 ;
  assign n43070 = n43069 ^ n17011 ^ 1'b0 ;
  assign n43071 = ~n456 & n8283 ;
  assign n43072 = ~n2230 & n43071 ;
  assign n43073 = n4375 & ~n41588 ;
  assign n43074 = n24770 ^ n12668 ^ 1'b0 ;
  assign n43075 = n7294 & ~n43074 ;
  assign n43076 = ~n11573 & n13846 ;
  assign n43077 = n43076 ^ n33617 ^ 1'b0 ;
  assign n43078 = n6064 | n28576 ;
  assign n43079 = n9553 & ~n43078 ;
  assign n43080 = n18050 ^ n13881 ^ x82 ;
  assign n43081 = n43080 ^ n24860 ^ n15374 ;
  assign n43082 = n14330 | n42854 ;
  assign n43083 = n11482 & n43082 ;
  assign n43084 = ~n6856 & n43083 ;
  assign n43085 = n3099 | n5931 ;
  assign n43086 = ~n6988 & n43085 ;
  assign n43087 = n43086 ^ n22574 ^ 1'b0 ;
  assign n43088 = n16567 ^ n7083 ^ 1'b0 ;
  assign n43089 = n16233 & n43088 ;
  assign n43090 = ~n3282 & n43089 ;
  assign n43091 = n2380 ^ n1342 ^ 1'b0 ;
  assign n43092 = n10617 & n43091 ;
  assign n43093 = n43092 ^ n7661 ^ 1'b0 ;
  assign n43094 = n24913 ^ n22346 ^ 1'b0 ;
  assign n43095 = n27586 ^ n3904 ^ 1'b0 ;
  assign n43096 = n35481 ^ n25567 ^ n4306 ;
  assign n43097 = ( n2486 & n21711 ) | ( n2486 & ~n43096 ) | ( n21711 & ~n43096 ) ;
  assign n43098 = n31969 ^ n25747 ^ n8996 ;
  assign n43099 = n1760 & n17468 ;
  assign n43100 = n21793 & ~n35819 ;
  assign n43101 = ~n12894 & n20079 ;
  assign n43102 = ~n27879 & n37841 ;
  assign n43103 = n41641 ^ n7969 ^ 1'b0 ;
  assign n43104 = n30664 & ~n43103 ;
  assign n43105 = n3610 & n28132 ;
  assign n43106 = ~n31238 & n43105 ;
  assign n43107 = n34702 ^ n8340 ^ 1'b0 ;
  assign n43108 = ~n22549 & n31555 ;
  assign n43109 = n43108 ^ n8058 ^ 1'b0 ;
  assign n43110 = ( ~n258 & n4207 ) | ( ~n258 & n4317 ) | ( n4207 & n4317 ) ;
  assign n43111 = n18462 & ~n37886 ;
  assign n43112 = n8932 | n18713 ;
  assign n43113 = n43112 ^ n8662 ^ 1'b0 ;
  assign n43114 = n43113 ^ n9757 ^ n4361 ;
  assign n43115 = ( n6381 & n19758 ) | ( n6381 & ~n43114 ) | ( n19758 & ~n43114 ) ;
  assign n43116 = n33581 ^ n25682 ^ 1'b0 ;
  assign n43117 = n1940 & n18555 ;
  assign n43118 = n6458 & ~n11633 ;
  assign n43119 = n17432 ^ n9423 ^ 1'b0 ;
  assign n43120 = n39961 & n43119 ;
  assign n43121 = ~n7839 & n18610 ;
  assign n43122 = n24354 & ~n31475 ;
  assign n43123 = n43122 ^ n5350 ^ 1'b0 ;
  assign n43124 = ( n29559 & ~n33642 ) | ( n29559 & n43123 ) | ( ~n33642 & n43123 ) ;
  assign n43125 = n18408 ^ n16657 ^ 1'b0 ;
  assign n43126 = n34128 & n43125 ;
  assign n43127 = n43126 ^ n22410 ^ n7556 ;
  assign n43128 = n19481 ^ n991 ^ 1'b0 ;
  assign n43129 = n22638 & ~n43128 ;
  assign n43130 = ( ~n13460 & n16018 ) | ( ~n13460 & n43129 ) | ( n16018 & n43129 ) ;
  assign n43131 = ( ~n22529 & n24258 ) | ( ~n22529 & n43130 ) | ( n24258 & n43130 ) ;
  assign n43133 = ( n4954 & ~n9271 ) | ( n4954 & n9942 ) | ( ~n9271 & n9942 ) ;
  assign n43132 = n31440 & n34969 ;
  assign n43134 = n43133 ^ n43132 ^ 1'b0 ;
  assign n43135 = n12057 ^ n9483 ^ 1'b0 ;
  assign n43136 = n527 | n7512 ;
  assign n43137 = n43136 ^ n25599 ^ 1'b0 ;
  assign n43138 = n25381 | n43137 ;
  assign n43139 = n4487 ^ n1275 ^ 1'b0 ;
  assign n43140 = n5534 | n43139 ;
  assign n43141 = n10027 ^ n2680 ^ 1'b0 ;
  assign n43142 = n16171 & n43141 ;
  assign n43143 = ~n12651 & n27642 ;
  assign n43144 = n43142 | n43143 ;
  assign n43145 = n2777 ^ n1486 ^ 1'b0 ;
  assign n43146 = n39910 ^ n20803 ^ 1'b0 ;
  assign n43147 = n43145 & n43146 ;
  assign n43148 = n18101 | n22826 ;
  assign n43149 = n28319 ^ n15130 ^ 1'b0 ;
  assign n43150 = ( n17700 & n18296 ) | ( n17700 & ~n37117 ) | ( n18296 & ~n37117 ) ;
  assign n43151 = n11115 & ~n43150 ;
  assign n43152 = ~n43149 & n43151 ;
  assign n43154 = n3542 ^ n3435 ^ 1'b0 ;
  assign n43153 = n12278 | n18653 ;
  assign n43155 = n43154 ^ n43153 ^ 1'b0 ;
  assign n43156 = n1703 ^ x231 ^ 1'b0 ;
  assign n43157 = n37477 ^ n15663 ^ 1'b0 ;
  assign n43158 = ( n541 & ~n43156 ) | ( n541 & n43157 ) | ( ~n43156 & n43157 ) ;
  assign n43159 = n14437 ^ n4080 ^ 1'b0 ;
  assign n43161 = n15412 ^ n14133 ^ 1'b0 ;
  assign n43162 = ~n15621 & n43161 ;
  assign n43160 = n5678 & n33226 ;
  assign n43163 = n43162 ^ n43160 ^ 1'b0 ;
  assign n43164 = n9767 & ~n31588 ;
  assign n43165 = n5144 ^ n1520 ^ 1'b0 ;
  assign n43166 = n43164 & n43165 ;
  assign n43167 = n3119 ^ n3084 ^ 1'b0 ;
  assign n43168 = n25096 & ~n43167 ;
  assign n43169 = n20227 ^ n3947 ^ n3746 ;
  assign n43170 = n43169 ^ n5387 ^ 1'b0 ;
  assign n43171 = n7600 & ~n11384 ;
  assign n43172 = n16841 & n43171 ;
  assign n43173 = n5286 | n43172 ;
  assign n43174 = n43173 ^ n38491 ^ 1'b0 ;
  assign n43175 = n43174 ^ n12635 ^ 1'b0 ;
  assign n43176 = n19249 ^ n4654 ^ 1'b0 ;
  assign n43177 = n38892 ^ n24972 ^ 1'b0 ;
  assign n43178 = n5512 | n11905 ;
  assign n43179 = ~n7611 & n43178 ;
  assign n43180 = n15747 & n30549 ;
  assign n43181 = n15240 ^ n5144 ^ 1'b0 ;
  assign n43182 = n2454 | n27589 ;
  assign n43183 = ( n11434 & n43181 ) | ( n11434 & ~n43182 ) | ( n43181 & ~n43182 ) ;
  assign n43184 = ( n32715 & n34113 ) | ( n32715 & n43183 ) | ( n34113 & n43183 ) ;
  assign n43185 = n14787 & n43184 ;
  assign n43186 = n2574 & n5763 ;
  assign n43187 = n7538 & n43186 ;
  assign n43188 = n31846 | n35299 ;
  assign n43189 = n43187 & ~n43188 ;
  assign n43190 = ~n867 & n6198 ;
  assign n43191 = n43190 ^ n8801 ^ 1'b0 ;
  assign n43192 = n3193 & ~n23592 ;
  assign n43193 = n43192 ^ n27795 ^ 1'b0 ;
  assign n43194 = ~n28109 & n43193 ;
  assign n43195 = n2897 & n27283 ;
  assign n43196 = n1645 & n43195 ;
  assign n43197 = n8039 | n31338 ;
  assign n43198 = n2178 & ~n43197 ;
  assign n43199 = n16424 & ~n43198 ;
  assign n43200 = n6912 & n43199 ;
  assign n43201 = n13863 ^ n856 ^ 1'b0 ;
  assign n43202 = n11004 & n37676 ;
  assign n43203 = n43202 ^ n10991 ^ 1'b0 ;
  assign n43204 = n43203 ^ n10316 ^ 1'b0 ;
  assign n43205 = ~n10751 & n43204 ;
  assign n43206 = ( n5495 & n9128 ) | ( n5495 & n43205 ) | ( n9128 & n43205 ) ;
  assign n43207 = n13157 | n21841 ;
  assign n43208 = n11117 & n43207 ;
  assign n43209 = n30043 ^ n20879 ^ 1'b0 ;
  assign n43210 = n15992 ^ n6409 ^ 1'b0 ;
  assign n43211 = n40637 ^ n3697 ^ 1'b0 ;
  assign n43212 = n38349 ^ n13555 ^ 1'b0 ;
  assign n43213 = n6501 & ~n39260 ;
  assign n43214 = ( n5864 & ~n10131 ) | ( n5864 & n15295 ) | ( ~n10131 & n15295 ) ;
  assign n43215 = n5422 & ~n13650 ;
  assign n43216 = ~n17200 & n43215 ;
  assign n43217 = ( n19982 & n43214 ) | ( n19982 & ~n43216 ) | ( n43214 & ~n43216 ) ;
  assign n43218 = n43217 ^ n30026 ^ n2682 ;
  assign n43219 = ~n6506 & n13297 ;
  assign n43220 = n35871 ^ n26137 ^ 1'b0 ;
  assign n43221 = n31426 ^ n26528 ^ n14095 ;
  assign n43222 = n4758 & ~n32029 ;
  assign n43223 = ~n19943 & n43222 ;
  assign n43224 = n15434 ^ n11317 ^ 1'b0 ;
  assign n43225 = n27470 & ~n28130 ;
  assign n43226 = n22122 & n43225 ;
  assign n43227 = n36398 ^ n1203 ^ 1'b0 ;
  assign n43228 = x116 & ~n43227 ;
  assign n43229 = n43228 ^ n17949 ^ 1'b0 ;
  assign n43230 = n42456 ^ n34849 ^ 1'b0 ;
  assign n43231 = ~n7844 & n8830 ;
  assign n43232 = n43231 ^ n13223 ^ 1'b0 ;
  assign n43233 = n516 & n43232 ;
  assign n43234 = n24780 ^ n1348 ^ 1'b0 ;
  assign n43235 = n17800 | n43234 ;
  assign n43236 = n43233 & ~n43235 ;
  assign n43237 = n2553 & ~n8113 ;
  assign n43238 = ~n4347 & n43237 ;
  assign n43239 = n43238 ^ n12389 ^ 1'b0 ;
  assign n43240 = n11222 ^ n5230 ^ 1'b0 ;
  assign n43241 = n19946 | n43240 ;
  assign n43242 = n808 & n43241 ;
  assign n43243 = ~n35068 & n43242 ;
  assign n43244 = n30609 & ~n43243 ;
  assign n43245 = n32397 & n43244 ;
  assign n43246 = ~n6588 & n37082 ;
  assign n43247 = n43246 ^ n24276 ^ 1'b0 ;
  assign n43248 = n17725 ^ n6297 ^ 1'b0 ;
  assign n43249 = ~n19543 & n28155 ;
  assign n43250 = ~n4606 & n4664 ;
  assign n43251 = n33953 & n43250 ;
  assign n43252 = n1997 | n18432 ;
  assign n43253 = n42188 ^ n447 ^ 1'b0 ;
  assign n43254 = n35822 & ~n43253 ;
  assign n43255 = ~n706 & n43254 ;
  assign n43256 = n30826 ^ x58 ^ 1'b0 ;
  assign n43257 = n40655 ^ n22364 ^ 1'b0 ;
  assign n43258 = x7 & n43257 ;
  assign n43259 = n4306 | n13628 ;
  assign n43260 = n43259 ^ n28845 ^ 1'b0 ;
  assign n43261 = n12317 & ~n30633 ;
  assign n43262 = ~n42623 & n43261 ;
  assign n43263 = ~n6421 & n25455 ;
  assign n43264 = n1235 & ~n3150 ;
  assign n43265 = n3150 & n43264 ;
  assign n43266 = n4544 & ~n43265 ;
  assign n43267 = n43265 & n43266 ;
  assign n43268 = n4538 | n43267 ;
  assign n43269 = n43268 ^ n30217 ^ 1'b0 ;
  assign n43270 = n5775 | n11458 ;
  assign n43271 = ( n1307 & n43269 ) | ( n1307 & ~n43270 ) | ( n43269 & ~n43270 ) ;
  assign n43273 = n13868 ^ n13366 ^ 1'b0 ;
  assign n43274 = ~n1521 & n43273 ;
  assign n43275 = n26519 & ~n43274 ;
  assign n43272 = ( n1667 & n8837 ) | ( n1667 & n28501 ) | ( n8837 & n28501 ) ;
  assign n43276 = n43275 ^ n43272 ^ 1'b0 ;
  assign n43277 = n43276 ^ n32674 ^ 1'b0 ;
  assign n43280 = n20304 | n20873 ;
  assign n43281 = n43280 ^ n14253 ^ 1'b0 ;
  assign n43279 = n5910 & ~n17982 ;
  assign n43282 = n43281 ^ n43279 ^ 1'b0 ;
  assign n43278 = x111 & n13861 ;
  assign n43283 = n43282 ^ n43278 ^ 1'b0 ;
  assign n43284 = n4398 & ~n15229 ;
  assign n43285 = n43284 ^ n6001 ^ 1'b0 ;
  assign n43286 = n24168 ^ n3404 ^ 1'b0 ;
  assign n43287 = ~n19301 & n43286 ;
  assign n43288 = n35345 ^ n9362 ^ n1259 ;
  assign n43289 = n13518 | n32735 ;
  assign n43290 = n4957 | n28872 ;
  assign n43291 = n21556 ^ n395 ^ 1'b0 ;
  assign n43292 = ~n1735 & n43291 ;
  assign n43293 = n14116 & n43292 ;
  assign n43294 = ~n16124 & n17231 ;
  assign n43295 = n17526 ^ n12515 ^ n2774 ;
  assign n43296 = ~n3360 & n26941 ;
  assign n43297 = n18823 ^ n9075 ^ 1'b0 ;
  assign n43298 = n19808 ^ n4425 ^ 1'b0 ;
  assign n43299 = n5380 & n19060 ;
  assign n43300 = ~n38313 & n43299 ;
  assign n43301 = ~x232 & n1298 ;
  assign n43302 = n43301 ^ n13046 ^ 1'b0 ;
  assign n43303 = n17395 ^ n7381 ^ 1'b0 ;
  assign n43304 = n43303 ^ n34797 ^ n24114 ;
  assign n43305 = ~n18338 & n34018 ;
  assign n43306 = n43305 ^ n21095 ^ 1'b0 ;
  assign n43307 = n29105 | n39179 ;
  assign n43308 = n43306 & ~n43307 ;
  assign n43309 = n9032 ^ n1037 ^ 1'b0 ;
  assign n43310 = n8447 ^ n2067 ^ 1'b0 ;
  assign n43311 = ~n8217 & n38310 ;
  assign n43312 = ~n43310 & n43311 ;
  assign n43313 = n10011 ^ n8545 ^ 1'b0 ;
  assign n43314 = ( ~n274 & n41614 ) | ( ~n274 & n43313 ) | ( n41614 & n43313 ) ;
  assign n43315 = ( n4995 & n7764 ) | ( n4995 & ~n36926 ) | ( n7764 & ~n36926 ) ;
  assign n43316 = n17578 ^ n12007 ^ 1'b0 ;
  assign n43317 = ~n33413 & n43316 ;
  assign n43318 = n4872 | n39115 ;
  assign n43319 = n1708 & n14220 ;
  assign n43320 = n674 & ~n3770 ;
  assign n43321 = n43319 & n43320 ;
  assign n43322 = ~n1486 & n6682 ;
  assign n43323 = n43322 ^ n14175 ^ 1'b0 ;
  assign n43324 = ~n29247 & n43323 ;
  assign n43325 = n43324 ^ n13262 ^ 1'b0 ;
  assign n43326 = ~n1208 & n5378 ;
  assign n43327 = n43326 ^ n12018 ^ 1'b0 ;
  assign n43328 = ( n10707 & ~n29909 ) | ( n10707 & n43327 ) | ( ~n29909 & n43327 ) ;
  assign n43329 = ~n2547 & n3056 ;
  assign n43330 = ~n16761 & n43329 ;
  assign n43332 = n9436 & n34702 ;
  assign n43333 = ~n9436 & n43332 ;
  assign n43334 = n11164 & ~n43333 ;
  assign n43335 = ~n21317 & n24514 ;
  assign n43336 = n11278 & n43335 ;
  assign n43337 = ( n29988 & n43334 ) | ( n29988 & n43336 ) | ( n43334 & n43336 ) ;
  assign n43331 = n25467 ^ n21230 ^ n19909 ;
  assign n43338 = n43337 ^ n43331 ^ 1'b0 ;
  assign n43339 = ( n9583 & n43330 ) | ( n9583 & ~n43338 ) | ( n43330 & ~n43338 ) ;
  assign n43340 = n21912 ^ n12590 ^ n9539 ;
  assign n43341 = n6448 & ~n10193 ;
  assign n43342 = n43341 ^ n4754 ^ 1'b0 ;
  assign n43343 = n31585 ^ n24623 ^ 1'b0 ;
  assign n43344 = n43342 & ~n43343 ;
  assign n43345 = n43344 ^ n38859 ^ 1'b0 ;
  assign n43346 = n41451 & n43345 ;
  assign n43347 = n13637 ^ n6979 ^ n351 ;
  assign n43348 = n10200 | n43347 ;
  assign n43354 = n29246 ^ n3422 ^ 1'b0 ;
  assign n43355 = ~n21523 & n24839 ;
  assign n43356 = n43354 & n43355 ;
  assign n43349 = ~n19163 & n21785 ;
  assign n43350 = n30559 & n43349 ;
  assign n43351 = n6366 ^ n559 ^ 1'b0 ;
  assign n43352 = ~n43350 & n43351 ;
  assign n43353 = n11368 & n43352 ;
  assign n43357 = n43356 ^ n43353 ^ 1'b0 ;
  assign n43358 = ~n26124 & n41524 ;
  assign n43359 = n43358 ^ n31205 ^ 1'b0 ;
  assign n43360 = ~n6630 & n30885 ;
  assign n43361 = n31846 ^ n10990 ^ 1'b0 ;
  assign n43362 = n12002 & n22413 ;
  assign n43363 = n43362 ^ n5079 ^ 1'b0 ;
  assign n43364 = n38789 | n43363 ;
  assign n43365 = n7839 | n35657 ;
  assign n43366 = n20010 & ~n43365 ;
  assign n43367 = n35582 ^ n8437 ^ 1'b0 ;
  assign n43368 = n15542 & n43367 ;
  assign n43369 = n15136 | n43368 ;
  assign n43370 = n26624 ^ n20858 ^ 1'b0 ;
  assign n43371 = n20339 | n43370 ;
  assign n43373 = ~n2791 & n37685 ;
  assign n43372 = n2266 | n40655 ;
  assign n43374 = n43373 ^ n43372 ^ 1'b0 ;
  assign n43375 = ( n5961 & n17501 ) | ( n5961 & ~n40645 ) | ( n17501 & ~n40645 ) ;
  assign n43376 = n27642 ^ n23360 ^ n10525 ;
  assign n43377 = n9776 ^ n3776 ^ 1'b0 ;
  assign n43378 = n31821 ^ n25173 ^ n5965 ;
  assign n43379 = x82 & n43378 ;
  assign n43380 = ~n645 & n43379 ;
  assign n43381 = n43380 ^ n32308 ^ 1'b0 ;
  assign n43382 = ~n723 & n9962 ;
  assign n43383 = n663 | n24060 ;
  assign n43384 = n21697 & ~n43383 ;
  assign n43385 = n37029 ^ n14536 ^ 1'b0 ;
  assign n43386 = n4917 | n9731 ;
  assign n43387 = n16247 ^ n7497 ^ 1'b0 ;
  assign n43388 = n43386 & n43387 ;
  assign n43389 = n3466 & n7049 ;
  assign n43390 = n43389 ^ n14557 ^ 1'b0 ;
  assign n43391 = n18103 & n43390 ;
  assign n43392 = n43391 ^ n9582 ^ 1'b0 ;
  assign n43393 = n43388 & n43392 ;
  assign n43394 = n8088 ^ n2124 ^ n1822 ;
  assign n43395 = n604 & n43394 ;
  assign n43396 = ( n20137 & ~n21012 ) | ( n20137 & n26524 ) | ( ~n21012 & n26524 ) ;
  assign n43397 = ( n9718 & n21338 ) | ( n9718 & ~n27496 ) | ( n21338 & ~n27496 ) ;
  assign n43398 = n43396 & ~n43397 ;
  assign n43399 = ( n9598 & n14536 ) | ( n9598 & n43398 ) | ( n14536 & n43398 ) ;
  assign n43400 = n24194 ^ n727 ^ n711 ;
  assign n43401 = n12203 & ~n43400 ;
  assign n43402 = n6041 & n7950 ;
  assign n43403 = ~n32022 & n43402 ;
  assign n43404 = n43403 ^ n5963 ^ 1'b0 ;
  assign n43405 = n13287 & ~n16419 ;
  assign n43406 = n28704 & ~n42063 ;
  assign n43407 = ~n43405 & n43406 ;
  assign n43408 = n3854 | n23546 ;
  assign n43409 = n42471 ^ n8921 ^ n4200 ;
  assign n43410 = ( ~n5549 & n20574 ) | ( ~n5549 & n43409 ) | ( n20574 & n43409 ) ;
  assign n43411 = n11465 & n26617 ;
  assign n43412 = ~n13487 & n43411 ;
  assign n43413 = n38897 ^ n37088 ^ n13161 ;
  assign n43414 = n890 & ~n15341 ;
  assign n43417 = n12799 & ~n31164 ;
  assign n43418 = n614 | n3721 ;
  assign n43419 = n43417 | n43418 ;
  assign n43415 = n36916 ^ n20686 ^ 1'b0 ;
  assign n43416 = n18460 & n43415 ;
  assign n43420 = n43419 ^ n43416 ^ 1'b0 ;
  assign n43421 = n29080 ^ n6868 ^ 1'b0 ;
  assign n43422 = n32959 & n43060 ;
  assign n43423 = n23403 ^ n2887 ^ 1'b0 ;
  assign n43424 = n2698 ^ n743 ^ 1'b0 ;
  assign n43425 = n43424 ^ n28927 ^ n8564 ;
  assign n43426 = n4145 & ~n34123 ;
  assign n43427 = n43426 ^ n5010 ^ n2659 ;
  assign n43428 = n43427 ^ n32690 ^ 1'b0 ;
  assign n43429 = n5489 | n17178 ;
  assign n43430 = n43429 ^ n20793 ^ 1'b0 ;
  assign n43431 = n16362 ^ n12343 ^ 1'b0 ;
  assign n43432 = n11114 & ~n22769 ;
  assign n43433 = n43432 ^ n37450 ^ 1'b0 ;
  assign n43434 = n24510 | n43433 ;
  assign n43435 = n16691 ^ n5646 ^ 1'b0 ;
  assign n43436 = n13805 & ~n43435 ;
  assign n43437 = n20692 | n39114 ;
  assign n43438 = n43437 ^ n40436 ^ 1'b0 ;
  assign n43439 = n10402 & n30675 ;
  assign n43440 = n43439 ^ n41158 ^ 1'b0 ;
  assign n43441 = n42968 ^ n7154 ^ 1'b0 ;
  assign n43442 = n24835 | n43441 ;
  assign n43443 = n8923 | n15443 ;
  assign n43444 = n43443 ^ n2959 ^ 1'b0 ;
  assign n43445 = ( n12435 & ~n22348 ) | ( n12435 & n43444 ) | ( ~n22348 & n43444 ) ;
  assign n43446 = n7965 | n22035 ;
  assign n43447 = n27575 & ~n43446 ;
  assign n43448 = n28051 & n42124 ;
  assign n43449 = n9152 & n36522 ;
  assign n43450 = n43449 ^ n19850 ^ 1'b0 ;
  assign n43451 = n7857 | n15736 ;
  assign n43452 = n2596 & n29052 ;
  assign n43453 = ~n4518 & n20044 ;
  assign n43454 = n43453 ^ n12651 ^ 1'b0 ;
  assign n43455 = n26362 & ~n39868 ;
  assign n43456 = ~n24723 & n32860 ;
  assign n43457 = n43456 ^ n33368 ^ 1'b0 ;
  assign n43458 = n25986 ^ n677 ^ 1'b0 ;
  assign n43459 = n27831 ^ n5691 ^ 1'b0 ;
  assign n43460 = ( ~n14610 & n35476 ) | ( ~n14610 & n43459 ) | ( n35476 & n43459 ) ;
  assign n43461 = ~n3047 & n12443 ;
  assign n43462 = ( n1944 & n16143 ) | ( n1944 & ~n43461 ) | ( n16143 & ~n43461 ) ;
  assign n43463 = ( n7916 & n16808 ) | ( n7916 & ~n36527 ) | ( n16808 & ~n36527 ) ;
  assign n43464 = ~n6627 & n37301 ;
  assign n43465 = n43464 ^ n41952 ^ 1'b0 ;
  assign n43466 = n10563 ^ n10088 ^ 1'b0 ;
  assign n43467 = ~n13827 & n27563 ;
  assign n43468 = n26079 & n43467 ;
  assign n43469 = ( ~n25694 & n43466 ) | ( ~n25694 & n43468 ) | ( n43466 & n43468 ) ;
  assign n43470 = n10214 | n43469 ;
  assign n43471 = n6430 & ~n20087 ;
  assign n43472 = ~n27525 & n43471 ;
  assign n43473 = n9105 | n21711 ;
  assign n43474 = n8930 & ~n43473 ;
  assign n43475 = n10396 & n11488 ;
  assign n43476 = n9287 | n41777 ;
  assign n43477 = ~n13593 & n21573 ;
  assign n43478 = ~n32251 & n43477 ;
  assign n43479 = ( x179 & n7978 ) | ( x179 & n38273 ) | ( n7978 & n38273 ) ;
  assign n43480 = n714 | n29741 ;
  assign n43481 = n296 | n43480 ;
  assign n43482 = n22478 ^ n10757 ^ 1'b0 ;
  assign n43483 = n25607 & ~n43482 ;
  assign n43484 = ~n16686 & n43483 ;
  assign n43485 = n43484 ^ n10863 ^ 1'b0 ;
  assign n43486 = n7143 & n11584 ;
  assign n43487 = n43486 ^ n17495 ^ 1'b0 ;
  assign n43488 = n22465 & n43487 ;
  assign n43489 = ~n2483 & n43488 ;
  assign n43490 = n25298 ^ n770 ^ 1'b0 ;
  assign n43491 = n19538 & n35910 ;
  assign n43492 = n43491 ^ n3366 ^ 1'b0 ;
  assign n43496 = n7308 & ~n28417 ;
  assign n43493 = n2248 & ~n7411 ;
  assign n43494 = ~n1622 & n43493 ;
  assign n43495 = n14047 & ~n43494 ;
  assign n43497 = n43496 ^ n43495 ^ 1'b0 ;
  assign n43498 = n43497 ^ n3161 ^ 1'b0 ;
  assign n43499 = n30524 ^ n1946 ^ 1'b0 ;
  assign n43500 = n35305 & ~n43499 ;
  assign n43501 = n648 & n13754 ;
  assign n43502 = n43501 ^ n21255 ^ 1'b0 ;
  assign n43503 = ~n514 & n4272 ;
  assign n43504 = ~n8623 & n43503 ;
  assign n43505 = n43504 ^ n26087 ^ n18589 ;
  assign n43506 = n3531 | n43505 ;
  assign n43507 = n10474 & n43506 ;
  assign n43508 = n16381 & ~n22364 ;
  assign n43509 = n23617 ^ n17437 ^ n16078 ;
  assign n43510 = n22914 | n41139 ;
  assign n43511 = n43510 ^ n13741 ^ 1'b0 ;
  assign n43512 = ( n29012 & ~n39845 ) | ( n29012 & n43511 ) | ( ~n39845 & n43511 ) ;
  assign n43513 = ~n16654 & n18172 ;
  assign n43514 = n43513 ^ n13196 ^ 1'b0 ;
  assign n43515 = n16714 & n24967 ;
  assign n43516 = ~n2702 & n43515 ;
  assign n43517 = n11844 | n19386 ;
  assign n43518 = ( n24284 & n29174 ) | ( n24284 & ~n40198 ) | ( n29174 & ~n40198 ) ;
  assign n43519 = n15723 & n18871 ;
  assign n43520 = n43518 & n43519 ;
  assign n43521 = ~n17226 & n34102 ;
  assign n43522 = n43520 & n43521 ;
  assign n43523 = n40220 & ~n40556 ;
  assign n43524 = n20159 & n24136 ;
  assign n43525 = ~n43523 & n43524 ;
  assign n43526 = ~n9222 & n22905 ;
  assign n43527 = ~n11667 & n43526 ;
  assign n43528 = n21358 & n31240 ;
  assign n43529 = ~n13920 & n43528 ;
  assign n43530 = n8377 & ~n43529 ;
  assign n43531 = n27597 & n43530 ;
  assign n43532 = n25602 ^ n1708 ^ 1'b0 ;
  assign n43533 = ~n27660 & n43532 ;
  assign n43534 = ( n4934 & n28198 ) | ( n4934 & ~n31132 ) | ( n28198 & ~n31132 ) ;
  assign n43535 = n2816 | n8260 ;
  assign n43536 = n40323 ^ n22040 ^ n4331 ;
  assign n43539 = n2937 & ~n17007 ;
  assign n43540 = n43539 ^ n824 ^ 1'b0 ;
  assign n43537 = n14983 & ~n22042 ;
  assign n43538 = ~n32419 & n43537 ;
  assign n43541 = n43540 ^ n43538 ^ 1'b0 ;
  assign n43542 = n1136 | n43541 ;
  assign n43543 = n8250 & ~n11908 ;
  assign n43544 = ~n3642 & n43543 ;
  assign n43545 = n3196 & n4721 ;
  assign n43546 = ~n42116 & n43545 ;
  assign n43547 = n22665 & ~n39346 ;
  assign n43548 = n26016 & n43547 ;
  assign n43549 = ( n19374 & n25215 ) | ( n19374 & ~n33920 ) | ( n25215 & ~n33920 ) ;
  assign n43550 = n3272 & n11900 ;
  assign n43551 = ~n759 & n43550 ;
  assign n43552 = ( n10701 & n12776 ) | ( n10701 & n43551 ) | ( n12776 & n43551 ) ;
  assign n43553 = n2058 & ~n6348 ;
  assign n43554 = n43553 ^ n30404 ^ n4654 ;
  assign n43555 = n5683 & n6796 ;
  assign n43556 = ~n23797 & n43555 ;
  assign n43557 = n7871 | n20414 ;
  assign n43558 = n4990 | n35060 ;
  assign n43559 = n4765 | n43558 ;
  assign n43560 = n10737 & n43559 ;
  assign n43561 = n43560 ^ n4404 ^ 1'b0 ;
  assign n43562 = n29836 & ~n37404 ;
  assign n43563 = n43562 ^ n36472 ^ 1'b0 ;
  assign n43564 = ~n8964 & n10994 ;
  assign n43565 = n3604 | n43462 ;
  assign n43566 = n33313 ^ n12612 ^ 1'b0 ;
  assign n43567 = n3052 & n6409 ;
  assign n43568 = n43567 ^ n4971 ^ 1'b0 ;
  assign n43569 = n43568 ^ n41994 ^ 1'b0 ;
  assign n43570 = n36483 ^ n23221 ^ 1'b0 ;
  assign n43571 = n43569 & n43570 ;
  assign n43572 = n9219 & n27807 ;
  assign n43573 = n34990 & n43572 ;
  assign n43574 = ~n3894 & n40730 ;
  assign n43575 = ~n41324 & n43574 ;
  assign n43576 = n32279 & n41460 ;
  assign n43577 = ~x17 & n858 ;
  assign n43578 = n21276 ^ n6036 ^ 1'b0 ;
  assign n43579 = n2836 & n43578 ;
  assign n43580 = ( n7378 & n25005 ) | ( n7378 & n43579 ) | ( n25005 & n43579 ) ;
  assign n43581 = n7629 & n37553 ;
  assign n43582 = ~n32044 & n39066 ;
  assign n43583 = ~n43581 & n43582 ;
  assign n43589 = ~n1639 & n22629 ;
  assign n43584 = n2689 & ~n19081 ;
  assign n43585 = n43584 ^ n15616 ^ 1'b0 ;
  assign n43586 = n15808 | n43585 ;
  assign n43587 = n43586 ^ n4845 ^ 1'b0 ;
  assign n43588 = n1801 | n43587 ;
  assign n43590 = n43589 ^ n43588 ^ 1'b0 ;
  assign n43591 = n43590 ^ n6885 ^ 1'b0 ;
  assign n43592 = ~n34350 & n43591 ;
  assign n43593 = ~n875 & n43592 ;
  assign n43594 = ~n645 & n39627 ;
  assign n43595 = n12350 | n21673 ;
  assign n43596 = n43595 ^ n7559 ^ 1'b0 ;
  assign n43597 = n43596 ^ n24208 ^ 1'b0 ;
  assign n43598 = n7499 | n43597 ;
  assign n43599 = n2298 & n31904 ;
  assign n43600 = n43599 ^ n12317 ^ 1'b0 ;
  assign n43601 = n43600 ^ n5099 ^ 1'b0 ;
  assign n43602 = n35831 & n43601 ;
  assign n43603 = n13305 & ~n35968 ;
  assign n43604 = ( n2680 & ~n15535 ) | ( n2680 & n27222 ) | ( ~n15535 & n27222 ) ;
  assign n43605 = n43604 ^ n38165 ^ 1'b0 ;
  assign n43606 = n34691 ^ n30227 ^ n28872 ;
  assign n43608 = n17128 & ~n26873 ;
  assign n43607 = ~n12786 & n35183 ;
  assign n43609 = n43608 ^ n43607 ^ n10121 ;
  assign n43610 = n31587 ^ n16812 ^ 1'b0 ;
  assign n43611 = ~n12231 & n43610 ;
  assign n43612 = ~n456 & n22836 ;
  assign n43613 = n43612 ^ n40115 ^ 1'b0 ;
  assign n43614 = n8458 ^ n6279 ^ 1'b0 ;
  assign n43615 = n43614 ^ n43419 ^ n15403 ;
  assign n43616 = n39974 | n43615 ;
  assign n43617 = n20156 & ~n43616 ;
  assign n43618 = n24831 ^ n16238 ^ 1'b0 ;
  assign n43619 = n28531 & n43618 ;
  assign n43620 = n27647 & n43619 ;
  assign n43621 = n21084 ^ n11770 ^ n2768 ;
  assign n43622 = n6931 & ~n43621 ;
  assign n43623 = ~n987 & n43622 ;
  assign n43627 = ( n524 & ~n7980 ) | ( n524 & n36609 ) | ( ~n7980 & n36609 ) ;
  assign n43624 = n23571 | n32566 ;
  assign n43625 = n24175 & n43624 ;
  assign n43626 = n20979 & n43625 ;
  assign n43628 = n43627 ^ n43626 ^ n25291 ;
  assign n43629 = n6184 & ~n6432 ;
  assign n43630 = n43629 ^ n8902 ^ 1'b0 ;
  assign n43631 = n8029 | n19609 ;
  assign n43632 = n15459 | n22753 ;
  assign n43633 = n43632 ^ n25340 ^ 1'b0 ;
  assign n43634 = ~n1030 & n23513 ;
  assign n43635 = ~n8651 & n32774 ;
  assign n43636 = ~n8999 & n43635 ;
  assign n43637 = n43634 & ~n43636 ;
  assign n43638 = ~n5235 & n19298 ;
  assign n43639 = n9201 & n23282 ;
  assign n43640 = n38461 & n43639 ;
  assign n43641 = ~n43638 & n43640 ;
  assign n43642 = n8266 | n16402 ;
  assign n43643 = n2829 & ~n43642 ;
  assign n43644 = n17504 | n41487 ;
  assign n43645 = n43644 ^ n18997 ^ 1'b0 ;
  assign n43646 = n11658 | n43645 ;
  assign n43647 = n38340 & ~n43646 ;
  assign n43648 = ( ~x170 & n853 ) | ( ~x170 & n26880 ) | ( n853 & n26880 ) ;
  assign n43649 = n9625 ^ n7014 ^ 1'b0 ;
  assign n43650 = n42193 ^ n29789 ^ 1'b0 ;
  assign n43651 = ( ~n1635 & n9648 ) | ( ~n1635 & n9820 ) | ( n9648 & n9820 ) ;
  assign n43652 = n19911 & n43651 ;
  assign n43653 = n43652 ^ n5592 ^ 1'b0 ;
  assign n43654 = n24347 ^ n20946 ^ 1'b0 ;
  assign n43655 = n1543 & ~n14366 ;
  assign n43656 = n7535 & ~n16078 ;
  assign n43657 = n43656 ^ n13571 ^ 1'b0 ;
  assign n43659 = n2444 & n33550 ;
  assign n43658 = n3443 & ~n43047 ;
  assign n43660 = n43659 ^ n43658 ^ 1'b0 ;
  assign n43661 = n2201 & ~n36950 ;
  assign n43662 = n43661 ^ n4410 ^ 1'b0 ;
  assign n43663 = n17845 ^ n10326 ^ 1'b0 ;
  assign n43664 = ~n15284 & n17867 ;
  assign n43665 = n43663 & n43664 ;
  assign n43666 = n15695 | n43665 ;
  assign n43667 = n43662 | n43666 ;
  assign n43668 = n21791 & ~n31084 ;
  assign n43669 = ~n28378 & n43668 ;
  assign n43670 = ( ~n18549 & n18551 ) | ( ~n18549 & n18660 ) | ( n18551 & n18660 ) ;
  assign n43671 = n43670 ^ n25752 ^ 1'b0 ;
  assign n43672 = n34825 & n43671 ;
  assign n43673 = n24268 | n43577 ;
  assign n43674 = n20832 & ~n43673 ;
  assign n43675 = n11083 ^ n3389 ^ 1'b0 ;
  assign n43676 = n6795 ^ n1967 ^ 1'b0 ;
  assign n43677 = ~n13589 & n43676 ;
  assign n43678 = n27914 ^ n7280 ^ 1'b0 ;
  assign n43679 = n16379 | n43678 ;
  assign n43680 = n43677 & n43679 ;
  assign n43681 = ~n43675 & n43680 ;
  assign n43682 = n39631 ^ n6577 ^ 1'b0 ;
  assign n43683 = n23272 ^ n3781 ^ 1'b0 ;
  assign n43684 = n12836 | n27315 ;
  assign n43685 = ~n12078 & n29188 ;
  assign n43686 = n43685 ^ n2337 ^ 1'b0 ;
  assign n43687 = n643 & n43686 ;
  assign n43688 = n43687 ^ n29678 ^ 1'b0 ;
  assign n43689 = n4852 | n25990 ;
  assign n43690 = n5211 | n43689 ;
  assign n43691 = n36853 & n43690 ;
  assign n43692 = n43691 ^ n29778 ^ 1'b0 ;
  assign n43693 = n29106 ^ n988 ^ 1'b0 ;
  assign n43694 = n28480 & ~n43693 ;
  assign n43695 = n3554 & n24793 ;
  assign n43696 = n36206 & ~n43695 ;
  assign n43697 = n6766 & ~n38821 ;
  assign n43698 = ~n11709 & n43697 ;
  assign n43699 = n12497 & ~n27936 ;
  assign n43700 = ~n806 & n43699 ;
  assign n43701 = n43700 ^ n14049 ^ 1'b0 ;
  assign n43702 = n1156 | n18775 ;
  assign n43703 = n9490 ^ n5793 ^ 1'b0 ;
  assign n43704 = n26723 & n37740 ;
  assign n43706 = ~n12310 & n18817 ;
  assign n43705 = ~n20957 & n27309 ;
  assign n43707 = n43706 ^ n43705 ^ 1'b0 ;
  assign n43708 = ~n26373 & n43707 ;
  assign n43709 = x210 & n21190 ;
  assign n43710 = n9363 | n43709 ;
  assign n43711 = n5837 ^ n620 ^ 1'b0 ;
  assign n43712 = ( n24328 & ~n30814 ) | ( n24328 & n43711 ) | ( ~n30814 & n43711 ) ;
  assign n43713 = n9170 | n25488 ;
  assign n43714 = n1760 & n9091 ;
  assign n43715 = n14269 & n43714 ;
  assign n43716 = ~n22994 & n30639 ;
  assign n43717 = n43716 ^ n3363 ^ 1'b0 ;
  assign n43718 = ~n31541 & n42650 ;
  assign n43719 = n11258 & n43718 ;
  assign n43720 = n13151 ^ n1715 ^ 1'b0 ;
  assign n43721 = ~n23095 & n43720 ;
  assign n43722 = n21949 ^ n3142 ^ 1'b0 ;
  assign n43723 = n2530 | n43722 ;
  assign n43724 = n7099 & ~n43723 ;
  assign n43725 = n40497 ^ n6870 ^ 1'b0 ;
  assign n43726 = n17634 ^ n14434 ^ n4010 ;
  assign n43727 = n43726 ^ n3903 ^ n2180 ;
  assign n43728 = n22729 ^ n12213 ^ 1'b0 ;
  assign n43729 = ~n36219 & n43728 ;
  assign n43730 = n43729 ^ n14239 ^ 1'b0 ;
  assign n43732 = n1212 & ~n9525 ;
  assign n43731 = n21100 | n33482 ;
  assign n43733 = n43732 ^ n43731 ^ 1'b0 ;
  assign n43734 = n29639 ^ n22722 ^ 1'b0 ;
  assign n43735 = n43733 & n43734 ;
  assign n43736 = n14002 ^ n4746 ^ 1'b0 ;
  assign n43737 = ~n15624 & n43736 ;
  assign n43738 = n16480 & n43737 ;
  assign n43739 = n13458 & ~n14165 ;
  assign n43740 = n10314 ^ n3908 ^ 1'b0 ;
  assign n43741 = n3257 ^ n547 ^ 1'b0 ;
  assign n43742 = n38721 ^ n12956 ^ 1'b0 ;
  assign n43743 = n30299 | n43742 ;
  assign n43744 = n33902 & ~n43743 ;
  assign n43745 = n15025 & ~n20150 ;
  assign n43746 = n9461 ^ n2441 ^ 1'b0 ;
  assign n43747 = n43746 ^ n35677 ^ n28181 ;
  assign n43748 = n2224 | n36652 ;
  assign n43749 = n14636 & ~n30338 ;
  assign n43750 = n30250 ^ n1030 ^ 1'b0 ;
  assign n43751 = n13347 | n43750 ;
  assign n43752 = n2937 & n20850 ;
  assign n43753 = n1419 & n43752 ;
  assign n43754 = n12601 | n43753 ;
  assign n43755 = n9099 & ~n43754 ;
  assign n43756 = n24083 & n28634 ;
  assign n43757 = n43756 ^ n4509 ^ 1'b0 ;
  assign n43761 = n30529 ^ n8781 ^ n5143 ;
  assign n43760 = n6825 & n9559 ;
  assign n43758 = n15985 ^ n6488 ^ 1'b0 ;
  assign n43759 = ~n41573 & n43758 ;
  assign n43762 = n43761 ^ n43760 ^ n43759 ;
  assign n43763 = ~x228 & n5996 ;
  assign n43764 = n13765 & n25039 ;
  assign n43765 = n21874 & n43764 ;
  assign n43766 = n21071 | n43765 ;
  assign n43767 = n43766 ^ n25300 ^ 1'b0 ;
  assign n43768 = n3361 | n43767 ;
  assign n43769 = ~n1574 & n20030 ;
  assign n43770 = n43769 ^ n42761 ^ 1'b0 ;
  assign n43771 = n43770 ^ n42253 ^ 1'b0 ;
  assign n43772 = n28810 & ~n39344 ;
  assign n43773 = n9835 & ~n14116 ;
  assign n43774 = ~n1706 & n11328 ;
  assign n43775 = ~n12002 & n43774 ;
  assign n43776 = n43775 ^ n2686 ^ 1'b0 ;
  assign n43777 = n43776 ^ n2995 ^ 1'b0 ;
  assign n43778 = ~n3891 & n43777 ;
  assign n43779 = n15141 ^ n13659 ^ n11075 ;
  assign n43780 = n5699 & n19325 ;
  assign n43781 = ( n2699 & n25018 ) | ( n2699 & ~n43780 ) | ( n25018 & ~n43780 ) ;
  assign n43782 = ( ~n10188 & n18265 ) | ( ~n10188 & n18317 ) | ( n18265 & n18317 ) ;
  assign n43783 = n6954 & ~n8773 ;
  assign n43784 = n12350 & n43783 ;
  assign n43785 = n14027 | n43784 ;
  assign n43786 = n14219 | n43785 ;
  assign n43787 = n43782 & n43786 ;
  assign n43788 = n5903 | n13040 ;
  assign n43789 = n28995 ^ n5550 ^ 1'b0 ;
  assign n43790 = n5807 & n43789 ;
  assign n43791 = n18222 & n43790 ;
  assign n43792 = n13146 | n23349 ;
  assign n43793 = n15183 & ~n43792 ;
  assign n43794 = n21984 | n43793 ;
  assign n43795 = n27914 | n43794 ;
  assign n43796 = n14242 ^ n11261 ^ 1'b0 ;
  assign n43797 = n30924 | n43796 ;
  assign n43798 = n10724 & ~n43797 ;
  assign n43799 = n18410 ^ n13009 ^ 1'b0 ;
  assign n43800 = n9610 & ~n43799 ;
  assign n43801 = n43800 ^ n37580 ^ n20335 ;
  assign n43802 = n11997 & n29188 ;
  assign n43803 = n21788 ^ n13889 ^ 1'b0 ;
  assign n43804 = ( ~n5176 & n43802 ) | ( ~n5176 & n43803 ) | ( n43802 & n43803 ) ;
  assign n43805 = ~n13650 & n43804 ;
  assign n43806 = ~n3773 & n27056 ;
  assign n43807 = n21025 ^ x178 ^ 1'b0 ;
  assign n43808 = n21223 & ~n30085 ;
  assign n43809 = n30602 ^ n9496 ^ 1'b0 ;
  assign n43810 = n22030 & n43809 ;
  assign n43811 = ~n23815 & n43810 ;
  assign n43812 = n43811 ^ n31498 ^ 1'b0 ;
  assign n43813 = n14813 ^ n3709 ^ n1998 ;
  assign n43814 = n31058 ^ n11915 ^ 1'b0 ;
  assign n43815 = n2448 & ~n43814 ;
  assign n43816 = n43815 ^ n8340 ^ 1'b0 ;
  assign n43817 = n13556 & ~n43816 ;
  assign n43818 = ( ~n31789 & n43813 ) | ( ~n31789 & n43817 ) | ( n43813 & n43817 ) ;
  assign n43819 = ( n11227 & n11312 ) | ( n11227 & n41614 ) | ( n11312 & n41614 ) ;
  assign n43820 = ~n6737 & n11863 ;
  assign n43821 = n43820 ^ n18037 ^ 1'b0 ;
  assign n43822 = n19978 ^ n13413 ^ n4831 ;
  assign n43823 = n31062 ^ n8138 ^ n5876 ;
  assign n43824 = n15242 & n43823 ;
  assign n43825 = n19733 ^ n2675 ^ 1'b0 ;
  assign n43826 = ~n19665 & n43825 ;
  assign n43827 = n40912 ^ n8503 ^ n6484 ;
  assign n43828 = ~n19578 & n43827 ;
  assign n43829 = ( n7485 & n9914 ) | ( n7485 & n43828 ) | ( n9914 & n43828 ) ;
  assign n43830 = n3627 ^ n527 ^ 1'b0 ;
  assign n43831 = n24403 & ~n43830 ;
  assign n43832 = n43831 ^ n849 ^ 1'b0 ;
  assign n43833 = n43832 ^ n33823 ^ n5131 ;
  assign n43834 = n4996 & n13146 ;
  assign n43835 = ( n1509 & ~n17430 ) | ( n1509 & n23153 ) | ( ~n17430 & n23153 ) ;
  assign n43836 = n43835 ^ n18585 ^ 1'b0 ;
  assign n43837 = ~n4002 & n7605 ;
  assign n43838 = ( n3404 & ~n15930 ) | ( n3404 & n34815 ) | ( ~n15930 & n34815 ) ;
  assign n43839 = n43837 & n43838 ;
  assign n43840 = n43839 ^ n3883 ^ 1'b0 ;
  assign n43841 = n34404 ^ n19021 ^ n14129 ;
  assign n43842 = n43841 ^ n2345 ^ 1'b0 ;
  assign n43843 = ~n3552 & n43842 ;
  assign n43844 = n11650 ^ n3340 ^ 1'b0 ;
  assign n43845 = n16149 & n43844 ;
  assign n43846 = n23784 ^ n13623 ^ 1'b0 ;
  assign n43847 = ( n890 & n8789 ) | ( n890 & n23512 ) | ( n8789 & n23512 ) ;
  assign n43848 = n353 | n7925 ;
  assign n43849 = n43848 ^ n38008 ^ n15227 ;
  assign n43850 = n3439 & n9403 ;
  assign n43851 = n12663 & n43850 ;
  assign n43852 = n25461 & ~n43851 ;
  assign n43853 = n3981 & n5896 ;
  assign n43854 = n15465 & n43853 ;
  assign n43855 = n38433 ^ n7776 ^ 1'b0 ;
  assign n43856 = n9979 & ~n43855 ;
  assign n43857 = n19278 & n28173 ;
  assign n43858 = n32272 | n34072 ;
  assign n43859 = n42987 ^ n10827 ^ 1'b0 ;
  assign n43860 = ~n43858 & n43859 ;
  assign n43861 = n1291 ^ n704 ^ 1'b0 ;
  assign n43862 = n33798 ^ n5057 ^ n2915 ;
  assign n43863 = n31911 & n43862 ;
  assign n43864 = ~n7428 & n27099 ;
  assign n43865 = n43864 ^ n23937 ^ n21697 ;
  assign n43866 = ( ~n12355 & n41716 ) | ( ~n12355 & n43865 ) | ( n41716 & n43865 ) ;
  assign n43867 = x139 & ~n26201 ;
  assign n43868 = n43867 ^ n791 ^ 1'b0 ;
  assign n43869 = n43868 ^ n39812 ^ n29742 ;
  assign n43870 = x175 & n33397 ;
  assign n43871 = x22 & n43870 ;
  assign n43872 = n43871 ^ n2149 ^ 1'b0 ;
  assign n43873 = n36866 & n43872 ;
  assign n43874 = n14450 ^ n10926 ^ n2114 ;
  assign n43875 = n5851 | n37272 ;
  assign n43876 = n15770 ^ n14605 ^ n12822 ;
  assign n43877 = n43140 ^ n13195 ^ 1'b0 ;
  assign n43878 = n7544 | n11158 ;
  assign n43879 = n759 & ~n13373 ;
  assign n43880 = ~n43878 & n43879 ;
  assign n43881 = ( ~n36740 & n43877 ) | ( ~n36740 & n43880 ) | ( n43877 & n43880 ) ;
  assign n43882 = n19982 ^ n10510 ^ 1'b0 ;
  assign n43883 = n24757 ^ n4099 ^ 1'b0 ;
  assign n43884 = n12595 | n26744 ;
  assign n43885 = ~n21151 & n23336 ;
  assign n43886 = n43885 ^ n835 ^ 1'b0 ;
  assign n43887 = n9445 | n43886 ;
  assign n43888 = n43884 | n43887 ;
  assign n43889 = n8787 ^ n6271 ^ 1'b0 ;
  assign n43890 = n20578 & ~n43889 ;
  assign n43891 = n38573 ^ n14178 ^ 1'b0 ;
  assign n43892 = n24084 & n43891 ;
  assign n43893 = n26091 ^ n15533 ^ 1'b0 ;
  assign n43894 = ~n9422 & n17230 ;
  assign n43895 = n30079 & n43894 ;
  assign n43896 = n20323 ^ n7418 ^ 1'b0 ;
  assign n43897 = ( n43893 & n43895 ) | ( n43893 & ~n43896 ) | ( n43895 & ~n43896 ) ;
  assign n43898 = n29731 ^ n20974 ^ 1'b0 ;
  assign n43899 = ~n24318 & n35802 ;
  assign n43900 = n43899 ^ n22256 ^ 1'b0 ;
  assign n43901 = ~n4120 & n15861 ;
  assign n43902 = n43901 ^ n13644 ^ 1'b0 ;
  assign n43903 = n31832 ^ n5910 ^ 1'b0 ;
  assign n43904 = ~n1233 & n9607 ;
  assign n43905 = ( ~n7073 & n22189 ) | ( ~n7073 & n43904 ) | ( n22189 & n43904 ) ;
  assign n43906 = x133 & n38090 ;
  assign n43907 = n43905 & n43906 ;
  assign n43908 = ~n9353 & n22613 ;
  assign n43909 = n15829 & ~n30901 ;
  assign n43910 = n995 | n14496 ;
  assign n43911 = ( ~n3210 & n23886 ) | ( ~n3210 & n43910 ) | ( n23886 & n43910 ) ;
  assign n43912 = n12876 & ~n43911 ;
  assign n43913 = n16332 & n43912 ;
  assign n43914 = n38790 & ~n43913 ;
  assign n43915 = n4783 | n21717 ;
  assign n43916 = ( n26334 & ~n31412 ) | ( n26334 & n43915 ) | ( ~n31412 & n43915 ) ;
  assign n43917 = n1013 & ~n26531 ;
  assign n43918 = n3814 | n43917 ;
  assign n43919 = n16492 | n43918 ;
  assign n43920 = n2006 & ~n2965 ;
  assign n43921 = n43920 ^ n886 ^ 1'b0 ;
  assign n43922 = n43921 ^ n10850 ^ 1'b0 ;
  assign n43923 = n9860 & ~n43922 ;
  assign n43924 = ( n28085 & ~n43919 ) | ( n28085 & n43923 ) | ( ~n43919 & n43923 ) ;
  assign n43925 = n32146 ^ n19178 ^ 1'b0 ;
  assign n43926 = n10859 & ~n43925 ;
  assign n43927 = n8005 | n43926 ;
  assign n43928 = ~n23755 & n35084 ;
  assign n43929 = n23672 | n43928 ;
  assign n43930 = n24119 & ~n43929 ;
  assign n43931 = n14408 ^ n11950 ^ 1'b0 ;
  assign n43932 = n27324 & ~n43931 ;
  assign n43933 = n14071 & ~n19794 ;
  assign n43934 = n5338 & n43933 ;
  assign n43935 = n11930 | n36198 ;
  assign n43936 = n11171 & n11543 ;
  assign n43937 = n43936 ^ n31742 ^ n28932 ;
  assign n43938 = n19138 & ~n43937 ;
  assign n43939 = n8556 & n8934 ;
  assign n43940 = n43939 ^ n40543 ^ 1'b0 ;
  assign n43941 = n29604 & n43940 ;
  assign n43942 = ( ~n7029 & n8902 ) | ( ~n7029 & n43941 ) | ( n8902 & n43941 ) ;
  assign n43943 = n27022 ^ n3909 ^ 1'b0 ;
  assign n43944 = n13217 ^ n10183 ^ 1'b0 ;
  assign n43945 = ( n5065 & ~n15585 ) | ( n5065 & n21498 ) | ( ~n15585 & n21498 ) ;
  assign n43946 = n43945 ^ n20514 ^ n15758 ;
  assign n43947 = n43944 & n43946 ;
  assign n43952 = ~n13640 & n23614 ;
  assign n43953 = n15772 & n43952 ;
  assign n43954 = ~x220 & n43953 ;
  assign n43949 = n14954 ^ n1274 ^ 1'b0 ;
  assign n43948 = ~n10856 & n11772 ;
  assign n43950 = n43949 ^ n43948 ^ 1'b0 ;
  assign n43951 = n29536 | n43950 ;
  assign n43955 = n43954 ^ n43951 ^ 1'b0 ;
  assign n43956 = n936 & ~n22547 ;
  assign n43957 = n43956 ^ n5719 ^ 1'b0 ;
  assign n43958 = n32122 & ~n39827 ;
  assign n43959 = n38229 ^ n9577 ^ 1'b0 ;
  assign n43960 = n9752 & n43959 ;
  assign n43961 = ~n33489 & n35732 ;
  assign n43962 = ~n13906 & n33990 ;
  assign n43963 = n10168 & n43962 ;
  assign n43964 = n43963 ^ n15618 ^ n418 ;
  assign n43966 = n41800 ^ n26621 ^ n14498 ;
  assign n43965 = ~n9676 & n14352 ;
  assign n43967 = n43966 ^ n43965 ^ n15806 ;
  assign n43968 = ~n17184 & n18894 ;
  assign n43969 = ~n13715 & n43968 ;
  assign n43970 = n6814 | n17392 ;
  assign n43971 = ~n32056 & n43970 ;
  assign n43972 = ~n26541 & n43971 ;
  assign n43973 = n3015 & n3493 ;
  assign n43974 = n22715 ^ n2898 ^ 1'b0 ;
  assign n43975 = ~n43973 & n43974 ;
  assign n43976 = n10925 ^ n2042 ^ 1'b0 ;
  assign n43977 = ~n4880 & n43976 ;
  assign n43978 = n43977 ^ n13380 ^ 1'b0 ;
  assign n43979 = ~n393 & n43978 ;
  assign n43980 = n20070 ^ n3905 ^ 1'b0 ;
  assign n43981 = n11655 | n26852 ;
  assign n43982 = n3425 | n25319 ;
  assign n43983 = n13413 | n27456 ;
  assign n43984 = n43983 ^ n12229 ^ 1'b0 ;
  assign n43985 = n43984 ^ n7135 ^ n4646 ;
  assign n43986 = ~n25353 & n29842 ;
  assign n43987 = n17324 ^ n3910 ^ 1'b0 ;
  assign n43988 = x81 | n43987 ;
  assign n43989 = n18383 ^ n3104 ^ 1'b0 ;
  assign n43990 = n43988 | n43989 ;
  assign n43991 = n43990 ^ n7359 ^ 1'b0 ;
  assign n43992 = n18257 & ~n21288 ;
  assign n43993 = n25381 & n43992 ;
  assign n43994 = n23490 ^ n10779 ^ 1'b0 ;
  assign n43995 = n1635 | n16052 ;
  assign n43996 = n37638 ^ n12546 ^ 1'b0 ;
  assign n43997 = n43995 | n43996 ;
  assign n43998 = n508 & ~n3433 ;
  assign n43999 = n7567 & ~n43998 ;
  assign n44000 = n43999 ^ n34473 ^ 1'b0 ;
  assign n44001 = ~n9172 & n13122 ;
  assign n44002 = n9350 & n44001 ;
  assign n44003 = n35845 ^ n7764 ^ 1'b0 ;
  assign n44006 = n28318 & ~n37220 ;
  assign n44007 = n44006 ^ n33807 ^ 1'b0 ;
  assign n44004 = n4647 & n6605 ;
  assign n44005 = ( n12624 & n14395 ) | ( n12624 & ~n44004 ) | ( n14395 & ~n44004 ) ;
  assign n44008 = n44007 ^ n44005 ^ n35360 ;
  assign n44009 = n10643 ^ n7431 ^ 1'b0 ;
  assign n44010 = n14382 & n44009 ;
  assign n44011 = n21523 | n24829 ;
  assign n44012 = ~n1998 & n8752 ;
  assign n44013 = n3326 & n19374 ;
  assign n44014 = ~n20439 & n44013 ;
  assign n44015 = n783 & ~n1474 ;
  assign n44016 = n15978 & n22066 ;
  assign n44017 = ~n44015 & n44016 ;
  assign n44018 = n44017 ^ n6754 ^ 1'b0 ;
  assign n44019 = ~n23484 & n44018 ;
  assign n44020 = ~n2305 & n20546 ;
  assign n44021 = n17366 & n20519 ;
  assign n44022 = ~n33539 & n44021 ;
  assign n44023 = n34154 & ~n44022 ;
  assign n44024 = n40226 ^ n10338 ^ 1'b0 ;
  assign n44025 = n32705 | n44024 ;
  assign n44026 = n30051 ^ n19876 ^ 1'b0 ;
  assign n44027 = ~n26979 & n43089 ;
  assign n44028 = n44027 ^ n31877 ^ 1'b0 ;
  assign n44029 = ~n8033 & n27404 ;
  assign n44030 = n44029 ^ n11486 ^ 1'b0 ;
  assign n44031 = n511 & n44030 ;
  assign n44032 = n11442 & ~n29923 ;
  assign n44033 = n1561 | n2067 ;
  assign n44034 = n23936 & ~n44033 ;
  assign n44035 = n44034 ^ n8022 ^ n6352 ;
  assign n44039 = x81 | n966 ;
  assign n44036 = n8189 | n25381 ;
  assign n44037 = n14877 | n44036 ;
  assign n44038 = n44037 ^ n42086 ^ n13605 ;
  assign n44040 = n44039 ^ n44038 ^ n39163 ;
  assign n44041 = n12763 & n30689 ;
  assign n44042 = n44041 ^ n25387 ^ 1'b0 ;
  assign n44043 = n1826 & ~n14112 ;
  assign n44044 = ~n15372 & n44043 ;
  assign n44045 = n19934 ^ n19438 ^ 1'b0 ;
  assign n44046 = ~n44044 & n44045 ;
  assign n44047 = n4390 ^ n4194 ^ 1'b0 ;
  assign n44048 = n2137 | n29361 ;
  assign n44049 = n2733 | n17788 ;
  assign n44050 = n44049 ^ n12359 ^ 1'b0 ;
  assign n44051 = n44050 ^ n18594 ^ 1'b0 ;
  assign n44052 = n21757 ^ n11316 ^ n9612 ;
  assign n44053 = ~n5269 & n43010 ;
  assign n44054 = n37225 & n44053 ;
  assign n44055 = n16100 ^ n7992 ^ n6375 ;
  assign n44056 = x180 & n44055 ;
  assign n44057 = n8420 & n44056 ;
  assign n44058 = ~n5676 & n44057 ;
  assign n44059 = n41989 ^ n11165 ^ 1'b0 ;
  assign n44060 = n6451 | n44059 ;
  assign n44061 = ~n10767 & n34633 ;
  assign n44062 = n29808 & n44061 ;
  assign n44063 = n3742 | n12044 ;
  assign n44064 = n44063 ^ n39751 ^ 1'b0 ;
  assign n44065 = ( ~n2168 & n40120 ) | ( ~n2168 & n44064 ) | ( n40120 & n44064 ) ;
  assign n44066 = n2513 & ~n39105 ;
  assign n44067 = ~n44065 & n44066 ;
  assign n44068 = n8190 & n27445 ;
  assign n44069 = n44068 ^ n11515 ^ 1'b0 ;
  assign n44070 = n31471 & ~n44069 ;
  assign n44071 = ( ~n3448 & n28069 ) | ( ~n3448 & n31653 ) | ( n28069 & n31653 ) ;
  assign n44072 = n25412 | n44071 ;
  assign n44073 = n44072 ^ n40473 ^ 1'b0 ;
  assign n44074 = n41514 ^ n26281 ^ n23634 ;
  assign n44075 = ( n25115 & n40335 ) | ( n25115 & n44074 ) | ( n40335 & n44074 ) ;
  assign n44076 = n23883 ^ n1085 ^ 1'b0 ;
  assign n44077 = n3008 & ~n24928 ;
  assign n44078 = n12901 | n44077 ;
  assign n44079 = n22276 | n44078 ;
  assign n44080 = n44079 ^ n25018 ^ n11568 ;
  assign n44081 = n11706 ^ n10218 ^ 1'b0 ;
  assign n44082 = n44080 | n44081 ;
  assign n44083 = n32006 ^ n21214 ^ 1'b0 ;
  assign n44084 = n20805 | n44083 ;
  assign n44085 = n44084 ^ n14286 ^ 1'b0 ;
  assign n44086 = ~n2676 & n10764 ;
  assign n44087 = ( ~n867 & n14487 ) | ( ~n867 & n17628 ) | ( n14487 & n17628 ) ;
  assign n44088 = ~n31298 & n44087 ;
  assign n44089 = ( n376 & ~n44086 ) | ( n376 & n44088 ) | ( ~n44086 & n44088 ) ;
  assign n44090 = n7317 & ~n9836 ;
  assign n44091 = ( n8819 & n29693 ) | ( n8819 & n44090 ) | ( n29693 & n44090 ) ;
  assign n44092 = x144 & ~n44091 ;
  assign n44093 = n39805 ^ n26051 ^ 1'b0 ;
  assign n44094 = ~n9498 & n44093 ;
  assign n44095 = n11486 ^ n4179 ^ 1'b0 ;
  assign n44096 = ~n17051 & n44095 ;
  assign n44097 = n17420 & n44096 ;
  assign n44098 = n10181 & n44097 ;
  assign n44099 = n19481 ^ n7732 ^ 1'b0 ;
  assign n44100 = n7471 | n44099 ;
  assign n44101 = n44098 & ~n44100 ;
  assign n44102 = n19118 & n33709 ;
  assign n44103 = ~n9562 & n44102 ;
  assign n44104 = n24602 | n33880 ;
  assign n44105 = n44104 ^ n14517 ^ 1'b0 ;
  assign n44106 = n1073 | n3232 ;
  assign n44107 = n2807 & ~n44106 ;
  assign n44108 = n44107 ^ n3746 ^ 1'b0 ;
  assign n44109 = n44108 ^ n25573 ^ 1'b0 ;
  assign n44110 = ~n2073 & n44109 ;
  assign n44112 = n11524 | n12974 ;
  assign n44113 = n44112 ^ n956 ^ 1'b0 ;
  assign n44114 = n8780 & n14886 ;
  assign n44115 = n19399 & n44114 ;
  assign n44116 = ( n12327 & ~n44113 ) | ( n12327 & n44115 ) | ( ~n44113 & n44115 ) ;
  assign n44111 = n13013 | n20824 ;
  assign n44117 = n44116 ^ n44111 ^ 1'b0 ;
  assign n44118 = ( n4585 & n21112 ) | ( n4585 & ~n36657 ) | ( n21112 & ~n36657 ) ;
  assign n44119 = ( n17271 & n19885 ) | ( n17271 & n24914 ) | ( n19885 & n24914 ) ;
  assign n44120 = n28652 ^ n28140 ^ 1'b0 ;
  assign n44121 = n28550 ^ n7431 ^ 1'b0 ;
  assign n44122 = n395 & ~n20366 ;
  assign n44123 = n44122 ^ n41229 ^ 1'b0 ;
  assign n44124 = n32204 | n44123 ;
  assign n44125 = n44124 ^ n5623 ^ 1'b0 ;
  assign n44126 = ~n10747 & n15328 ;
  assign n44127 = n23642 ^ n17614 ^ 1'b0 ;
  assign n44128 = n1575 & n44127 ;
  assign n44129 = n44128 ^ n24533 ^ 1'b0 ;
  assign n44130 = n10582 | n44129 ;
  assign n44131 = n39092 ^ n8453 ^ n6808 ;
  assign n44132 = n38790 ^ n30774 ^ n23932 ;
  assign n44133 = n24902 & ~n31804 ;
  assign n44134 = n44133 ^ n5740 ^ 1'b0 ;
  assign n44135 = n43936 ^ n27693 ^ 1'b0 ;
  assign n44136 = ~n8169 & n12019 ;
  assign n44137 = n12090 | n29988 ;
  assign n44138 = ( n2406 & n44136 ) | ( n2406 & n44137 ) | ( n44136 & n44137 ) ;
  assign n44139 = n29727 ^ n28392 ^ 1'b0 ;
  assign n44140 = ~n44138 & n44139 ;
  assign n44141 = n9542 & n16923 ;
  assign n44142 = ~n24701 & n44141 ;
  assign n44143 = n18432 ^ n4157 ^ 1'b0 ;
  assign n44144 = n314 & n34881 ;
  assign n44145 = n44144 ^ n33771 ^ 1'b0 ;
  assign n44146 = n37622 ^ n22373 ^ 1'b0 ;
  assign n44147 = ~n7349 & n9093 ;
  assign n44148 = n33639 ^ n2847 ^ 1'b0 ;
  assign n44149 = ~n25734 & n44148 ;
  assign n44150 = n44149 ^ n34591 ^ 1'b0 ;
  assign n44151 = n3545 | n11821 ;
  assign n44152 = ( ~n10138 & n15941 ) | ( ~n10138 & n19303 ) | ( n15941 & n19303 ) ;
  assign n44153 = n44152 ^ n3848 ^ 1'b0 ;
  assign n44154 = n1313 & n44153 ;
  assign n44155 = n16331 & n16411 ;
  assign n44156 = n44155 ^ n26060 ^ n5934 ;
  assign n44157 = n36704 & ~n44156 ;
  assign n44158 = n6257 & n14046 ;
  assign n44159 = ( n17665 & n21673 ) | ( n17665 & n30944 ) | ( n21673 & n30944 ) ;
  assign n44160 = n44159 ^ n20756 ^ 1'b0 ;
  assign n44161 = n44160 ^ n33769 ^ n4931 ;
  assign n44162 = n44161 ^ n31746 ^ 1'b0 ;
  assign n44163 = n6588 & n6904 ;
  assign n44164 = n37937 ^ n14756 ^ n3118 ;
  assign n44165 = n13056 & ~n19046 ;
  assign n44166 = n19820 & n33301 ;
  assign n44167 = ~n19303 & n44166 ;
  assign n44168 = ~n36488 & n44167 ;
  assign n44169 = ~n18173 & n22998 ;
  assign n44170 = n44169 ^ n8073 ^ 1'b0 ;
  assign n44171 = n44170 ^ n27524 ^ 1'b0 ;
  assign n44172 = n44064 ^ n17572 ^ n2896 ;
  assign n44173 = n43468 & ~n44172 ;
  assign n44174 = ~n12118 & n28706 ;
  assign n44175 = n44174 ^ n6375 ^ 1'b0 ;
  assign n44176 = ~n23479 & n44175 ;
  assign n44177 = n5054 | n11014 ;
  assign n44178 = n44177 ^ n1327 ^ 1'b0 ;
  assign n44179 = ( n23552 & n29326 ) | ( n23552 & n44178 ) | ( n29326 & n44178 ) ;
  assign n44180 = n35872 | n37276 ;
  assign n44181 = n31389 & ~n44180 ;
  assign n44182 = ~x155 & n44181 ;
  assign n44183 = n8443 & ~n44182 ;
  assign n44189 = n11475 & ~n17384 ;
  assign n44184 = x187 & n5090 ;
  assign n44185 = n44184 ^ n4959 ^ 1'b0 ;
  assign n44186 = ~n4744 & n44185 ;
  assign n44187 = n44186 ^ n950 ^ 1'b0 ;
  assign n44188 = n7930 | n44187 ;
  assign n44190 = n44189 ^ n44188 ^ n9990 ;
  assign n44191 = n43518 ^ n19631 ^ 1'b0 ;
  assign n44192 = n22545 & ~n44191 ;
  assign n44193 = n34355 ^ n12171 ^ 1'b0 ;
  assign n44194 = n18091 ^ n15825 ^ n5489 ;
  assign n44195 = n31848 & n44194 ;
  assign n44196 = n44195 ^ n35012 ^ 1'b0 ;
  assign n44197 = n44196 ^ n23674 ^ 1'b0 ;
  assign n44198 = n26392 & ~n44197 ;
  assign n44199 = n33781 ^ n22343 ^ 1'b0 ;
  assign n44200 = ( n7571 & ~n29249 ) | ( n7571 & n36262 ) | ( ~n29249 & n36262 ) ;
  assign n44201 = n4428 & n18335 ;
  assign n44202 = n34353 | n34815 ;
  assign n44203 = n44202 ^ n20678 ^ 1'b0 ;
  assign n44204 = n9432 | n26122 ;
  assign n44205 = ~n16238 & n26519 ;
  assign n44206 = n4911 ^ n4027 ^ 1'b0 ;
  assign n44207 = n44206 ^ n22429 ^ n2885 ;
  assign n44208 = n23407 ^ n20218 ^ n8058 ;
  assign n44209 = n12518 | n13225 ;
  assign n44210 = n44209 ^ n9297 ^ 1'b0 ;
  assign n44211 = n34355 | n44210 ;
  assign n44212 = n6819 & ~n8325 ;
  assign n44213 = n44212 ^ n13581 ^ 1'b0 ;
  assign n44214 = n15657 | n40866 ;
  assign n44215 = n27949 | n29138 ;
  assign n44216 = n32567 | n44215 ;
  assign n44217 = n6196 & ~n32240 ;
  assign n44218 = n44217 ^ n2661 ^ 1'b0 ;
  assign n44219 = n15561 & n36469 ;
  assign n44220 = ~n9833 & n21274 ;
  assign n44221 = n39158 ^ n8531 ^ 1'b0 ;
  assign n44222 = n6019 | n11518 ;
  assign n44223 = n2690 & n15222 ;
  assign n44224 = ~n14690 & n44223 ;
  assign n44225 = ~n12125 & n19393 ;
  assign n44226 = n24657 ^ n3554 ^ n2949 ;
  assign n44227 = n3205 & ~n44226 ;
  assign n44228 = ( n16322 & ~n22391 ) | ( n16322 & n44227 ) | ( ~n22391 & n44227 ) ;
  assign n44229 = n526 | n44228 ;
  assign n44230 = n15909 ^ n15403 ^ 1'b0 ;
  assign n44231 = n41553 ^ n41116 ^ n21993 ;
  assign n44232 = n37973 ^ n35400 ^ n11103 ;
  assign n44233 = n41034 ^ n16954 ^ 1'b0 ;
  assign n44234 = n579 & n3708 ;
  assign n44235 = n41231 ^ n11040 ^ 1'b0 ;
  assign n44236 = n15430 ^ n15404 ^ 1'b0 ;
  assign n44237 = ~n44235 & n44236 ;
  assign n44238 = n44237 ^ n21867 ^ 1'b0 ;
  assign n44239 = n3315 | n44238 ;
  assign n44240 = ~n11421 & n39353 ;
  assign n44241 = ~n10344 & n44240 ;
  assign n44242 = n7879 | n37502 ;
  assign n44243 = n18731 & ~n44242 ;
  assign n44244 = n23442 ^ n13926 ^ n2941 ;
  assign n44247 = n19025 ^ n7298 ^ n1040 ;
  assign n44245 = n7670 & n7843 ;
  assign n44246 = n44245 ^ n18797 ^ 1'b0 ;
  assign n44248 = n44247 ^ n44246 ^ n4016 ;
  assign n44249 = n2450 | n8912 ;
  assign n44250 = n36713 | n44249 ;
  assign n44251 = n19780 & n27653 ;
  assign n44252 = n44250 & n44251 ;
  assign n44253 = n37700 ^ n1228 ^ 1'b0 ;
  assign n44254 = n906 & ~n39257 ;
  assign n44255 = ~n36882 & n44254 ;
  assign n44256 = n27800 ^ n288 ^ 1'b0 ;
  assign n44257 = ~n23055 & n44256 ;
  assign n44258 = n2071 & n12806 ;
  assign n44259 = n44258 ^ n24932 ^ 1'b0 ;
  assign n44260 = n36527 ^ n24310 ^ n4205 ;
  assign n44261 = n9212 & n32299 ;
  assign n44262 = n44261 ^ n1285 ^ 1'b0 ;
  assign n44263 = ( ~n17625 & n43675 ) | ( ~n17625 & n44262 ) | ( n43675 & n44262 ) ;
  assign n44264 = ( ~n9621 & n31240 ) | ( ~n9621 & n32680 ) | ( n31240 & n32680 ) ;
  assign n44265 = n37550 ^ n27404 ^ 1'b0 ;
  assign n44266 = n2103 | n44265 ;
  assign n44267 = n37955 ^ n16954 ^ 1'b0 ;
  assign n44268 = n11857 | n44267 ;
  assign n44269 = n4247 & ~n5739 ;
  assign n44270 = n34254 ^ n5154 ^ 1'b0 ;
  assign n44271 = n5449 & ~n44270 ;
  assign n44272 = ~n44269 & n44271 ;
  assign n44273 = ~n531 & n11389 ;
  assign n44274 = n35622 ^ n19860 ^ n17948 ;
  assign n44275 = n29217 & n40806 ;
  assign n44276 = ~n947 & n44275 ;
  assign n44277 = n2692 ^ n2481 ^ 1'b0 ;
  assign n44278 = n6485 & ~n44277 ;
  assign n44279 = n29275 ^ n14604 ^ 1'b0 ;
  assign n44280 = n2883 | n44279 ;
  assign n44281 = n39952 & ~n44280 ;
  assign n44282 = n10292 & n18183 ;
  assign n44283 = ~n8886 & n44282 ;
  assign n44284 = n1574 | n8113 ;
  assign n44285 = ( n17589 & ~n41727 ) | ( n17589 & n44284 ) | ( ~n41727 & n44284 ) ;
  assign n44286 = n36568 | n39829 ;
  assign n44287 = n23981 ^ n8159 ^ n4643 ;
  assign n44288 = n44287 ^ n21232 ^ 1'b0 ;
  assign n44289 = n17684 & n44288 ;
  assign n44290 = n44289 ^ n5367 ^ n4152 ;
  assign n44291 = ~n5081 & n16711 ;
  assign n44292 = n13246 & n44291 ;
  assign n44293 = ~n15865 & n17687 ;
  assign n44294 = ~n10309 & n19710 ;
  assign n44295 = n44293 & n44294 ;
  assign n44296 = n43314 ^ n26435 ^ 1'b0 ;
  assign n44297 = n20126 ^ n13861 ^ n3360 ;
  assign n44298 = n7905 & ~n22351 ;
  assign n44299 = ~n14941 & n44298 ;
  assign n44300 = ~n11645 & n44299 ;
  assign n44301 = ( ~n11092 & n44297 ) | ( ~n11092 & n44300 ) | ( n44297 & n44300 ) ;
  assign n44302 = n289 & ~n14427 ;
  assign n44303 = n44302 ^ n20761 ^ 1'b0 ;
  assign n44304 = n44303 ^ n4867 ^ n4703 ;
  assign n44305 = n2723 & n8356 ;
  assign n44306 = ~n26640 & n44305 ;
  assign n44307 = ( n34867 & n37682 ) | ( n34867 & ~n41156 ) | ( n37682 & ~n41156 ) ;
  assign n44308 = n44307 ^ n11483 ^ 1'b0 ;
  assign n44309 = n8527 & n44308 ;
  assign n44310 = ( n6757 & n7481 ) | ( n6757 & ~n17109 ) | ( n7481 & ~n17109 ) ;
  assign n44311 = ~n17714 & n44310 ;
  assign n44312 = n17873 & ~n29047 ;
  assign n44313 = ~n26461 & n44312 ;
  assign n44314 = ~n18634 & n21385 ;
  assign n44315 = n20038 ^ n17392 ^ n14422 ;
  assign n44320 = n20781 ^ n16986 ^ 1'b0 ;
  assign n44316 = ~n4832 & n25578 ;
  assign n44317 = ~n333 & n44316 ;
  assign n44318 = ~n4236 & n44317 ;
  assign n44319 = n44318 ^ n32666 ^ n6884 ;
  assign n44321 = n44320 ^ n44319 ^ n32718 ;
  assign n44322 = n37983 ^ n30349 ^ 1'b0 ;
  assign n44323 = n26702 & n44322 ;
  assign n44324 = n10066 | n15608 ;
  assign n44325 = n1366 & ~n44324 ;
  assign n44326 = n17780 | n19029 ;
  assign n44327 = n14615 | n44326 ;
  assign n44330 = n10479 & ~n42219 ;
  assign n44328 = n15322 & ~n34350 ;
  assign n44329 = ~n2963 & n44328 ;
  assign n44331 = n44330 ^ n44329 ^ 1'b0 ;
  assign n44332 = n44331 ^ n9352 ^ 1'b0 ;
  assign n44333 = n34313 ^ n33443 ^ n15693 ;
  assign n44334 = ( ~n2376 & n9201 ) | ( ~n2376 & n22976 ) | ( n9201 & n22976 ) ;
  assign n44335 = n35682 ^ n1509 ^ 1'b0 ;
  assign n44336 = n18492 & ~n39113 ;
  assign n44337 = n10387 & ~n14009 ;
  assign n44338 = n44337 ^ n597 ^ 1'b0 ;
  assign n44339 = n44338 ^ n26053 ^ 1'b0 ;
  assign n44340 = n15387 & n44339 ;
  assign n44341 = ( n11812 & n22016 ) | ( n11812 & n24559 ) | ( n22016 & n24559 ) ;
  assign n44342 = n17373 & n44341 ;
  assign n44343 = n44342 ^ n17752 ^ 1'b0 ;
  assign n44344 = n44343 ^ n13826 ^ 1'b0 ;
  assign n44347 = ~n835 & n41716 ;
  assign n44345 = n30422 ^ n29193 ^ 1'b0 ;
  assign n44346 = n6998 & ~n44345 ;
  assign n44348 = n44347 ^ n44346 ^ 1'b0 ;
  assign n44349 = n34102 ^ n22090 ^ 1'b0 ;
  assign n44350 = n10236 & ~n44349 ;
  assign n44351 = n44350 ^ n25250 ^ n6881 ;
  assign n44352 = n31685 & ~n40819 ;
  assign n44353 = n16647 ^ n5984 ^ 1'b0 ;
  assign n44354 = n5947 & ~n44353 ;
  assign n44355 = ( n22962 & n44352 ) | ( n22962 & n44354 ) | ( n44352 & n44354 ) ;
  assign n44356 = ~n14356 & n23917 ;
  assign n44357 = n44356 ^ n38207 ^ 1'b0 ;
  assign n44358 = n44357 ^ n20841 ^ n10236 ;
  assign n44359 = ( n9023 & n36722 ) | ( n9023 & n44358 ) | ( n36722 & n44358 ) ;
  assign n44360 = n7137 ^ n6917 ^ 1'b0 ;
  assign n44361 = n26689 & n44360 ;
  assign n44362 = n1943 | n34376 ;
  assign n44363 = n33651 | n44362 ;
  assign n44364 = n4975 | n36600 ;
  assign n44365 = n28484 ^ n17514 ^ 1'b0 ;
  assign n44366 = x121 & n44365 ;
  assign n44367 = n31287 & n44366 ;
  assign n44368 = n44367 ^ n15096 ^ 1'b0 ;
  assign n44369 = ( x187 & n13574 ) | ( x187 & n44368 ) | ( n13574 & n44368 ) ;
  assign n44370 = n12517 ^ n11326 ^ n7362 ;
  assign n44371 = n43933 ^ n12739 ^ 1'b0 ;
  assign n44372 = n31646 ^ n26130 ^ 1'b0 ;
  assign n44373 = ~n11990 & n33744 ;
  assign n44374 = n8630 & n44373 ;
  assign n44375 = n42530 & n44374 ;
  assign n44376 = n32202 ^ n31446 ^ 1'b0 ;
  assign n44377 = n8899 & n44376 ;
  assign n44378 = n6507 | n41785 ;
  assign n44379 = n4976 & ~n9689 ;
  assign n44380 = n39829 ^ n36481 ^ 1'b0 ;
  assign n44381 = ~n3642 & n44380 ;
  assign n44382 = n40115 ^ n37502 ^ n31746 ;
  assign n44383 = n9267 ^ n6276 ^ 1'b0 ;
  assign n44384 = n982 | n10436 ;
  assign n44385 = n44384 ^ n10071 ^ 1'b0 ;
  assign n44386 = n44385 ^ n39846 ^ 1'b0 ;
  assign n44387 = n24498 ^ n12011 ^ n10151 ;
  assign n44388 = n44387 ^ n27547 ^ 1'b0 ;
  assign n44389 = ~n1851 & n12907 ;
  assign n44390 = ~n908 & n11608 ;
  assign n44391 = n44390 ^ n25014 ^ 1'b0 ;
  assign n44392 = n5175 & ~n12639 ;
  assign n44393 = n21377 ^ n597 ^ 1'b0 ;
  assign n44394 = n13907 | n44393 ;
  assign n44395 = n44394 ^ n43728 ^ n24264 ;
  assign n44396 = n11335 & n32010 ;
  assign n44397 = n44396 ^ n40677 ^ n35831 ;
  assign n44398 = ( n811 & n16868 ) | ( n811 & n40657 ) | ( n16868 & n40657 ) ;
  assign n44399 = n8781 & n19235 ;
  assign n44400 = n911 & ~n18009 ;
  assign n44401 = n38124 & n44400 ;
  assign n44402 = n44401 ^ n18622 ^ 1'b0 ;
  assign n44403 = n29744 ^ n26244 ^ 1'b0 ;
  assign n44404 = ~n44402 & n44403 ;
  assign n44405 = n44404 ^ n11087 ^ 1'b0 ;
  assign n44406 = ~n4508 & n36767 ;
  assign n44407 = ~n11479 & n44406 ;
  assign n44408 = n4468 ^ n2573 ^ 1'b0 ;
  assign n44409 = n43753 | n44408 ;
  assign n44411 = n12399 & n26594 ;
  assign n44410 = n22486 & n23810 ;
  assign n44412 = n44411 ^ n44410 ^ 1'b0 ;
  assign n44413 = n39284 ^ n22088 ^ n13384 ;
  assign n44414 = n6704 & ~n26806 ;
  assign n44415 = n14837 | n44414 ;
  assign n44416 = n44415 ^ n28492 ^ 1'b0 ;
  assign n44417 = ( ~n559 & n28280 ) | ( ~n559 & n44416 ) | ( n28280 & n44416 ) ;
  assign n44418 = n8683 & ~n12989 ;
  assign n44419 = n36604 ^ n27560 ^ 1'b0 ;
  assign n44420 = n29862 & n44419 ;
  assign n44421 = n9483 & ~n17573 ;
  assign n44422 = n44421 ^ n26829 ^ 1'b0 ;
  assign n44423 = n31775 ^ n24947 ^ n12145 ;
  assign n44424 = n44423 ^ n8271 ^ 1'b0 ;
  assign n44425 = n20161 & n44424 ;
  assign n44426 = n2916 | n41959 ;
  assign n44427 = x254 & ~n3732 ;
  assign n44428 = n44427 ^ n10679 ^ 1'b0 ;
  assign n44429 = n44428 ^ n10511 ^ 1'b0 ;
  assign n44430 = n4286 ^ n606 ^ x187 ;
  assign n44431 = ~n1495 & n18340 ;
  assign n44432 = n44431 ^ n38902 ^ 1'b0 ;
  assign n44433 = n44432 ^ n32502 ^ n28886 ;
  assign n44434 = n37604 ^ n21977 ^ 1'b0 ;
  assign n44435 = n30382 ^ n17426 ^ 1'b0 ;
  assign n44436 = n5807 & n5865 ;
  assign n44437 = n24490 | n25099 ;
  assign n44438 = n18514 & ~n44437 ;
  assign n44439 = ( n9179 & ~n12625 ) | ( n9179 & n44438 ) | ( ~n12625 & n44438 ) ;
  assign n44440 = ( n4410 & n4521 ) | ( n4410 & n25210 ) | ( n4521 & n25210 ) ;
  assign n44441 = n44440 ^ n33097 ^ n24818 ;
  assign n44442 = n20665 ^ n7897 ^ n4957 ;
  assign n44443 = n18317 | n44442 ;
  assign n44444 = n16642 & ~n44443 ;
  assign n44445 = n31827 ^ n26797 ^ 1'b0 ;
  assign n44446 = ~n37008 & n44445 ;
  assign n44447 = n12723 | n44446 ;
  assign n44448 = ~n9230 & n9687 ;
  assign n44449 = n10532 & n44448 ;
  assign n44450 = n12355 | n44449 ;
  assign n44451 = n6172 | n22604 ;
  assign n44452 = n44451 ^ n21607 ^ 1'b0 ;
  assign n44453 = n44450 & n44452 ;
  assign n44454 = n15551 ^ n10076 ^ 1'b0 ;
  assign n44455 = n32533 ^ n2057 ^ 1'b0 ;
  assign n44456 = n31061 ^ n9870 ^ 1'b0 ;
  assign n44457 = n3422 | n44456 ;
  assign n44458 = n44457 ^ n32237 ^ 1'b0 ;
  assign n44459 = ( n5780 & n9078 ) | ( n5780 & ~n24017 ) | ( n9078 & ~n24017 ) ;
  assign n44460 = n25099 ^ n6888 ^ 1'b0 ;
  assign n44461 = n35200 | n44460 ;
  assign n44462 = n44461 ^ n31927 ^ 1'b0 ;
  assign n44463 = n12712 ^ n6622 ^ 1'b0 ;
  assign n44464 = n24531 | n44463 ;
  assign n44465 = ( n9103 & n25061 ) | ( n9103 & ~n44464 ) | ( n25061 & ~n44464 ) ;
  assign n44466 = n793 | n1188 ;
  assign n44467 = n44466 ^ n36888 ^ 1'b0 ;
  assign n44468 = n17956 | n33032 ;
  assign n44469 = n16766 & ~n31317 ;
  assign n44470 = n6871 & n43250 ;
  assign n44471 = n13441 & n19134 ;
  assign n44472 = n44471 ^ n37661 ^ 1'b0 ;
  assign n44473 = n25199 & n32875 ;
  assign n44474 = ( n28934 & ~n33560 ) | ( n28934 & n35071 ) | ( ~n33560 & n35071 ) ;
  assign n44475 = ( n33788 & ~n44473 ) | ( n33788 & n44474 ) | ( ~n44473 & n44474 ) ;
  assign n44476 = n16725 | n27600 ;
  assign n44477 = n44476 ^ n11407 ^ 1'b0 ;
  assign n44478 = n26358 ^ n11163 ^ 1'b0 ;
  assign n44479 = n11747 | n25686 ;
  assign n44480 = n981 | n44479 ;
  assign n44482 = ~n5974 & n6382 ;
  assign n44483 = ~n7196 & n44482 ;
  assign n44484 = n11338 & n11847 ;
  assign n44485 = n44483 & n44484 ;
  assign n44481 = ~n1213 & n10573 ;
  assign n44486 = n44485 ^ n44481 ^ 1'b0 ;
  assign n44487 = n377 | n31209 ;
  assign n44488 = n44486 | n44487 ;
  assign n44489 = n30247 ^ n25931 ^ 1'b0 ;
  assign n44490 = n16002 & n44489 ;
  assign n44491 = ( x65 & ~n3626 ) | ( x65 & n21201 ) | ( ~n3626 & n21201 ) ;
  assign n44492 = n10262 & ~n14057 ;
  assign n44493 = n21055 & n21549 ;
  assign n44494 = ~n20784 & n44493 ;
  assign n44495 = ~n44492 & n44494 ;
  assign n44496 = n7174 | n29483 ;
  assign n44497 = n10965 & ~n44496 ;
  assign n44498 = ( n20952 & n43538 ) | ( n20952 & ~n44497 ) | ( n43538 & ~n44497 ) ;
  assign n44499 = n27295 ^ n21740 ^ n18360 ;
  assign n44500 = x46 & n18857 ;
  assign n44501 = n44500 ^ n33841 ^ 1'b0 ;
  assign n44502 = ( n11885 & ~n44499 ) | ( n11885 & n44501 ) | ( ~n44499 & n44501 ) ;
  assign n44503 = n37819 & ~n44502 ;
  assign n44504 = n44503 ^ n6977 ^ 1'b0 ;
  assign n44505 = n15290 & n22163 ;
  assign n44506 = n20864 ^ n3480 ^ 1'b0 ;
  assign n44507 = ~n44505 & n44506 ;
  assign n44508 = n44507 ^ n8319 ^ 1'b0 ;
  assign n44509 = n4119 & ~n21875 ;
  assign n44510 = n13928 & n44509 ;
  assign n44511 = n6268 | n44510 ;
  assign n44512 = n44511 ^ n13643 ^ 1'b0 ;
  assign n44513 = n44512 ^ n19125 ^ 1'b0 ;
  assign n44514 = n29577 & ~n44513 ;
  assign n44515 = ~n11564 & n38454 ;
  assign n44516 = ~n5788 & n6700 ;
  assign n44517 = n22160 ^ n7053 ^ n397 ;
  assign n44518 = ( n5850 & ~n26888 ) | ( n5850 & n42081 ) | ( ~n26888 & n42081 ) ;
  assign n44520 = n1897 | n9461 ;
  assign n44519 = ( n7310 & n8762 ) | ( n7310 & ~n33041 ) | ( n8762 & ~n33041 ) ;
  assign n44521 = n44520 ^ n44519 ^ n8438 ;
  assign n44522 = n15307 ^ n1779 ^ 1'b0 ;
  assign n44523 = n12780 & n26606 ;
  assign n44524 = n12142 & n44523 ;
  assign n44525 = n7718 ^ n5064 ^ 1'b0 ;
  assign n44526 = n597 & n44525 ;
  assign n44527 = n26092 | n44526 ;
  assign n44529 = ~n5277 & n9408 ;
  assign n44528 = n16972 | n19303 ;
  assign n44530 = n44529 ^ n44528 ^ 1'b0 ;
  assign n44531 = n15091 | n44530 ;
  assign n44532 = ~n3879 & n29851 ;
  assign n44533 = n5170 & n44532 ;
  assign n44534 = n6216 & ~n12019 ;
  assign n44535 = n44533 & n44534 ;
  assign n44536 = n25429 | n44535 ;
  assign n44537 = n1365 & n3843 ;
  assign n44538 = n44537 ^ n35351 ^ 1'b0 ;
  assign n44539 = ( ~n9106 & n22354 ) | ( ~n9106 & n24450 ) | ( n22354 & n24450 ) ;
  assign n44542 = n28680 ^ n7764 ^ n1885 ;
  assign n44540 = n19166 & ~n20998 ;
  assign n44541 = n44540 ^ n3540 ^ 1'b0 ;
  assign n44543 = n44542 ^ n44541 ^ n13527 ;
  assign n44544 = n16004 & ~n18222 ;
  assign n44545 = n3283 & ~n28015 ;
  assign n44546 = n31230 ^ n14540 ^ 1'b0 ;
  assign n44547 = n15996 ^ n4007 ^ 1'b0 ;
  assign n44548 = n17602 & ~n44547 ;
  assign n44549 = n9512 & n44548 ;
  assign n44550 = n30767 & n44549 ;
  assign n44551 = n6967 ^ n2475 ^ 1'b0 ;
  assign n44552 = ~n21777 & n44551 ;
  assign n44553 = n4762 | n44552 ;
  assign n44554 = n11960 & ~n12145 ;
  assign n44555 = x60 | n29395 ;
  assign n44556 = n44555 ^ n6440 ^ 1'b0 ;
  assign n44557 = n9694 & ~n24975 ;
  assign n44558 = n16655 ^ n4183 ^ 1'b0 ;
  assign n44559 = ~n2519 & n14366 ;
  assign n44560 = ~n12678 & n18523 ;
  assign n44561 = n44560 ^ n25737 ^ 1'b0 ;
  assign n44562 = n35971 ^ n32176 ^ 1'b0 ;
  assign n44563 = ~n6867 & n28435 ;
  assign n44564 = n44563 ^ n31913 ^ 1'b0 ;
  assign n44566 = n30695 ^ n15629 ^ 1'b0 ;
  assign n44567 = n21508 | n44566 ;
  assign n44565 = n6726 & n25391 ;
  assign n44568 = n44567 ^ n44565 ^ 1'b0 ;
  assign n44569 = ( n1811 & n8721 ) | ( n1811 & ~n29483 ) | ( n8721 & ~n29483 ) ;
  assign n44570 = n14677 & ~n43711 ;
  assign n44571 = n31557 & n44570 ;
  assign n44572 = ~n23760 & n26482 ;
  assign n44573 = n616 & n44572 ;
  assign n44574 = ~n31169 & n38062 ;
  assign n44575 = n19799 & n44574 ;
  assign n44576 = n44575 ^ n35111 ^ 1'b0 ;
  assign n44577 = ( n529 & ~n14273 ) | ( n529 & n18465 ) | ( ~n14273 & n18465 ) ;
  assign n44578 = n36053 ^ n22381 ^ 1'b0 ;
  assign n44579 = n44577 | n44578 ;
  assign n44580 = ~n5070 & n20230 ;
  assign n44581 = ~n6953 & n44580 ;
  assign n44583 = n20357 & ~n21853 ;
  assign n44584 = n44583 ^ n13392 ^ 1'b0 ;
  assign n44582 = n2804 & ~n5243 ;
  assign n44585 = n44584 ^ n44582 ^ 1'b0 ;
  assign n44586 = n40366 ^ n18560 ^ n4729 ;
  assign n44587 = n30928 ^ n16235 ^ 1'b0 ;
  assign n44588 = n20531 ^ n6002 ^ 1'b0 ;
  assign n44589 = n3586 & ~n6309 ;
  assign n44590 = n32647 & n44589 ;
  assign n44591 = ~n28573 & n37450 ;
  assign n44592 = n33417 & n44591 ;
  assign n44593 = n24310 ^ n5626 ^ 1'b0 ;
  assign n44594 = ~n2274 & n4397 ;
  assign n44595 = ( n8589 & ~n28509 ) | ( n8589 & n44594 ) | ( ~n28509 & n44594 ) ;
  assign n44596 = n3988 ^ n3066 ^ 1'b0 ;
  assign n44597 = ~n22019 & n44596 ;
  assign n44598 = n44597 ^ n38400 ^ n35118 ;
  assign n44599 = n4405 & ~n19132 ;
  assign n44600 = ~n32484 & n44599 ;
  assign n44604 = x50 | n11302 ;
  assign n44601 = n5843 & ~n10928 ;
  assign n44602 = n44601 ^ n3785 ^ 1'b0 ;
  assign n44603 = ~n23477 & n44602 ;
  assign n44605 = n44604 ^ n44603 ^ 1'b0 ;
  assign n44606 = n13765 ^ n1270 ^ n397 ;
  assign n44607 = n16466 ^ n12343 ^ n11176 ;
  assign n44608 = ~x159 & n4552 ;
  assign n44609 = n44608 ^ n25093 ^ 1'b0 ;
  assign n44611 = n3384 ^ x237 ^ 1'b0 ;
  assign n44610 = n17794 & ~n33012 ;
  assign n44612 = n44611 ^ n44610 ^ 1'b0 ;
  assign n44613 = n24311 ^ n22064 ^ 1'b0 ;
  assign n44614 = n2142 & ~n44613 ;
  assign n44617 = n16168 ^ n9371 ^ 1'b0 ;
  assign n44615 = n29344 ^ n4009 ^ 1'b0 ;
  assign n44616 = n25129 | n44615 ;
  assign n44618 = n44617 ^ n44616 ^ 1'b0 ;
  assign n44619 = n36933 ^ n19820 ^ 1'b0 ;
  assign n44620 = n44618 & n44619 ;
  assign n44621 = n24855 ^ n10187 ^ n5211 ;
  assign n44622 = n24044 | n44621 ;
  assign n44623 = n44622 ^ n3520 ^ 1'b0 ;
  assign n44624 = n33617 ^ n5491 ^ 1'b0 ;
  assign n44625 = n1758 & ~n20946 ;
  assign n44626 = n44625 ^ n10509 ^ 1'b0 ;
  assign n44627 = ( n3912 & n9208 ) | ( n3912 & n29507 ) | ( n9208 & n29507 ) ;
  assign n44628 = n4966 & n17694 ;
  assign n44629 = n44628 ^ n32680 ^ 1'b0 ;
  assign n44630 = ~n6249 & n44629 ;
  assign n44631 = n41875 ^ n8825 ^ 1'b0 ;
  assign n44632 = n4950 & ~n33106 ;
  assign n44633 = n44632 ^ n24537 ^ 1'b0 ;
  assign n44634 = n5121 & ~n23028 ;
  assign n44635 = n6912 & n44634 ;
  assign n44636 = n8517 & n34607 ;
  assign n44637 = n10221 & n11803 ;
  assign n44638 = ~n7564 & n11854 ;
  assign n44639 = n44638 ^ n21073 ^ n6859 ;
  assign n44640 = ( n1453 & n21359 ) | ( n1453 & ~n44639 ) | ( n21359 & ~n44639 ) ;
  assign n44641 = n5896 | n7786 ;
  assign n44642 = ~n25820 & n44641 ;
  assign n44643 = n39727 ^ n4243 ^ 1'b0 ;
  assign n44644 = n29984 | n44643 ;
  assign n44645 = n17350 & ~n39953 ;
  assign n44646 = n2299 & ~n9117 ;
  assign n44647 = n44646 ^ n2419 ^ 1'b0 ;
  assign n44648 = n12547 & n44647 ;
  assign n44649 = n44648 ^ n19975 ^ 1'b0 ;
  assign n44650 = n16338 ^ n12285 ^ n9810 ;
  assign n44651 = n44650 ^ n36443 ^ n35221 ;
  assign n44655 = n36130 ^ n30813 ^ 1'b0 ;
  assign n44656 = n9529 & ~n44655 ;
  assign n44652 = n12762 | n27034 ;
  assign n44653 = n10658 & ~n44652 ;
  assign n44654 = n44653 ^ n25277 ^ n9773 ;
  assign n44657 = n44656 ^ n44654 ^ 1'b0 ;
  assign n44658 = n1347 | n22749 ;
  assign n44659 = n8810 & ~n44658 ;
  assign n44660 = n44659 ^ n26297 ^ n6608 ;
  assign n44662 = n6661 ^ n4340 ^ 1'b0 ;
  assign n44663 = n29207 & n44662 ;
  assign n44661 = n16719 & ~n26631 ;
  assign n44664 = n44663 ^ n44661 ^ 1'b0 ;
  assign n44665 = ~n13542 & n14454 ;
  assign n44666 = n4037 & ~n18485 ;
  assign n44667 = n44666 ^ n20317 ^ 1'b0 ;
  assign n44668 = n6868 | n23784 ;
  assign n44669 = n4027 & ~n44668 ;
  assign n44671 = ( n1564 & ~n15018 ) | ( n1564 & n31187 ) | ( ~n15018 & n31187 ) ;
  assign n44670 = n8945 & ~n23883 ;
  assign n44672 = n44671 ^ n44670 ^ 1'b0 ;
  assign n44673 = n26489 ^ n5726 ^ 1'b0 ;
  assign n44674 = n1922 & n44673 ;
  assign n44675 = n17631 ^ n4135 ^ n315 ;
  assign n44676 = n44675 ^ n20508 ^ n1988 ;
  assign n44677 = n38310 ^ n20575 ^ 1'b0 ;
  assign n44678 = n36828 & n44677 ;
  assign n44679 = n44678 ^ n18260 ^ n10612 ;
  assign n44680 = n5536 & ~n23209 ;
  assign n44681 = n44680 ^ n13391 ^ 1'b0 ;
  assign n44682 = n44681 ^ n21010 ^ 1'b0 ;
  assign n44683 = n44682 ^ n25111 ^ 1'b0 ;
  assign n44684 = ( ~n482 & n3872 ) | ( ~n482 & n13243 ) | ( n3872 & n13243 ) ;
  assign n44685 = n23603 | n44684 ;
  assign n44686 = n44685 ^ n38786 ^ 1'b0 ;
  assign n44687 = n10949 & ~n38834 ;
  assign n44688 = n36481 ^ n14340 ^ 1'b0 ;
  assign n44689 = ~n26438 & n44688 ;
  assign n44690 = n44689 ^ n21709 ^ n14697 ;
  assign n44691 = n10421 & ~n13183 ;
  assign n44692 = ( n3709 & n8461 ) | ( n3709 & ~n25515 ) | ( n8461 & ~n25515 ) ;
  assign n44693 = n28616 | n31404 ;
  assign n44695 = n13921 ^ n7637 ^ n2225 ;
  assign n44694 = n10120 & ~n29649 ;
  assign n44696 = n44695 ^ n44694 ^ 1'b0 ;
  assign n44697 = n7947 | n30845 ;
  assign n44698 = n20809 & ~n44697 ;
  assign n44699 = n10288 | n44698 ;
  assign n44700 = n15903 & ~n44699 ;
  assign n44701 = n9860 & n18953 ;
  assign n44702 = n44701 ^ n6119 ^ 1'b0 ;
  assign n44703 = ~n34382 & n42181 ;
  assign n44705 = ~n10183 & n21664 ;
  assign n44704 = n18455 & ~n26671 ;
  assign n44706 = n44705 ^ n44704 ^ 1'b0 ;
  assign n44707 = n19772 ^ n1093 ^ 1'b0 ;
  assign n44708 = ( n2276 & n36511 ) | ( n2276 & ~n44707 ) | ( n36511 & ~n44707 ) ;
  assign n44709 = ~n25669 & n43459 ;
  assign n44710 = ~x170 & n7824 ;
  assign n44711 = n6908 & ~n44710 ;
  assign n44712 = ~n17816 & n31021 ;
  assign n44713 = n18451 | n36138 ;
  assign n44714 = n44712 & ~n44713 ;
  assign n44716 = ( n4232 & ~n19722 ) | ( n4232 & n25820 ) | ( ~n19722 & n25820 ) ;
  assign n44715 = n21170 | n25125 ;
  assign n44717 = n44716 ^ n44715 ^ 1'b0 ;
  assign n44718 = n23915 ^ n15707 ^ 1'b0 ;
  assign n44719 = ~n29324 & n44718 ;
  assign n44720 = n7664 & n13596 ;
  assign n44721 = n21981 & ~n44720 ;
  assign n44722 = ~n5255 & n29229 ;
  assign n44723 = ( n413 & ~n29914 ) | ( n413 & n43804 ) | ( ~n29914 & n43804 ) ;
  assign n44724 = n6191 & ~n40440 ;
  assign n44725 = ( x4 & n24546 ) | ( x4 & n44724 ) | ( n24546 & n44724 ) ;
  assign n44726 = n16427 & ~n40344 ;
  assign n44727 = ~x133 & n44726 ;
  assign n44728 = ~n6555 & n11873 ;
  assign n44729 = n3330 | n25552 ;
  assign n44732 = n22195 ^ n19212 ^ 1'b0 ;
  assign n44733 = n7584 & ~n44732 ;
  assign n44734 = ( n5112 & n38362 ) | ( n5112 & ~n44733 ) | ( n38362 & ~n44733 ) ;
  assign n44730 = n31342 ^ n12727 ^ 1'b0 ;
  assign n44731 = n27838 & n44730 ;
  assign n44735 = n44734 ^ n44731 ^ 1'b0 ;
  assign n44736 = n1526 | n9849 ;
  assign n44737 = n5359 | n44736 ;
  assign n44738 = n11196 | n22645 ;
  assign n44739 = ~n17143 & n25965 ;
  assign n44740 = n44738 & n44739 ;
  assign n44741 = n44740 ^ n1230 ^ 1'b0 ;
  assign n44742 = ~n2426 & n42621 ;
  assign n44743 = n31475 & n40475 ;
  assign n44744 = n719 | n3986 ;
  assign n44745 = n44744 ^ n2054 ^ 1'b0 ;
  assign n44746 = ~n5330 & n9524 ;
  assign n44747 = ~n12548 & n44746 ;
  assign n44748 = n1455 & ~n7372 ;
  assign n44749 = n5415 & ~n11948 ;
  assign n44750 = n44748 & n44749 ;
  assign n44751 = ( n44745 & n44747 ) | ( n44745 & ~n44750 ) | ( n44747 & ~n44750 ) ;
  assign n44752 = n14412 & n25576 ;
  assign n44753 = n1875 & ~n12329 ;
  assign n44754 = n44752 & n44753 ;
  assign n44755 = n2553 & n9166 ;
  assign n44756 = n791 ^ n585 ^ 1'b0 ;
  assign n44757 = n15930 & n44756 ;
  assign n44758 = n31259 & ~n34492 ;
  assign n44759 = n2981 | n44758 ;
  assign n44762 = ( n8411 & n17235 ) | ( n8411 & ~n21993 ) | ( n17235 & ~n21993 ) ;
  assign n44760 = n15113 & ~n19616 ;
  assign n44761 = n29395 & n44760 ;
  assign n44763 = n44762 ^ n44761 ^ n14962 ;
  assign n44764 = n35410 ^ n16133 ^ n11887 ;
  assign n44765 = n44764 ^ n21044 ^ 1'b0 ;
  assign n44766 = n44763 | n44765 ;
  assign n44767 = n2824 | n24865 ;
  assign n44768 = n1499 & n20035 ;
  assign n44769 = ~n24450 & n44768 ;
  assign n44770 = n44769 ^ n21128 ^ 1'b0 ;
  assign n44771 = n30192 ^ n22059 ^ x82 ;
  assign n44772 = ~n2959 & n7443 ;
  assign n44773 = n20759 & ~n33312 ;
  assign n44774 = ~n10230 & n44773 ;
  assign n44775 = n10071 & n38067 ;
  assign n44776 = n33839 ^ n15246 ^ 1'b0 ;
  assign n44777 = n12713 & n44776 ;
  assign n44778 = n44777 ^ n24284 ^ 1'b0 ;
  assign n44779 = n4552 & ~n44778 ;
  assign n44780 = n40635 ^ n19303 ^ 1'b0 ;
  assign n44781 = ~n24708 & n44780 ;
  assign n44782 = ~n4312 & n44781 ;
  assign n44783 = n33978 ^ n30886 ^ 1'b0 ;
  assign n44784 = ( n2462 & n7468 ) | ( n2462 & ~n11694 ) | ( n7468 & ~n11694 ) ;
  assign n44785 = n15664 & ~n44784 ;
  assign n44786 = ~n6352 & n44785 ;
  assign n44787 = n44786 ^ n13406 ^ 1'b0 ;
  assign n44788 = ~n10827 & n18060 ;
  assign n44789 = ~n18060 & n44788 ;
  assign n44790 = n6824 & ~n32519 ;
  assign n44791 = ( ~n19210 & n44789 ) | ( ~n19210 & n44790 ) | ( n44789 & n44790 ) ;
  assign n44792 = n5669 | n25936 ;
  assign n44793 = ( n5569 & n13757 ) | ( n5569 & ~n26664 ) | ( n13757 & ~n26664 ) ;
  assign n44794 = n42469 | n44793 ;
  assign n44795 = n12722 & ~n44794 ;
  assign n44796 = ( ~n5855 & n30051 ) | ( ~n5855 & n44795 ) | ( n30051 & n44795 ) ;
  assign n44797 = n44161 ^ n6993 ^ 1'b0 ;
  assign n44798 = ~n44796 & n44797 ;
  assign n44799 = n18171 & n22188 ;
  assign n44800 = ( n40149 & ~n44050 ) | ( n40149 & n44799 ) | ( ~n44050 & n44799 ) ;
  assign n44801 = n26405 ^ n11246 ^ 1'b0 ;
  assign n44802 = n8038 | n44801 ;
  assign n44803 = n44802 ^ n5029 ^ n3570 ;
  assign n44804 = n29983 ^ n29472 ^ n706 ;
  assign n44805 = n7453 & n21827 ;
  assign n44806 = n44804 & n44805 ;
  assign n44807 = ( n21210 & n33575 ) | ( n21210 & n44806 ) | ( n33575 & n44806 ) ;
  assign n44808 = x241 ^ x152 ^ 1'b0 ;
  assign n44809 = n16184 | n44808 ;
  assign n44810 = n44809 ^ n44538 ^ 1'b0 ;
  assign n44811 = n14382 ^ n5556 ^ 1'b0 ;
  assign n44812 = n28739 & n44811 ;
  assign n44813 = n37062 ^ n1024 ^ 1'b0 ;
  assign n44814 = n633 & n6063 ;
  assign n44815 = n7740 & n44814 ;
  assign n44816 = n21929 & ~n44815 ;
  assign n44817 = n9112 & n44816 ;
  assign n44818 = n44813 & n44817 ;
  assign n44819 = ( n18964 & n22795 ) | ( n18964 & ~n34262 ) | ( n22795 & ~n34262 ) ;
  assign n44820 = ~n6648 & n44819 ;
  assign n44821 = n34955 ^ n2652 ^ 1'b0 ;
  assign n44822 = n9651 & n44821 ;
  assign n44823 = n44822 ^ n27427 ^ 1'b0 ;
  assign n44824 = n39482 ^ n9144 ^ n4703 ;
  assign n44825 = n7155 | n39916 ;
  assign n44826 = n11284 & ~n24071 ;
  assign n44827 = n44826 ^ n32445 ^ n3474 ;
  assign n44828 = n36855 ^ n17684 ^ n8490 ;
  assign n44829 = n36263 ^ n451 ^ 1'b0 ;
  assign n44830 = n3803 & n44829 ;
  assign n44831 = n2991 | n15093 ;
  assign n44832 = n44831 ^ n22671 ^ 1'b0 ;
  assign n44833 = ~n35582 & n36373 ;
  assign n44834 = n43607 & n44833 ;
  assign n44835 = ~n704 & n30076 ;
  assign n44836 = n44835 ^ n7068 ^ 1'b0 ;
  assign n44837 = n21398 ^ n15012 ^ 1'b0 ;
  assign n44838 = ~n23626 & n44837 ;
  assign n44839 = n13754 & n42863 ;
  assign n44840 = n44839 ^ n905 ^ 1'b0 ;
  assign n44841 = n23637 ^ n9962 ^ 1'b0 ;
  assign n44842 = ( n2158 & n2368 ) | ( n2158 & n31187 ) | ( n2368 & n31187 ) ;
  assign n44843 = ~n10332 & n44842 ;
  assign n44844 = ( n30520 & ~n36829 ) | ( n30520 & n44843 ) | ( ~n36829 & n44843 ) ;
  assign n44845 = n29179 ^ n4853 ^ n575 ;
  assign n44846 = n44845 ^ n11298 ^ 1'b0 ;
  assign n44847 = n3129 & ~n8567 ;
  assign n44848 = n26178 & n44847 ;
  assign n44849 = ~n5812 & n44848 ;
  assign n44850 = n7095 ^ n1489 ^ 1'b0 ;
  assign n44851 = n44850 ^ n9529 ^ n4419 ;
  assign n44852 = ~n24608 & n44851 ;
  assign n44853 = n15491 ^ n7527 ^ 1'b0 ;
  assign n44854 = n14983 ^ n6700 ^ 1'b0 ;
  assign n44855 = n44853 | n44854 ;
  assign n44856 = ~n6064 & n13380 ;
  assign n44857 = ~n5354 & n44856 ;
  assign n44858 = ~n471 & n44857 ;
  assign n44859 = n37833 & n44858 ;
  assign n44860 = n7723 ^ n7475 ^ 1'b0 ;
  assign n44861 = ~n44859 & n44860 ;
  assign n44862 = n37192 ^ n17523 ^ 1'b0 ;
  assign n44863 = n11157 ^ n1387 ^ 1'b0 ;
  assign n44864 = n9311 | n37119 ;
  assign n44865 = n21165 & ~n44864 ;
  assign n44866 = n10203 | n18693 ;
  assign n44867 = n42377 ^ n23763 ^ 1'b0 ;
  assign n44868 = n13589 ^ n2868 ^ 1'b0 ;
  assign n44869 = ~n29982 & n44868 ;
  assign n44871 = n6018 ^ n5481 ^ 1'b0 ;
  assign n44872 = ~n6369 & n44871 ;
  assign n44870 = n3306 | n10525 ;
  assign n44873 = n44872 ^ n44870 ^ 1'b0 ;
  assign n44874 = n44873 ^ n27390 ^ 1'b0 ;
  assign n44875 = ( n24063 & n40052 ) | ( n24063 & ~n44874 ) | ( n40052 & ~n44874 ) ;
  assign n44876 = ~n5370 & n44875 ;
  assign n44877 = ~n44869 & n44876 ;
  assign n44879 = n24768 & n40879 ;
  assign n44880 = n44879 ^ n21067 ^ 1'b0 ;
  assign n44878 = n15107 & n44782 ;
  assign n44881 = n44880 ^ n44878 ^ 1'b0 ;
  assign n44882 = n36800 | n43537 ;
  assign n44883 = n5837 | n44882 ;
  assign n44884 = n4957 | n7799 ;
  assign n44885 = n2601 | n44884 ;
  assign n44886 = n44885 ^ n37833 ^ n8284 ;
  assign n44887 = n19475 & ~n44886 ;
  assign n44888 = ~n8634 & n44887 ;
  assign n44889 = n44888 ^ n30727 ^ 1'b0 ;
  assign n44890 = n6830 | n32610 ;
  assign n44891 = n30026 | n44890 ;
  assign n44892 = ~n1758 & n4463 ;
  assign n44893 = n44892 ^ n7726 ^ 1'b0 ;
  assign n44894 = n32329 ^ n25702 ^ 1'b0 ;
  assign n44895 = n1291 | n44894 ;
  assign n44896 = ( ~n11526 & n13081 ) | ( ~n11526 & n44895 ) | ( n13081 & n44895 ) ;
  assign n44897 = n29373 ^ n25813 ^ 1'b0 ;
  assign n44898 = n7952 ^ n1483 ^ 1'b0 ;
  assign n44899 = n5075 & n44898 ;
  assign n44900 = n42148 ^ n28734 ^ n22453 ;
  assign n44901 = n32447 | n44900 ;
  assign n44902 = n44901 ^ n8281 ^ 1'b0 ;
  assign n44903 = ~n516 & n8622 ;
  assign n44904 = n25900 & ~n44903 ;
  assign n44905 = n40953 ^ n30415 ^ 1'b0 ;
  assign n44906 = n23514 & ~n44905 ;
  assign n44907 = n7035 | n13185 ;
  assign n44908 = ~n11932 & n14422 ;
  assign n44909 = n37569 ^ n34681 ^ n31871 ;
  assign n44910 = n5562 ^ n4676 ^ n1991 ;
  assign n44911 = ~n1769 & n44910 ;
  assign n44912 = n5954 & n17954 ;
  assign n44913 = n908 & n1731 ;
  assign n44914 = n14551 ^ n8284 ^ 1'b0 ;
  assign n44915 = n6632 | n27652 ;
  assign n44916 = n10324 & ~n44915 ;
  assign n44917 = n17620 ^ n16579 ^ 1'b0 ;
  assign n44918 = ~n44916 & n44917 ;
  assign n44919 = ( n2955 & ~n17689 ) | ( n2955 & n23691 ) | ( ~n17689 & n23691 ) ;
  assign n44920 = ~n7048 & n20061 ;
  assign n44921 = ( ~n3304 & n12142 ) | ( ~n3304 & n44920 ) | ( n12142 & n44920 ) ;
  assign n44922 = n8702 ^ n4810 ^ 1'b0 ;
  assign n44923 = n2376 & n44922 ;
  assign n44926 = ( n14786 & n26347 ) | ( n14786 & n28678 ) | ( n26347 & n28678 ) ;
  assign n44924 = n14856 ^ n7584 ^ n555 ;
  assign n44925 = n3676 & n44924 ;
  assign n44927 = n44926 ^ n44925 ^ 1'b0 ;
  assign n44928 = n6723 & n20575 ;
  assign n44929 = ~n1324 & n44928 ;
  assign n44931 = ~n9324 & n40177 ;
  assign n44930 = n9493 | n15919 ;
  assign n44932 = n44931 ^ n44930 ^ 1'b0 ;
  assign n44933 = n37592 ^ n27098 ^ 1'b0 ;
  assign n44935 = n5967 | n8592 ;
  assign n44934 = n15536 | n23356 ;
  assign n44936 = n44935 ^ n44934 ^ 1'b0 ;
  assign n44937 = ( n8257 & n8773 ) | ( n8257 & ~n10631 ) | ( n8773 & ~n10631 ) ;
  assign n44938 = n44937 ^ n34034 ^ 1'b0 ;
  assign n44939 = n44936 & n44938 ;
  assign n44940 = n8632 ^ n1713 ^ 1'b0 ;
  assign n44941 = ~n14388 & n44940 ;
  assign n44942 = ~n31710 & n44941 ;
  assign n44943 = n44939 & n44942 ;
  assign n44944 = n3882 | n13899 ;
  assign n44945 = n3882 & ~n44944 ;
  assign n44946 = n44945 ^ n43319 ^ n42947 ;
  assign n44947 = n10284 ^ n5039 ^ 1'b0 ;
  assign n44948 = ~n4058 & n44947 ;
  assign n44949 = ( n33670 & ~n42881 ) | ( n33670 & n44948 ) | ( ~n42881 & n44948 ) ;
  assign n44951 = n12185 & ~n34713 ;
  assign n44952 = n44951 ^ n17094 ^ 1'b0 ;
  assign n44953 = n14793 | n44952 ;
  assign n44950 = n21584 ^ n8112 ^ 1'b0 ;
  assign n44954 = n44953 ^ n44950 ^ n44347 ;
  assign n44955 = n21777 & n31973 ;
  assign n44956 = n8630 ^ n3685 ^ 1'b0 ;
  assign n44957 = n3295 | n44956 ;
  assign n44958 = n44957 ^ n22554 ^ 1'b0 ;
  assign n44959 = n37938 | n44958 ;
  assign n44960 = ( n3615 & ~n6174 ) | ( n3615 & n10504 ) | ( ~n6174 & n10504 ) ;
  assign n44961 = n44960 ^ n34577 ^ n28340 ;
  assign n44962 = n19852 & n44961 ;
  assign n44963 = ~n2224 & n11842 ;
  assign n44964 = ~n11842 & n44963 ;
  assign n44965 = x61 & n2979 ;
  assign n44966 = ~x61 & n44965 ;
  assign n44967 = n44964 | n44966 ;
  assign n44968 = n44964 & ~n44967 ;
  assign n44969 = ( n5455 & n6030 ) | ( n5455 & n44968 ) | ( n6030 & n44968 ) ;
  assign n44970 = n10783 & n44969 ;
  assign n44971 = n16767 & n44970 ;
  assign n44972 = n23530 | n30918 ;
  assign n44973 = n1368 | n33685 ;
  assign n44974 = n9201 ^ n3013 ^ 1'b0 ;
  assign n44975 = ( ~n10125 & n20778 ) | ( ~n10125 & n39141 ) | ( n20778 & n39141 ) ;
  assign n44976 = n22362 ^ n15944 ^ 1'b0 ;
  assign n44977 = ~n5699 & n44976 ;
  assign n44978 = n44977 ^ n41641 ^ n31329 ;
  assign n44980 = n38174 ^ n15002 ^ 1'b0 ;
  assign n44979 = n7721 & n44037 ;
  assign n44981 = n44980 ^ n44979 ^ 1'b0 ;
  assign n44982 = n44981 ^ n1396 ^ 1'b0 ;
  assign n44983 = n43123 ^ n1988 ^ 1'b0 ;
  assign n44984 = n13382 ^ n2022 ^ 1'b0 ;
  assign n44985 = ~n44983 & n44984 ;
  assign n44986 = n18289 | n42355 ;
  assign n44987 = n15862 | n22246 ;
  assign n44988 = ~n1304 & n43254 ;
  assign n44989 = n44988 ^ n25612 ^ 1'b0 ;
  assign n44990 = n44989 ^ n15692 ^ 1'b0 ;
  assign n44991 = n41237 ^ n13153 ^ n11009 ;
  assign n44992 = n18258 & ~n22661 ;
  assign n44993 = n44992 ^ n30978 ^ 1'b0 ;
  assign n44994 = ~n44077 & n44993 ;
  assign n44995 = ~n24121 & n44994 ;
  assign n44996 = n5178 | n44995 ;
  assign n44997 = n15802 ^ n3632 ^ 1'b0 ;
  assign n44998 = n15077 | n24485 ;
  assign n44999 = n44998 ^ n35638 ^ 1'b0 ;
  assign n45000 = n44999 ^ n7489 ^ 1'b0 ;
  assign n45001 = n45000 ^ n3343 ^ 1'b0 ;
  assign n45002 = n11745 & ~n45001 ;
  assign n45003 = n19399 & n22598 ;
  assign n45004 = n8216 & n45003 ;
  assign n45005 = n2082 & n6361 ;
  assign n45006 = n20941 & n45005 ;
  assign n45007 = n44857 ^ n35385 ^ n10653 ;
  assign n45008 = n31708 ^ n12895 ^ 1'b0 ;
  assign n45009 = n2512 | n45008 ;
  assign n45010 = ~n15040 & n27020 ;
  assign n45011 = n45010 ^ n2684 ^ 1'b0 ;
  assign n45012 = n30174 & ~n45011 ;
  assign n45013 = n45012 ^ n31437 ^ 1'b0 ;
  assign n45014 = ~n45009 & n45013 ;
  assign n45015 = ( n13469 & n18886 ) | ( n13469 & n20731 ) | ( n18886 & n20731 ) ;
  assign n45016 = n1164 | n45015 ;
  assign n45017 = n4907 ^ n4471 ^ 1'b0 ;
  assign n45018 = ~n45016 & n45017 ;
  assign n45019 = n36547 ^ n35531 ^ 1'b0 ;
  assign n45020 = ~n3573 & n5452 ;
  assign n45021 = n12083 & n36469 ;
  assign n45022 = n45021 ^ n18749 ^ 1'b0 ;
  assign n45024 = ~n9891 & n14618 ;
  assign n45023 = ~n4124 & n22883 ;
  assign n45025 = n45024 ^ n45023 ^ n26671 ;
  assign n45026 = ~n20587 & n41199 ;
  assign n45027 = n10953 ^ n5399 ^ 1'b0 ;
  assign n45028 = n4532 & ~n45027 ;
  assign n45029 = n45028 ^ n31336 ^ 1'b0 ;
  assign n45030 = ~n2506 & n14258 ;
  assign n45031 = n18376 & n24914 ;
  assign n45032 = n45031 ^ n16239 ^ 1'b0 ;
  assign n45033 = ~n37317 & n45032 ;
  assign n45034 = n13937 ^ n10351 ^ n9196 ;
  assign n45035 = n45034 ^ n25551 ^ x14 ;
  assign n45036 = n37668 ^ n14154 ^ 1'b0 ;
  assign n45037 = n13075 & ~n45036 ;
  assign n45038 = n45037 ^ n22665 ^ 1'b0 ;
  assign n45039 = n15637 ^ n4855 ^ 1'b0 ;
  assign n45040 = ~n8588 & n45039 ;
  assign n45041 = ~n12917 & n45040 ;
  assign n45042 = n45041 ^ n17184 ^ 1'b0 ;
  assign n45043 = n45042 ^ n22269 ^ 1'b0 ;
  assign n45044 = ( n15027 & ~n29724 ) | ( n15027 & n45043 ) | ( ~n29724 & n45043 ) ;
  assign n45045 = n13056 & n28656 ;
  assign n45046 = n16584 & n30316 ;
  assign n45047 = ~n4142 & n45046 ;
  assign n45048 = ( n22665 & n45045 ) | ( n22665 & n45047 ) | ( n45045 & n45047 ) ;
  assign n45049 = n6784 & n8137 ;
  assign n45050 = ~n45048 & n45049 ;
  assign n45051 = ( n3622 & n5550 ) | ( n3622 & ~n12080 ) | ( n5550 & ~n12080 ) ;
  assign n45052 = n4754 | n45051 ;
  assign n45053 = n10872 | n45052 ;
  assign n45054 = n13568 ^ n8477 ^ 1'b0 ;
  assign n45055 = n14248 & n45054 ;
  assign n45056 = n714 | n18070 ;
  assign n45057 = n45056 ^ n20046 ^ 1'b0 ;
  assign n45058 = ~x235 & n13181 ;
  assign n45059 = x14 & x79 ;
  assign n45060 = n45059 ^ n7932 ^ 1'b0 ;
  assign n45061 = n45060 ^ n22390 ^ n2689 ;
  assign n45062 = ~n4831 & n5070 ;
  assign n45063 = n45062 ^ n39712 ^ n2020 ;
  assign n45064 = n21865 ^ n6069 ^ 1'b0 ;
  assign n45065 = n3278 & ~n17595 ;
  assign n45066 = n38994 ^ n6950 ^ 1'b0 ;
  assign n45067 = ~n4126 & n45066 ;
  assign n45068 = n7182 & ~n8936 ;
  assign n45069 = n5586 & n45068 ;
  assign n45070 = ~n3363 & n10855 ;
  assign n45071 = n45069 & n45070 ;
  assign n45072 = ~n4421 & n37036 ;
  assign n45076 = n2955 & ~n22669 ;
  assign n45073 = ~n557 & n9638 ;
  assign n45074 = ~n27329 & n45073 ;
  assign n45075 = n4491 | n45074 ;
  assign n45077 = n45076 ^ n45075 ^ n6417 ;
  assign n45079 = n8634 & ~n25175 ;
  assign n45078 = n326 | n27581 ;
  assign n45080 = n45079 ^ n45078 ^ 1'b0 ;
  assign n45081 = ( n8477 & n32790 ) | ( n8477 & ~n45080 ) | ( n32790 & ~n45080 ) ;
  assign n45082 = n16239 ^ n8417 ^ 1'b0 ;
  assign n45083 = ~n5751 & n36450 ;
  assign n45085 = n36913 & n38504 ;
  assign n45084 = n18275 & n29324 ;
  assign n45086 = n45085 ^ n45084 ^ 1'b0 ;
  assign n45087 = n25501 ^ n17447 ^ 1'b0 ;
  assign n45088 = ( n8329 & n38654 ) | ( n8329 & ~n41094 ) | ( n38654 & ~n41094 ) ;
  assign n45090 = ~n19019 & n20471 ;
  assign n45089 = n2120 & ~n10271 ;
  assign n45091 = n45090 ^ n45089 ^ 1'b0 ;
  assign n45092 = n45088 & ~n45091 ;
  assign n45093 = ~n19729 & n41549 ;
  assign n45094 = n19847 | n23142 ;
  assign n45095 = n45094 ^ n25890 ^ 1'b0 ;
  assign n45096 = n11956 | n25360 ;
  assign n45097 = n23974 & ~n45096 ;
  assign n45098 = n9289 & ~n45097 ;
  assign n45099 = n5200 & ~n37027 ;
  assign n45100 = n45099 ^ n16045 ^ 1'b0 ;
  assign n45101 = n45100 ^ n21446 ^ n18449 ;
  assign n45102 = n39719 ^ n29982 ^ 1'b0 ;
  assign n45103 = ~n15820 & n19512 ;
  assign n45104 = n37863 & n45103 ;
  assign n45105 = n15734 ^ x94 ^ 1'b0 ;
  assign n45106 = n9998 & ~n45105 ;
  assign n45107 = n7495 & n16234 ;
  assign n45108 = n45107 ^ n35375 ^ 1'b0 ;
  assign n45109 = n39195 ^ n8620 ^ 1'b0 ;
  assign n45110 = n38457 | n45109 ;
  assign n45111 = n45110 ^ n36979 ^ 1'b0 ;
  assign n45112 = ~n16189 & n22452 ;
  assign n45113 = n42188 & n45112 ;
  assign n45114 = n8791 ^ n4902 ^ n1213 ;
  assign n45115 = ~n45113 & n45114 ;
  assign n45116 = ~n34291 & n45115 ;
  assign n45117 = n2234 & n6516 ;
  assign n45118 = ( ~n12210 & n34789 ) | ( ~n12210 & n45117 ) | ( n34789 & n45117 ) ;
  assign n45119 = ( n10332 & n32164 ) | ( n10332 & ~n45118 ) | ( n32164 & ~n45118 ) ;
  assign n45120 = n13547 ^ n5956 ^ n1433 ;
  assign n45121 = n45120 ^ n22527 ^ 1'b0 ;
  assign n45123 = n35652 & ~n39886 ;
  assign n45124 = n45123 ^ n16257 ^ 1'b0 ;
  assign n45122 = ~n2661 & n33087 ;
  assign n45125 = n45124 ^ n45122 ^ 1'b0 ;
  assign n45126 = n18344 & ~n38715 ;
  assign n45127 = ~n15994 & n45126 ;
  assign n45128 = ~n9934 & n23366 ;
  assign n45129 = ~n5915 & n45128 ;
  assign n45130 = n9224 & n42014 ;
  assign n45131 = n3144 ^ x7 ^ 1'b0 ;
  assign n45132 = n599 & n45131 ;
  assign n45133 = n45132 ^ n17084 ^ 1'b0 ;
  assign n45134 = ( n5243 & ~n17820 ) | ( n5243 & n23513 ) | ( ~n17820 & n23513 ) ;
  assign n45135 = n13272 ^ n13140 ^ 1'b0 ;
  assign n45136 = n8531 & n27174 ;
  assign n45137 = ~n5040 & n45136 ;
  assign n45138 = n6563 ^ n1805 ^ 1'b0 ;
  assign n45139 = ~n14371 & n45138 ;
  assign n45140 = n41067 ^ n643 ^ 1'b0 ;
  assign n45141 = ( n37406 & n37502 ) | ( n37406 & ~n45140 ) | ( n37502 & ~n45140 ) ;
  assign n45142 = x109 & ~n45141 ;
  assign n45143 = n18775 ^ x30 ^ 1'b0 ;
  assign n45144 = n45142 | n45143 ;
  assign n45145 = n5230 & ~n7756 ;
  assign n45146 = n34994 & n45145 ;
  assign n45147 = ~n40688 & n45146 ;
  assign n45148 = n12978 & n45147 ;
  assign n45149 = n6537 & n14963 ;
  assign n45150 = ~n29484 & n45149 ;
  assign n45151 = n24696 & ~n45150 ;
  assign n45152 = n45151 ^ n34356 ^ 1'b0 ;
  assign n45153 = n34078 ^ n26111 ^ 1'b0 ;
  assign n45154 = n19994 | n45153 ;
  assign n45155 = n13939 & ~n26581 ;
  assign n45156 = ~n17772 & n24261 ;
  assign n45157 = n5413 ^ n1347 ^ n471 ;
  assign n45158 = n22344 & ~n45157 ;
  assign n45159 = ~n590 & n45158 ;
  assign n45160 = ~n3127 & n44370 ;
  assign n45161 = n36818 & n45160 ;
  assign n45162 = n22713 ^ n797 ^ 1'b0 ;
  assign n45163 = n11516 ^ n7834 ^ n2552 ;
  assign n45165 = n33136 ^ n27759 ^ n5775 ;
  assign n45166 = n23960 ^ n8125 ^ 1'b0 ;
  assign n45167 = ~n45165 & n45166 ;
  assign n45164 = n3394 & ~n7824 ;
  assign n45168 = n45167 ^ n45164 ^ 1'b0 ;
  assign n45170 = n14352 ^ n4561 ^ 1'b0 ;
  assign n45171 = n45170 ^ n25094 ^ 1'b0 ;
  assign n45172 = n14012 & n45171 ;
  assign n45173 = n14562 | n25405 ;
  assign n45174 = n45173 ^ n40689 ^ 1'b0 ;
  assign n45175 = n45172 & n45174 ;
  assign n45169 = ( n4569 & n13801 ) | ( n4569 & ~n21515 ) | ( n13801 & ~n21515 ) ;
  assign n45176 = n45175 ^ n45169 ^ 1'b0 ;
  assign n45177 = n25659 ^ n25160 ^ 1'b0 ;
  assign n45178 = n42645 ^ n4415 ^ 1'b0 ;
  assign n45179 = ~n45177 & n45178 ;
  assign n45180 = ( n3834 & ~n9489 ) | ( n3834 & n45179 ) | ( ~n9489 & n45179 ) ;
  assign n45182 = n4405 ^ n2422 ^ n1499 ;
  assign n45183 = ~n21198 & n45182 ;
  assign n45184 = n45183 ^ n13360 ^ 1'b0 ;
  assign n45181 = n39723 ^ n3481 ^ 1'b0 ;
  assign n45185 = n45184 ^ n45181 ^ n29473 ;
  assign n45188 = n11989 ^ n4741 ^ 1'b0 ;
  assign n45190 = ~n12700 & n16043 ;
  assign n45191 = ~n34286 & n45190 ;
  assign n45192 = n45191 ^ n12647 ^ 1'b0 ;
  assign n45189 = n5603 & n13760 ;
  assign n45193 = n45192 ^ n45189 ^ 1'b0 ;
  assign n45194 = n45188 | n45193 ;
  assign n45186 = n26422 | n27449 ;
  assign n45187 = n13646 & ~n45186 ;
  assign n45195 = n45194 ^ n45187 ^ 1'b0 ;
  assign n45196 = n1519 & n8503 ;
  assign n45197 = n45196 ^ n27896 ^ n27578 ;
  assign n45198 = n13372 | n45197 ;
  assign n45199 = n45198 ^ n16625 ^ 1'b0 ;
  assign n45200 = n5448 & ~n38889 ;
  assign n45201 = n36269 ^ n27025 ^ 1'b0 ;
  assign n45202 = n960 & n33301 ;
  assign n45203 = n39465 ^ n24849 ^ 1'b0 ;
  assign n45204 = n12483 ^ n1855 ^ 1'b0 ;
  assign n45205 = n1027 & n45204 ;
  assign n45206 = n45205 ^ n14474 ^ 1'b0 ;
  assign n45207 = n21365 ^ n3806 ^ 1'b0 ;
  assign n45208 = n29567 & n45207 ;
  assign n45209 = ~n10289 & n26611 ;
  assign n45210 = n460 | n14175 ;
  assign n45211 = n45210 ^ n18771 ^ 1'b0 ;
  assign n45212 = n45211 ^ n9261 ^ 1'b0 ;
  assign n45213 = n17182 & ~n45212 ;
  assign n45214 = n14605 & n34639 ;
  assign n45215 = ~n45213 & n45214 ;
  assign n45216 = n13469 ^ n8293 ^ 1'b0 ;
  assign n45217 = n13533 & ~n45216 ;
  assign n45225 = n5853 ^ n688 ^ 1'b0 ;
  assign n45221 = n17738 ^ n11885 ^ 1'b0 ;
  assign n45222 = ~n13873 & n45221 ;
  assign n45223 = n45222 ^ n15849 ^ 1'b0 ;
  assign n45224 = n25989 & n45223 ;
  assign n45218 = n8889 | n16642 ;
  assign n45219 = n45218 ^ n2169 ^ 1'b0 ;
  assign n45220 = n13873 | n45219 ;
  assign n45226 = n45225 ^ n45224 ^ n45220 ;
  assign n45227 = n11287 & ~n18879 ;
  assign n45228 = n45227 ^ n34503 ^ 1'b0 ;
  assign n45229 = n6781 | n45228 ;
  assign n45230 = n2528 & n12448 ;
  assign n45231 = n20223 | n29657 ;
  assign n45232 = n16597 ^ n4493 ^ 1'b0 ;
  assign n45233 = n18616 ^ n2182 ^ 1'b0 ;
  assign n45234 = ~n45232 & n45233 ;
  assign n45235 = ~n5637 & n7023 ;
  assign n45236 = n12994 & n23998 ;
  assign n45237 = ~n45235 & n45236 ;
  assign n45238 = n24934 | n27694 ;
  assign n45239 = n45238 ^ n3472 ^ 1'b0 ;
  assign n45240 = ~n6510 & n10060 ;
  assign n45241 = n35686 ^ n4207 ^ 1'b0 ;
  assign n45242 = n23332 ^ n10504 ^ n9298 ;
  assign n45243 = n38647 & n43817 ;
  assign n45244 = ( ~n17571 & n17634 ) | ( ~n17571 & n39206 ) | ( n17634 & n39206 ) ;
  assign n45245 = n593 & ~n45244 ;
  assign n45246 = n3568 | n6483 ;
  assign n45247 = n3321 | n45246 ;
  assign n45248 = n37090 & n45247 ;
  assign n45249 = n45248 ^ n357 ^ 1'b0 ;
  assign n45250 = n3002 & ~n8779 ;
  assign n45251 = n9869 & n39425 ;
  assign n45252 = n45250 & n45251 ;
  assign n45253 = n1557 & n30103 ;
  assign n45254 = n32628 & n45253 ;
  assign n45255 = n8477 | n16610 ;
  assign n45256 = n4442 & ~n19741 ;
  assign n45257 = n3958 & n45256 ;
  assign n45258 = ( n33711 & ~n41961 ) | ( n33711 & n45257 ) | ( ~n41961 & n45257 ) ;
  assign n45259 = n29544 & ~n40160 ;
  assign n45260 = n45259 ^ n11529 ^ 1'b0 ;
  assign n45261 = ~n4898 & n10798 ;
  assign n45263 = n11559 | n11885 ;
  assign n45262 = ~n14669 & n44892 ;
  assign n45264 = n45263 ^ n45262 ^ 1'b0 ;
  assign n45265 = n22001 ^ n20450 ^ 1'b0 ;
  assign n45266 = ~n13640 & n45265 ;
  assign n45267 = n35420 ^ n6225 ^ 1'b0 ;
  assign n45268 = n17707 & n25493 ;
  assign n45269 = n583 & ~n17254 ;
  assign n45270 = n3365 & n45269 ;
  assign n45271 = n45270 ^ n10128 ^ 1'b0 ;
  assign n45272 = ( ~n38936 & n45268 ) | ( ~n38936 & n45271 ) | ( n45268 & n45271 ) ;
  assign n45273 = n11075 ^ n3574 ^ 1'b0 ;
  assign n45274 = n2501 ^ n2455 ^ 1'b0 ;
  assign n45275 = n15453 | n26338 ;
  assign n45276 = n45275 ^ n27198 ^ 1'b0 ;
  assign n45277 = n24341 ^ n7739 ^ 1'b0 ;
  assign n45278 = ~n2509 & n30341 ;
  assign n45279 = ~n20190 & n45278 ;
  assign n45280 = n45279 ^ n32327 ^ 1'b0 ;
  assign n45281 = x108 & ~n30845 ;
  assign n45282 = n16865 ^ n7686 ^ 1'b0 ;
  assign n45283 = ~n29422 & n39398 ;
  assign n45284 = ~n19596 & n45283 ;
  assign n45285 = n19198 ^ n10209 ^ 1'b0 ;
  assign n45286 = n3119 & n45285 ;
  assign n45287 = n45286 ^ n2422 ^ 1'b0 ;
  assign n45288 = n27288 | n45287 ;
  assign n45289 = n22861 & ~n30929 ;
  assign n45290 = ~n9192 & n45289 ;
  assign n45291 = n28501 ^ n21199 ^ 1'b0 ;
  assign n45292 = n28604 & ~n45291 ;
  assign n45293 = n5129 & ~n23260 ;
  assign n45294 = ( n3183 & ~n34766 ) | ( n3183 & n45293 ) | ( ~n34766 & n45293 ) ;
  assign n45295 = n15020 ^ n2326 ^ 1'b0 ;
  assign n45296 = ~n9790 & n45295 ;
  assign n45297 = n45296 ^ n24328 ^ n10761 ;
  assign n45298 = n26249 ^ n14192 ^ 1'b0 ;
  assign n45299 = n16464 & n22145 ;
  assign n45300 = n7409 | n8075 ;
  assign n45301 = n45300 ^ n9506 ^ 1'b0 ;
  assign n45302 = n27534 & ~n29731 ;
  assign n45303 = ~n45301 & n45302 ;
  assign n45304 = n4550 & n23581 ;
  assign n45305 = n25929 ^ n3158 ^ 1'b0 ;
  assign n45306 = n45304 & ~n45305 ;
  assign n45307 = ( n2221 & n10440 ) | ( n2221 & n29422 ) | ( n10440 & n29422 ) ;
  assign n45308 = n21370 ^ n21017 ^ 1'b0 ;
  assign n45309 = n4292 | n45308 ;
  assign n45310 = ( n40050 & n45307 ) | ( n40050 & n45309 ) | ( n45307 & n45309 ) ;
  assign n45311 = n28565 ^ n7756 ^ 1'b0 ;
  assign n45312 = n8594 & n45311 ;
  assign n45315 = n3754 | n4909 ;
  assign n45316 = n45315 ^ x206 ^ 1'b0 ;
  assign n45317 = n27696 & n45316 ;
  assign n45313 = ( n4426 & n7963 ) | ( n4426 & ~n9178 ) | ( n7963 & ~n9178 ) ;
  assign n45314 = n3687 & ~n45313 ;
  assign n45318 = n45317 ^ n45314 ^ n40768 ;
  assign n45320 = ~n8680 & n28692 ;
  assign n45321 = n45320 ^ n10696 ^ 1'b0 ;
  assign n45322 = ( ~n10801 & n29050 ) | ( ~n10801 & n45321 ) | ( n29050 & n45321 ) ;
  assign n45319 = n411 & ~n22742 ;
  assign n45323 = n45322 ^ n45319 ^ n37424 ;
  assign n45324 = n9993 | n25818 ;
  assign n45325 = n29158 & ~n45324 ;
  assign n45326 = n20926 | n21846 ;
  assign n45327 = n8497 & ~n45326 ;
  assign n45328 = n45325 & n45327 ;
  assign n45329 = n45328 ^ n15219 ^ 1'b0 ;
  assign n45330 = n19396 & ~n22244 ;
  assign n45331 = n418 | n19326 ;
  assign n45332 = n45331 ^ n39514 ^ 1'b0 ;
  assign n45333 = ~n16534 & n27343 ;
  assign n45334 = n19191 ^ n8811 ^ 1'b0 ;
  assign n45335 = n33739 & ~n45334 ;
  assign n45336 = n1311 & n10677 ;
  assign n45337 = n13452 | n24611 ;
  assign n45338 = x65 | n45337 ;
  assign n45339 = ~n23851 & n45338 ;
  assign n45340 = x185 | n3287 ;
  assign n45341 = n20120 | n33971 ;
  assign n45342 = ~n23609 & n45341 ;
  assign n45343 = n16534 & ~n35506 ;
  assign n45344 = n3659 | n5059 ;
  assign n45345 = n45343 | n45344 ;
  assign n45346 = n20261 | n32625 ;
  assign n45347 = n23317 & ~n28987 ;
  assign n45348 = n45347 ^ n42126 ^ 1'b0 ;
  assign n45349 = n3172 & n45348 ;
  assign n45350 = n2440 ^ n1232 ^ 1'b0 ;
  assign n45351 = ~n14362 & n45350 ;
  assign n45352 = ( n1829 & ~n33720 ) | ( n1829 & n45351 ) | ( ~n33720 & n45351 ) ;
  assign n45353 = ( n3562 & ~n19033 ) | ( n3562 & n29351 ) | ( ~n19033 & n29351 ) ;
  assign n45354 = n45353 ^ n37653 ^ n1404 ;
  assign n45355 = n39708 ^ n4775 ^ 1'b0 ;
  assign n45356 = n45355 ^ n9581 ^ 1'b0 ;
  assign n45357 = n1850 & n14449 ;
  assign n45358 = n45357 ^ x41 ^ 1'b0 ;
  assign n45359 = ( n10070 & ~n17324 ) | ( n10070 & n45358 ) | ( ~n17324 & n45358 ) ;
  assign n45360 = ( n24228 & n37073 ) | ( n24228 & ~n45359 ) | ( n37073 & ~n45359 ) ;
  assign n45361 = n43806 | n45360 ;
  assign n45362 = n45361 ^ n32713 ^ 1'b0 ;
  assign n45363 = n21877 | n24924 ;
  assign n45364 = n45363 ^ n19738 ^ 1'b0 ;
  assign n45365 = n14673 ^ n1981 ^ 1'b0 ;
  assign n45366 = n25018 ^ n19677 ^ 1'b0 ;
  assign n45367 = n45366 ^ n23370 ^ 1'b0 ;
  assign n45368 = n29538 ^ n16490 ^ 1'b0 ;
  assign n45369 = n1975 | n45368 ;
  assign n45370 = n42623 ^ n7987 ^ n6375 ;
  assign n45371 = n12850 ^ n1024 ^ 1'b0 ;
  assign n45372 = n1346 | n7714 ;
  assign n45373 = n8345 & ~n16409 ;
  assign n45374 = ~n33487 & n45373 ;
  assign n45375 = n3261 & n19425 ;
  assign n45376 = n8622 & ~n20058 ;
  assign n45377 = ~n20987 & n45376 ;
  assign n45378 = n45377 ^ n11213 ^ 1'b0 ;
  assign n45379 = ~n45375 & n45378 ;
  assign n45380 = n38006 ^ n9843 ^ 1'b0 ;
  assign n45381 = n3738 & ~n45380 ;
  assign n45382 = n27450 ^ n6881 ^ 1'b0 ;
  assign n45383 = ~n17845 & n45382 ;
  assign n45384 = n8048 & ~n11143 ;
  assign n45385 = ~n4458 & n45384 ;
  assign n45386 = n20721 ^ n16133 ^ n8453 ;
  assign n45387 = n39841 ^ n2127 ^ 1'b0 ;
  assign n45388 = n3815 | n19326 ;
  assign n45389 = n45388 ^ n7322 ^ 1'b0 ;
  assign n45390 = ( n23736 & n39570 ) | ( n23736 & ~n45389 ) | ( n39570 & ~n45389 ) ;
  assign n45391 = ( n7750 & n17495 ) | ( n7750 & n45390 ) | ( n17495 & n45390 ) ;
  assign n45396 = n20285 | n28576 ;
  assign n45392 = n23280 & ~n34200 ;
  assign n45393 = n45392 ^ n6774 ^ 1'b0 ;
  assign n45394 = n17739 & ~n45393 ;
  assign n45395 = n33726 | n45394 ;
  assign n45397 = n45396 ^ n45395 ^ 1'b0 ;
  assign n45398 = n45397 ^ n36111 ^ 1'b0 ;
  assign n45399 = n8066 & n45398 ;
  assign n45400 = n8086 ^ n7901 ^ 1'b0 ;
  assign n45401 = n18360 & n45400 ;
  assign n45402 = n1999 & ~n5637 ;
  assign n45403 = n45402 ^ n17467 ^ 1'b0 ;
  assign n45404 = n45403 ^ n18271 ^ 1'b0 ;
  assign n45405 = n16547 & ~n25686 ;
  assign n45406 = n38226 & n45405 ;
  assign n45407 = n9425 ^ n2434 ^ 1'b0 ;
  assign n45408 = n45407 ^ n20527 ^ n12790 ;
  assign n45409 = ( n1233 & n10218 ) | ( n1233 & ~n45408 ) | ( n10218 & ~n45408 ) ;
  assign n45410 = ( ~n5843 & n20027 ) | ( ~n5843 & n28579 ) | ( n20027 & n28579 ) ;
  assign n45411 = ( n9486 & ~n20958 ) | ( n9486 & n21895 ) | ( ~n20958 & n21895 ) ;
  assign n45412 = n23560 ^ n11548 ^ 1'b0 ;
  assign n45413 = ~n1728 & n45412 ;
  assign n45414 = ~n41365 & n45413 ;
  assign n45415 = n42977 ^ n18934 ^ 1'b0 ;
  assign n45416 = ~n36256 & n45415 ;
  assign n45417 = n17420 & ~n18490 ;
  assign n45418 = ~n45416 & n45417 ;
  assign n45419 = n10066 | n10231 ;
  assign n45420 = n45419 ^ n31999 ^ 1'b0 ;
  assign n45421 = x30 & ~n45420 ;
  assign n45422 = n45421 ^ n6322 ^ 1'b0 ;
  assign n45423 = ( ~n3579 & n7435 ) | ( ~n3579 & n12455 ) | ( n7435 & n12455 ) ;
  assign n45424 = n45423 ^ n32022 ^ n10913 ;
  assign n45425 = n42058 & n45424 ;
  assign n45426 = n45425 ^ n24468 ^ 1'b0 ;
  assign n45430 = n17302 ^ n15580 ^ 1'b0 ;
  assign n45431 = n3791 & n45430 ;
  assign n45432 = n14285 & n45431 ;
  assign n45429 = ~n21559 & n27586 ;
  assign n45427 = n3011 | n14773 ;
  assign n45428 = n45427 ^ n25778 ^ 1'b0 ;
  assign n45433 = n45432 ^ n45429 ^ n45428 ;
  assign n45434 = n38423 ^ n30072 ^ 1'b0 ;
  assign n45435 = x61 & n3804 ;
  assign n45436 = ( n27031 & n40352 ) | ( n27031 & n40388 ) | ( n40352 & n40388 ) ;
  assign n45437 = n45436 ^ n40618 ^ 1'b0 ;
  assign n45438 = n26858 & ~n45437 ;
  assign n45439 = n3493 | n18205 ;
  assign n45440 = n10292 | n32848 ;
  assign n45441 = n23050 ^ n5632 ^ 1'b0 ;
  assign n45442 = ~n7788 & n11252 ;
  assign n45443 = n24700 & n45442 ;
  assign n45444 = n33097 ^ n31686 ^ 1'b0 ;
  assign n45445 = n27947 & n30414 ;
  assign n45446 = n45444 & n45445 ;
  assign n45447 = ~n14027 & n26625 ;
  assign n45448 = n11342 & n45447 ;
  assign n45449 = n41551 ^ n9156 ^ 1'b0 ;
  assign n45450 = ~n45448 & n45449 ;
  assign n45451 = n42139 ^ n16870 ^ n2728 ;
  assign n45452 = n30618 ^ n3897 ^ 1'b0 ;
  assign n45453 = n16512 & ~n39911 ;
  assign n45454 = ~n6971 & n21949 ;
  assign n45455 = n39504 ^ n19232 ^ 1'b0 ;
  assign n45456 = n41162 | n45455 ;
  assign n45457 = n7485 | n45456 ;
  assign n45458 = n45454 & ~n45457 ;
  assign n45459 = n19352 ^ n13574 ^ 1'b0 ;
  assign n45460 = n45459 ^ n7925 ^ n2617 ;
  assign n45461 = n44064 & ~n45460 ;
  assign n45462 = n35638 ^ n14310 ^ n12629 ;
  assign n45463 = n45461 | n45462 ;
  assign n45464 = n30788 ^ n18594 ^ 1'b0 ;
  assign n45465 = ~n18778 & n39349 ;
  assign n45466 = ~n10886 & n45465 ;
  assign n45467 = n20542 & n20578 ;
  assign n45468 = n45467 ^ n14784 ^ 1'b0 ;
  assign n45469 = n972 | n33094 ;
  assign n45470 = ~n13505 & n45469 ;
  assign n45471 = n31260 & n41609 ;
  assign n45472 = ~n42691 & n45471 ;
  assign n45473 = ( n4626 & n29171 ) | ( n4626 & ~n45472 ) | ( n29171 & ~n45472 ) ;
  assign n45474 = n18899 ^ n13080 ^ 1'b0 ;
  assign n45475 = ~n28166 & n45474 ;
  assign n45476 = n19267 & n45475 ;
  assign n45477 = n15430 ^ n5865 ^ 1'b0 ;
  assign n45478 = ~n15930 & n45477 ;
  assign n45479 = x0 & ~n18396 ;
  assign n45480 = n357 | n45479 ;
  assign n45481 = n1036 | n23628 ;
  assign n45482 = n15002 & n15621 ;
  assign n45483 = n35126 | n45482 ;
  assign n45484 = ( n21388 & n26556 ) | ( n21388 & n43157 ) | ( n26556 & n43157 ) ;
  assign n45485 = n41408 & ~n45484 ;
  assign n45486 = n13354 ^ n3242 ^ 1'b0 ;
  assign n45487 = n12971 & n45486 ;
  assign n45488 = n31634 & n34715 ;
  assign n45489 = ~n45487 & n45488 ;
  assign n45490 = n11713 ^ n3283 ^ 1'b0 ;
  assign n45491 = n1783 & ~n45490 ;
  assign n45492 = n45491 ^ n28280 ^ 1'b0 ;
  assign n45493 = n21771 & n45492 ;
  assign n45494 = n4435 ^ n4331 ^ 1'b0 ;
  assign n45495 = n4659 & ~n45494 ;
  assign n45496 = n3501 & ~n32817 ;
  assign n45497 = n45496 ^ n19960 ^ 1'b0 ;
  assign n45498 = n19668 | n45497 ;
  assign n45499 = n45495 | n45498 ;
  assign n45503 = n8781 ^ n5999 ^ 1'b0 ;
  assign n45504 = n40623 & ~n45503 ;
  assign n45500 = ( ~n2855 & n21349 ) | ( ~n2855 & n32690 ) | ( n21349 & n32690 ) ;
  assign n45501 = n6180 & ~n45500 ;
  assign n45502 = n1457 & n45501 ;
  assign n45505 = n45504 ^ n45502 ^ 1'b0 ;
  assign n45506 = n31031 ^ n19894 ^ 1'b0 ;
  assign n45507 = n31164 ^ n11696 ^ n1184 ;
  assign n45508 = ~n8325 & n45507 ;
  assign n45509 = n17518 & n45508 ;
  assign n45510 = n36968 ^ n21053 ^ n9983 ;
  assign n45511 = n4931 & n12579 ;
  assign n45512 = ~n45510 & n45511 ;
  assign n45513 = n9416 ^ n6833 ^ n3253 ;
  assign n45514 = n23019 ^ n2317 ^ 1'b0 ;
  assign n45515 = n7838 | n45514 ;
  assign n45516 = n45515 ^ n19895 ^ 1'b0 ;
  assign n45517 = n19536 ^ n16820 ^ 1'b0 ;
  assign n45518 = ~n19147 & n45517 ;
  assign n45519 = n28200 ^ x134 ^ 1'b0 ;
  assign n45520 = n14264 & ~n45519 ;
  assign n45521 = ~n7333 & n8130 ;
  assign n45522 = n45521 ^ n19998 ^ 1'b0 ;
  assign n45523 = n19941 & ~n21584 ;
  assign n45524 = n15946 & ~n16131 ;
  assign n45525 = n8919 | n28270 ;
  assign n45526 = n8266 | n45525 ;
  assign n45527 = n16165 ^ n14304 ^ 1'b0 ;
  assign n45528 = n17387 | n45527 ;
  assign n45529 = n45528 ^ n35927 ^ 1'b0 ;
  assign n45530 = n6322 ^ n1611 ^ 1'b0 ;
  assign n45531 = n37729 & ~n45530 ;
  assign n45532 = n30551 ^ n1553 ^ 1'b0 ;
  assign n45533 = n9170 | n45532 ;
  assign n45534 = x243 & n27040 ;
  assign n45536 = ( ~n861 & n9029 ) | ( ~n861 & n14340 ) | ( n9029 & n14340 ) ;
  assign n45535 = ~n20007 & n29247 ;
  assign n45537 = n45536 ^ n45535 ^ n25552 ;
  assign n45538 = n24016 | n44438 ;
  assign n45539 = n45537 | n45538 ;
  assign n45540 = n12637 & n29505 ;
  assign n45541 = ( n577 & n6874 ) | ( n577 & ~n45540 ) | ( n6874 & ~n45540 ) ;
  assign n45542 = n38828 ^ n21797 ^ 1'b0 ;
  assign n45543 = n5623 & n45542 ;
  assign n45544 = n45543 ^ n32849 ^ 1'b0 ;
  assign n45545 = n45541 & ~n45544 ;
  assign n45546 = n39223 ^ n33025 ^ 1'b0 ;
  assign n45547 = n36283 & ~n45546 ;
  assign n45548 = ( n1340 & n17707 ) | ( n1340 & ~n45547 ) | ( n17707 & ~n45547 ) ;
  assign n45549 = n4036 & ~n18805 ;
  assign n45550 = n8605 | n42136 ;
  assign n45551 = n42136 & ~n45550 ;
  assign n45552 = n301 | n45551 ;
  assign n45553 = n752 | n45552 ;
  assign n45554 = n45553 ^ n24551 ^ 1'b0 ;
  assign n45555 = n23284 ^ n23244 ^ 1'b0 ;
  assign n45556 = n10412 & ~n32791 ;
  assign n45557 = ~n27022 & n43409 ;
  assign n45558 = n44531 ^ n34938 ^ 1'b0 ;
  assign n45559 = n4174 & ~n45558 ;
  assign n45560 = n2234 & ~n18307 ;
  assign n45561 = n22126 & ~n27949 ;
  assign n45562 = n45561 ^ n8011 ^ 1'b0 ;
  assign n45563 = n45562 ^ n10196 ^ 1'b0 ;
  assign n45564 = ~n4772 & n7130 ;
  assign n45565 = n45564 ^ n19669 ^ 1'b0 ;
  assign n45566 = n11050 | n45565 ;
  assign n45567 = n26911 ^ n20245 ^ n3072 ;
  assign n45568 = ~n7995 & n34818 ;
  assign n45569 = ( ~n31171 & n36403 ) | ( ~n31171 & n45568 ) | ( n36403 & n45568 ) ;
  assign n45570 = n44350 ^ n4211 ^ 1'b0 ;
  assign n45571 = n4741 ^ n1253 ^ 1'b0 ;
  assign n45572 = n8233 & n39218 ;
  assign n45573 = n45571 & n45572 ;
  assign n45574 = n8577 & n32669 ;
  assign n45575 = n25059 & n30300 ;
  assign n45576 = n45575 ^ n1811 ^ 1'b0 ;
  assign n45577 = n23829 ^ n14226 ^ 1'b0 ;
  assign n45578 = n31710 ^ n31290 ^ n25340 ;
  assign n45579 = n36667 ^ n516 ^ 1'b0 ;
  assign n45580 = n3112 & n21565 ;
  assign n45581 = n45580 ^ n7307 ^ 1'b0 ;
  assign n45582 = n7521 & ~n45581 ;
  assign n45583 = n17808 ^ n17471 ^ 1'b0 ;
  assign n45584 = n45582 & ~n45583 ;
  assign n45585 = ~n3043 & n45584 ;
  assign n45586 = ~n32403 & n45585 ;
  assign n45587 = n11658 & n41122 ;
  assign n45588 = n10682 ^ n10078 ^ 1'b0 ;
  assign n45589 = ~n16118 & n45588 ;
  assign n45590 = n11859 ^ n5469 ^ n4161 ;
  assign n45591 = n23429 ^ n21559 ^ 1'b0 ;
  assign n45592 = n45590 & n45591 ;
  assign n45593 = ~n13606 & n26489 ;
  assign n45596 = n13452 ^ n8123 ^ 1'b0 ;
  assign n45595 = n24281 ^ n5511 ^ 1'b0 ;
  assign n45594 = n2836 & ~n15990 ;
  assign n45597 = n45596 ^ n45595 ^ n45594 ;
  assign n45598 = n5657 & ~n39518 ;
  assign n45599 = n43802 ^ n6272 ^ 1'b0 ;
  assign n45600 = n15563 ^ n8772 ^ 1'b0 ;
  assign n45601 = n2401 | n45600 ;
  assign n45602 = n32504 & ~n45601 ;
  assign n45603 = n13906 & n45602 ;
  assign n45604 = n30355 ^ n1707 ^ 1'b0 ;
  assign n45605 = ~n4540 & n41170 ;
  assign n45606 = n7490 & n45605 ;
  assign n45607 = n5509 | n34233 ;
  assign n45608 = n36206 & ~n45607 ;
  assign n45609 = n41441 ^ n14427 ^ 1'b0 ;
  assign n45610 = n12405 & ~n45609 ;
  assign n45611 = n45610 ^ n39149 ^ 1'b0 ;
  assign n45612 = n32695 ^ n10582 ^ 1'b0 ;
  assign n45613 = n36584 & ~n40019 ;
  assign n45614 = ~n14873 & n43030 ;
  assign n45615 = n3604 | n39181 ;
  assign n45616 = n10312 & ~n45615 ;
  assign n45617 = n30208 ^ n903 ^ 1'b0 ;
  assign n45618 = n23079 ^ n21756 ^ 1'b0 ;
  assign n45619 = n18348 ^ n1033 ^ 1'b0 ;
  assign n45620 = ~n37049 & n45152 ;
  assign n45621 = n42942 & ~n43035 ;
  assign n45622 = ~n12114 & n45621 ;
  assign n45623 = n8035 & ~n12341 ;
  assign n45624 = n7360 & n45623 ;
  assign n45625 = n45624 ^ n8964 ^ 1'b0 ;
  assign n45626 = n4513 & ~n27274 ;
  assign n45627 = n45626 ^ n19724 ^ 1'b0 ;
  assign n45628 = n45627 ^ n9578 ^ 1'b0 ;
  assign n45629 = n16088 ^ n12118 ^ 1'b0 ;
  assign n45630 = n45629 ^ n17435 ^ n4493 ;
  assign n45631 = n30245 ^ n11981 ^ 1'b0 ;
  assign n45632 = n22395 & ~n45631 ;
  assign n45633 = n12402 & n21025 ;
  assign n45634 = n38555 & n45633 ;
  assign n45635 = ~n294 & n45634 ;
  assign n45636 = n6512 ^ n1967 ^ 1'b0 ;
  assign n45637 = n14623 & n45636 ;
  assign n45638 = n10338 & ~n29254 ;
  assign n45639 = ~n45637 & n45638 ;
  assign n45640 = ~n5496 & n15427 ;
  assign n45641 = n45640 ^ n34592 ^ 1'b0 ;
  assign n45642 = n28281 | n33375 ;
  assign n45643 = n45642 ^ n19825 ^ 1'b0 ;
  assign n45646 = n9181 & ~n12219 ;
  assign n45644 = n9610 & n16652 ;
  assign n45645 = n45644 ^ n26124 ^ 1'b0 ;
  assign n45647 = n45646 ^ n45645 ^ n21585 ;
  assign n45648 = n20319 ^ n3854 ^ 1'b0 ;
  assign n45649 = n21983 & ~n45648 ;
  assign n45650 = n45649 ^ n22978 ^ 1'b0 ;
  assign n45651 = ( n5352 & n15680 ) | ( n5352 & n45650 ) | ( n15680 & n45650 ) ;
  assign n45652 = ~n16143 & n21495 ;
  assign n45653 = n1235 & ~n30504 ;
  assign n45654 = n38504 & n45653 ;
  assign n45655 = n1486 & ~n45654 ;
  assign n45656 = n1697 | n31932 ;
  assign n45657 = n1777 | n45656 ;
  assign n45658 = n45657 ^ n1946 ^ 1'b0 ;
  assign n45659 = n14655 ^ n3772 ^ 1'b0 ;
  assign n45660 = n8016 & ~n45659 ;
  assign n45661 = ~n3050 & n16651 ;
  assign n45662 = n8271 & ~n13209 ;
  assign n45663 = ~n45661 & n45662 ;
  assign n45664 = n16407 | n25777 ;
  assign n45665 = n45663 & ~n45664 ;
  assign n45666 = n45665 ^ n12167 ^ n8337 ;
  assign n45667 = ( n15102 & n43782 ) | ( n15102 & ~n45666 ) | ( n43782 & ~n45666 ) ;
  assign n45668 = n41053 ^ n27863 ^ 1'b0 ;
  assign n45669 = n16417 & ~n45668 ;
  assign n45670 = n35597 & n45669 ;
  assign n45671 = n5707 & n11168 ;
  assign n45672 = ( n7035 & ~n29257 ) | ( n7035 & n45671 ) | ( ~n29257 & n45671 ) ;
  assign n45673 = n4571 & n30003 ;
  assign n45674 = n16687 | n27390 ;
  assign n45675 = n29724 & ~n45674 ;
  assign n45676 = n17657 ^ n16221 ^ n2849 ;
  assign n45677 = n36026 | n45676 ;
  assign n45678 = n697 & n9152 ;
  assign n45679 = n45678 ^ n23565 ^ 1'b0 ;
  assign n45680 = n4773 & ~n27506 ;
  assign n45681 = n5471 & n45680 ;
  assign n45682 = n1298 & n45681 ;
  assign n45683 = n16381 | n19790 ;
  assign n45684 = n18661 ^ n294 ^ 1'b0 ;
  assign n45685 = n45683 & ~n45684 ;
  assign n45686 = n30367 ^ n11124 ^ 1'b0 ;
  assign n45687 = n5425 & n12152 ;
  assign n45688 = n27524 & n45687 ;
  assign n45689 = n4363 & ~n27806 ;
  assign n45690 = n45689 ^ n286 ^ 1'b0 ;
  assign n45691 = n22511 & ~n31294 ;
  assign n45692 = n7172 & n45691 ;
  assign n45693 = n8245 & ~n14870 ;
  assign n45694 = n29202 ^ n744 ^ 1'b0 ;
  assign n45695 = ~n45693 & n45694 ;
  assign n45696 = n11684 & ~n29984 ;
  assign n45697 = n45696 ^ n30079 ^ 1'b0 ;
  assign n45698 = n6808 | n21626 ;
  assign n45699 = n33200 ^ n28049 ^ 1'b0 ;
  assign n45700 = n45698 & n45699 ;
  assign n45701 = n20395 & n29289 ;
  assign n45702 = ( n6232 & n40104 ) | ( n6232 & n41780 ) | ( n40104 & n41780 ) ;
  assign n45703 = n45702 ^ n16352 ^ n1998 ;
  assign n45704 = ~n307 & n1975 ;
  assign n45705 = n16974 | n28987 ;
  assign n45706 = n45705 ^ n4980 ^ 1'b0 ;
  assign n45707 = n45706 ^ n21732 ^ 1'b0 ;
  assign n45708 = ( n6337 & ~n45704 ) | ( n6337 & n45707 ) | ( ~n45704 & n45707 ) ;
  assign n45709 = n17677 ^ n14306 ^ 1'b0 ;
  assign n45710 = n18399 & n44084 ;
  assign n45711 = ~n11824 & n17158 ;
  assign n45712 = n45711 ^ n6546 ^ 1'b0 ;
  assign n45713 = n21589 ^ n685 ^ 1'b0 ;
  assign n45714 = n45712 | n45713 ;
  assign n45715 = n37290 ^ n6628 ^ 1'b0 ;
  assign n45716 = ~n3671 & n16622 ;
  assign n45717 = n45715 & n45716 ;
  assign n45718 = n27623 ^ n2864 ^ 1'b0 ;
  assign n45719 = n12571 & ~n19317 ;
  assign n45720 = n27153 ^ n18973 ^ n3417 ;
  assign n45721 = n13884 & ~n30122 ;
  assign n45722 = ~n3543 & n43163 ;
  assign n45723 = n15365 & n16494 ;
  assign n45725 = n23620 ^ n11667 ^ 1'b0 ;
  assign n45726 = n37105 & n45725 ;
  assign n45724 = n24000 | n36199 ;
  assign n45727 = n45726 ^ n45724 ^ 1'b0 ;
  assign n45728 = ~n713 & n9273 ;
  assign n45729 = n45728 ^ n18410 ^ 1'b0 ;
  assign n45730 = n25996 ^ n15550 ^ 1'b0 ;
  assign n45731 = n29824 & ~n45730 ;
  assign n45732 = ~n45729 & n45731 ;
  assign n45733 = x41 | n28432 ;
  assign n45734 = n45733 ^ n10935 ^ 1'b0 ;
  assign n45735 = n29135 ^ n2751 ^ 1'b0 ;
  assign n45736 = n39220 & n45735 ;
  assign n45737 = n23849 & n45736 ;
  assign n45738 = ~n10947 & n45737 ;
  assign n45739 = n45738 ^ n34793 ^ n33535 ;
  assign n45740 = n14339 & ~n33375 ;
  assign n45741 = n3431 & n30161 ;
  assign n45742 = ~n11107 & n45741 ;
  assign n45743 = n45742 ^ n44387 ^ 1'b0 ;
  assign n45749 = n29065 ^ n3334 ^ 1'b0 ;
  assign n45750 = n3460 & n45749 ;
  assign n45751 = n45750 ^ n28069 ^ n7306 ;
  assign n45747 = n8751 ^ n6998 ^ 1'b0 ;
  assign n45748 = n40341 | n45747 ;
  assign n45752 = n45751 ^ n45748 ^ n33524 ;
  assign n45744 = n3376 & n38043 ;
  assign n45745 = ~n22072 & n45744 ;
  assign n45746 = n21538 | n45745 ;
  assign n45753 = n45752 ^ n45746 ^ 1'b0 ;
  assign n45754 = n45448 ^ n14610 ^ n13604 ;
  assign n45755 = n33583 ^ n27098 ^ 1'b0 ;
  assign n45757 = n20591 ^ n6651 ^ 1'b0 ;
  assign n45756 = ~n7750 & n18473 ;
  assign n45758 = n45757 ^ n45756 ^ n28200 ;
  assign n45759 = ~n35348 & n40866 ;
  assign n45760 = n1409 & ~n4580 ;
  assign n45761 = n27706 | n42898 ;
  assign n45762 = n45761 ^ n6592 ^ 1'b0 ;
  assign n45763 = n22549 | n45762 ;
  assign n45764 = n35645 ^ n4672 ^ 1'b0 ;
  assign n45765 = n7330 & n45764 ;
  assign n45766 = ( n5443 & n16830 ) | ( n5443 & ~n42488 ) | ( n16830 & ~n42488 ) ;
  assign n45767 = ( n11332 & n24530 ) | ( n11332 & ~n30494 ) | ( n24530 & ~n30494 ) ;
  assign n45768 = n28856 & n45767 ;
  assign n45769 = n4985 | n45027 ;
  assign n45770 = n16477 & n20614 ;
  assign n45771 = n11769 ^ n5989 ^ 1'b0 ;
  assign n45772 = ~n32554 & n45771 ;
  assign n45773 = n13972 & ~n17894 ;
  assign n45774 = n11046 & n45773 ;
  assign n45775 = n30484 | n45774 ;
  assign n45776 = n45775 ^ n18895 ^ 1'b0 ;
  assign n45777 = n30482 ^ n7023 ^ 1'b0 ;
  assign n45778 = n13015 & ~n37481 ;
  assign n45779 = ~n42650 & n45778 ;
  assign n45780 = n16118 ^ n10391 ^ 1'b0 ;
  assign n45782 = n27787 ^ n7518 ^ 1'b0 ;
  assign n45783 = ~n13695 & n45782 ;
  assign n45781 = n20684 ^ n16996 ^ n6776 ;
  assign n45784 = n45783 ^ n45781 ^ n20159 ;
  assign n45785 = n45018 ^ n27144 ^ 1'b0 ;
  assign n45786 = ~n3922 & n8027 ;
  assign n45787 = n45786 ^ n10073 ^ 1'b0 ;
  assign n45788 = x24 & ~n13452 ;
  assign n45789 = ~n11328 & n45788 ;
  assign n45790 = n45789 ^ n3508 ^ 1'b0 ;
  assign n45791 = n45787 | n45790 ;
  assign n45792 = ~n27299 & n38369 ;
  assign n45793 = n45792 ^ n36525 ^ 1'b0 ;
  assign n45794 = ~n4306 & n16503 ;
  assign n45795 = n18974 ^ n16432 ^ 1'b0 ;
  assign n45796 = n45794 & n45795 ;
  assign n45797 = x190 & n45796 ;
  assign n45798 = n45797 ^ n23696 ^ 1'b0 ;
  assign n45799 = n13189 ^ n8675 ^ 1'b0 ;
  assign n45800 = n16218 & ~n45799 ;
  assign n45801 = n45800 ^ n7339 ^ 1'b0 ;
  assign n45802 = n36182 ^ n29262 ^ n13744 ;
  assign n45803 = ~n45801 & n45802 ;
  assign n45804 = n21252 ^ n2842 ^ 1'b0 ;
  assign n45805 = n12256 & ~n20734 ;
  assign n45806 = ~n35295 & n45805 ;
  assign n45807 = n27365 ^ n10236 ^ 1'b0 ;
  assign n45808 = ~n45806 & n45807 ;
  assign n45809 = n45808 ^ n28697 ^ 1'b0 ;
  assign n45810 = n4447 & n23997 ;
  assign n45811 = n21462 & n45810 ;
  assign n45812 = ~n29566 & n45811 ;
  assign n45813 = ( x178 & n14472 ) | ( x178 & ~n17352 ) | ( n14472 & ~n17352 ) ;
  assign n45814 = ~n5909 & n44762 ;
  assign n45815 = n6589 ^ n1620 ^ 1'b0 ;
  assign n45816 = n11435 | n23649 ;
  assign n45817 = n12591 & ~n45816 ;
  assign n45818 = n40623 ^ n12330 ^ n6223 ;
  assign n45819 = ( n26119 & ~n31576 ) | ( n26119 & n36022 ) | ( ~n31576 & n36022 ) ;
  assign n45820 = ~n6648 & n17175 ;
  assign n45821 = n21010 & ~n38422 ;
  assign n45822 = n19763 & n23612 ;
  assign n45823 = ~n23612 & n45822 ;
  assign n45824 = n4241 | n45823 ;
  assign n45825 = n45824 ^ n10411 ^ 1'b0 ;
  assign n45826 = n45825 ^ n42076 ^ 1'b0 ;
  assign n45827 = n11770 ^ n11474 ^ n6768 ;
  assign n45828 = ~x228 & n38814 ;
  assign n45829 = ~n27307 & n45828 ;
  assign n45830 = n9900 | n31157 ;
  assign n45831 = x43 & ~n45830 ;
  assign n45832 = n45831 ^ n6330 ^ 1'b0 ;
  assign n45833 = n24542 & ~n36256 ;
  assign n45834 = n29242 | n45833 ;
  assign n45835 = ~n5421 & n41779 ;
  assign n45836 = n2853 & ~n11784 ;
  assign n45837 = n22951 ^ n4478 ^ 1'b0 ;
  assign n45838 = n45837 ^ n607 ^ n495 ;
  assign n45839 = n12968 | n14322 ;
  assign n45840 = n14253 & ~n45839 ;
  assign n45841 = n45840 ^ n37898 ^ n16409 ;
  assign n45842 = n21590 | n32305 ;
  assign n45843 = n29473 ^ n4855 ^ 1'b0 ;
  assign n45844 = n45843 ^ n10625 ^ n10275 ;
  assign n45845 = n7277 & n15818 ;
  assign n45846 = ~n45844 & n45845 ;
  assign n45847 = ~n9867 & n33742 ;
  assign n45848 = ~n427 & n45847 ;
  assign n45849 = n34561 ^ n8076 ^ 1'b0 ;
  assign n45850 = n4784 & ~n22966 ;
  assign n45851 = n45850 ^ n19963 ^ 1'b0 ;
  assign n45852 = n45851 ^ n20721 ^ 1'b0 ;
  assign n45854 = n21846 | n34491 ;
  assign n45853 = n14088 & n25105 ;
  assign n45855 = n45854 ^ n45853 ^ 1'b0 ;
  assign n45856 = ( n21756 & ~n45852 ) | ( n21756 & n45855 ) | ( ~n45852 & n45855 ) ;
  assign n45857 = n45856 ^ n20502 ^ 1'b0 ;
  assign n45858 = n7172 | n45857 ;
  assign n45859 = n38887 ^ n15366 ^ 1'b0 ;
  assign n45860 = n2991 & ~n14970 ;
  assign n45861 = n45860 ^ n26179 ^ 1'b0 ;
  assign n45862 = n45861 ^ n13666 ^ 1'b0 ;
  assign n45863 = ( ~n18816 & n27890 ) | ( ~n18816 & n34892 ) | ( n27890 & n34892 ) ;
  assign n45864 = ~n17992 & n26099 ;
  assign n45865 = ~n11413 & n32099 ;
  assign n45866 = n34040 & n45865 ;
  assign n45867 = n12357 & n45024 ;
  assign n45868 = n45867 ^ n1048 ^ 1'b0 ;
  assign n45869 = n23223 ^ n2434 ^ 1'b0 ;
  assign n45870 = n45868 | n45869 ;
  assign n45871 = n11986 ^ n9802 ^ 1'b0 ;
  assign n45872 = ~n7253 & n45871 ;
  assign n45873 = n2765 | n11690 ;
  assign n45874 = n45873 ^ n22827 ^ 1'b0 ;
  assign n45875 = n12384 ^ n9661 ^ 1'b0 ;
  assign n45876 = n45874 & ~n45875 ;
  assign n45877 = ( ~n4910 & n8717 ) | ( ~n4910 & n45876 ) | ( n8717 & n45876 ) ;
  assign n45878 = ~n774 & n45877 ;
  assign n45879 = ~n45872 & n45878 ;
  assign n45880 = n26832 | n38485 ;
  assign n45881 = n45880 ^ n23502 ^ 1'b0 ;
  assign n45882 = n1347 & ~n4467 ;
  assign n45883 = n5157 ^ n2194 ^ 1'b0 ;
  assign n45884 = n11070 | n14543 ;
  assign n45885 = ~n5921 & n45884 ;
  assign n45886 = n2041 & ~n14520 ;
  assign n45887 = n45886 ^ n18832 ^ 1'b0 ;
  assign n45888 = n28488 | n45887 ;
  assign n45889 = n45888 ^ n21487 ^ 1'b0 ;
  assign n45890 = n7323 ^ n441 ^ 1'b0 ;
  assign n45891 = ~n45889 & n45890 ;
  assign n45892 = n45891 ^ n25189 ^ n9390 ;
  assign n45893 = ( n2982 & n5260 ) | ( n2982 & n7569 ) | ( n5260 & n7569 ) ;
  assign n45894 = n30395 & ~n45893 ;
  assign n45895 = ~n2000 & n21808 ;
  assign n45896 = n45895 ^ x161 ^ 1'b0 ;
  assign n45897 = n18222 ^ n11819 ^ 1'b0 ;
  assign n45898 = n39163 | n45897 ;
  assign n45899 = n45896 | n45898 ;
  assign n45900 = n5485 & n9694 ;
  assign n45901 = ~n12019 & n45900 ;
  assign n45902 = n45901 ^ n33138 ^ 1'b0 ;
  assign n45903 = n9257 | n16142 ;
  assign n45904 = n45903 ^ n22166 ^ 1'b0 ;
  assign n45905 = n25018 & n45904 ;
  assign n45906 = n45902 & n45905 ;
  assign n45907 = n524 & ~n45906 ;
  assign n45908 = ~n4758 & n45907 ;
  assign n45909 = n45908 ^ n40134 ^ 1'b0 ;
  assign n45910 = n41485 ^ n20300 ^ n7506 ;
  assign n45911 = n42422 ^ n35060 ^ 1'b0 ;
  assign n45912 = n45910 | n45911 ;
  assign n45913 = n24049 & n33769 ;
  assign n45914 = n5448 & ~n45913 ;
  assign n45915 = ( n13941 & n30055 ) | ( n13941 & n32058 ) | ( n30055 & n32058 ) ;
  assign n45916 = ( n8610 & n21931 ) | ( n8610 & n36312 ) | ( n21931 & n36312 ) ;
  assign n45917 = n5965 & ~n43156 ;
  assign n45918 = n45917 ^ n18442 ^ 1'b0 ;
  assign n45919 = n36622 ^ n18034 ^ 1'b0 ;
  assign n45920 = ( n8274 & n22856 ) | ( n8274 & n45919 ) | ( n22856 & n45919 ) ;
  assign n45921 = n16839 & ~n45920 ;
  assign n45922 = n45921 ^ n23592 ^ 1'b0 ;
  assign n45923 = n20126 ^ n9375 ^ 1'b0 ;
  assign n45924 = ~n17854 & n45923 ;
  assign n45925 = n45924 ^ n22001 ^ 1'b0 ;
  assign n45926 = n3751 & n29861 ;
  assign n45927 = n45926 ^ n2791 ^ 1'b0 ;
  assign n45928 = n16884 ^ n8884 ^ 1'b0 ;
  assign n45929 = n22945 | n45928 ;
  assign n45930 = n45929 ^ x61 ^ 1'b0 ;
  assign n45931 = ~n42182 & n45066 ;
  assign n45932 = n11124 | n14992 ;
  assign n45933 = ( n19276 & n24056 ) | ( n19276 & ~n33617 ) | ( n24056 & ~n33617 ) ;
  assign n45934 = n2066 & ~n13744 ;
  assign n45935 = n39584 & n45934 ;
  assign n45936 = n21041 ^ n6260 ^ n4347 ;
  assign n45937 = n6491 ^ n4339 ^ 1'b0 ;
  assign n45938 = n7680 & ~n39603 ;
  assign n45941 = n7519 & n12927 ;
  assign n45939 = n15622 & n22182 ;
  assign n45940 = n7918 & n45939 ;
  assign n45942 = n45941 ^ n45940 ^ 1'b0 ;
  assign n45943 = n40533 ^ n16928 ^ 1'b0 ;
  assign n45944 = n25570 & ~n45943 ;
  assign n45945 = ~n5050 & n20790 ;
  assign n45946 = n45945 ^ n10940 ^ 1'b0 ;
  assign n45947 = n18714 | n45946 ;
  assign n45948 = n45947 ^ n12350 ^ 1'b0 ;
  assign n45949 = n45576 ^ n18660 ^ 1'b0 ;
  assign n45950 = n41379 & ~n45949 ;
  assign n45951 = ~n2477 & n5666 ;
  assign n45952 = ~n8301 & n13246 ;
  assign n45953 = ~n5055 & n45952 ;
  assign n45954 = n45953 ^ n42639 ^ n19099 ;
  assign n45955 = n17053 | n20625 ;
  assign n45956 = n13802 & ~n45955 ;
  assign n45957 = n45956 ^ n19027 ^ 1'b0 ;
  assign n45958 = n45957 ^ n33952 ^ n33296 ;
  assign n45959 = n45900 ^ n9518 ^ 1'b0 ;
  assign n45960 = ~n27153 & n45959 ;
  assign n45961 = n17453 ^ n4931 ^ 1'b0 ;
  assign n45962 = n38068 & n45961 ;
  assign n45963 = n45962 ^ n17118 ^ 1'b0 ;
  assign n45964 = n6749 | n43432 ;
  assign n45965 = n1400 & ~n45964 ;
  assign n45968 = ~n11564 & n12253 ;
  assign n45969 = ~n20581 & n45968 ;
  assign n45966 = n10761 & ~n35183 ;
  assign n45967 = ~n10686 & n45966 ;
  assign n45970 = n45969 ^ n45967 ^ 1'b0 ;
  assign n45971 = n3960 | n23532 ;
  assign n45972 = n19205 & ~n45971 ;
  assign n45973 = n23209 ^ n13086 ^ n4604 ;
  assign n45974 = n16147 ^ n10541 ^ 1'b0 ;
  assign n45975 = n42810 ^ n24937 ^ n8500 ;
  assign n45976 = n6975 & n39283 ;
  assign n45977 = n45976 ^ n43748 ^ 1'b0 ;
  assign n45978 = n5888 | n40974 ;
  assign n45979 = n704 & ~n45978 ;
  assign n45980 = n4182 & n14629 ;
  assign n45981 = n45980 ^ n15258 ^ 1'b0 ;
  assign n45982 = n21153 ^ n14184 ^ 1'b0 ;
  assign n45983 = n13171 | n26624 ;
  assign n45984 = n45983 ^ n9157 ^ 1'b0 ;
  assign n45989 = n20883 ^ n7387 ^ n5055 ;
  assign n45985 = n45893 ^ n13921 ^ n3051 ;
  assign n45986 = n45985 ^ n2544 ^ 1'b0 ;
  assign n45987 = n4865 & n24173 ;
  assign n45988 = n45986 & n45987 ;
  assign n45990 = n45989 ^ n45988 ^ n20426 ;
  assign n45997 = n3667 | n12744 ;
  assign n45998 = n45997 ^ n1886 ^ 1'b0 ;
  assign n45996 = n39130 ^ n7175 ^ 1'b0 ;
  assign n45992 = n36469 ^ n7465 ^ 1'b0 ;
  assign n45993 = n19639 & ~n45992 ;
  assign n45994 = n32625 & ~n45993 ;
  assign n45991 = ~n575 & n7495 ;
  assign n45995 = n45994 ^ n45991 ^ 1'b0 ;
  assign n45999 = n45998 ^ n45996 ^ n45995 ;
  assign n46004 = ~n2382 & n6683 ;
  assign n46005 = n46004 ^ n5868 ^ 1'b0 ;
  assign n46000 = n9385 & n21618 ;
  assign n46001 = n20127 & n46000 ;
  assign n46002 = n46001 ^ n8931 ^ 1'b0 ;
  assign n46003 = n46002 ^ n2281 ^ 1'b0 ;
  assign n46006 = n46005 ^ n46003 ^ n12957 ;
  assign n46007 = n34272 ^ n17207 ^ 1'b0 ;
  assign n46008 = n3183 & ~n46007 ;
  assign n46010 = ~n23760 & n27652 ;
  assign n46009 = n8823 | n12918 ;
  assign n46011 = n46010 ^ n46009 ^ 1'b0 ;
  assign n46012 = n37506 ^ n11703 ^ 1'b0 ;
  assign n46013 = ~n13363 & n28652 ;
  assign n46014 = n36424 ^ n13695 ^ 1'b0 ;
  assign n46015 = ( ~n10882 & n34851 ) | ( ~n10882 & n46014 ) | ( n34851 & n46014 ) ;
  assign n46016 = ( ~n950 & n14025 ) | ( ~n950 & n20487 ) | ( n14025 & n20487 ) ;
  assign n46017 = n8934 ^ n1800 ^ n1319 ;
  assign n46018 = n36196 & ~n46017 ;
  assign n46019 = n21309 ^ n5075 ^ 1'b0 ;
  assign n46020 = n26350 ^ n17124 ^ 1'b0 ;
  assign n46021 = n26207 ^ n16338 ^ 1'b0 ;
  assign n46022 = n10490 ^ x169 ^ 1'b0 ;
  assign n46023 = ~n34891 & n46022 ;
  assign n46024 = n4768 ^ n4177 ^ 1'b0 ;
  assign n46025 = n33633 ^ n18839 ^ 1'b0 ;
  assign n46026 = n24984 ^ n16221 ^ n9222 ;
  assign n46027 = n12266 & ~n22760 ;
  assign n46028 = n45117 ^ n21806 ^ 1'b0 ;
  assign n46029 = n10885 ^ n5558 ^ 1'b0 ;
  assign n46030 = n11906 & n46029 ;
  assign n46031 = n311 & ~n22830 ;
  assign n46032 = n46031 ^ n9614 ^ 1'b0 ;
  assign n46033 = n8961 ^ n2914 ^ 1'b0 ;
  assign n46034 = n24937 & n46033 ;
  assign n46035 = n8090 | n28976 ;
  assign n46036 = n13574 & ~n46035 ;
  assign n46037 = n1533 | n4657 ;
  assign n46038 = n13630 | n46037 ;
  assign n46039 = n29533 & ~n33556 ;
  assign n46040 = n29902 ^ n14784 ^ n751 ;
  assign n46041 = n4038 & ~n30898 ;
  assign n46042 = ~n15027 & n46041 ;
  assign n46043 = ( n20774 & ~n27584 ) | ( n20774 & n46042 ) | ( ~n27584 & n46042 ) ;
  assign n46044 = ( n6296 & n11689 ) | ( n6296 & n46043 ) | ( n11689 & n46043 ) ;
  assign n46045 = n12460 ^ n4306 ^ 1'b0 ;
  assign n46046 = n18529 & n46045 ;
  assign n46047 = n25999 ^ n24709 ^ n14528 ;
  assign n46048 = n34484 | n46047 ;
  assign n46049 = n46048 ^ n1671 ^ 1'b0 ;
  assign n46050 = n1162 | n3454 ;
  assign n46051 = n46050 ^ n5408 ^ 1'b0 ;
  assign n46052 = n1807 & ~n46051 ;
  assign n46053 = n46052 ^ n9692 ^ n9553 ;
  assign n46055 = n28426 ^ n10102 ^ 1'b0 ;
  assign n46054 = n286 | n43742 ;
  assign n46056 = n46055 ^ n46054 ^ 1'b0 ;
  assign n46057 = n12864 | n22346 ;
  assign n46058 = n5107 & ~n15197 ;
  assign n46059 = n35068 & n46058 ;
  assign n46060 = n28436 & ~n36798 ;
  assign n46061 = n25534 & n46060 ;
  assign n46062 = n18600 | n46061 ;
  assign n46063 = n44055 ^ n34379 ^ n21286 ;
  assign n46068 = n16636 ^ n14523 ^ n12332 ;
  assign n46064 = n4907 & ~n23983 ;
  assign n46065 = n46064 ^ n14450 ^ 1'b0 ;
  assign n46066 = n46065 ^ n1665 ^ 1'b0 ;
  assign n46067 = n13436 & n46066 ;
  assign n46069 = n46068 ^ n46067 ^ n10548 ;
  assign n46070 = n7608 & ~n26776 ;
  assign n46071 = n46070 ^ n8765 ^ 1'b0 ;
  assign n46072 = ~x32 & n3611 ;
  assign n46073 = n8521 & ~n46072 ;
  assign n46074 = n46073 ^ n12382 ^ 1'b0 ;
  assign n46075 = n25167 ^ n11083 ^ 1'b0 ;
  assign n46076 = n14047 ^ n12888 ^ 1'b0 ;
  assign n46077 = n29153 ^ n4661 ^ 1'b0 ;
  assign n46078 = n23436 ^ n16796 ^ n2281 ;
  assign n46079 = n860 & ~n4160 ;
  assign n46080 = ( n4857 & ~n5670 ) | ( n4857 & n46079 ) | ( ~n5670 & n46079 ) ;
  assign n46081 = ~n10073 & n32111 ;
  assign n46082 = ~n23490 & n27583 ;
  assign n46083 = n46082 ^ n17424 ^ 1'b0 ;
  assign n46084 = ( n7844 & n12091 ) | ( n7844 & ~n30236 ) | ( n12091 & ~n30236 ) ;
  assign n46085 = n46084 ^ n7322 ^ 1'b0 ;
  assign n46086 = n45351 ^ n34001 ^ n577 ;
  assign n46087 = n46086 ^ n31182 ^ 1'b0 ;
  assign n46088 = n15181 ^ n9692 ^ 1'b0 ;
  assign n46089 = n10909 | n13511 ;
  assign n46090 = n38253 & ~n46089 ;
  assign n46091 = n33076 ^ n27350 ^ 1'b0 ;
  assign n46092 = n46091 ^ n24328 ^ 1'b0 ;
  assign n46093 = n26903 ^ n9804 ^ 1'b0 ;
  assign n46094 = ~n604 & n46093 ;
  assign n46095 = ( n8672 & n35730 ) | ( n8672 & n46094 ) | ( n35730 & n46094 ) ;
  assign n46096 = n16415 ^ n10171 ^ n1683 ;
  assign n46097 = n46096 ^ n19641 ^ 1'b0 ;
  assign n46098 = n46097 ^ n36241 ^ n35883 ;
  assign n46099 = n5637 & n23554 ;
  assign n46100 = n4342 & n46099 ;
  assign n46101 = n46100 ^ n18918 ^ n9406 ;
  assign n46102 = ~n1253 & n25933 ;
  assign n46103 = ~n5798 & n46102 ;
  assign n46104 = n3089 & n46103 ;
  assign n46105 = n10968 | n46104 ;
  assign n46106 = n46105 ^ n33941 ^ 1'b0 ;
  assign n46107 = n41656 & n46106 ;
  assign n46108 = n46107 ^ n11930 ^ 1'b0 ;
  assign n46110 = ( ~n15155 & n16058 ) | ( ~n15155 & n34037 ) | ( n16058 & n34037 ) ;
  assign n46109 = n3492 | n4832 ;
  assign n46111 = n46110 ^ n46109 ^ 1'b0 ;
  assign n46112 = n8282 & n10813 ;
  assign n46113 = n15530 & n40802 ;
  assign n46114 = n274 | n15812 ;
  assign n46115 = n35490 ^ n28424 ^ 1'b0 ;
  assign n46116 = ~n46114 & n46115 ;
  assign n46117 = ( ~n21506 & n40406 ) | ( ~n21506 & n45462 ) | ( n40406 & n45462 ) ;
  assign n46118 = ~n39106 & n45501 ;
  assign n46119 = n11667 & ~n12142 ;
  assign n46120 = n46119 ^ n25661 ^ 1'b0 ;
  assign n46121 = n46120 ^ n33658 ^ 1'b0 ;
  assign n46122 = n13626 & ~n46121 ;
  assign n46123 = n3517 & ~n18568 ;
  assign n46124 = n46123 ^ n16754 ^ 1'b0 ;
  assign n46125 = n24073 | n35933 ;
  assign n46126 = n46124 & ~n46125 ;
  assign n46127 = n22915 & ~n46126 ;
  assign n46128 = n46127 ^ n38816 ^ 1'b0 ;
  assign n46129 = ( n9833 & ~n35221 ) | ( n9833 & n38207 ) | ( ~n35221 & n38207 ) ;
  assign n46130 = n46129 ^ n27754 ^ 1'b0 ;
  assign n46131 = n5185 | n15551 ;
  assign n46132 = n17782 & ~n46131 ;
  assign n46133 = n45923 ^ n7262 ^ 1'b0 ;
  assign n46134 = n11434 | n46133 ;
  assign n46135 = ( n6502 & n37587 ) | ( n6502 & n43858 ) | ( n37587 & n43858 ) ;
  assign n46136 = n8886 | n46135 ;
  assign n46137 = n9518 & ~n12909 ;
  assign n46138 = n16631 ^ n6279 ^ 1'b0 ;
  assign n46139 = n1330 | n27251 ;
  assign n46140 = n14100 & ~n35623 ;
  assign n46141 = n46140 ^ n5980 ^ 1'b0 ;
  assign n46142 = n4538 | n38608 ;
  assign n46143 = n5977 & ~n46142 ;
  assign n46144 = ( ~n2228 & n20429 ) | ( ~n2228 & n24340 ) | ( n20429 & n24340 ) ;
  assign n46145 = n1270 & ~n46144 ;
  assign n46146 = n14458 & n46145 ;
  assign n46147 = n3241 & ~n7081 ;
  assign n46148 = n46147 ^ n23626 ^ 1'b0 ;
  assign n46149 = n3808 & ~n14648 ;
  assign n46150 = n46149 ^ n8374 ^ x126 ;
  assign n46151 = n23428 ^ n17853 ^ 1'b0 ;
  assign n46152 = ~n25291 & n46151 ;
  assign n46153 = n35904 ^ n31419 ^ 1'b0 ;
  assign n46154 = n14598 & n22932 ;
  assign n46155 = n14429 | n39536 ;
  assign n46156 = n46154 & ~n46155 ;
  assign n46157 = n18529 | n19413 ;
  assign n46158 = n46157 ^ n2078 ^ 1'b0 ;
  assign n46159 = ~n2129 & n26035 ;
  assign n46160 = n46159 ^ n34891 ^ 1'b0 ;
  assign n46161 = n12451 ^ n11910 ^ n1350 ;
  assign n46162 = n30816 & n46161 ;
  assign n46163 = n3376 ^ x220 ^ 1'b0 ;
  assign n46164 = n1536 & n6648 ;
  assign n46165 = n32848 & n46164 ;
  assign n46167 = ( n298 & ~n2054 ) | ( n298 & n15721 ) | ( ~n2054 & n15721 ) ;
  assign n46168 = n21252 ^ n9379 ^ 1'b0 ;
  assign n46169 = ~n46167 & n46168 ;
  assign n46170 = n46169 ^ n21242 ^ 1'b0 ;
  assign n46166 = n21012 ^ n733 ^ 1'b0 ;
  assign n46171 = n46170 ^ n46166 ^ n36924 ;
  assign n46172 = n33680 ^ n4464 ^ n1396 ;
  assign n46173 = n24977 ^ n16660 ^ n11357 ;
  assign n46174 = n30532 ^ n536 ^ 1'b0 ;
  assign n46175 = n15134 ^ x238 ^ 1'b0 ;
  assign n46176 = n34711 & n46175 ;
  assign n46177 = ~n15244 & n46176 ;
  assign n46178 = n46177 ^ n8768 ^ 1'b0 ;
  assign n46179 = ~n7027 & n39827 ;
  assign n46180 = n28856 | n34338 ;
  assign n46181 = n13021 | n24888 ;
  assign n46182 = n17175 ^ n2748 ^ 1'b0 ;
  assign n46183 = n46181 | n46182 ;
  assign n46184 = n46183 ^ n21882 ^ 1'b0 ;
  assign n46185 = n23905 | n28388 ;
  assign n46186 = n39961 | n46185 ;
  assign n46187 = n734 & ~n36376 ;
  assign n46188 = ~n7267 & n8794 ;
  assign n46189 = n2783 & n46188 ;
  assign n46190 = ( n5903 & n31603 ) | ( n5903 & ~n46189 ) | ( n31603 & ~n46189 ) ;
  assign n46191 = ~n6655 & n19307 ;
  assign n46192 = n3973 & n46191 ;
  assign n46193 = n11939 & n46192 ;
  assign n46194 = n46193 ^ n32671 ^ n25510 ;
  assign n46195 = ~n288 & n16207 ;
  assign n46196 = n10460 & n46195 ;
  assign n46197 = n11297 & n16581 ;
  assign n46198 = n46197 ^ n20788 ^ 1'b0 ;
  assign n46199 = n13943 ^ n9421 ^ n3523 ;
  assign n46200 = ~n46198 & n46199 ;
  assign n46201 = n29251 & n46200 ;
  assign n46203 = ~n18791 & n18889 ;
  assign n46204 = n11443 ^ n4132 ^ 1'b0 ;
  assign n46205 = ~n11083 & n46204 ;
  assign n46206 = ~n46203 & n46205 ;
  assign n46202 = n10383 | n44761 ;
  assign n46207 = n46206 ^ n46202 ^ 1'b0 ;
  assign n46208 = n46207 ^ n31346 ^ 1'b0 ;
  assign n46209 = n3720 & n26203 ;
  assign n46210 = n2715 & n23485 ;
  assign n46211 = ~n46209 & n46210 ;
  assign n46212 = n24329 | n42027 ;
  assign n46213 = n46211 & ~n46212 ;
  assign n46214 = n20346 ^ n6927 ^ 1'b0 ;
  assign n46215 = n29143 & n46214 ;
  assign n46216 = n46215 ^ n15594 ^ 1'b0 ;
  assign n46217 = ~n38599 & n46216 ;
  assign n46218 = n12497 ^ n4489 ^ 1'b0 ;
  assign n46219 = ~n1401 & n46218 ;
  assign n46220 = n2024 & n6317 ;
  assign n46221 = n16203 & n46220 ;
  assign n46222 = n5107 | n41917 ;
  assign n46223 = n24979 | n46222 ;
  assign y0 = x2 ;
  assign y1 = x8 ;
  assign y2 = x9 ;
  assign y3 = x15 ;
  assign y4 = x16 ;
  assign y5 = x21 ;
  assign y6 = x24 ;
  assign y7 = x30 ;
  assign y8 = x32 ;
  assign y9 = x33 ;
  assign y10 = x34 ;
  assign y11 = x40 ;
  assign y12 = x42 ;
  assign y13 = x45 ;
  assign y14 = x54 ;
  assign y15 = x62 ;
  assign y16 = x63 ;
  assign y17 = x66 ;
  assign y18 = x75 ;
  assign y19 = x84 ;
  assign y20 = x89 ;
  assign y21 = x93 ;
  assign y22 = x99 ;
  assign y23 = x102 ;
  assign y24 = x111 ;
  assign y25 = x114 ;
  assign y26 = x115 ;
  assign y27 = x116 ;
  assign y28 = x122 ;
  assign y29 = x134 ;
  assign y30 = x139 ;
  assign y31 = x163 ;
  assign y32 = x176 ;
  assign y33 = x183 ;
  assign y34 = x190 ;
  assign y35 = x197 ;
  assign y36 = x199 ;
  assign y37 = x201 ;
  assign y38 = x205 ;
  assign y39 = x208 ;
  assign y40 = x210 ;
  assign y41 = x211 ;
  assign y42 = x213 ;
  assign y43 = x216 ;
  assign y44 = x218 ;
  assign y45 = x219 ;
  assign y46 = x222 ;
  assign y47 = x223 ;
  assign y48 = x232 ;
  assign y49 = x237 ;
  assign y50 = x238 ;
  assign y51 = x240 ;
  assign y52 = x241 ;
  assign y53 = x245 ;
  assign y54 = n256 ;
  assign y55 = ~1'b0 ;
  assign y56 = ~n258 ;
  assign y57 = n259 ;
  assign y58 = ~1'b0 ;
  assign y59 = ~1'b0 ;
  assign y60 = ~n263 ;
  assign y61 = n265 ;
  assign y62 = ~n267 ;
  assign y63 = n269 ;
  assign y64 = ~n273 ;
  assign y65 = ~1'b0 ;
  assign y66 = n275 ;
  assign y67 = n277 ;
  assign y68 = ~n279 ;
  assign y69 = n281 ;
  assign y70 = ~1'b0 ;
  assign y71 = ~n283 ;
  assign y72 = ~n286 ;
  assign y73 = ~n288 ;
  assign y74 = n289 ;
  assign y75 = ~1'b0 ;
  assign y76 = ~n291 ;
  assign y77 = ~n292 ;
  assign y78 = ~n294 ;
  assign y79 = n299 ;
  assign y80 = ~n300 ;
  assign y81 = ~n301 ;
  assign y82 = ~1'b0 ;
  assign y83 = ~n302 ;
  assign y84 = ~n304 ;
  assign y85 = ~1'b0 ;
  assign y86 = ~n305 ;
  assign y87 = ~1'b0 ;
  assign y88 = ~1'b0 ;
  assign y89 = n306 ;
  assign y90 = n307 ;
  assign y91 = n314 ;
  assign y92 = ~n315 ;
  assign y93 = ~n319 ;
  assign y94 = ~n320 ;
  assign y95 = ~1'b0 ;
  assign y96 = ~n322 ;
  assign y97 = ~n323 ;
  assign y98 = ~n328 ;
  assign y99 = ~n331 ;
  assign y100 = ~n332 ;
  assign y101 = ~n333 ;
  assign y102 = ~n335 ;
  assign y103 = n338 ;
  assign y104 = n342 ;
  assign y105 = ~n349 ;
  assign y106 = ~n351 ;
  assign y107 = ~n354 ;
  assign y108 = ~n361 ;
  assign y109 = ~n366 ;
  assign y110 = ~1'b0 ;
  assign y111 = ~n371 ;
  assign y112 = ~n377 ;
  assign y113 = ~1'b0 ;
  assign y114 = n380 ;
  assign y115 = ~n381 ;
  assign y116 = ~n393 ;
  assign y117 = n395 ;
  assign y118 = ~1'b0 ;
  assign y119 = n397 ;
  assign y120 = n399 ;
  assign y121 = ~n400 ;
  assign y122 = ~n401 ;
  assign y123 = ~1'b0 ;
  assign y124 = ~n402 ;
  assign y125 = ~n405 ;
  assign y126 = ~n409 ;
  assign y127 = n412 ;
  assign y128 = ~n415 ;
  assign y129 = ~n417 ;
  assign y130 = ~n418 ;
  assign y131 = ~n431 ;
  assign y132 = ~n432 ;
  assign y133 = n433 ;
  assign y134 = ~n434 ;
  assign y135 = ~n436 ;
  assign y136 = n441 ;
  assign y137 = n446 ;
  assign y138 = n447 ;
  assign y139 = ~n453 ;
  assign y140 = n456 ;
  assign y141 = n459 ;
  assign y142 = ~n460 ;
  assign y143 = n462 ;
  assign y144 = n463 ;
  assign y145 = ~n467 ;
  assign y146 = n469 ;
  assign y147 = ~n471 ;
  assign y148 = ~1'b0 ;
  assign y149 = n473 ;
  assign y150 = ~1'b0 ;
  assign y151 = ~1'b0 ;
  assign y152 = ~n476 ;
  assign y153 = ~n478 ;
  assign y154 = n481 ;
  assign y155 = ~1'b0 ;
  assign y156 = ~n482 ;
  assign y157 = n484 ;
  assign y158 = n485 ;
  assign y159 = n488 ;
  assign y160 = n490 ;
  assign y161 = n491 ;
  assign y162 = n500 ;
  assign y163 = ~n504 ;
  assign y164 = ~1'b0 ;
  assign y165 = n505 ;
  assign y166 = n506 ;
  assign y167 = ~1'b0 ;
  assign y168 = ~1'b0 ;
  assign y169 = ~1'b0 ;
  assign y170 = ~n509 ;
  assign y171 = ~n511 ;
  assign y172 = n518 ;
  assign y173 = ~n522 ;
  assign y174 = ~x101 ;
  assign y175 = ~1'b0 ;
  assign y176 = n524 ;
  assign y177 = n526 ;
  assign y178 = ~n527 ;
  assign y179 = ~1'b0 ;
  assign y180 = ~n529 ;
  assign y181 = ~n541 ;
  assign y182 = ~1'b0 ;
  assign y183 = n546 ;
  assign y184 = ~n548 ;
  assign y185 = ~n550 ;
  assign y186 = ~1'b0 ;
  assign y187 = x7 ;
  assign y188 = ~1'b0 ;
  assign y189 = ~n552 ;
  assign y190 = ~n556 ;
  assign y191 = n558 ;
  assign y192 = n560 ;
  assign y193 = ~n563 ;
  assign y194 = ~n567 ;
  assign y195 = n571 ;
  assign y196 = ~n572 ;
  assign y197 = ~n575 ;
  assign y198 = ~n585 ;
  assign y199 = n591 ;
  assign y200 = ~1'b0 ;
  assign y201 = ~n592 ;
  assign y202 = n597 ;
  assign y203 = ~1'b0 ;
  assign y204 = n598 ;
  assign y205 = ~n600 ;
  assign y206 = ~1'b0 ;
  assign y207 = n606 ;
  assign y208 = ~n612 ;
  assign y209 = ~n617 ;
  assign y210 = n624 ;
  assign y211 = n634 ;
  assign y212 = x167 ;
  assign y213 = n636 ;
  assign y214 = ~1'b0 ;
  assign y215 = ~n642 ;
  assign y216 = ~1'b0 ;
  assign y217 = n643 ;
  assign y218 = n646 ;
  assign y219 = ~n648 ;
  assign y220 = ~n650 ;
  assign y221 = ~n653 ;
  assign y222 = n659 ;
  assign y223 = ~n365 ;
  assign y224 = ~n663 ;
  assign y225 = ~1'b0 ;
  assign y226 = ~1'b0 ;
  assign y227 = ~n665 ;
  assign y228 = ~x15 ;
  assign y229 = n666 ;
  assign y230 = n674 ;
  assign y231 = ~1'b0 ;
  assign y232 = n677 ;
  assign y233 = ~1'b0 ;
  assign y234 = ~1'b0 ;
  assign y235 = ~n685 ;
  assign y236 = ~1'b0 ;
  assign y237 = ~n692 ;
  assign y238 = ~n694 ;
  assign y239 = ~n698 ;
  assign y240 = ~n702 ;
  assign y241 = ~n706 ;
  assign y242 = n709 ;
  assign y243 = ~n711 ;
  assign y244 = ~n713 ;
  assign y245 = ~n714 ;
  assign y246 = n716 ;
  assign y247 = ~1'b0 ;
  assign y248 = ~1'b0 ;
  assign y249 = ~n718 ;
  assign y250 = ~n645 ;
  assign y251 = ~1'b0 ;
  assign y252 = ~1'b0 ;
  assign y253 = ~1'b0 ;
  assign y254 = ~n729 ;
  assign y255 = n732 ;
  assign y256 = ~n733 ;
  assign y257 = ~n735 ;
  assign y258 = ~n745 ;
  assign y259 = n749 ;
  assign y260 = ~1'b0 ;
  assign y261 = ~n752 ;
  assign y262 = n753 ;
  assign y263 = n755 ;
  assign y264 = ~n756 ;
  assign y265 = ~n758 ;
  assign y266 = ~n764 ;
  assign y267 = ~n766 ;
  assign y268 = ~n772 ;
  assign y269 = ~n774 ;
  assign y270 = ~1'b0 ;
  assign y271 = ~n535 ;
  assign y272 = n783 ;
  assign y273 = ~n789 ;
  assign y274 = n791 ;
  assign y275 = ~n795 ;
  assign y276 = ~n797 ;
  assign y277 = ~n798 ;
  assign y278 = n803 ;
  assign y279 = ~1'b0 ;
  assign y280 = n804 ;
  assign y281 = n808 ;
  assign y282 = ~n813 ;
  assign y283 = ~1'b0 ;
  assign y284 = ~n815 ;
  assign y285 = ~n818 ;
  assign y286 = ~n822 ;
  assign y287 = n826 ;
  assign y288 = ~1'b0 ;
  assign y289 = ~n835 ;
  assign y290 = n841 ;
  assign y291 = n845 ;
  assign y292 = n854 ;
  assign y293 = ~n861 ;
  assign y294 = ~1'b0 ;
  assign y295 = ~1'b0 ;
  assign y296 = ~n867 ;
  assign y297 = ~n872 ;
  assign y298 = n874 ;
  assign y299 = ~n878 ;
  assign y300 = ~1'b0 ;
  assign y301 = 1'b0 ;
  assign y302 = ~n880 ;
  assign y303 = ~n881 ;
  assign y304 = n887 ;
  assign y305 = ~n889 ;
  assign y306 = n890 ;
  assign y307 = n894 ;
  assign y308 = ~1'b0 ;
  assign y309 = n896 ;
  assign y310 = ~1'b0 ;
  assign y311 = n897 ;
  assign y312 = ~1'b0 ;
  assign y313 = ~1'b0 ;
  assign y314 = n902 ;
  assign y315 = ~n904 ;
  assign y316 = n906 ;
  assign y317 = ~1'b0 ;
  assign y318 = ~n908 ;
  assign y319 = n918 ;
  assign y320 = n921 ;
  assign y321 = ~1'b0 ;
  assign y322 = ~n928 ;
  assign y323 = n931 ;
  assign y324 = ~n940 ;
  assign y325 = ~1'b0 ;
  assign y326 = ~n952 ;
  assign y327 = n960 ;
  assign y328 = n961 ;
  assign y329 = ~n967 ;
  assign y330 = n968 ;
  assign y331 = ~1'b0 ;
  assign y332 = n976 ;
  assign y333 = n988 ;
  assign y334 = ~n989 ;
  assign y335 = ~n991 ;
  assign y336 = n995 ;
  assign y337 = ~n998 ;
  assign y338 = n1001 ;
  assign y339 = ~n1003 ;
  assign y340 = ~n1004 ;
  assign y341 = n1006 ;
  assign y342 = ~n1007 ;
  assign y343 = n1010 ;
  assign y344 = ~n1011 ;
  assign y345 = ~1'b0 ;
  assign y346 = n1021 ;
  assign y347 = ~n1023 ;
  assign y348 = n1024 ;
  assign y349 = ~n1026 ;
  assign y350 = n1030 ;
  assign y351 = n1034 ;
  assign y352 = n1040 ;
  assign y353 = ~n1041 ;
  assign y354 = ~1'b0 ;
  assign y355 = ~1'b0 ;
  assign y356 = n1042 ;
  assign y357 = ~1'b0 ;
  assign y358 = n1044 ;
  assign y359 = n1046 ;
  assign y360 = ~n1055 ;
  assign y361 = ~1'b0 ;
  assign y362 = ~n1058 ;
  assign y363 = n1060 ;
  assign y364 = ~n1063 ;
  assign y365 = ~n1068 ;
  assign y366 = n1070 ;
  assign y367 = ~n1073 ;
  assign y368 = ~n1077 ;
  assign y369 = ~1'b0 ;
  assign y370 = ~n1086 ;
  assign y371 = n1088 ;
  assign y372 = n1090 ;
  assign y373 = n1091 ;
  assign y374 = ~1'b0 ;
  assign y375 = ~1'b0 ;
  assign y376 = ~n1099 ;
  assign y377 = ~n1101 ;
  assign y378 = ~n1103 ;
  assign y379 = ~n1111 ;
  assign y380 = n1117 ;
  assign y381 = n1119 ;
  assign y382 = ~n1124 ;
  assign y383 = ~n1126 ;
  assign y384 = ~n1127 ;
  assign y385 = ~n1132 ;
  assign y386 = ~1'b0 ;
  assign y387 = ~n1134 ;
  assign y388 = ~n1137 ;
  assign y389 = n1138 ;
  assign y390 = ~n1139 ;
  assign y391 = ~n1148 ;
  assign y392 = ~n1152 ;
  assign y393 = n1160 ;
  assign y394 = ~n1162 ;
  assign y395 = ~n1173 ;
  assign y396 = ~n1186 ;
  assign y397 = ~1'b0 ;
  assign y398 = n1187 ;
  assign y399 = ~n1188 ;
  assign y400 = ~1'b0 ;
  assign y401 = ~1'b0 ;
  assign y402 = ~n1189 ;
  assign y403 = n1195 ;
  assign y404 = ~n1199 ;
  assign y405 = n1200 ;
  assign y406 = ~1'b0 ;
  assign y407 = ~n1201 ;
  assign y408 = n1203 ;
  assign y409 = ~n1208 ;
  assign y410 = ~n1212 ;
  assign y411 = n1213 ;
  assign y412 = n1214 ;
  assign y413 = n1218 ;
  assign y414 = n1220 ;
  assign y415 = ~1'b0 ;
  assign y416 = n1223 ;
  assign y417 = ~n1227 ;
  assign y418 = n1228 ;
  assign y419 = ~n1232 ;
  assign y420 = n1234 ;
  assign y421 = n1235 ;
  assign y422 = ~1'b0 ;
  assign y423 = ~1'b0 ;
  assign y424 = ~n1241 ;
  assign y425 = n1246 ;
  assign y426 = n1249 ;
  assign y427 = ~1'b0 ;
  assign y428 = ~n1255 ;
  assign y429 = n1256 ;
  assign y430 = ~n1264 ;
  assign y431 = n1265 ;
  assign y432 = ~1'b0 ;
  assign y433 = ~1'b0 ;
  assign y434 = ~1'b0 ;
  assign y435 = n1266 ;
  assign y436 = ~1'b0 ;
  assign y437 = n1270 ;
  assign y438 = ~n1271 ;
  assign y439 = ~1'b0 ;
  assign y440 = ~n1272 ;
  assign y441 = n1273 ;
  assign y442 = ~n1274 ;
  assign y443 = ~n1277 ;
  assign y444 = ~n1278 ;
  assign y445 = n1286 ;
  assign y446 = ~n1293 ;
  assign y447 = n1296 ;
  assign y448 = n1298 ;
  assign y449 = ~n1302 ;
  assign y450 = ~n1304 ;
  assign y451 = ~1'b0 ;
  assign y452 = n1010 ;
  assign y453 = ~n1308 ;
  assign y454 = n1310 ;
  assign y455 = ~n1313 ;
  assign y456 = ~1'b0 ;
  assign y457 = ~n1314 ;
  assign y458 = n405 ;
  assign y459 = ~1'b0 ;
  assign y460 = n1315 ;
  assign y461 = ~1'b0 ;
  assign y462 = ~n1321 ;
  assign y463 = ~n1325 ;
  assign y464 = ~1'b0 ;
  assign y465 = n1328 ;
  assign y466 = n1334 ;
  assign y467 = ~n1339 ;
  assign y468 = ~1'b0 ;
  assign y469 = n1348 ;
  assign y470 = n1349 ;
  assign y471 = ~1'b0 ;
  assign y472 = ~n1350 ;
  assign y473 = ~n1353 ;
  assign y474 = ~n634 ;
  assign y475 = ~n1356 ;
  assign y476 = n1362 ;
  assign y477 = ~n1365 ;
  assign y478 = ~n1368 ;
  assign y479 = ~n1370 ;
  assign y480 = ~n1373 ;
  assign y481 = ~n1378 ;
  assign y482 = n1380 ;
  assign y483 = ~n1381 ;
  assign y484 = ~n1384 ;
  assign y485 = n1386 ;
  assign y486 = n1388 ;
  assign y487 = ~n1390 ;
  assign y488 = n1392 ;
  assign y489 = ~1'b0 ;
  assign y490 = ~n1394 ;
  assign y491 = ~n1395 ;
  assign y492 = ~n1397 ;
  assign y493 = n1403 ;
  assign y494 = ~1'b0 ;
  assign y495 = ~n1411 ;
  assign y496 = ~n1425 ;
  assign y497 = ~1'b0 ;
  assign y498 = ~n1430 ;
  assign y499 = n1432 ;
  assign y500 = n1435 ;
  assign y501 = 1'b0 ;
  assign y502 = x83 ;
  assign y503 = ~n1442 ;
  assign y504 = ~n1444 ;
  assign y505 = ~n1451 ;
  assign y506 = ~1'b0 ;
  assign y507 = ~1'b0 ;
  assign y508 = ~1'b0 ;
  assign y509 = n1457 ;
  assign y510 = ~n1460 ;
  assign y511 = n1462 ;
  assign y512 = ~1'b0 ;
  assign y513 = ~1'b0 ;
  assign y514 = n1469 ;
  assign y515 = n1470 ;
  assign y516 = ~n593 ;
  assign y517 = n1471 ;
  assign y518 = ~1'b0 ;
  assign y519 = ~n1472 ;
  assign y520 = ~1'b0 ;
  assign y521 = ~n1480 ;
  assign y522 = n1484 ;
  assign y523 = ~n1488 ;
  assign y524 = ~1'b0 ;
  assign y525 = n1489 ;
  assign y526 = ~n432 ;
  assign y527 = ~n1493 ;
  assign y528 = n1499 ;
  assign y529 = n1509 ;
  assign y530 = ~n1515 ;
  assign y531 = n1518 ;
  assign y532 = n1519 ;
  assign y533 = ~1'b0 ;
  assign y534 = ~1'b0 ;
  assign y535 = ~1'b0 ;
  assign y536 = ~n1520 ;
  assign y537 = ~n1521 ;
  assign y538 = ~1'b0 ;
  assign y539 = ~1'b0 ;
  assign y540 = n1525 ;
  assign y541 = ~1'b0 ;
  assign y542 = n1528 ;
  assign y543 = ~n1530 ;
  assign y544 = ~n1532 ;
  assign y545 = ~n1533 ;
  assign y546 = ~1'b0 ;
  assign y547 = n1535 ;
  assign y548 = ~1'b0 ;
  assign y549 = ~1'b0 ;
  assign y550 = ~n1538 ;
  assign y551 = n1540 ;
  assign y552 = ~1'b0 ;
  assign y553 = ~n1546 ;
  assign y554 = n1547 ;
  assign y555 = ~n1553 ;
  assign y556 = n1557 ;
  assign y557 = ~n1561 ;
  assign y558 = ~n1563 ;
  assign y559 = ~n1564 ;
  assign y560 = n1565 ;
  assign y561 = n1567 ;
  assign y562 = n1587 ;
  assign y563 = ~n1595 ;
  assign y564 = ~1'b0 ;
  assign y565 = n1597 ;
  assign y566 = ~n1600 ;
  assign y567 = ~n1604 ;
  assign y568 = ~1'b0 ;
  assign y569 = ~1'b0 ;
  assign y570 = ~n1611 ;
  assign y571 = n1612 ;
  assign y572 = n395 ;
  assign y573 = ~n1613 ;
  assign y574 = n1618 ;
  assign y575 = n1619 ;
  assign y576 = n1626 ;
  assign y577 = ~1'b0 ;
  assign y578 = ~n1630 ;
  assign y579 = ~n1635 ;
  assign y580 = n1643 ;
  assign y581 = ~1'b0 ;
  assign y582 = ~n1646 ;
  assign y583 = ~n1648 ;
  assign y584 = n1651 ;
  assign y585 = ~1'b0 ;
  assign y586 = ~n1657 ;
  assign y587 = ~n1658 ;
  assign y588 = ~n1663 ;
  assign y589 = n1669 ;
  assign y590 = ~1'b0 ;
  assign y591 = ~x241 ;
  assign y592 = ~1'b0 ;
  assign y593 = ~n1673 ;
  assign y594 = n1679 ;
  assign y595 = n1688 ;
  assign y596 = n1690 ;
  assign y597 = ~n1693 ;
  assign y598 = ~n1694 ;
  assign y599 = ~1'b0 ;
  assign y600 = ~1'b0 ;
  assign y601 = ~n1695 ;
  assign y602 = n1701 ;
  assign y603 = ~n1703 ;
  assign y604 = ~n1706 ;
  assign y605 = ~n1713 ;
  assign y606 = ~1'b0 ;
  assign y607 = ~n1719 ;
  assign y608 = ~1'b0 ;
  assign y609 = ~1'b0 ;
  assign y610 = ~n1720 ;
  assign y611 = ~n1724 ;
  assign y612 = n1725 ;
  assign y613 = n1727 ;
  assign y614 = ~n1729 ;
  assign y615 = ~1'b0 ;
  assign y616 = n1730 ;
  assign y617 = n1731 ;
  assign y618 = ~x247 ;
  assign y619 = ~1'b0 ;
  assign y620 = n1733 ;
  assign y621 = ~1'b0 ;
  assign y622 = n1737 ;
  assign y623 = ~1'b0 ;
  assign y624 = n1233 ;
  assign y625 = ~1'b0 ;
  assign y626 = n1741 ;
  assign y627 = ~1'b0 ;
  assign y628 = n1742 ;
  assign y629 = ~n1744 ;
  assign y630 = n1746 ;
  assign y631 = ~1'b0 ;
  assign y632 = n1748 ;
  assign y633 = x22 ;
  assign y634 = ~n1757 ;
  assign y635 = n1758 ;
  assign y636 = n271 ;
  assign y637 = ~n1762 ;
  assign y638 = ~n1763 ;
  assign y639 = x121 ;
  assign y640 = n1764 ;
  assign y641 = n1775 ;
  assign y642 = n1776 ;
  assign y643 = ~n1777 ;
  assign y644 = ~1'b0 ;
  assign y645 = ~n1781 ;
  assign y646 = ~n1788 ;
  assign y647 = n1792 ;
  assign y648 = n1798 ;
  assign y649 = ~1'b0 ;
  assign y650 = ~n1804 ;
  assign y651 = ~n1805 ;
  assign y652 = ~n1806 ;
  assign y653 = n1807 ;
  assign y654 = ~1'b0 ;
  assign y655 = ~1'b0 ;
  assign y656 = ~n1816 ;
  assign y657 = ~n1819 ;
  assign y658 = n1826 ;
  assign y659 = n1827 ;
  assign y660 = ~n1830 ;
  assign y661 = n1831 ;
  assign y662 = n1835 ;
  assign y663 = ~n1836 ;
  assign y664 = n1838 ;
  assign y665 = n1843 ;
  assign y666 = ~1'b0 ;
  assign y667 = ~n1213 ;
  assign y668 = ~n1851 ;
  assign y669 = ~n1853 ;
  assign y670 = ~1'b0 ;
  assign y671 = ~1'b0 ;
  assign y672 = ~1'b0 ;
  assign y673 = ~1'b0 ;
  assign y674 = ~1'b0 ;
  assign y675 = n1855 ;
  assign y676 = n1860 ;
  assign y677 = ~1'b0 ;
  assign y678 = ~1'b0 ;
  assign y679 = ~n1863 ;
  assign y680 = n1866 ;
  assign y681 = ~1'b0 ;
  assign y682 = n791 ;
  assign y683 = n1868 ;
  assign y684 = ~1'b0 ;
  assign y685 = n1871 ;
  assign y686 = ~n1873 ;
  assign y687 = 1'b0 ;
  assign y688 = ~n1876 ;
  assign y689 = ~n1877 ;
  assign y690 = ~n1880 ;
  assign y691 = n1881 ;
  assign y692 = n1886 ;
  assign y693 = n1895 ;
  assign y694 = ~n1902 ;
  assign y695 = n1904 ;
  assign y696 = ~1'b0 ;
  assign y697 = ~n1907 ;
  assign y698 = n559 ;
  assign y699 = ~n1909 ;
  assign y700 = n1913 ;
  assign y701 = n1914 ;
  assign y702 = ~n1920 ;
  assign y703 = ~1'b0 ;
  assign y704 = n1926 ;
  assign y705 = n1935 ;
  assign y706 = ~1'b0 ;
  assign y707 = ~n793 ;
  assign y708 = ~1'b0 ;
  assign y709 = n1952 ;
  assign y710 = n1953 ;
  assign y711 = ~1'b0 ;
  assign y712 = ~1'b0 ;
  assign y713 = ~1'b0 ;
  assign y714 = n1955 ;
  assign y715 = ~n1960 ;
  assign y716 = n1963 ;
  assign y717 = ~1'b0 ;
  assign y718 = ~n1967 ;
  assign y719 = n1970 ;
  assign y720 = ~n1979 ;
  assign y721 = ~n1980 ;
  assign y722 = ~n1982 ;
  assign y723 = n1983 ;
  assign y724 = ~n1985 ;
  assign y725 = ~1'b0 ;
  assign y726 = n1995 ;
  assign y727 = n1999 ;
  assign y728 = n269 ;
  assign y729 = ~n1777 ;
  assign y730 = ~n2002 ;
  assign y731 = n2004 ;
  assign y732 = ~n2005 ;
  assign y733 = ~1'b0 ;
  assign y734 = ~n2008 ;
  assign y735 = ~n2010 ;
  assign y736 = ~1'b0 ;
  assign y737 = n2011 ;
  assign y738 = n2014 ;
  assign y739 = ~1'b0 ;
  assign y740 = ~n2015 ;
  assign y741 = ~1'b0 ;
  assign y742 = ~1'b0 ;
  assign y743 = ~1'b0 ;
  assign y744 = n2017 ;
  assign y745 = ~n2019 ;
  assign y746 = n2022 ;
  assign y747 = ~n1500 ;
  assign y748 = n2028 ;
  assign y749 = n2031 ;
  assign y750 = ~n2036 ;
  assign y751 = ~n2038 ;
  assign y752 = ~1'b0 ;
  assign y753 = n369 ;
  assign y754 = n2048 ;
  assign y755 = ~1'b0 ;
  assign y756 = ~n2051 ;
  assign y757 = n2053 ;
  assign y758 = n1255 ;
  assign y759 = ~n2055 ;
  assign y760 = n2057 ;
  assign y761 = 1'b0 ;
  assign y762 = ~n2064 ;
  assign y763 = ~n2065 ;
  assign y764 = ~1'b0 ;
  assign y765 = ~n2067 ;
  assign y766 = ~n2068 ;
  assign y767 = ~1'b0 ;
  assign y768 = ~n2070 ;
  assign y769 = ~n2074 ;
  assign y770 = n2075 ;
  assign y771 = ~n2076 ;
  assign y772 = n2082 ;
  assign y773 = ~n2087 ;
  assign y774 = ~1'b0 ;
  assign y775 = ~n2089 ;
  assign y776 = ~1'b0 ;
  assign y777 = n2091 ;
  assign y778 = ~n2095 ;
  assign y779 = ~1'b0 ;
  assign y780 = ~n2097 ;
  assign y781 = ~n2098 ;
  assign y782 = ~1'b0 ;
  assign y783 = ~n2099 ;
  assign y784 = ~1'b0 ;
  assign y785 = ~n2106 ;
  assign y786 = n2109 ;
  assign y787 = n2122 ;
  assign y788 = ~n2125 ;
  assign y789 = ~1'b0 ;
  assign y790 = ~n2129 ;
  assign y791 = ~1'b0 ;
  assign y792 = ~n2134 ;
  assign y793 = n2135 ;
  assign y794 = ~n2138 ;
  assign y795 = ~1'b0 ;
  assign y796 = n2140 ;
  assign y797 = n2141 ;
  assign y798 = ~n2148 ;
  assign y799 = ~n2149 ;
  assign y800 = n2151 ;
  assign y801 = n2153 ;
  assign y802 = ~n2158 ;
  assign y803 = ~n2161 ;
  assign y804 = ~1'b0 ;
  assign y805 = ~n2162 ;
  assign y806 = n2164 ;
  assign y807 = ~n2165 ;
  assign y808 = n1233 ;
  assign y809 = n2166 ;
  assign y810 = ~1'b0 ;
  assign y811 = ~n1851 ;
  assign y812 = ~n2171 ;
  assign y813 = n2173 ;
  assign y814 = 1'b0 ;
  assign y815 = n2178 ;
  assign y816 = ~1'b0 ;
  assign y817 = ~n2182 ;
  assign y818 = n2188 ;
  assign y819 = ~1'b0 ;
  assign y820 = ~1'b0 ;
  assign y821 = ~n2195 ;
  assign y822 = ~n2199 ;
  assign y823 = ~1'b0 ;
  assign y824 = ~n2203 ;
  assign y825 = ~n2214 ;
  assign y826 = n2217 ;
  assign y827 = n2221 ;
  assign y828 = n2224 ;
  assign y829 = n2225 ;
  assign y830 = ~n2231 ;
  assign y831 = ~1'b0 ;
  assign y832 = ~n2232 ;
  assign y833 = ~n2239 ;
  assign y834 = n2243 ;
  assign y835 = ~1'b0 ;
  assign y836 = n2244 ;
  assign y837 = ~n2246 ;
  assign y838 = 1'b0 ;
  assign y839 = ~n2247 ;
  assign y840 = n2250 ;
  assign y841 = n2252 ;
  assign y842 = ~n2266 ;
  assign y843 = ~n2267 ;
  assign y844 = ~n2274 ;
  assign y845 = ~n2275 ;
  assign y846 = ~n2277 ;
  assign y847 = x114 ;
  assign y848 = n2278 ;
  assign y849 = n2285 ;
  assign y850 = ~n2286 ;
  assign y851 = ~n2293 ;
  assign y852 = n2294 ;
  assign y853 = n2300 ;
  assign y854 = ~1'b0 ;
  assign y855 = n2302 ;
  assign y856 = ~1'b0 ;
  assign y857 = n2306 ;
  assign y858 = ~1'b0 ;
  assign y859 = ~n2307 ;
  assign y860 = n2309 ;
  assign y861 = ~n677 ;
  assign y862 = ~1'b0 ;
  assign y863 = n2311 ;
  assign y864 = n2313 ;
  assign y865 = n2314 ;
  assign y866 = n2317 ;
  assign y867 = n2318 ;
  assign y868 = n2326 ;
  assign y869 = ~n2338 ;
  assign y870 = ~n2342 ;
  assign y871 = ~n2345 ;
  assign y872 = ~n2349 ;
  assign y873 = n2353 ;
  assign y874 = ~1'b0 ;
  assign y875 = ~n2354 ;
  assign y876 = ~1'b0 ;
  assign y877 = n2355 ;
  assign y878 = n2357 ;
  assign y879 = n2358 ;
  assign y880 = n2359 ;
  assign y881 = ~n2360 ;
  assign y882 = ~1'b0 ;
  assign y883 = ~n2365 ;
  assign y884 = ~n2369 ;
  assign y885 = n2371 ;
  assign y886 = ~n2374 ;
  assign y887 = ~n2386 ;
  assign y888 = ~1'b0 ;
  assign y889 = ~n2389 ;
  assign y890 = n2390 ;
  assign y891 = n2394 ;
  assign y892 = ~n2395 ;
  assign y893 = n2397 ;
  assign y894 = ~n2401 ;
  assign y895 = ~n2406 ;
  assign y896 = ~n2407 ;
  assign y897 = ~n2409 ;
  assign y898 = ~1'b0 ;
  assign y899 = ~n781 ;
  assign y900 = ~1'b0 ;
  assign y901 = n1767 ;
  assign y902 = ~n2411 ;
  assign y903 = ~1'b0 ;
  assign y904 = n2413 ;
  assign y905 = ~1'b0 ;
  assign y906 = ~1'b0 ;
  assign y907 = ~n2414 ;
  assign y908 = ~1'b0 ;
  assign y909 = n2416 ;
  assign y910 = n2421 ;
  assign y911 = ~n2422 ;
  assign y912 = ~1'b0 ;
  assign y913 = ~n2425 ;
  assign y914 = ~n2430 ;
  assign y915 = ~n2433 ;
  assign y916 = ~n2438 ;
  assign y917 = 1'b0 ;
  assign y918 = ~n1073 ;
  assign y919 = ~n2440 ;
  assign y920 = ~n2441 ;
  assign y921 = n2442 ;
  assign y922 = n2444 ;
  assign y923 = n2449 ;
  assign y924 = ~n2450 ;
  assign y925 = ~n2452 ;
  assign y926 = ~n2454 ;
  assign y927 = n2459 ;
  assign y928 = ~1'b0 ;
  assign y929 = ~n2462 ;
  assign y930 = ~n2468 ;
  assign y931 = ~n2469 ;
  assign y932 = ~1'b0 ;
  assign y933 = n2470 ;
  assign y934 = ~n2473 ;
  assign y935 = ~n2475 ;
  assign y936 = ~n2476 ;
  assign y937 = n2489 ;
  assign y938 = n2490 ;
  assign y939 = ~n2493 ;
  assign y940 = ~1'b0 ;
  assign y941 = ~1'b0 ;
  assign y942 = ~n2495 ;
  assign y943 = ~1'b0 ;
  assign y944 = ~n2504 ;
  assign y945 = ~n2506 ;
  assign y946 = 1'b0 ;
  assign y947 = ~n2507 ;
  assign y948 = ~n2511 ;
  assign y949 = n2521 ;
  assign y950 = n2529 ;
  assign y951 = n2532 ;
  assign y952 = ~1'b0 ;
  assign y953 = n2534 ;
  assign y954 = n2536 ;
  assign y955 = ~1'b0 ;
  assign y956 = ~n2537 ;
  assign y957 = ~1'b0 ;
  assign y958 = ~n2538 ;
  assign y959 = ~1'b0 ;
  assign y960 = n2539 ;
  assign y961 = n2542 ;
  assign y962 = ~1'b0 ;
  assign y963 = n835 ;
  assign y964 = ~1'b0 ;
  assign y965 = ~1'b0 ;
  assign y966 = n2546 ;
  assign y967 = ~n2550 ;
  assign y968 = n2553 ;
  assign y969 = ~1'b0 ;
  assign y970 = ~n2057 ;
  assign y971 = n2556 ;
  assign y972 = ~n2561 ;
  assign y973 = ~n2564 ;
  assign y974 = ~1'b0 ;
  assign y975 = ~1'b0 ;
  assign y976 = ~n2566 ;
  assign y977 = n2567 ;
  assign y978 = ~n2571 ;
  assign y979 = ~1'b0 ;
  assign y980 = ~n2577 ;
  assign y981 = n2585 ;
  assign y982 = ~n2590 ;
  assign y983 = n2596 ;
  assign y984 = ~1'b0 ;
  assign y985 = n2603 ;
  assign y986 = ~n2610 ;
  assign y987 = ~1'b0 ;
  assign y988 = ~n2613 ;
  assign y989 = 1'b0 ;
  assign y990 = ~n2614 ;
  assign y991 = ~n2615 ;
  assign y992 = ~n2617 ;
  assign y993 = n2618 ;
  assign y994 = ~1'b0 ;
  assign y995 = ~1'b0 ;
  assign y996 = n2621 ;
  assign y997 = n2635 ;
  assign y998 = ~n2637 ;
  assign y999 = ~n2641 ;
  assign y1000 = ~n2644 ;
  assign y1001 = ~1'b0 ;
  assign y1002 = ~n2645 ;
  assign y1003 = ~n1762 ;
  assign y1004 = ~n2648 ;
  assign y1005 = ~n2650 ;
  assign y1006 = n2651 ;
  assign y1007 = ~1'b0 ;
  assign y1008 = ~1'b0 ;
  assign y1009 = ~n2652 ;
  assign y1010 = ~1'b0 ;
  assign y1011 = ~n2653 ;
  assign y1012 = n2654 ;
  assign y1013 = ~1'b0 ;
  assign y1014 = ~1'b0 ;
  assign y1015 = ~1'b0 ;
  assign y1016 = ~n2656 ;
  assign y1017 = ~1'b0 ;
  assign y1018 = n2658 ;
  assign y1019 = ~n2663 ;
  assign y1020 = ~x3 ;
  assign y1021 = n2670 ;
  assign y1022 = n2675 ;
  assign y1023 = n2678 ;
  assign y1024 = n2684 ;
  assign y1025 = ~1'b0 ;
  assign y1026 = ~n2688 ;
  assign y1027 = n2692 ;
  assign y1028 = ~n2696 ;
  assign y1029 = ~1'b0 ;
  assign y1030 = ~1'b0 ;
  assign y1031 = n2703 ;
  assign y1032 = ~n2704 ;
  assign y1033 = n2707 ;
  assign y1034 = ~n2712 ;
  assign y1035 = ~1'b0 ;
  assign y1036 = n2713 ;
  assign y1037 = ~1'b0 ;
  assign y1038 = ~n2714 ;
  assign y1039 = n2725 ;
  assign y1040 = ~1'b0 ;
  assign y1041 = ~n2727 ;
  assign y1042 = n2738 ;
  assign y1043 = ~1'b0 ;
  assign y1044 = n1000 ;
  assign y1045 = n2743 ;
  assign y1046 = ~n2752 ;
  assign y1047 = ~n2755 ;
  assign y1048 = n2756 ;
  assign y1049 = ~n514 ;
  assign y1050 = ~1'b0 ;
  assign y1051 = ~1'b0 ;
  assign y1052 = n2757 ;
  assign y1053 = ~n2761 ;
  assign y1054 = ~1'b0 ;
  assign y1055 = n2766 ;
  assign y1056 = n2774 ;
  assign y1057 = ~n2775 ;
  assign y1058 = n2778 ;
  assign y1059 = n2780 ;
  assign y1060 = ~n2783 ;
  assign y1061 = n2786 ;
  assign y1062 = ~n2787 ;
  assign y1063 = ~n2791 ;
  assign y1064 = ~1'b0 ;
  assign y1065 = n806 ;
  assign y1066 = n2796 ;
  assign y1067 = ~1'b0 ;
  assign y1068 = ~n2799 ;
  assign y1069 = ~n2800 ;
  assign y1070 = n2802 ;
  assign y1071 = ~1'b0 ;
  assign y1072 = ~n2806 ;
  assign y1073 = ~n2808 ;
  assign y1074 = ~n2810 ;
  assign y1075 = ~n2812 ;
  assign y1076 = ~n2817 ;
  assign y1077 = ~1'b0 ;
  assign y1078 = n2819 ;
  assign y1079 = ~n2826 ;
  assign y1080 = ~1'b0 ;
  assign y1081 = ~1'b0 ;
  assign y1082 = ~n2833 ;
  assign y1083 = n2841 ;
  assign y1084 = ~n2846 ;
  assign y1085 = 1'b0 ;
  assign y1086 = n2850 ;
  assign y1087 = n2853 ;
  assign y1088 = n2854 ;
  assign y1089 = ~n2860 ;
  assign y1090 = ~n2868 ;
  assign y1091 = ~n2873 ;
  assign y1092 = ~1'b0 ;
  assign y1093 = ~1'b0 ;
  assign y1094 = ~n2881 ;
  assign y1095 = n2882 ;
  assign y1096 = n538 ;
  assign y1097 = ~n2883 ;
  assign y1098 = n2884 ;
  assign y1099 = n2890 ;
  assign y1100 = ~n2892 ;
  assign y1101 = n2893 ;
  assign y1102 = n1155 ;
  assign y1103 = n2895 ;
  assign y1104 = n2897 ;
  assign y1105 = n2898 ;
  assign y1106 = n706 ;
  assign y1107 = n2899 ;
  assign y1108 = ~n2900 ;
  assign y1109 = ~1'b0 ;
  assign y1110 = ~1'b0 ;
  assign y1111 = ~n2081 ;
  assign y1112 = ~n2903 ;
  assign y1113 = n2907 ;
  assign y1114 = ~n2910 ;
  assign y1115 = ~n2916 ;
  assign y1116 = n2922 ;
  assign y1117 = n2925 ;
  assign y1118 = n2927 ;
  assign y1119 = ~n2932 ;
  assign y1120 = ~1'b0 ;
  assign y1121 = n2936 ;
  assign y1122 = ~1'b0 ;
  assign y1123 = n2937 ;
  assign y1124 = ~n2942 ;
  assign y1125 = ~n2946 ;
  assign y1126 = ~n2947 ;
  assign y1127 = ~n2952 ;
  assign y1128 = ~n2953 ;
  assign y1129 = ~1'b0 ;
  assign y1130 = n2957 ;
  assign y1131 = ~n2961 ;
  assign y1132 = ~n2968 ;
  assign y1133 = n2971 ;
  assign y1134 = ~n2973 ;
  assign y1135 = ~1'b0 ;
  assign y1136 = n2976 ;
  assign y1137 = n2982 ;
  assign y1138 = ~n2983 ;
  assign y1139 = n2984 ;
  assign y1140 = ~1'b0 ;
  assign y1141 = n2990 ;
  assign y1142 = n2993 ;
  assign y1143 = ~1'b0 ;
  assign y1144 = ~n2995 ;
  assign y1145 = ~n833 ;
  assign y1146 = n2996 ;
  assign y1147 = ~1'b0 ;
  assign y1148 = ~n2998 ;
  assign y1149 = ~n3001 ;
  assign y1150 = ~n3002 ;
  assign y1151 = ~n3005 ;
  assign y1152 = ~1'b0 ;
  assign y1153 = ~n3011 ;
  assign y1154 = ~1'b0 ;
  assign y1155 = ~n3029 ;
  assign y1156 = ~n3035 ;
  assign y1157 = ~1'b0 ;
  assign y1158 = ~1'b0 ;
  assign y1159 = ~n3040 ;
  assign y1160 = n3045 ;
  assign y1161 = ~n3048 ;
  assign y1162 = ~n3050 ;
  assign y1163 = ~n3051 ;
  assign y1164 = ~1'b0 ;
  assign y1165 = ~1'b0 ;
  assign y1166 = ~n1253 ;
  assign y1167 = n3052 ;
  assign y1168 = 1'b0 ;
  assign y1169 = n3056 ;
  assign y1170 = ~n3058 ;
  assign y1171 = ~1'b0 ;
  assign y1172 = ~n758 ;
  assign y1173 = n3060 ;
  assign y1174 = n3062 ;
  assign y1175 = n3064 ;
  assign y1176 = ~1'b0 ;
  assign y1177 = ~1'b0 ;
  assign y1178 = n3067 ;
  assign y1179 = n3068 ;
  assign y1180 = ~n3071 ;
  assign y1181 = n3074 ;
  assign y1182 = ~n2661 ;
  assign y1183 = ~n3078 ;
  assign y1184 = ~n3084 ;
  assign y1185 = ~n3085 ;
  assign y1186 = ~n3087 ;
  assign y1187 = n3090 ;
  assign y1188 = n3091 ;
  assign y1189 = ~n3093 ;
  assign y1190 = ~n3095 ;
  assign y1191 = ~x17 ;
  assign y1192 = ~n3100 ;
  assign y1193 = ~1'b0 ;
  assign y1194 = ~1'b0 ;
  assign y1195 = ~n3104 ;
  assign y1196 = ~1'b0 ;
  assign y1197 = 1'b0 ;
  assign y1198 = n3106 ;
  assign y1199 = ~n3109 ;
  assign y1200 = ~1'b0 ;
  assign y1201 = n2108 ;
  assign y1202 = n3111 ;
  assign y1203 = n3112 ;
  assign y1204 = n3115 ;
  assign y1205 = n3116 ;
  assign y1206 = ~1'b0 ;
  assign y1207 = ~n2547 ;
  assign y1208 = ~1'b0 ;
  assign y1209 = ~1'b0 ;
  assign y1210 = n2680 ;
  assign y1211 = n3120 ;
  assign y1212 = n3121 ;
  assign y1213 = ~n3124 ;
  assign y1214 = n3129 ;
  assign y1215 = ~n3133 ;
  assign y1216 = n3134 ;
  assign y1217 = ~n1930 ;
  assign y1218 = ~n3141 ;
  assign y1219 = n3145 ;
  assign y1220 = ~n3153 ;
  assign y1221 = ~n3156 ;
  assign y1222 = n3158 ;
  assign y1223 = ~n3163 ;
  assign y1224 = ~n3164 ;
  assign y1225 = ~n3171 ;
  assign y1226 = ~1'b0 ;
  assign y1227 = n3176 ;
  assign y1228 = n3180 ;
  assign y1229 = n3187 ;
  assign y1230 = ~1'b0 ;
  assign y1231 = n3196 ;
  assign y1232 = ~n3199 ;
  assign y1233 = ~1'b0 ;
  assign y1234 = ~n3201 ;
  assign y1235 = n3203 ;
  assign y1236 = ~n3204 ;
  assign y1237 = ~n3207 ;
  assign y1238 = n3210 ;
  assign y1239 = n3213 ;
  assign y1240 = ~n3223 ;
  assign y1241 = n1225 ;
  assign y1242 = ~n2885 ;
  assign y1243 = ~n1571 ;
  assign y1244 = ~n1486 ;
  assign y1245 = n3230 ;
  assign y1246 = ~n3233 ;
  assign y1247 = n3235 ;
  assign y1248 = ~1'b0 ;
  assign y1249 = ~1'b0 ;
  assign y1250 = n3237 ;
  assign y1251 = ~n3240 ;
  assign y1252 = ~1'b0 ;
  assign y1253 = ~n3241 ;
  assign y1254 = n3249 ;
  assign y1255 = ~1'b0 ;
  assign y1256 = n3255 ;
  assign y1257 = ~1'b0 ;
  assign y1258 = ~n3256 ;
  assign y1259 = ~n3264 ;
  assign y1260 = ~1'b0 ;
  assign y1261 = n3265 ;
  assign y1262 = n3267 ;
  assign y1263 = n3272 ;
  assign y1264 = ~1'b0 ;
  assign y1265 = n3273 ;
  assign y1266 = n3274 ;
  assign y1267 = ~n3282 ;
  assign y1268 = n3289 ;
  assign y1269 = n3292 ;
  assign y1270 = ~n3294 ;
  assign y1271 = ~1'b0 ;
  assign y1272 = ~n3296 ;
  assign y1273 = n3297 ;
  assign y1274 = 1'b0 ;
  assign y1275 = n3302 ;
  assign y1276 = ~n3306 ;
  assign y1277 = ~1'b0 ;
  assign y1278 = ~n3308 ;
  assign y1279 = ~n3312 ;
  assign y1280 = n3313 ;
  assign y1281 = n3317 ;
  assign y1282 = ~n3318 ;
  assign y1283 = n3322 ;
  assign y1284 = ~n3324 ;
  assign y1285 = n3325 ;
  assign y1286 = ~n3326 ;
  assign y1287 = n3332 ;
  assign y1288 = ~n3334 ;
  assign y1289 = ~n3340 ;
  assign y1290 = ~1'b0 ;
  assign y1291 = ~n3342 ;
  assign y1292 = n3344 ;
  assign y1293 = ~n3348 ;
  assign y1294 = n3352 ;
  assign y1295 = ~n3354 ;
  assign y1296 = ~1'b0 ;
  assign y1297 = ~n3362 ;
  assign y1298 = ~n3366 ;
  assign y1299 = n3367 ;
  assign y1300 = ~n3369 ;
  assign y1301 = n3376 ;
  assign y1302 = ~1'b0 ;
  assign y1303 = n3378 ;
  assign y1304 = n3381 ;
  assign y1305 = ~n3382 ;
  assign y1306 = ~n3383 ;
  assign y1307 = ~n3391 ;
  assign y1308 = n3393 ;
  assign y1309 = n3394 ;
  assign y1310 = ~1'b0 ;
  assign y1311 = ~n3398 ;
  assign y1312 = n3401 ;
  assign y1313 = n3405 ;
  assign y1314 = ~1'b0 ;
  assign y1315 = n3410 ;
  assign y1316 = n3415 ;
  assign y1317 = n3421 ;
  assign y1318 = ~1'b0 ;
  assign y1319 = ~1'b0 ;
  assign y1320 = ~n3422 ;
  assign y1321 = ~1'b0 ;
  assign y1322 = n3423 ;
  assign y1323 = ~1'b0 ;
  assign y1324 = ~1'b0 ;
  assign y1325 = ~n3431 ;
  assign y1326 = ~n3433 ;
  assign y1327 = ~1'b0 ;
  assign y1328 = n3439 ;
  assign y1329 = n3443 ;
  assign y1330 = n3445 ;
  assign y1331 = n3447 ;
  assign y1332 = n3450 ;
  assign y1333 = ~n3451 ;
  assign y1334 = n3453 ;
  assign y1335 = n3462 ;
  assign y1336 = 1'b0 ;
  assign y1337 = ~1'b0 ;
  assign y1338 = n3465 ;
  assign y1339 = n3467 ;
  assign y1340 = ~1'b0 ;
  assign y1341 = n3473 ;
  assign y1342 = n3475 ;
  assign y1343 = n3476 ;
  assign y1344 = ~1'b0 ;
  assign y1345 = n3479 ;
  assign y1346 = ~n3486 ;
  assign y1347 = ~n3489 ;
  assign y1348 = ~n3493 ;
  assign y1349 = ~1'b0 ;
  assign y1350 = ~n3497 ;
  assign y1351 = ~n3498 ;
  assign y1352 = ~n3507 ;
  assign y1353 = n3508 ;
  assign y1354 = n3509 ;
  assign y1355 = ~1'b0 ;
  assign y1356 = ~1'b0 ;
  assign y1357 = ~n3511 ;
  assign y1358 = ~n3515 ;
  assign y1359 = ~n3521 ;
  assign y1360 = ~1'b0 ;
  assign y1361 = 1'b0 ;
  assign y1362 = n3524 ;
  assign y1363 = n3526 ;
  assign y1364 = ~n3538 ;
  assign y1365 = n3540 ;
  assign y1366 = ~1'b0 ;
  assign y1367 = ~1'b0 ;
  assign y1368 = n3546 ;
  assign y1369 = ~1'b0 ;
  assign y1370 = ~1'b0 ;
  assign y1371 = ~1'b0 ;
  assign y1372 = ~1'b0 ;
  assign y1373 = n3547 ;
  assign y1374 = n3550 ;
  assign y1375 = n3551 ;
  assign y1376 = ~n3552 ;
  assign y1377 = ~n3554 ;
  assign y1378 = ~n3558 ;
  assign y1379 = ~n3566 ;
  assign y1380 = ~n3576 ;
  assign y1381 = n3586 ;
  assign y1382 = ~1'b0 ;
  assign y1383 = n3587 ;
  assign y1384 = ~1'b0 ;
  assign y1385 = n3588 ;
  assign y1386 = n3596 ;
  assign y1387 = n3606 ;
  assign y1388 = n3610 ;
  assign y1389 = n3611 ;
  assign y1390 = ~n3618 ;
  assign y1391 = ~1'b0 ;
  assign y1392 = ~n3622 ;
  assign y1393 = ~n3627 ;
  assign y1394 = ~1'b0 ;
  assign y1395 = ~n3635 ;
  assign y1396 = ~1'b0 ;
  assign y1397 = ~n3600 ;
  assign y1398 = n3643 ;
  assign y1399 = ~n3645 ;
  assign y1400 = n3648 ;
  assign y1401 = ~n3651 ;
  assign y1402 = ~1'b0 ;
  assign y1403 = n3652 ;
  assign y1404 = ~1'b0 ;
  assign y1405 = 1'b0 ;
  assign y1406 = ~1'b0 ;
  assign y1407 = n3653 ;
  assign y1408 = ~n3654 ;
  assign y1409 = ~n610 ;
  assign y1410 = n3660 ;
  assign y1411 = n3664 ;
  assign y1412 = ~n3666 ;
  assign y1413 = ~n3667 ;
  assign y1414 = ~1'b0 ;
  assign y1415 = n3672 ;
  assign y1416 = ~1'b0 ;
  assign y1417 = ~n3673 ;
  assign y1418 = n3676 ;
  assign y1419 = ~n3680 ;
  assign y1420 = n3685 ;
  assign y1421 = ~1'b0 ;
  assign y1422 = n3686 ;
  assign y1423 = n3689 ;
  assign y1424 = ~n1110 ;
  assign y1425 = n3690 ;
  assign y1426 = ~n3691 ;
  assign y1427 = ~1'b0 ;
  assign y1428 = n3694 ;
  assign y1429 = ~n3697 ;
  assign y1430 = n3700 ;
  assign y1431 = n1913 ;
  assign y1432 = ~n3701 ;
  assign y1433 = n3706 ;
  assign y1434 = n3708 ;
  assign y1435 = ~n3714 ;
  assign y1436 = n3720 ;
  assign y1437 = ~n3721 ;
  assign y1438 = ~n3732 ;
  assign y1439 = ~1'b0 ;
  assign y1440 = n3734 ;
  assign y1441 = ~n3744 ;
  assign y1442 = n3746 ;
  assign y1443 = ~n3749 ;
  assign y1444 = n3750 ;
  assign y1445 = ~1'b0 ;
  assign y1446 = n3755 ;
  assign y1447 = ~n3759 ;
  assign y1448 = n1665 ;
  assign y1449 = ~1'b0 ;
  assign y1450 = ~n3761 ;
  assign y1451 = ~1'b0 ;
  assign y1452 = n3763 ;
  assign y1453 = n3765 ;
  assign y1454 = n3767 ;
  assign y1455 = n704 ;
  assign y1456 = ~1'b0 ;
  assign y1457 = n3769 ;
  assign y1458 = n3772 ;
  assign y1459 = n3782 ;
  assign y1460 = ~n3785 ;
  assign y1461 = ~1'b0 ;
  assign y1462 = ~n3786 ;
  assign y1463 = ~n3788 ;
  assign y1464 = n3793 ;
  assign y1465 = ~1'b0 ;
  assign y1466 = ~1'b0 ;
  assign y1467 = ~n3796 ;
  assign y1468 = ~1'b0 ;
  assign y1469 = ~n3798 ;
  assign y1470 = n3800 ;
  assign y1471 = ~n3806 ;
  assign y1472 = ~n3815 ;
  assign y1473 = ~1'b0 ;
  assign y1474 = n3817 ;
  assign y1475 = ~n3819 ;
  assign y1476 = n3822 ;
  assign y1477 = ~1'b0 ;
  assign y1478 = ~1'b0 ;
  assign y1479 = n3827 ;
  assign y1480 = ~1'b0 ;
  assign y1481 = n3831 ;
  assign y1482 = ~1'b0 ;
  assign y1483 = ~n1323 ;
  assign y1484 = ~1'b0 ;
  assign y1485 = ~1'b0 ;
  assign y1486 = ~n3833 ;
  assign y1487 = ~n3837 ;
  assign y1488 = n3841 ;
  assign y1489 = ~n3844 ;
  assign y1490 = ~n3847 ;
  assign y1491 = ~n3848 ;
  assign y1492 = ~1'b0 ;
  assign y1493 = n3853 ;
  assign y1494 = n3859 ;
  assign y1495 = n3864 ;
  assign y1496 = ~1'b0 ;
  assign y1497 = ~1'b0 ;
  assign y1498 = n3871 ;
  assign y1499 = n3874 ;
  assign y1500 = ~1'b0 ;
  assign y1501 = ~1'b0 ;
  assign y1502 = ~n3879 ;
  assign y1503 = n3880 ;
  assign y1504 = ~n3882 ;
  assign y1505 = ~n3884 ;
  assign y1506 = ~n3885 ;
  assign y1507 = n3887 ;
  assign y1508 = n2544 ;
  assign y1509 = n3889 ;
  assign y1510 = ~n3893 ;
  assign y1511 = ~1'b0 ;
  assign y1512 = ~n3894 ;
  assign y1513 = n3899 ;
  assign y1514 = ~1'b0 ;
  assign y1515 = ~n3901 ;
  assign y1516 = ~n3915 ;
  assign y1517 = ~n3921 ;
  assign y1518 = ~1'b0 ;
  assign y1519 = ~1'b0 ;
  assign y1520 = ~n3924 ;
  assign y1521 = n3938 ;
  assign y1522 = n3940 ;
  assign y1523 = ~1'b0 ;
  assign y1524 = ~1'b0 ;
  assign y1525 = ~n3946 ;
  assign y1526 = n3947 ;
  assign y1527 = ~n3951 ;
  assign y1528 = n3953 ;
  assign y1529 = n3955 ;
  assign y1530 = ~n3958 ;
  assign y1531 = ~n3960 ;
  assign y1532 = ~1'b0 ;
  assign y1533 = n3962 ;
  assign y1534 = ~n3965 ;
  assign y1535 = n3968 ;
  assign y1536 = ~1'b0 ;
  assign y1537 = ~n3973 ;
  assign y1538 = ~n3975 ;
  assign y1539 = n3981 ;
  assign y1540 = ~1'b0 ;
  assign y1541 = ~1'b0 ;
  assign y1542 = ~n3983 ;
  assign y1543 = ~1'b0 ;
  assign y1544 = ~n3985 ;
  assign y1545 = ~1'b0 ;
  assign y1546 = ~n3986 ;
  assign y1547 = n3997 ;
  assign y1548 = ~n4000 ;
  assign y1549 = ~n4001 ;
  assign y1550 = n4004 ;
  assign y1551 = n4007 ;
  assign y1552 = ~n4020 ;
  assign y1553 = ~n4029 ;
  assign y1554 = ~n4035 ;
  assign y1555 = ~n4037 ;
  assign y1556 = n4038 ;
  assign y1557 = ~1'b0 ;
  assign y1558 = ~1'b0 ;
  assign y1559 = ~n4039 ;
  assign y1560 = ~n4046 ;
  assign y1561 = ~n4048 ;
  assign y1562 = ~n4055 ;
  assign y1563 = n4056 ;
  assign y1564 = 1'b0 ;
  assign y1565 = n4059 ;
  assign y1566 = n4062 ;
  assign y1567 = n4063 ;
  assign y1568 = ~1'b0 ;
  assign y1569 = ~1'b0 ;
  assign y1570 = ~n4068 ;
  assign y1571 = ~1'b0 ;
  assign y1572 = ~n4076 ;
  assign y1573 = ~n4086 ;
  assign y1574 = n4087 ;
  assign y1575 = ~n4093 ;
  assign y1576 = ~1'b0 ;
  assign y1577 = ~n4095 ;
  assign y1578 = ~n4099 ;
  assign y1579 = ~n4104 ;
  assign y1580 = ~n4114 ;
  assign y1581 = n4120 ;
  assign y1582 = n4129 ;
  assign y1583 = ~1'b0 ;
  assign y1584 = n4136 ;
  assign y1585 = ~1'b0 ;
  assign y1586 = n4144 ;
  assign y1587 = ~1'b0 ;
  assign y1588 = ~n4146 ;
  assign y1589 = ~n4147 ;
  assign y1590 = ~n4152 ;
  assign y1591 = n4153 ;
  assign y1592 = n4158 ;
  assign y1593 = ~n4160 ;
  assign y1594 = ~n4167 ;
  assign y1595 = ~n4169 ;
  assign y1596 = ~n4172 ;
  assign y1597 = ~n4173 ;
  assign y1598 = n4180 ;
  assign y1599 = n4186 ;
  assign y1600 = ~n4187 ;
  assign y1601 = n4193 ;
  assign y1602 = n4194 ;
  assign y1603 = n4195 ;
  assign y1604 = ~n4198 ;
  assign y1605 = ~n4203 ;
  assign y1606 = ~n4210 ;
  assign y1607 = ~n4211 ;
  assign y1608 = ~n4228 ;
  assign y1609 = ~1'b0 ;
  assign y1610 = ~n4229 ;
  assign y1611 = n4235 ;
  assign y1612 = ~n4246 ;
  assign y1613 = n4247 ;
  assign y1614 = n4253 ;
  assign y1615 = ~n2907 ;
  assign y1616 = ~n4256 ;
  assign y1617 = ~1'b0 ;
  assign y1618 = n4257 ;
  assign y1619 = n4258 ;
  assign y1620 = n4259 ;
  assign y1621 = ~n4263 ;
  assign y1622 = ~n4267 ;
  assign y1623 = ~1'b0 ;
  assign y1624 = ~1'b0 ;
  assign y1625 = ~n4275 ;
  assign y1626 = ~1'b0 ;
  assign y1627 = n4279 ;
  assign y1628 = n4283 ;
  assign y1629 = n4290 ;
  assign y1630 = ~n4292 ;
  assign y1631 = n4296 ;
  assign y1632 = ~1'b0 ;
  assign y1633 = ~n4303 ;
  assign y1634 = ~n512 ;
  assign y1635 = ~n4306 ;
  assign y1636 = ~1'b0 ;
  assign y1637 = 1'b0 ;
  assign y1638 = n4308 ;
  assign y1639 = n4309 ;
  assign y1640 = ~n4310 ;
  assign y1641 = ~1'b0 ;
  assign y1642 = ~n4312 ;
  assign y1643 = ~1'b0 ;
  assign y1644 = ~n4315 ;
  assign y1645 = n4323 ;
  assign y1646 = n4328 ;
  assign y1647 = ~n4334 ;
  assign y1648 = ~1'b0 ;
  assign y1649 = ~n4340 ;
  assign y1650 = n4346 ;
  assign y1651 = n4347 ;
  assign y1652 = ~n4352 ;
  assign y1653 = ~n4354 ;
  assign y1654 = n4359 ;
  assign y1655 = ~1'b0 ;
  assign y1656 = ~1'b0 ;
  assign y1657 = ~1'b0 ;
  assign y1658 = n4364 ;
  assign y1659 = ~n4368 ;
  assign y1660 = ~n4369 ;
  assign y1661 = ~n4371 ;
  assign y1662 = ~1'b0 ;
  assign y1663 = ~1'b0 ;
  assign y1664 = ~1'b0 ;
  assign y1665 = ~1'b0 ;
  assign y1666 = n4375 ;
  assign y1667 = ~1'b0 ;
  assign y1668 = ~n4379 ;
  assign y1669 = n1930 ;
  assign y1670 = ~n4383 ;
  assign y1671 = ~n4391 ;
  assign y1672 = n4396 ;
  assign y1673 = ~n4402 ;
  assign y1674 = ~1'b0 ;
  assign y1675 = ~n4405 ;
  assign y1676 = n4406 ;
  assign y1677 = ~1'b0 ;
  assign y1678 = n4407 ;
  assign y1679 = ~n4415 ;
  assign y1680 = ~1'b0 ;
  assign y1681 = n4418 ;
  assign y1682 = ~n4421 ;
  assign y1683 = 1'b0 ;
  assign y1684 = ~n4425 ;
  assign y1685 = ~1'b0 ;
  assign y1686 = ~1'b0 ;
  assign y1687 = ~1'b0 ;
  assign y1688 = n4426 ;
  assign y1689 = ~n4432 ;
  assign y1690 = n4433 ;
  assign y1691 = ~1'b0 ;
  assign y1692 = n4442 ;
  assign y1693 = n4445 ;
  assign y1694 = ~n4450 ;
  assign y1695 = ~1'b0 ;
  assign y1696 = ~n4452 ;
  assign y1697 = ~n4454 ;
  assign y1698 = ~n4455 ;
  assign y1699 = n4457 ;
  assign y1700 = n4196 ;
  assign y1701 = ~n4466 ;
  assign y1702 = ~1'b0 ;
  assign y1703 = ~n4467 ;
  assign y1704 = ~n4468 ;
  assign y1705 = ~n4473 ;
  assign y1706 = ~1'b0 ;
  assign y1707 = ~n4474 ;
  assign y1708 = n4477 ;
  assign y1709 = ~n4479 ;
  assign y1710 = ~n4483 ;
  assign y1711 = n4485 ;
  assign y1712 = ~n4487 ;
  assign y1713 = ~n4488 ;
  assign y1714 = n4491 ;
  assign y1715 = ~1'b0 ;
  assign y1716 = ~n4495 ;
  assign y1717 = ~1'b0 ;
  assign y1718 = ~1'b0 ;
  assign y1719 = n4496 ;
  assign y1720 = n4497 ;
  assign y1721 = ~n4498 ;
  assign y1722 = n4501 ;
  assign y1723 = n4503 ;
  assign y1724 = ~n4507 ;
  assign y1725 = ~1'b0 ;
  assign y1726 = ~n4508 ;
  assign y1727 = n4511 ;
  assign y1728 = ~1'b0 ;
  assign y1729 = n4520 ;
  assign y1730 = ~n4528 ;
  assign y1731 = ~n4529 ;
  assign y1732 = ~n4531 ;
  assign y1733 = n4532 ;
  assign y1734 = ~n4534 ;
  assign y1735 = n4537 ;
  assign y1736 = ~n4540 ;
  assign y1737 = ~n4545 ;
  assign y1738 = ~1'b0 ;
  assign y1739 = ~n4548 ;
  assign y1740 = n4549 ;
  assign y1741 = n4550 ;
  assign y1742 = n4553 ;
  assign y1743 = ~1'b0 ;
  assign y1744 = ~n4556 ;
  assign y1745 = ~n4557 ;
  assign y1746 = ~1'b0 ;
  assign y1747 = n4561 ;
  assign y1748 = n4567 ;
  assign y1749 = n4576 ;
  assign y1750 = ~1'b0 ;
  assign y1751 = ~n4579 ;
  assign y1752 = ~n4580 ;
  assign y1753 = n2922 ;
  assign y1754 = ~n4582 ;
  assign y1755 = ~n4583 ;
  assign y1756 = ~n4584 ;
  assign y1757 = n4587 ;
  assign y1758 = ~1'b0 ;
  assign y1759 = ~n4590 ;
  assign y1760 = n4593 ;
  assign y1761 = n4595 ;
  assign y1762 = ~1'b0 ;
  assign y1763 = ~1'b0 ;
  assign y1764 = n4599 ;
  assign y1765 = n4600 ;
  assign y1766 = n4602 ;
  assign y1767 = ~n4607 ;
  assign y1768 = ~n4611 ;
  assign y1769 = ~n4614 ;
  assign y1770 = ~1'b0 ;
  assign y1771 = ~n4616 ;
  assign y1772 = ~n4622 ;
  assign y1773 = ~n4627 ;
  assign y1774 = ~n4630 ;
  assign y1775 = n4634 ;
  assign y1776 = x142 ;
  assign y1777 = n4643 ;
  assign y1778 = 1'b0 ;
  assign y1779 = ~1'b0 ;
  assign y1780 = ~1'b0 ;
  assign y1781 = n4648 ;
  assign y1782 = ~n4650 ;
  assign y1783 = n4651 ;
  assign y1784 = ~n4658 ;
  assign y1785 = n4666 ;
  assign y1786 = 1'b0 ;
  assign y1787 = ~n2213 ;
  assign y1788 = ~n4672 ;
  assign y1789 = ~n4673 ;
  assign y1790 = n4674 ;
  assign y1791 = n4681 ;
  assign y1792 = ~n4684 ;
  assign y1793 = ~n4691 ;
  assign y1794 = n4693 ;
  assign y1795 = ~1'b0 ;
  assign y1796 = ~1'b0 ;
  assign y1797 = ~n4696 ;
  assign y1798 = n4705 ;
  assign y1799 = ~n4707 ;
  assign y1800 = ~1'b0 ;
  assign y1801 = n4711 ;
  assign y1802 = ~n4713 ;
  assign y1803 = ~n4714 ;
  assign y1804 = ~1'b0 ;
  assign y1805 = ~1'b0 ;
  assign y1806 = n4716 ;
  assign y1807 = ~n4719 ;
  assign y1808 = n4722 ;
  assign y1809 = ~1'b0 ;
  assign y1810 = 1'b0 ;
  assign y1811 = 1'b0 ;
  assign y1812 = ~1'b0 ;
  assign y1813 = n4723 ;
  assign y1814 = n1254 ;
  assign y1815 = n4731 ;
  assign y1816 = n648 ;
  assign y1817 = ~n4736 ;
  assign y1818 = n4741 ;
  assign y1819 = n4742 ;
  assign y1820 = ~n4744 ;
  assign y1821 = ~1'b0 ;
  assign y1822 = ~n4749 ;
  assign y1823 = ~n4751 ;
  assign y1824 = ~n2495 ;
  assign y1825 = ~n4752 ;
  assign y1826 = ~1'b0 ;
  assign y1827 = ~1'b0 ;
  assign y1828 = ~n4754 ;
  assign y1829 = ~n4762 ;
  assign y1830 = ~1'b0 ;
  assign y1831 = ~n4767 ;
  assign y1832 = n4774 ;
  assign y1833 = ~1'b0 ;
  assign y1834 = ~1'b0 ;
  assign y1835 = ~n4775 ;
  assign y1836 = ~1'b0 ;
  assign y1837 = ~n1930 ;
  assign y1838 = ~n2651 ;
  assign y1839 = n4778 ;
  assign y1840 = n4783 ;
  assign y1841 = n4790 ;
  assign y1842 = n4792 ;
  assign y1843 = ~1'b0 ;
  assign y1844 = n4797 ;
  assign y1845 = ~1'b0 ;
  assign y1846 = ~n4800 ;
  assign y1847 = ~1'b0 ;
  assign y1848 = n4803 ;
  assign y1849 = n4806 ;
  assign y1850 = ~1'b0 ;
  assign y1851 = n4810 ;
  assign y1852 = ~1'b0 ;
  assign y1853 = n4812 ;
  assign y1854 = ~n4815 ;
  assign y1855 = n4818 ;
  assign y1856 = ~n4820 ;
  assign y1857 = n3915 ;
  assign y1858 = ~n4826 ;
  assign y1859 = ~1'b0 ;
  assign y1860 = n4830 ;
  assign y1861 = ~1'b0 ;
  assign y1862 = ~n4832 ;
  assign y1863 = ~n4840 ;
  assign y1864 = n4842 ;
  assign y1865 = ~n4844 ;
  assign y1866 = ~n4846 ;
  assign y1867 = ~n3587 ;
  assign y1868 = n4849 ;
  assign y1869 = ~1'b0 ;
  assign y1870 = ~1'b0 ;
  assign y1871 = n4850 ;
  assign y1872 = n4858 ;
  assign y1873 = n4865 ;
  assign y1874 = ~1'b0 ;
  assign y1875 = n4868 ;
  assign y1876 = ~1'b0 ;
  assign y1877 = n4870 ;
  assign y1878 = n4873 ;
  assign y1879 = ~n4880 ;
  assign y1880 = n4881 ;
  assign y1881 = ~n4882 ;
  assign y1882 = ~n4890 ;
  assign y1883 = n4900 ;
  assign y1884 = n4905 ;
  assign y1885 = ~n4907 ;
  assign y1886 = ~n4912 ;
  assign y1887 = n4913 ;
  assign y1888 = ~n4915 ;
  assign y1889 = ~n4925 ;
  assign y1890 = n4927 ;
  assign y1891 = n4929 ;
  assign y1892 = n4937 ;
  assign y1893 = ~n4945 ;
  assign y1894 = ~n4950 ;
  assign y1895 = ~n4951 ;
  assign y1896 = ~1'b0 ;
  assign y1897 = ~1'b0 ;
  assign y1898 = ~n4954 ;
  assign y1899 = ~n4960 ;
  assign y1900 = ~1'b0 ;
  assign y1901 = n4969 ;
  assign y1902 = ~1'b0 ;
  assign y1903 = ~n4971 ;
  assign y1904 = n4977 ;
  assign y1905 = n4978 ;
  assign y1906 = ~n2002 ;
  assign y1907 = n4982 ;
  assign y1908 = ~x153 ;
  assign y1909 = n4991 ;
  assign y1910 = ~n4994 ;
  assign y1911 = n4995 ;
  assign y1912 = n4999 ;
  assign y1913 = ~n5001 ;
  assign y1914 = n5003 ;
  assign y1915 = ~n5006 ;
  assign y1916 = n5009 ;
  assign y1917 = ~1'b0 ;
  assign y1918 = ~1'b0 ;
  assign y1919 = ~1'b0 ;
  assign y1920 = n5011 ;
  assign y1921 = n5017 ;
  assign y1922 = ~1'b0 ;
  assign y1923 = n5020 ;
  assign y1924 = n5021 ;
  assign y1925 = ~1'b0 ;
  assign y1926 = ~n5022 ;
  assign y1927 = n5023 ;
  assign y1928 = ~n5027 ;
  assign y1929 = ~n5029 ;
  assign y1930 = ~1'b0 ;
  assign y1931 = n5031 ;
  assign y1932 = ~n2080 ;
  assign y1933 = n5036 ;
  assign y1934 = n5039 ;
  assign y1935 = ~1'b0 ;
  assign y1936 = ~n5045 ;
  assign y1937 = ~n4580 ;
  assign y1938 = ~n1585 ;
  assign y1939 = n5046 ;
  assign y1940 = ~1'b0 ;
  assign y1941 = n5047 ;
  assign y1942 = ~1'b0 ;
  assign y1943 = ~n5048 ;
  assign y1944 = ~n5050 ;
  assign y1945 = n5052 ;
  assign y1946 = n5053 ;
  assign y1947 = ~n5054 ;
  assign y1948 = n5056 ;
  assign y1949 = ~n5057 ;
  assign y1950 = ~n5061 ;
  assign y1951 = ~n5063 ;
  assign y1952 = n5064 ;
  assign y1953 = ~n5067 ;
  assign y1954 = ~1'b0 ;
  assign y1955 = ~n3814 ;
  assign y1956 = ~n5068 ;
  assign y1957 = ~n5070 ;
  assign y1958 = n5072 ;
  assign y1959 = ~n5074 ;
  assign y1960 = ~n5075 ;
  assign y1961 = ~n5081 ;
  assign y1962 = ~1'b0 ;
  assign y1963 = n5084 ;
  assign y1964 = ~n5090 ;
  assign y1965 = ~n5091 ;
  assign y1966 = n5092 ;
  assign y1967 = n5093 ;
  assign y1968 = ~1'b0 ;
  assign y1969 = n5099 ;
  assign y1970 = ~n5102 ;
  assign y1971 = n5105 ;
  assign y1972 = ~1'b0 ;
  assign y1973 = ~n4462 ;
  assign y1974 = n5110 ;
  assign y1975 = ~1'b0 ;
  assign y1976 = ~n5113 ;
  assign y1977 = ~n5116 ;
  assign y1978 = n5117 ;
  assign y1979 = 1'b0 ;
  assign y1980 = n5124 ;
  assign y1981 = ~1'b0 ;
  assign y1982 = ~n3624 ;
  assign y1983 = ~1'b0 ;
  assign y1984 = ~n5131 ;
  assign y1985 = ~n5133 ;
  assign y1986 = n5134 ;
  assign y1987 = n5139 ;
  assign y1988 = ~1'b0 ;
  assign y1989 = ~1'b0 ;
  assign y1990 = ~n5141 ;
  assign y1991 = ~n5142 ;
  assign y1992 = n5143 ;
  assign y1993 = ~1'b0 ;
  assign y1994 = n5145 ;
  assign y1995 = n5150 ;
  assign y1996 = n5154 ;
  assign y1997 = n4460 ;
  assign y1998 = ~1'b0 ;
  assign y1999 = ~n5160 ;
  assign y2000 = ~n5164 ;
  assign y2001 = n5167 ;
  assign y2002 = ~n5172 ;
  assign y2003 = n5173 ;
  assign y2004 = n5176 ;
  assign y2005 = ~n5178 ;
  assign y2006 = ~1'b0 ;
  assign y2007 = ~n5185 ;
  assign y2008 = ~1'b0 ;
  assign y2009 = ~1'b0 ;
  assign y2010 = ~n5190 ;
  assign y2011 = n5200 ;
  assign y2012 = n5203 ;
  assign y2013 = ~n5205 ;
  assign y2014 = n5208 ;
  assign y2015 = ~n5216 ;
  assign y2016 = n5223 ;
  assign y2017 = ~1'b0 ;
  assign y2018 = ~n5225 ;
  assign y2019 = ~1'b0 ;
  assign y2020 = ~n5230 ;
  assign y2021 = ~1'b0 ;
  assign y2022 = n5231 ;
  assign y2023 = ~n5235 ;
  assign y2024 = ~1'b0 ;
  assign y2025 = ~1'b0 ;
  assign y2026 = n5244 ;
  assign y2027 = n5248 ;
  assign y2028 = n5252 ;
  assign y2029 = ~n5253 ;
  assign y2030 = ~1'b0 ;
  assign y2031 = ~n5255 ;
  assign y2032 = n5256 ;
  assign y2033 = ~1'b0 ;
  assign y2034 = ~n5259 ;
  assign y2035 = ~n5266 ;
  assign y2036 = ~n4300 ;
  assign y2037 = ~n5269 ;
  assign y2038 = n5276 ;
  assign y2039 = n5282 ;
  assign y2040 = ~n5283 ;
  assign y2041 = n5285 ;
  assign y2042 = ~1'b0 ;
  assign y2043 = ~n5286 ;
  assign y2044 = ~n5292 ;
  assign y2045 = n5296 ;
  assign y2046 = n5298 ;
  assign y2047 = ~1'b0 ;
  assign y2048 = n5303 ;
  assign y2049 = n5304 ;
  assign y2050 = ~n5310 ;
  assign y2051 = ~1'b0 ;
  assign y2052 = ~1'b0 ;
  assign y2053 = n5317 ;
  assign y2054 = ~n5319 ;
  assign y2055 = n5324 ;
  assign y2056 = n5329 ;
  assign y2057 = ~1'b0 ;
  assign y2058 = n5339 ;
  assign y2059 = n5356 ;
  assign y2060 = ~n5361 ;
  assign y2061 = ~1'b0 ;
  assign y2062 = n5363 ;
  assign y2063 = ~n5369 ;
  assign y2064 = ~n5370 ;
  assign y2065 = n5372 ;
  assign y2066 = ~1'b0 ;
  assign y2067 = ~n5376 ;
  assign y2068 = n5380 ;
  assign y2069 = ~n5381 ;
  assign y2070 = n5385 ;
  assign y2071 = n5386 ;
  assign y2072 = n1553 ;
  assign y2073 = n5387 ;
  assign y2074 = n5391 ;
  assign y2075 = ~n5398 ;
  assign y2076 = ~n5400 ;
  assign y2077 = ~n5402 ;
  assign y2078 = ~n5406 ;
  assign y2079 = n5408 ;
  assign y2080 = n5412 ;
  assign y2081 = ~1'b0 ;
  assign y2082 = n5413 ;
  assign y2083 = n5414 ;
  assign y2084 = ~n5417 ;
  assign y2085 = n5421 ;
  assign y2086 = ~1'b0 ;
  assign y2087 = ~n3104 ;
  assign y2088 = ~n5426 ;
  assign y2089 = n5430 ;
  assign y2090 = ~n5437 ;
  assign y2091 = n5439 ;
  assign y2092 = ~n5445 ;
  assign y2093 = ~n4194 ;
  assign y2094 = n5446 ;
  assign y2095 = n5448 ;
  assign y2096 = n5449 ;
  assign y2097 = n5451 ;
  assign y2098 = ~1'b0 ;
  assign y2099 = n5455 ;
  assign y2100 = ~1'b0 ;
  assign y2101 = ~n5461 ;
  assign y2102 = 1'b0 ;
  assign y2103 = ~n5468 ;
  assign y2104 = n5478 ;
  assign y2105 = ~1'b0 ;
  assign y2106 = ~1'b0 ;
  assign y2107 = n5479 ;
  assign y2108 = n5483 ;
  assign y2109 = n5493 ;
  assign y2110 = ~n5497 ;
  assign y2111 = ~n5499 ;
  assign y2112 = n5501 ;
  assign y2113 = ~1'b0 ;
  assign y2114 = ~1'b0 ;
  assign y2115 = ~1'b0 ;
  assign y2116 = ~1'b0 ;
  assign y2117 = n5502 ;
  assign y2118 = n5504 ;
  assign y2119 = ~1'b0 ;
  assign y2120 = n5510 ;
  assign y2121 = n5511 ;
  assign y2122 = ~n5514 ;
  assign y2123 = ~1'b0 ;
  assign y2124 = ~n5518 ;
  assign y2125 = ~1'b0 ;
  assign y2126 = ~1'b0 ;
  assign y2127 = n5522 ;
  assign y2128 = ~n5523 ;
  assign y2129 = ~n5525 ;
  assign y2130 = n5528 ;
  assign y2131 = ~n5529 ;
  assign y2132 = ~n5531 ;
  assign y2133 = ~1'b0 ;
  assign y2134 = ~1'b0 ;
  assign y2135 = ~1'b0 ;
  assign y2136 = ~n5535 ;
  assign y2137 = n5536 ;
  assign y2138 = ~1'b0 ;
  assign y2139 = ~1'b0 ;
  assign y2140 = ~1'b0 ;
  assign y2141 = ~n5537 ;
  assign y2142 = ~n5541 ;
  assign y2143 = ~1'b0 ;
  assign y2144 = x244 ;
  assign y2145 = ~1'b0 ;
  assign y2146 = ~1'b0 ;
  assign y2147 = ~n5552 ;
  assign y2148 = ~1'b0 ;
  assign y2149 = n5556 ;
  assign y2150 = ~1'b0 ;
  assign y2151 = 1'b0 ;
  assign y2152 = ~1'b0 ;
  assign y2153 = ~1'b0 ;
  assign y2154 = ~n5558 ;
  assign y2155 = ~n5560 ;
  assign y2156 = ~1'b0 ;
  assign y2157 = n5567 ;
  assign y2158 = ~1'b0 ;
  assign y2159 = ~1'b0 ;
  assign y2160 = ~1'b0 ;
  assign y2161 = ~n5568 ;
  assign y2162 = ~1'b0 ;
  assign y2163 = ~n5569 ;
  assign y2164 = ~n5573 ;
  assign y2165 = n5576 ;
  assign y2166 = n2074 ;
  assign y2167 = ~n5577 ;
  assign y2168 = n5578 ;
  assign y2169 = ~1'b0 ;
  assign y2170 = ~n5581 ;
  assign y2171 = n5582 ;
  assign y2172 = ~n5583 ;
  assign y2173 = ~n5589 ;
  assign y2174 = n5590 ;
  assign y2175 = ~1'b0 ;
  assign y2176 = n5596 ;
  assign y2177 = ~1'b0 ;
  assign y2178 = ~n5598 ;
  assign y2179 = n5599 ;
  assign y2180 = n5601 ;
  assign y2181 = ~1'b0 ;
  assign y2182 = ~1'b0 ;
  assign y2183 = ~1'b0 ;
  assign y2184 = n5607 ;
  assign y2185 = ~n5608 ;
  assign y2186 = n5617 ;
  assign y2187 = n5618 ;
  assign y2188 = ~n5620 ;
  assign y2189 = n780 ;
  assign y2190 = n5621 ;
  assign y2191 = ~1'b0 ;
  assign y2192 = n5636 ;
  assign y2193 = n5637 ;
  assign y2194 = ~n5638 ;
  assign y2195 = ~1'b0 ;
  assign y2196 = ~1'b0 ;
  assign y2197 = ~n5639 ;
  assign y2198 = n5643 ;
  assign y2199 = ~n5647 ;
  assign y2200 = ~n5648 ;
  assign y2201 = n5649 ;
  assign y2202 = n5655 ;
  assign y2203 = ~1'b0 ;
  assign y2204 = ~1'b0 ;
  assign y2205 = ~1'b0 ;
  assign y2206 = n5660 ;
  assign y2207 = ~n5667 ;
  assign y2208 = ~1'b0 ;
  assign y2209 = ~n5669 ;
  assign y2210 = ~n5672 ;
  assign y2211 = ~n5673 ;
  assign y2212 = ~1'b0 ;
  assign y2213 = ~n5674 ;
  assign y2214 = n5676 ;
  assign y2215 = ~n5677 ;
  assign y2216 = n5678 ;
  assign y2217 = ~n2539 ;
  assign y2218 = ~n5680 ;
  assign y2219 = n5681 ;
  assign y2220 = ~n5683 ;
  assign y2221 = n5685 ;
  assign y2222 = n5688 ;
  assign y2223 = ~1'b0 ;
  assign y2224 = n5690 ;
  assign y2225 = n5691 ;
  assign y2226 = ~n5698 ;
  assign y2227 = ~1'b0 ;
  assign y2228 = ~1'b0 ;
  assign y2229 = ~1'b0 ;
  assign y2230 = ~1'b0 ;
  assign y2231 = n5699 ;
  assign y2232 = ~1'b0 ;
  assign y2233 = n5701 ;
  assign y2234 = n5703 ;
  assign y2235 = ~n5705 ;
  assign y2236 = ~n5710 ;
  assign y2237 = ~n5716 ;
  assign y2238 = ~1'b0 ;
  assign y2239 = n5718 ;
  assign y2240 = ~1'b0 ;
  assign y2241 = ~1'b0 ;
  assign y2242 = ~n5720 ;
  assign y2243 = n5721 ;
  assign y2244 = n5726 ;
  assign y2245 = ~n5738 ;
  assign y2246 = ~1'b0 ;
  assign y2247 = n5741 ;
  assign y2248 = ~1'b0 ;
  assign y2249 = ~n5742 ;
  assign y2250 = n5750 ;
  assign y2251 = n5751 ;
  assign y2252 = n5752 ;
  assign y2253 = n5755 ;
  assign y2254 = ~n880 ;
  assign y2255 = ~1'b0 ;
  assign y2256 = n5759 ;
  assign y2257 = n5760 ;
  assign y2258 = n5767 ;
  assign y2259 = ~n5768 ;
  assign y2260 = ~1'b0 ;
  assign y2261 = ~n5772 ;
  assign y2262 = n5773 ;
  assign y2263 = ~n5775 ;
  assign y2264 = n5778 ;
  assign y2265 = ~n5786 ;
  assign y2266 = ~n5788 ;
  assign y2267 = n5791 ;
  assign y2268 = ~1'b0 ;
  assign y2269 = ~n5793 ;
  assign y2270 = n5795 ;
  assign y2271 = ~n1813 ;
  assign y2272 = ~n5797 ;
  assign y2273 = ~n5798 ;
  assign y2274 = ~n5800 ;
  assign y2275 = ~n5801 ;
  assign y2276 = n5802 ;
  assign y2277 = ~n5806 ;
  assign y2278 = ~n5812 ;
  assign y2279 = ~1'b0 ;
  assign y2280 = ~n5813 ;
  assign y2281 = n5814 ;
  assign y2282 = ~n5818 ;
  assign y2283 = ~n5820 ;
  assign y2284 = ~n5824 ;
  assign y2285 = ~n3043 ;
  assign y2286 = ~n5826 ;
  assign y2287 = ~n5830 ;
  assign y2288 = n5832 ;
  assign y2289 = ~n5833 ;
  assign y2290 = ~n5834 ;
  assign y2291 = ~1'b0 ;
  assign y2292 = n5839 ;
  assign y2293 = ~1'b0 ;
  assign y2294 = n5550 ;
  assign y2295 = ~1'b0 ;
  assign y2296 = ~1'b0 ;
  assign y2297 = ~n5840 ;
  assign y2298 = n2698 ;
  assign y2299 = n5841 ;
  assign y2300 = ~n5846 ;
  assign y2301 = ~n5849 ;
  assign y2302 = ~n5851 ;
  assign y2303 = n5852 ;
  assign y2304 = n1932 ;
  assign y2305 = ~n5855 ;
  assign y2306 = ~n5865 ;
  assign y2307 = ~n5866 ;
  assign y2308 = ~1'b0 ;
  assign y2309 = ~n5868 ;
  assign y2310 = n5869 ;
  assign y2311 = ~1'b0 ;
  assign y2312 = n5870 ;
  assign y2313 = ~1'b0 ;
  assign y2314 = ~n5874 ;
  assign y2315 = n4719 ;
  assign y2316 = ~1'b0 ;
  assign y2317 = ~1'b0 ;
  assign y2318 = n5876 ;
  assign y2319 = ~1'b0 ;
  assign y2320 = ~n5884 ;
  assign y2321 = ~1'b0 ;
  assign y2322 = ~n5888 ;
  assign y2323 = ~n5895 ;
  assign y2324 = ~n5899 ;
  assign y2325 = n5901 ;
  assign y2326 = ~1'b0 ;
  assign y2327 = ~1'b0 ;
  assign y2328 = ~n5909 ;
  assign y2329 = ~1'b0 ;
  assign y2330 = n5910 ;
  assign y2331 = ~n5916 ;
  assign y2332 = n5918 ;
  assign y2333 = n5920 ;
  assign y2334 = ~1'b0 ;
  assign y2335 = ~1'b0 ;
  assign y2336 = ~n5921 ;
  assign y2337 = n5923 ;
  assign y2338 = ~n5926 ;
  assign y2339 = n5927 ;
  assign y2340 = ~1'b0 ;
  assign y2341 = n5929 ;
  assign y2342 = ~n5941 ;
  assign y2343 = ~n5943 ;
  assign y2344 = n5945 ;
  assign y2345 = ~n5954 ;
  assign y2346 = ~n5956 ;
  assign y2347 = ~1'b0 ;
  assign y2348 = n5960 ;
  assign y2349 = ~n2995 ;
  assign y2350 = ~n5963 ;
  assign y2351 = n5965 ;
  assign y2352 = n5966 ;
  assign y2353 = n5971 ;
  assign y2354 = ~1'b0 ;
  assign y2355 = ~1'b0 ;
  assign y2356 = n5973 ;
  assign y2357 = ~n5974 ;
  assign y2358 = n5230 ;
  assign y2359 = n5976 ;
  assign y2360 = n5978 ;
  assign y2361 = ~n5981 ;
  assign y2362 = ~n5984 ;
  assign y2363 = n5985 ;
  assign y2364 = ~n5988 ;
  assign y2365 = ~1'b0 ;
  assign y2366 = ~n5989 ;
  assign y2367 = n5999 ;
  assign y2368 = ~1'b0 ;
  assign y2369 = n6003 ;
  assign y2370 = ~n6012 ;
  assign y2371 = ~1'b0 ;
  assign y2372 = n4509 ;
  assign y2373 = n6021 ;
  assign y2374 = ~n5884 ;
  assign y2375 = ~n2230 ;
  assign y2376 = ~n6025 ;
  assign y2377 = n6030 ;
  assign y2378 = ~1'b0 ;
  assign y2379 = ~n6033 ;
  assign y2380 = ~n6034 ;
  assign y2381 = ~n6035 ;
  assign y2382 = n6038 ;
  assign y2383 = n6042 ;
  assign y2384 = ~1'b0 ;
  assign y2385 = n6044 ;
  assign y2386 = n6054 ;
  assign y2387 = n6058 ;
  assign y2388 = ~n6060 ;
  assign y2389 = ~1'b0 ;
  assign y2390 = n6061 ;
  assign y2391 = n6063 ;
  assign y2392 = ~n6064 ;
  assign y2393 = ~n1024 ;
  assign y2394 = ~n6066 ;
  assign y2395 = ~n6072 ;
  assign y2396 = ~1'b0 ;
  assign y2397 = ~1'b0 ;
  assign y2398 = n6074 ;
  assign y2399 = n6084 ;
  assign y2400 = n6085 ;
  assign y2401 = ~n6088 ;
  assign y2402 = n6091 ;
  assign y2403 = ~1'b0 ;
  assign y2404 = ~n6092 ;
  assign y2405 = ~n6096 ;
  assign y2406 = ~1'b0 ;
  assign y2407 = ~n6101 ;
  assign y2408 = ~n6103 ;
  assign y2409 = n6114 ;
  assign y2410 = ~n6121 ;
  assign y2411 = ~n6122 ;
  assign y2412 = ~n6123 ;
  assign y2413 = ~1'b0 ;
  assign y2414 = n6127 ;
  assign y2415 = n6129 ;
  assign y2416 = ~n6131 ;
  assign y2417 = n6134 ;
  assign y2418 = n6139 ;
  assign y2419 = n6141 ;
  assign y2420 = n6146 ;
  assign y2421 = ~n6149 ;
  assign y2422 = ~1'b0 ;
  assign y2423 = ~1'b0 ;
  assign y2424 = ~1'b0 ;
  assign y2425 = ~1'b0 ;
  assign y2426 = ~1'b0 ;
  assign y2427 = ~n6150 ;
  assign y2428 = n6158 ;
  assign y2429 = n6161 ;
  assign y2430 = n6164 ;
  assign y2431 = ~n6167 ;
  assign y2432 = ~n6169 ;
  assign y2433 = ~1'b0 ;
  assign y2434 = ~n6170 ;
  assign y2435 = ~n6172 ;
  assign y2436 = n6176 ;
  assign y2437 = n6179 ;
  assign y2438 = ~n6180 ;
  assign y2439 = ~1'b0 ;
  assign y2440 = n6182 ;
  assign y2441 = ~1'b0 ;
  assign y2442 = n6184 ;
  assign y2443 = ~n6186 ;
  assign y2444 = ~n6189 ;
  assign y2445 = n6196 ;
  assign y2446 = n432 ;
  assign y2447 = ~n286 ;
  assign y2448 = ~n6200 ;
  assign y2449 = ~n6203 ;
  assign y2450 = ~n6204 ;
  assign y2451 = ~1'b0 ;
  assign y2452 = n6206 ;
  assign y2453 = n6207 ;
  assign y2454 = ~1'b0 ;
  assign y2455 = ~n6212 ;
  assign y2456 = ~1'b0 ;
  assign y2457 = n6213 ;
  assign y2458 = ~1'b0 ;
  assign y2459 = ~n6215 ;
  assign y2460 = ~1'b0 ;
  assign y2461 = 1'b0 ;
  assign y2462 = ~1'b0 ;
  assign y2463 = n6216 ;
  assign y2464 = n6220 ;
  assign y2465 = n6221 ;
  assign y2466 = n6227 ;
  assign y2467 = n6230 ;
  assign y2468 = ~1'b0 ;
  assign y2469 = n6232 ;
  assign y2470 = n6234 ;
  assign y2471 = n6238 ;
  assign y2472 = n6242 ;
  assign y2473 = ~n6255 ;
  assign y2474 = ~n6257 ;
  assign y2475 = ~n6258 ;
  assign y2476 = ~n6259 ;
  assign y2477 = n6264 ;
  assign y2478 = ~n6267 ;
  assign y2479 = ~n6268 ;
  assign y2480 = n6270 ;
  assign y2481 = ~n6271 ;
  assign y2482 = ~1'b0 ;
  assign y2483 = ~n6272 ;
  assign y2484 = ~1'b0 ;
  assign y2485 = n6276 ;
  assign y2486 = n6284 ;
  assign y2487 = ~n6286 ;
  assign y2488 = n6287 ;
  assign y2489 = ~n6288 ;
  assign y2490 = n6291 ;
  assign y2491 = n6294 ;
  assign y2492 = n6295 ;
  assign y2493 = ~1'b0 ;
  assign y2494 = ~n6300 ;
  assign y2495 = ~n6305 ;
  assign y2496 = n6307 ;
  assign y2497 = n6312 ;
  assign y2498 = n5304 ;
  assign y2499 = n6313 ;
  assign y2500 = ~1'b0 ;
  assign y2501 = ~n6314 ;
  assign y2502 = n6318 ;
  assign y2503 = ~n6319 ;
  assign y2504 = ~n6325 ;
  assign y2505 = ~n6327 ;
  assign y2506 = ~n6330 ;
  assign y2507 = ~n6331 ;
  assign y2508 = n6332 ;
  assign y2509 = ~n6336 ;
  assign y2510 = n6346 ;
  assign y2511 = ~1'b0 ;
  assign y2512 = n6348 ;
  assign y2513 = n674 ;
  assign y2514 = ~n6350 ;
  assign y2515 = ~n6351 ;
  assign y2516 = ~1'b0 ;
  assign y2517 = n6353 ;
  assign y2518 = ~1'b0 ;
  assign y2519 = ~n6357 ;
  assign y2520 = 1'b0 ;
  assign y2521 = n6362 ;
  assign y2522 = ~n6363 ;
  assign y2523 = ~1'b0 ;
  assign y2524 = n6365 ;
  assign y2525 = ~1'b0 ;
  assign y2526 = ~n6370 ;
  assign y2527 = ~n6371 ;
  assign y2528 = ~1'b0 ;
  assign y2529 = ~n6373 ;
  assign y2530 = ~1'b0 ;
  assign y2531 = ~1'b0 ;
  assign y2532 = 1'b0 ;
  assign y2533 = ~n6377 ;
  assign y2534 = ~n6379 ;
  assign y2535 = n6383 ;
  assign y2536 = ~n6384 ;
  assign y2537 = ~n6388 ;
  assign y2538 = n6390 ;
  assign y2539 = n6398 ;
  assign y2540 = n1297 ;
  assign y2541 = ~1'b0 ;
  assign y2542 = ~1'b0 ;
  assign y2543 = ~n6400 ;
  assign y2544 = ~n6402 ;
  assign y2545 = ~1'b0 ;
  assign y2546 = ~n6405 ;
  assign y2547 = ~1'b0 ;
  assign y2548 = n6406 ;
  assign y2549 = n6409 ;
  assign y2550 = n6420 ;
  assign y2551 = ~1'b0 ;
  assign y2552 = n6421 ;
  assign y2553 = ~1'b0 ;
  assign y2554 = ~n6423 ;
  assign y2555 = n1324 ;
  assign y2556 = n6428 ;
  assign y2557 = 1'b0 ;
  assign y2558 = n6429 ;
  assign y2559 = n6436 ;
  assign y2560 = n6438 ;
  assign y2561 = n6442 ;
  assign y2562 = ~n6444 ;
  assign y2563 = ~n6445 ;
  assign y2564 = ~1'b0 ;
  assign y2565 = n6448 ;
  assign y2566 = n6450 ;
  assign y2567 = ~1'b0 ;
  assign y2568 = n6453 ;
  assign y2569 = n6455 ;
  assign y2570 = n6456 ;
  assign y2571 = ~n6462 ;
  assign y2572 = ~n6464 ;
  assign y2573 = n6466 ;
  assign y2574 = n5775 ;
  assign y2575 = ~1'b0 ;
  assign y2576 = ~1'b0 ;
  assign y2577 = n6467 ;
  assign y2578 = n6469 ;
  assign y2579 = ~n6472 ;
  assign y2580 = ~n6483 ;
  assign y2581 = ~1'b0 ;
  assign y2582 = ~n6491 ;
  assign y2583 = ~1'b0 ;
  assign y2584 = ~n6493 ;
  assign y2585 = ~n6494 ;
  assign y2586 = ~n6498 ;
  assign y2587 = ~n6500 ;
  assign y2588 = ~n6506 ;
  assign y2589 = ~n6507 ;
  assign y2590 = ~1'b0 ;
  assign y2591 = ~1'b0 ;
  assign y2592 = n6513 ;
  assign y2593 = n6514 ;
  assign y2594 = ~n6515 ;
  assign y2595 = n6516 ;
  assign y2596 = ~n6518 ;
  assign y2597 = n6525 ;
  assign y2598 = ~n6533 ;
  assign y2599 = ~n6541 ;
  assign y2600 = n6542 ;
  assign y2601 = n6543 ;
  assign y2602 = ~n6555 ;
  assign y2603 = ~n6565 ;
  assign y2604 = n6567 ;
  assign y2605 = n6573 ;
  assign y2606 = ~n6574 ;
  assign y2607 = ~1'b0 ;
  assign y2608 = n6575 ;
  assign y2609 = ~n6578 ;
  assign y2610 = n6589 ;
  assign y2611 = n6590 ;
  assign y2612 = n6196 ;
  assign y2613 = n6591 ;
  assign y2614 = ~n6592 ;
  assign y2615 = ~n6595 ;
  assign y2616 = x178 ;
  assign y2617 = n6596 ;
  assign y2618 = ~n6597 ;
  assign y2619 = ~1'b0 ;
  assign y2620 = n6605 ;
  assign y2621 = ~n6606 ;
  assign y2622 = 1'b0 ;
  assign y2623 = n6607 ;
  assign y2624 = ~1'b0 ;
  assign y2625 = n4750 ;
  assign y2626 = ~1'b0 ;
  assign y2627 = ~n6610 ;
  assign y2628 = n6615 ;
  assign y2629 = n6618 ;
  assign y2630 = n6623 ;
  assign y2631 = ~n6632 ;
  assign y2632 = ~1'b0 ;
  assign y2633 = n6640 ;
  assign y2634 = ~1'b0 ;
  assign y2635 = n3551 ;
  assign y2636 = n6646 ;
  assign y2637 = ~n6655 ;
  assign y2638 = ~1'b0 ;
  assign y2639 = ~n6658 ;
  assign y2640 = ~n6668 ;
  assign y2641 = ~1'b0 ;
  assign y2642 = ~n6672 ;
  assign y2643 = ~n6676 ;
  assign y2644 = n6677 ;
  assign y2645 = ~n6679 ;
  assign y2646 = n6683 ;
  assign y2647 = n6684 ;
  assign y2648 = ~n6686 ;
  assign y2649 = ~n6688 ;
  assign y2650 = n6693 ;
  assign y2651 = ~n6700 ;
  assign y2652 = n6703 ;
  assign y2653 = ~1'b0 ;
  assign y2654 = n6704 ;
  assign y2655 = n6705 ;
  assign y2656 = n6709 ;
  assign y2657 = n6711 ;
  assign y2658 = n6715 ;
  assign y2659 = ~n6719 ;
  assign y2660 = ~n6724 ;
  assign y2661 = n6726 ;
  assign y2662 = ~1'b0 ;
  assign y2663 = ~n6727 ;
  assign y2664 = n6730 ;
  assign y2665 = ~n6734 ;
  assign y2666 = ~1'b0 ;
  assign y2667 = n6739 ;
  assign y2668 = n6743 ;
  assign y2669 = ~n6747 ;
  assign y2670 = ~n6748 ;
  assign y2671 = ~n6749 ;
  assign y2672 = ~n6760 ;
  assign y2673 = ~1'b0 ;
  assign y2674 = n6762 ;
  assign y2675 = ~n6770 ;
  assign y2676 = n6771 ;
  assign y2677 = ~n6772 ;
  assign y2678 = ~n6773 ;
  assign y2679 = ~1'b0 ;
  assign y2680 = n6777 ;
  assign y2681 = ~n6780 ;
  assign y2682 = n650 ;
  assign y2683 = ~n6787 ;
  assign y2684 = n4962 ;
  assign y2685 = ~n6790 ;
  assign y2686 = ~1'b0 ;
  assign y2687 = ~n6795 ;
  assign y2688 = n6797 ;
  assign y2689 = ~1'b0 ;
  assign y2690 = ~n6801 ;
  assign y2691 = ~1'b0 ;
  assign y2692 = ~n6808 ;
  assign y2693 = n6810 ;
  assign y2694 = ~n6815 ;
  assign y2695 = n6816 ;
  assign y2696 = ~1'b0 ;
  assign y2697 = ~n6818 ;
  assign y2698 = ~n6820 ;
  assign y2699 = ~n6822 ;
  assign y2700 = ~n6676 ;
  assign y2701 = ~n6824 ;
  assign y2702 = n6825 ;
  assign y2703 = ~n6828 ;
  assign y2704 = ~1'b0 ;
  assign y2705 = ~n6830 ;
  assign y2706 = ~n6831 ;
  assign y2707 = ~n6834 ;
  assign y2708 = n6840 ;
  assign y2709 = ~1'b0 ;
  assign y2710 = n6841 ;
  assign y2711 = ~n6846 ;
  assign y2712 = n681 ;
  assign y2713 = n6849 ;
  assign y2714 = n6850 ;
  assign y2715 = n6851 ;
  assign y2716 = n6852 ;
  assign y2717 = ~n6853 ;
  assign y2718 = ~n6854 ;
  assign y2719 = n6866 ;
  assign y2720 = ~n6867 ;
  assign y2721 = ~n6868 ;
  assign y2722 = ~1'b0 ;
  assign y2723 = 1'b0 ;
  assign y2724 = ~n6869 ;
  assign y2725 = ~n6873 ;
  assign y2726 = ~n6877 ;
  assign y2727 = ~n6882 ;
  assign y2728 = ~n4518 ;
  assign y2729 = ~n6885 ;
  assign y2730 = n6889 ;
  assign y2731 = ~1'b0 ;
  assign y2732 = x247 ;
  assign y2733 = ~1'b0 ;
  assign y2734 = ~n6894 ;
  assign y2735 = n6898 ;
  assign y2736 = ~n6901 ;
  assign y2737 = n6903 ;
  assign y2738 = ~n6911 ;
  assign y2739 = n6914 ;
  assign y2740 = ~1'b0 ;
  assign y2741 = ~1'b0 ;
  assign y2742 = n6915 ;
  assign y2743 = n6920 ;
  assign y2744 = ~1'b0 ;
  assign y2745 = ~n6923 ;
  assign y2746 = n6931 ;
  assign y2747 = n5051 ;
  assign y2748 = ~n6934 ;
  assign y2749 = n6936 ;
  assign y2750 = ~1'b0 ;
  assign y2751 = n6938 ;
  assign y2752 = n6940 ;
  assign y2753 = ~n6949 ;
  assign y2754 = n6950 ;
  assign y2755 = ~n6952 ;
  assign y2756 = n6954 ;
  assign y2757 = n6955 ;
  assign y2758 = n6956 ;
  assign y2759 = ~n6958 ;
  assign y2760 = ~1'b0 ;
  assign y2761 = ~n6962 ;
  assign y2762 = n6966 ;
  assign y2763 = n6968 ;
  assign y2764 = ~n6969 ;
  assign y2765 = ~1'b0 ;
  assign y2766 = ~1'b0 ;
  assign y2767 = n6976 ;
  assign y2768 = ~n6979 ;
  assign y2769 = n6982 ;
  assign y2770 = ~1'b0 ;
  assign y2771 = n6984 ;
  assign y2772 = ~1'b0 ;
  assign y2773 = ~n6985 ;
  assign y2774 = ~n6986 ;
  assign y2775 = n6987 ;
  assign y2776 = ~1'b0 ;
  assign y2777 = ~n6988 ;
  assign y2778 = ~n6993 ;
  assign y2779 = ~1'b0 ;
  assign y2780 = ~n6994 ;
  assign y2781 = n6998 ;
  assign y2782 = ~n7003 ;
  assign y2783 = ~1'b0 ;
  assign y2784 = ~n7007 ;
  assign y2785 = ~n7008 ;
  assign y2786 = ~1'b0 ;
  assign y2787 = ~1'b0 ;
  assign y2788 = n5726 ;
  assign y2789 = n7013 ;
  assign y2790 = n6338 ;
  assign y2791 = n7016 ;
  assign y2792 = ~1'b0 ;
  assign y2793 = n7017 ;
  assign y2794 = ~n7019 ;
  assign y2795 = n7026 ;
  assign y2796 = ~n7027 ;
  assign y2797 = ~n7033 ;
  assign y2798 = ~1'b0 ;
  assign y2799 = 1'b0 ;
  assign y2800 = ~n7035 ;
  assign y2801 = ~n7036 ;
  assign y2802 = n7038 ;
  assign y2803 = n7039 ;
  assign y2804 = ~n7043 ;
  assign y2805 = n7046 ;
  assign y2806 = n7047 ;
  assign y2807 = n3088 ;
  assign y2808 = n1760 ;
  assign y2809 = n7049 ;
  assign y2810 = ~1'b0 ;
  assign y2811 = n7055 ;
  assign y2812 = n7058 ;
  assign y2813 = n7062 ;
  assign y2814 = ~1'b0 ;
  assign y2815 = ~1'b0 ;
  assign y2816 = ~n7068 ;
  assign y2817 = n7070 ;
  assign y2818 = ~n7071 ;
  assign y2819 = n7072 ;
  assign y2820 = n7074 ;
  assign y2821 = n7078 ;
  assign y2822 = ~1'b0 ;
  assign y2823 = ~n7081 ;
  assign y2824 = ~1'b0 ;
  assign y2825 = ~n7083 ;
  assign y2826 = ~n7086 ;
  assign y2827 = n7089 ;
  assign y2828 = ~1'b0 ;
  assign y2829 = n7090 ;
  assign y2830 = n7091 ;
  assign y2831 = n7102 ;
  assign y2832 = n7105 ;
  assign y2833 = n7113 ;
  assign y2834 = ~n7114 ;
  assign y2835 = ~n7118 ;
  assign y2836 = n7119 ;
  assign y2837 = ~1'b0 ;
  assign y2838 = ~n7122 ;
  assign y2839 = n7123 ;
  assign y2840 = n7126 ;
  assign y2841 = ~1'b0 ;
  assign y2842 = ~n7127 ;
  assign y2843 = n7130 ;
  assign y2844 = n7132 ;
  assign y2845 = ~n7135 ;
  assign y2846 = ~1'b0 ;
  assign y2847 = n7137 ;
  assign y2848 = n6068 ;
  assign y2849 = n7144 ;
  assign y2850 = n7145 ;
  assign y2851 = n7149 ;
  assign y2852 = ~n7154 ;
  assign y2853 = ~1'b0 ;
  assign y2854 = n7156 ;
  assign y2855 = n7160 ;
  assign y2856 = ~n7167 ;
  assign y2857 = n7169 ;
  assign y2858 = ~1'b0 ;
  assign y2859 = ~n7171 ;
  assign y2860 = ~n7174 ;
  assign y2861 = n7178 ;
  assign y2862 = ~1'b0 ;
  assign y2863 = ~1'b0 ;
  assign y2864 = n6768 ;
  assign y2865 = n4719 ;
  assign y2866 = ~1'b0 ;
  assign y2867 = n7184 ;
  assign y2868 = n7185 ;
  assign y2869 = n3791 ;
  assign y2870 = ~n7191 ;
  assign y2871 = ~1'b0 ;
  assign y2872 = n7196 ;
  assign y2873 = ~1'b0 ;
  assign y2874 = n7204 ;
  assign y2875 = n7209 ;
  assign y2876 = ~1'b0 ;
  assign y2877 = ~1'b0 ;
  assign y2878 = ~1'b0 ;
  assign y2879 = ~1'b0 ;
  assign y2880 = ~n7211 ;
  assign y2881 = ~1'b0 ;
  assign y2882 = n7216 ;
  assign y2883 = n7217 ;
  assign y2884 = ~n7225 ;
  assign y2885 = ~n7227 ;
  assign y2886 = ~n7233 ;
  assign y2887 = n7235 ;
  assign y2888 = n7241 ;
  assign y2889 = n1030 ;
  assign y2890 = n7246 ;
  assign y2891 = n7247 ;
  assign y2892 = ~n7252 ;
  assign y2893 = n7257 ;
  assign y2894 = n7258 ;
  assign y2895 = n7259 ;
  assign y2896 = ~1'b0 ;
  assign y2897 = ~n7262 ;
  assign y2898 = ~n7263 ;
  assign y2899 = ~n7265 ;
  assign y2900 = n7271 ;
  assign y2901 = n7274 ;
  assign y2902 = n7277 ;
  assign y2903 = ~n7278 ;
  assign y2904 = ~n7281 ;
  assign y2905 = ~1'b0 ;
  assign y2906 = ~n7282 ;
  assign y2907 = ~1'b0 ;
  assign y2908 = ~n7283 ;
  assign y2909 = ~n7291 ;
  assign y2910 = n7296 ;
  assign y2911 = n7297 ;
  assign y2912 = ~n7298 ;
  assign y2913 = ~n7300 ;
  assign y2914 = n7307 ;
  assign y2915 = n7308 ;
  assign y2916 = n7313 ;
  assign y2917 = ~1'b0 ;
  assign y2918 = ~1'b0 ;
  assign y2919 = ~n7314 ;
  assign y2920 = ~1'b0 ;
  assign y2921 = ~n7315 ;
  assign y2922 = ~1'b0 ;
  assign y2923 = n7318 ;
  assign y2924 = n7321 ;
  assign y2925 = n7327 ;
  assign y2926 = ~n7331 ;
  assign y2927 = ~n7335 ;
  assign y2928 = ~n7336 ;
  assign y2929 = ~n7341 ;
  assign y2930 = ~n7344 ;
  assign y2931 = ~1'b0 ;
  assign y2932 = ~n7346 ;
  assign y2933 = n7352 ;
  assign y2934 = n7360 ;
  assign y2935 = n7363 ;
  assign y2936 = ~n7365 ;
  assign y2937 = n7369 ;
  assign y2938 = ~n7370 ;
  assign y2939 = ~n7374 ;
  assign y2940 = ~1'b0 ;
  assign y2941 = ~n7376 ;
  assign y2942 = ~1'b0 ;
  assign y2943 = n7377 ;
  assign y2944 = ~1'b0 ;
  assign y2945 = ~n7380 ;
  assign y2946 = ~1'b0 ;
  assign y2947 = n7385 ;
  assign y2948 = ~n7390 ;
  assign y2949 = ~1'b0 ;
  assign y2950 = ~n7391 ;
  assign y2951 = ~n7394 ;
  assign y2952 = n7396 ;
  assign y2953 = n7399 ;
  assign y2954 = ~n7400 ;
  assign y2955 = ~n7403 ;
  assign y2956 = ~1'b0 ;
  assign y2957 = ~1'b0 ;
  assign y2958 = ~1'b0 ;
  assign y2959 = n7405 ;
  assign y2960 = ~n7409 ;
  assign y2961 = ~n7411 ;
  assign y2962 = n7415 ;
  assign y2963 = ~1'b0 ;
  assign y2964 = ~1'b0 ;
  assign y2965 = ~n7420 ;
  assign y2966 = ~n7423 ;
  assign y2967 = ~n7424 ;
  assign y2968 = n7426 ;
  assign y2969 = n7428 ;
  assign y2970 = ~1'b0 ;
  assign y2971 = n7429 ;
  assign y2972 = n7431 ;
  assign y2973 = ~n7436 ;
  assign y2974 = ~1'b0 ;
  assign y2975 = n7439 ;
  assign y2976 = ~n7445 ;
  assign y2977 = n7448 ;
  assign y2978 = ~1'b0 ;
  assign y2979 = ~n7450 ;
  assign y2980 = ~1'b0 ;
  assign y2981 = ~n7452 ;
  assign y2982 = ~1'b0 ;
  assign y2983 = n7453 ;
  assign y2984 = ~n7457 ;
  assign y2985 = ~1'b0 ;
  assign y2986 = ~1'b0 ;
  assign y2987 = ~1'b0 ;
  assign y2988 = ~n7463 ;
  assign y2989 = ~n7464 ;
  assign y2990 = ~n7465 ;
  assign y2991 = ~n1007 ;
  assign y2992 = ~n7471 ;
  assign y2993 = ~1'b0 ;
  assign y2994 = ~1'b0 ;
  assign y2995 = ~1'b0 ;
  assign y2996 = n7476 ;
  assign y2997 = n7480 ;
  assign y2998 = ~n7484 ;
  assign y2999 = ~1'b0 ;
  assign y3000 = ~n7485 ;
  assign y3001 = ~1'b0 ;
  assign y3002 = ~n7489 ;
  assign y3003 = ~n7500 ;
  assign y3004 = ~n7505 ;
  assign y3005 = n7507 ;
  assign y3006 = ~n7512 ;
  assign y3007 = n7518 ;
  assign y3008 = n7521 ;
  assign y3009 = ~1'b0 ;
  assign y3010 = ~1'b0 ;
  assign y3011 = ~n7522 ;
  assign y3012 = ~n7525 ;
  assign y3013 = n7530 ;
  assign y3014 = n6643 ;
  assign y3015 = ~n7534 ;
  assign y3016 = n7535 ;
  assign y3017 = ~n7538 ;
  assign y3018 = ~1'b0 ;
  assign y3019 = 1'b0 ;
  assign y3020 = n7542 ;
  assign y3021 = n7546 ;
  assign y3022 = n7558 ;
  assign y3023 = n7560 ;
  assign y3024 = n2963 ;
  assign y3025 = ~1'b0 ;
  assign y3026 = n7568 ;
  assign y3027 = ~1'b0 ;
  assign y3028 = n7570 ;
  assign y3029 = n7572 ;
  assign y3030 = n7575 ;
  assign y3031 = ~n7576 ;
  assign y3032 = n7581 ;
  assign y3033 = n3439 ;
  assign y3034 = n7583 ;
  assign y3035 = n7585 ;
  assign y3036 = ~1'b0 ;
  assign y3037 = ~1'b0 ;
  assign y3038 = ~n7601 ;
  assign y3039 = n7602 ;
  assign y3040 = ~n7604 ;
  assign y3041 = 1'b0 ;
  assign y3042 = n7609 ;
  assign y3043 = ~n7619 ;
  assign y3044 = n7622 ;
  assign y3045 = ~1'b0 ;
  assign y3046 = n7627 ;
  assign y3047 = ~1'b0 ;
  assign y3048 = n4442 ;
  assign y3049 = n7630 ;
  assign y3050 = n7633 ;
  assign y3051 = n5278 ;
  assign y3052 = ~n7645 ;
  assign y3053 = ~n7647 ;
  assign y3054 = ~1'b0 ;
  assign y3055 = ~1'b0 ;
  assign y3056 = ~n7650 ;
  assign y3057 = ~n7656 ;
  assign y3058 = ~1'b0 ;
  assign y3059 = ~n7663 ;
  assign y3060 = ~n7664 ;
  assign y3061 = ~n7667 ;
  assign y3062 = ~n7671 ;
  assign y3063 = n7677 ;
  assign y3064 = ~n7679 ;
  assign y3065 = n7680 ;
  assign y3066 = ~n7682 ;
  assign y3067 = n7683 ;
  assign y3068 = ~n7688 ;
  assign y3069 = ~1'b0 ;
  assign y3070 = n7694 ;
  assign y3071 = n7696 ;
  assign y3072 = ~1'b0 ;
  assign y3073 = ~1'b0 ;
  assign y3074 = ~n7700 ;
  assign y3075 = n7701 ;
  assign y3076 = ~n7706 ;
  assign y3077 = ~n7710 ;
  assign y3078 = ~n7711 ;
  assign y3079 = ~n7713 ;
  assign y3080 = n7714 ;
  assign y3081 = n7715 ;
  assign y3082 = ~n7716 ;
  assign y3083 = ~n7718 ;
  assign y3084 = n7719 ;
  assign y3085 = ~1'b0 ;
  assign y3086 = n7723 ;
  assign y3087 = n7727 ;
  assign y3088 = ~1'b0 ;
  assign y3089 = ~1'b0 ;
  assign y3090 = ~1'b0 ;
  assign y3091 = ~n7729 ;
  assign y3092 = ~n7732 ;
  assign y3093 = n7735 ;
  assign y3094 = n7737 ;
  assign y3095 = ~n7739 ;
  assign y3096 = ~n7741 ;
  assign y3097 = ~n7746 ;
  assign y3098 = n7749 ;
  assign y3099 = ~n7750 ;
  assign y3100 = ~n7753 ;
  assign y3101 = ~n7758 ;
  assign y3102 = ~n7761 ;
  assign y3103 = ~1'b0 ;
  assign y3104 = ~n7765 ;
  assign y3105 = n7766 ;
  assign y3106 = n7771 ;
  assign y3107 = ~1'b0 ;
  assign y3108 = ~n7776 ;
  assign y3109 = n7777 ;
  assign y3110 = ~n7786 ;
  assign y3111 = n7790 ;
  assign y3112 = ~n7791 ;
  assign y3113 = n7793 ;
  assign y3114 = ~n7794 ;
  assign y3115 = ~n7795 ;
  assign y3116 = n7798 ;
  assign y3117 = ~n7806 ;
  assign y3118 = n7813 ;
  assign y3119 = ~1'b0 ;
  assign y3120 = ~n7814 ;
  assign y3121 = ~n7822 ;
  assign y3122 = ~n7831 ;
  assign y3123 = ~n7846 ;
  assign y3124 = n7853 ;
  assign y3125 = n7854 ;
  assign y3126 = n7864 ;
  assign y3127 = ~n7866 ;
  assign y3128 = x97 ;
  assign y3129 = n7870 ;
  assign y3130 = ~n7873 ;
  assign y3131 = ~n7876 ;
  assign y3132 = ~n7879 ;
  assign y3133 = ~1'b0 ;
  assign y3134 = n7883 ;
  assign y3135 = ~1'b0 ;
  assign y3136 = n5850 ;
  assign y3137 = ~n7886 ;
  assign y3138 = x241 ;
  assign y3139 = ~1'b0 ;
  assign y3140 = ~1'b0 ;
  assign y3141 = ~n7887 ;
  assign y3142 = ~1'b0 ;
  assign y3143 = ~n7895 ;
  assign y3144 = ~1'b0 ;
  assign y3145 = ~1'b0 ;
  assign y3146 = n7899 ;
  assign y3147 = ~1'b0 ;
  assign y3148 = n7901 ;
  assign y3149 = n7903 ;
  assign y3150 = n7905 ;
  assign y3151 = ~1'b0 ;
  assign y3152 = ~1'b0 ;
  assign y3153 = ~n7906 ;
  assign y3154 = ~1'b0 ;
  assign y3155 = ~n7912 ;
  assign y3156 = n7915 ;
  assign y3157 = ~1'b0 ;
  assign y3158 = n7918 ;
  assign y3159 = ~1'b0 ;
  assign y3160 = n7921 ;
  assign y3161 = ~n7922 ;
  assign y3162 = ~n7924 ;
  assign y3163 = ~n7928 ;
  assign y3164 = ~n7932 ;
  assign y3165 = ~n7935 ;
  assign y3166 = ~1'b0 ;
  assign y3167 = ~n7936 ;
  assign y3168 = ~n7940 ;
  assign y3169 = ~n7941 ;
  assign y3170 = n7944 ;
  assign y3171 = ~1'b0 ;
  assign y3172 = n7954 ;
  assign y3173 = n7957 ;
  assign y3174 = n7958 ;
  assign y3175 = ~1'b0 ;
  assign y3176 = ~n952 ;
  assign y3177 = ~1'b0 ;
  assign y3178 = ~1'b0 ;
  assign y3179 = ~1'b0 ;
  assign y3180 = ~n4917 ;
  assign y3181 = n7962 ;
  assign y3182 = ~n7969 ;
  assign y3183 = ~n7970 ;
  assign y3184 = n7971 ;
  assign y3185 = n7972 ;
  assign y3186 = ~n7975 ;
  assign y3187 = n7983 ;
  assign y3188 = n7986 ;
  assign y3189 = n1524 ;
  assign y3190 = n7999 ;
  assign y3191 = ~n8000 ;
  assign y3192 = ~1'b0 ;
  assign y3193 = ~n8005 ;
  assign y3194 = ~1'b0 ;
  assign y3195 = ~1'b0 ;
  assign y3196 = ~n8009 ;
  assign y3197 = ~n8014 ;
  assign y3198 = n8017 ;
  assign y3199 = ~1'b0 ;
  assign y3200 = n8018 ;
  assign y3201 = ~n727 ;
  assign y3202 = n8024 ;
  assign y3203 = n8027 ;
  assign y3204 = n8030 ;
  assign y3205 = ~n8038 ;
  assign y3206 = ~n8039 ;
  assign y3207 = ~n8040 ;
  assign y3208 = ~n8041 ;
  assign y3209 = ~n8042 ;
  assign y3210 = n8044 ;
  assign y3211 = ~n8046 ;
  assign y3212 = n8048 ;
  assign y3213 = ~1'b0 ;
  assign y3214 = ~n8052 ;
  assign y3215 = ~1'b0 ;
  assign y3216 = ~n8054 ;
  assign y3217 = ~1'b0 ;
  assign y3218 = n8060 ;
  assign y3219 = ~n8064 ;
  assign y3220 = ~1'b0 ;
  assign y3221 = n8071 ;
  assign y3222 = ~n8076 ;
  assign y3223 = ~n8080 ;
  assign y3224 = ~n8081 ;
  assign y3225 = ~n8084 ;
  assign y3226 = n8085 ;
  assign y3227 = ~1'b0 ;
  assign y3228 = n8087 ;
  assign y3229 = ~n8088 ;
  assign y3230 = ~n8090 ;
  assign y3231 = n8091 ;
  assign y3232 = n8100 ;
  assign y3233 = ~n8107 ;
  assign y3234 = ~n8112 ;
  assign y3235 = ~1'b0 ;
  assign y3236 = n8114 ;
  assign y3237 = ~n8118 ;
  assign y3238 = n8120 ;
  assign y3239 = ~1'b0 ;
  assign y3240 = ~n8121 ;
  assign y3241 = ~n8122 ;
  assign y3242 = ~n8123 ;
  assign y3243 = ~n8124 ;
  assign y3244 = n8130 ;
  assign y3245 = n8137 ;
  assign y3246 = n8138 ;
  assign y3247 = n8139 ;
  assign y3248 = ~n8140 ;
  assign y3249 = ~x237 ;
  assign y3250 = ~1'b0 ;
  assign y3251 = ~n8144 ;
  assign y3252 = ~1'b0 ;
  assign y3253 = ~n8149 ;
  assign y3254 = n6153 ;
  assign y3255 = ~1'b0 ;
  assign y3256 = n8153 ;
  assign y3257 = n8154 ;
  assign y3258 = n8158 ;
  assign y3259 = ~n8161 ;
  assign y3260 = ~n8163 ;
  assign y3261 = n8165 ;
  assign y3262 = n8171 ;
  assign y3263 = n8173 ;
  assign y3264 = n8176 ;
  assign y3265 = ~1'b0 ;
  assign y3266 = 1'b0 ;
  assign y3267 = ~1'b0 ;
  assign y3268 = ~1'b0 ;
  assign y3269 = n6683 ;
  assign y3270 = n8190 ;
  assign y3271 = n8194 ;
  assign y3272 = ~1'b0 ;
  assign y3273 = n8195 ;
  assign y3274 = n8198 ;
  assign y3275 = n8203 ;
  assign y3276 = ~1'b0 ;
  assign y3277 = n8216 ;
  assign y3278 = ~n8217 ;
  assign y3279 = n8218 ;
  assign y3280 = ~1'b0 ;
  assign y3281 = n8219 ;
  assign y3282 = ~n8220 ;
  assign y3283 = n8227 ;
  assign y3284 = n8233 ;
  assign y3285 = n8243 ;
  assign y3286 = 1'b0 ;
  assign y3287 = ~n8244 ;
  assign y3288 = n8246 ;
  assign y3289 = ~n6754 ;
  assign y3290 = ~1'b0 ;
  assign y3291 = n8251 ;
  assign y3292 = ~n8253 ;
  assign y3293 = ~1'b0 ;
  assign y3294 = ~n8257 ;
  assign y3295 = ~n8261 ;
  assign y3296 = n8262 ;
  assign y3297 = ~1'b0 ;
  assign y3298 = ~n8265 ;
  assign y3299 = n8271 ;
  assign y3300 = n8275 ;
  assign y3301 = ~1'b0 ;
  assign y3302 = n8276 ;
  assign y3303 = ~1'b0 ;
  assign y3304 = n8282 ;
  assign y3305 = ~n8283 ;
  assign y3306 = ~1'b0 ;
  assign y3307 = ~n8284 ;
  assign y3308 = n8287 ;
  assign y3309 = ~1'b0 ;
  assign y3310 = ~1'b0 ;
  assign y3311 = n8293 ;
  assign y3312 = ~n674 ;
  assign y3313 = ~n8294 ;
  assign y3314 = ~n8298 ;
  assign y3315 = ~1'b0 ;
  assign y3316 = n8299 ;
  assign y3317 = n5415 ;
  assign y3318 = ~1'b0 ;
  assign y3319 = ~1'b0 ;
  assign y3320 = ~n8301 ;
  assign y3321 = ~n8302 ;
  assign y3322 = ~1'b0 ;
  assign y3323 = 1'b0 ;
  assign y3324 = n8303 ;
  assign y3325 = 1'b0 ;
  assign y3326 = n8307 ;
  assign y3327 = ~n8311 ;
  assign y3328 = ~n8314 ;
  assign y3329 = ~n8316 ;
  assign y3330 = ~n8319 ;
  assign y3331 = n4797 ;
  assign y3332 = n8320 ;
  assign y3333 = ~n8321 ;
  assign y3334 = ~1'b0 ;
  assign y3335 = ~n8323 ;
  assign y3336 = ~n8324 ;
  assign y3337 = ~n8325 ;
  assign y3338 = ~1'b0 ;
  assign y3339 = n8327 ;
  assign y3340 = ~n8329 ;
  assign y3341 = n8336 ;
  assign y3342 = ~1'b0 ;
  assign y3343 = 1'b0 ;
  assign y3344 = ~1'b0 ;
  assign y3345 = n8339 ;
  assign y3346 = ~n8340 ;
  assign y3347 = ~1'b0 ;
  assign y3348 = ~1'b0 ;
  assign y3349 = n8345 ;
  assign y3350 = n8346 ;
  assign y3351 = n8350 ;
  assign y3352 = ~n8352 ;
  assign y3353 = n4828 ;
  assign y3354 = ~n8358 ;
  assign y3355 = ~n8362 ;
  assign y3356 = ~n8364 ;
  assign y3357 = n8367 ;
  assign y3358 = n2249 ;
  assign y3359 = ~n8369 ;
  assign y3360 = ~n8376 ;
  assign y3361 = ~1'b0 ;
  assign y3362 = n8377 ;
  assign y3363 = ~n8378 ;
  assign y3364 = n8382 ;
  assign y3365 = n8384 ;
  assign y3366 = ~1'b0 ;
  assign y3367 = ~1'b0 ;
  assign y3368 = n8387 ;
  assign y3369 = n8390 ;
  assign y3370 = n8391 ;
  assign y3371 = ~n8393 ;
  assign y3372 = ~n8395 ;
  assign y3373 = ~n8399 ;
  assign y3374 = n8408 ;
  assign y3375 = ~n8409 ;
  assign y3376 = n8411 ;
  assign y3377 = ~1'b0 ;
  assign y3378 = 1'b0 ;
  assign y3379 = ~1'b0 ;
  assign y3380 = ~n8419 ;
  assign y3381 = n8420 ;
  assign y3382 = ~n8423 ;
  assign y3383 = ~1'b0 ;
  assign y3384 = n8424 ;
  assign y3385 = n8428 ;
  assign y3386 = ~1'b0 ;
  assign y3387 = n8432 ;
  assign y3388 = n8433 ;
  assign y3389 = ~n8435 ;
  assign y3390 = ~1'b0 ;
  assign y3391 = ~n8445 ;
  assign y3392 = ~n8450 ;
  assign y3393 = n8451 ;
  assign y3394 = ~1'b0 ;
  assign y3395 = n8457 ;
  assign y3396 = ~n8463 ;
  assign y3397 = n8468 ;
  assign y3398 = ~n3659 ;
  assign y3399 = n7532 ;
  assign y3400 = ~n8470 ;
  assign y3401 = ~1'b0 ;
  assign y3402 = n8478 ;
  assign y3403 = ~1'b0 ;
  assign y3404 = n8481 ;
  assign y3405 = n8482 ;
  assign y3406 = ~n8493 ;
  assign y3407 = n8494 ;
  assign y3408 = n8496 ;
  assign y3409 = n8497 ;
  assign y3410 = n8501 ;
  assign y3411 = n8505 ;
  assign y3412 = ~1'b0 ;
  assign y3413 = n8509 ;
  assign y3414 = n8510 ;
  assign y3415 = n8513 ;
  assign y3416 = ~1'b0 ;
  assign y3417 = ~n8517 ;
  assign y3418 = n8521 ;
  assign y3419 = ~1'b0 ;
  assign y3420 = ~n8524 ;
  assign y3421 = n8526 ;
  assign y3422 = ~n8528 ;
  assign y3423 = ~1'b0 ;
  assign y3424 = n8542 ;
  assign y3425 = ~n8548 ;
  assign y3426 = ~n8550 ;
  assign y3427 = ~n8557 ;
  assign y3428 = ~n8558 ;
  assign y3429 = ~1'b0 ;
  assign y3430 = n8560 ;
  assign y3431 = ~n8567 ;
  assign y3432 = ~n8570 ;
  assign y3433 = ~n8575 ;
  assign y3434 = n8577 ;
  assign y3435 = ~n8578 ;
  assign y3436 = n8581 ;
  assign y3437 = ~n8583 ;
  assign y3438 = ~1'b0 ;
  assign y3439 = ~n8584 ;
  assign y3440 = ~n8585 ;
  assign y3441 = ~1'b0 ;
  assign y3442 = n8587 ;
  assign y3443 = ~n8592 ;
  assign y3444 = ~n8602 ;
  assign y3445 = ~n8605 ;
  assign y3446 = ~n8610 ;
  assign y3447 = n8614 ;
  assign y3448 = n8621 ;
  assign y3449 = ~1'b0 ;
  assign y3450 = ~1'b0 ;
  assign y3451 = ~n8623 ;
  assign y3452 = ~n8635 ;
  assign y3453 = n8636 ;
  assign y3454 = ~n8637 ;
  assign y3455 = n8639 ;
  assign y3456 = ~1'b0 ;
  assign y3457 = ~n563 ;
  assign y3458 = n8642 ;
  assign y3459 = ~n8643 ;
  assign y3460 = ~n8651 ;
  assign y3461 = n8653 ;
  assign y3462 = n8655 ;
  assign y3463 = ~n8657 ;
  assign y3464 = 1'b0 ;
  assign y3465 = n8659 ;
  assign y3466 = ~1'b0 ;
  assign y3467 = x65 ;
  assign y3468 = n8664 ;
  assign y3469 = n8669 ;
  assign y3470 = n8674 ;
  assign y3471 = n8677 ;
  assign y3472 = n8678 ;
  assign y3473 = ~n8680 ;
  assign y3474 = ~1'b0 ;
  assign y3475 = ~n8684 ;
  assign y3476 = ~n8686 ;
  assign y3477 = ~n8691 ;
  assign y3478 = ~n8692 ;
  assign y3479 = ~n8694 ;
  assign y3480 = ~1'b0 ;
  assign y3481 = ~n8696 ;
  assign y3482 = ~1'b0 ;
  assign y3483 = n8697 ;
  assign y3484 = ~n8699 ;
  assign y3485 = ~1'b0 ;
  assign y3486 = ~n8704 ;
  assign y3487 = ~n8705 ;
  assign y3488 = ~1'b0 ;
  assign y3489 = ~n8708 ;
  assign y3490 = n8709 ;
  assign y3491 = ~n8712 ;
  assign y3492 = n8716 ;
  assign y3493 = n8720 ;
  assign y3494 = n1304 ;
  assign y3495 = ~n8739 ;
  assign y3496 = ~n8746 ;
  assign y3497 = n8752 ;
  assign y3498 = ~1'b0 ;
  assign y3499 = ~n8754 ;
  assign y3500 = n8762 ;
  assign y3501 = ~n8769 ;
  assign y3502 = ~n8772 ;
  assign y3503 = ~n8775 ;
  assign y3504 = ~1'b0 ;
  assign y3505 = 1'b0 ;
  assign y3506 = n8780 ;
  assign y3507 = n8782 ;
  assign y3508 = n8787 ;
  assign y3509 = n8790 ;
  assign y3510 = ~n8793 ;
  assign y3511 = n8799 ;
  assign y3512 = 1'b0 ;
  assign y3513 = ~n8802 ;
  assign y3514 = ~n5988 ;
  assign y3515 = n8805 ;
  assign y3516 = ~n8807 ;
  assign y3517 = n8808 ;
  assign y3518 = n1440 ;
  assign y3519 = 1'b0 ;
  assign y3520 = ~n8811 ;
  assign y3521 = n8817 ;
  assign y3522 = n8819 ;
  assign y3523 = ~1'b0 ;
  assign y3524 = n8820 ;
  assign y3525 = n8824 ;
  assign y3526 = ~n8825 ;
  assign y3527 = n8826 ;
  assign y3528 = n8834 ;
  assign y3529 = n8836 ;
  assign y3530 = n8839 ;
  assign y3531 = ~1'b0 ;
  assign y3532 = ~n8844 ;
  assign y3533 = n8845 ;
  assign y3534 = n8848 ;
  assign y3535 = ~n8855 ;
  assign y3536 = ~1'b0 ;
  assign y3537 = ~1'b0 ;
  assign y3538 = ~1'b0 ;
  assign y3539 = ~1'b0 ;
  assign y3540 = ~n8856 ;
  assign y3541 = ~n8862 ;
  assign y3542 = ~1'b0 ;
  assign y3543 = ~n8865 ;
  assign y3544 = ~n8877 ;
  assign y3545 = n8880 ;
  assign y3546 = n8882 ;
  assign y3547 = n8884 ;
  assign y3548 = n8888 ;
  assign y3549 = ~1'b0 ;
  assign y3550 = ~1'b0 ;
  assign y3551 = ~n8889 ;
  assign y3552 = ~1'b0 ;
  assign y3553 = n8892 ;
  assign y3554 = n8894 ;
  assign y3555 = n8895 ;
  assign y3556 = ~1'b0 ;
  assign y3557 = n8901 ;
  assign y3558 = n8903 ;
  assign y3559 = ~1'b0 ;
  assign y3560 = ~1'b0 ;
  assign y3561 = ~n8906 ;
  assign y3562 = ~n8911 ;
  assign y3563 = ~1'b0 ;
  assign y3564 = ~n8914 ;
  assign y3565 = ~n8923 ;
  assign y3566 = n8927 ;
  assign y3567 = ~1'b0 ;
  assign y3568 = ~n8929 ;
  assign y3569 = n8931 ;
  assign y3570 = ~n7962 ;
  assign y3571 = ~n8932 ;
  assign y3572 = ~n8936 ;
  assign y3573 = ~1'b0 ;
  assign y3574 = n8940 ;
  assign y3575 = n8941 ;
  assign y3576 = ~n8944 ;
  assign y3577 = n8945 ;
  assign y3578 = n8948 ;
  assign y3579 = ~n8951 ;
  assign y3580 = ~n8956 ;
  assign y3581 = ~n8959 ;
  assign y3582 = ~n8961 ;
  assign y3583 = ~n8963 ;
  assign y3584 = n8965 ;
  assign y3585 = ~1'b0 ;
  assign y3586 = n8966 ;
  assign y3587 = ~1'b0 ;
  assign y3588 = n8974 ;
  assign y3589 = n8977 ;
  assign y3590 = ~n8988 ;
  assign y3591 = ~1'b0 ;
  assign y3592 = ~1'b0 ;
  assign y3593 = n1582 ;
  assign y3594 = ~1'b0 ;
  assign y3595 = ~n8990 ;
  assign y3596 = ~n8993 ;
  assign y3597 = n8994 ;
  assign y3598 = n8995 ;
  assign y3599 = ~n8998 ;
  assign y3600 = n3229 ;
  assign y3601 = ~1'b0 ;
  assign y3602 = ~n9001 ;
  assign y3603 = ~n9002 ;
  assign y3604 = ~1'b0 ;
  assign y3605 = ~n9014 ;
  assign y3606 = ~n9015 ;
  assign y3607 = n9020 ;
  assign y3608 = ~n9024 ;
  assign y3609 = n9027 ;
  assign y3610 = ~1'b0 ;
  assign y3611 = ~n9030 ;
  assign y3612 = n9033 ;
  assign y3613 = ~n9034 ;
  assign y3614 = ~1'b0 ;
  assign y3615 = ~n9035 ;
  assign y3616 = n9040 ;
  assign y3617 = ~1'b0 ;
  assign y3618 = ~1'b0 ;
  assign y3619 = n9044 ;
  assign y3620 = n9047 ;
  assign y3621 = n9048 ;
  assign y3622 = ~n9051 ;
  assign y3623 = ~n9052 ;
  assign y3624 = ~n9054 ;
  assign y3625 = n9056 ;
  assign y3626 = ~n9057 ;
  assign y3627 = n9058 ;
  assign y3628 = ~1'b0 ;
  assign y3629 = n9059 ;
  assign y3630 = n9062 ;
  assign y3631 = n9064 ;
  assign y3632 = ~n9065 ;
  assign y3633 = n9066 ;
  assign y3634 = n9069 ;
  assign y3635 = ~n9070 ;
  assign y3636 = ~1'b0 ;
  assign y3637 = ~n9075 ;
  assign y3638 = ~n9081 ;
  assign y3639 = n8386 ;
  assign y3640 = n9083 ;
  assign y3641 = n9087 ;
  assign y3642 = n9094 ;
  assign y3643 = ~n9096 ;
  assign y3644 = ~n9104 ;
  assign y3645 = ~n9105 ;
  assign y3646 = ~1'b0 ;
  assign y3647 = n9110 ;
  assign y3648 = n9111 ;
  assign y3649 = ~1'b0 ;
  assign y3650 = ~1'b0 ;
  assign y3651 = ~1'b0 ;
  assign y3652 = n9112 ;
  assign y3653 = ~n9119 ;
  assign y3654 = n9121 ;
  assign y3655 = ~n9130 ;
  assign y3656 = ~n9132 ;
  assign y3657 = n6302 ;
  assign y3658 = ~n9134 ;
  assign y3659 = ~n9137 ;
  assign y3660 = ~n9141 ;
  assign y3661 = n9144 ;
  assign y3662 = n9146 ;
  assign y3663 = n9151 ;
  assign y3664 = n9152 ;
  assign y3665 = ~n9153 ;
  assign y3666 = ~n9154 ;
  assign y3667 = ~n9155 ;
  assign y3668 = n9156 ;
  assign y3669 = ~1'b0 ;
  assign y3670 = ~1'b0 ;
  assign y3671 = n9164 ;
  assign y3672 = n9169 ;
  assign y3673 = n9170 ;
  assign y3674 = ~1'b0 ;
  assign y3675 = ~n9172 ;
  assign y3676 = ~1'b0 ;
  assign y3677 = ~1'b0 ;
  assign y3678 = ~n9174 ;
  assign y3679 = ~n9187 ;
  assign y3680 = ~n9194 ;
  assign y3681 = ~n9195 ;
  assign y3682 = ~n9204 ;
  assign y3683 = n9209 ;
  assign y3684 = n9212 ;
  assign y3685 = n9213 ;
  assign y3686 = ~n9214 ;
  assign y3687 = 1'b0 ;
  assign y3688 = n5914 ;
  assign y3689 = n9217 ;
  assign y3690 = ~1'b0 ;
  assign y3691 = ~n3922 ;
  assign y3692 = ~1'b0 ;
  assign y3693 = ~1'b0 ;
  assign y3694 = n9219 ;
  assign y3695 = n7785 ;
  assign y3696 = ~1'b0 ;
  assign y3697 = ~1'b0 ;
  assign y3698 = ~1'b0 ;
  assign y3699 = ~1'b0 ;
  assign y3700 = n9233 ;
  assign y3701 = n319 ;
  assign y3702 = n9234 ;
  assign y3703 = n9239 ;
  assign y3704 = n9242 ;
  assign y3705 = n9245 ;
  assign y3706 = ~n9249 ;
  assign y3707 = ~1'b0 ;
  assign y3708 = ~n9251 ;
  assign y3709 = ~1'b0 ;
  assign y3710 = ~n9252 ;
  assign y3711 = ~n9257 ;
  assign y3712 = ~n9261 ;
  assign y3713 = ~n9269 ;
  assign y3714 = n9274 ;
  assign y3715 = ~1'b0 ;
  assign y3716 = ~1'b0 ;
  assign y3717 = n9278 ;
  assign y3718 = n9282 ;
  assign y3719 = ~n9287 ;
  assign y3720 = n867 ;
  assign y3721 = ~n9292 ;
  assign y3722 = n6232 ;
  assign y3723 = n9293 ;
  assign y3724 = n9296 ;
  assign y3725 = ~n9297 ;
  assign y3726 = ~n9300 ;
  assign y3727 = ~1'b0 ;
  assign y3728 = n9305 ;
  assign y3729 = n9309 ;
  assign y3730 = ~n9313 ;
  assign y3731 = n9318 ;
  assign y3732 = 1'b0 ;
  assign y3733 = ~n9324 ;
  assign y3734 = ~1'b0 ;
  assign y3735 = ~1'b0 ;
  assign y3736 = ~1'b0 ;
  assign y3737 = n2829 ;
  assign y3738 = ~1'b0 ;
  assign y3739 = ~n9327 ;
  assign y3740 = ~1'b0 ;
  assign y3741 = ~n9329 ;
  assign y3742 = ~n9333 ;
  assign y3743 = n9340 ;
  assign y3744 = n9345 ;
  assign y3745 = ~1'b0 ;
  assign y3746 = ~n9347 ;
  assign y3747 = ~n9349 ;
  assign y3748 = ~n9356 ;
  assign y3749 = ~n9359 ;
  assign y3750 = ~n9361 ;
  assign y3751 = n9362 ;
  assign y3752 = ~n9363 ;
  assign y3753 = ~1'b0 ;
  assign y3754 = n9366 ;
  assign y3755 = 1'b0 ;
  assign y3756 = ~n9367 ;
  assign y3757 = n9369 ;
  assign y3758 = ~1'b0 ;
  assign y3759 = n9373 ;
  assign y3760 = n9381 ;
  assign y3761 = n9385 ;
  assign y3762 = ~n9387 ;
  assign y3763 = ~1'b0 ;
  assign y3764 = n9394 ;
  assign y3765 = n9401 ;
  assign y3766 = n9402 ;
  assign y3767 = ~1'b0 ;
  assign y3768 = n9404 ;
  assign y3769 = n9409 ;
  assign y3770 = ~1'b0 ;
  assign y3771 = ~n9418 ;
  assign y3772 = ~n9420 ;
  assign y3773 = ~n9421 ;
  assign y3774 = ~n9422 ;
  assign y3775 = ~n9423 ;
  assign y3776 = n9427 ;
  assign y3777 = n9429 ;
  assign y3778 = ~n9431 ;
  assign y3779 = ~n9437 ;
  assign y3780 = ~1'b0 ;
  assign y3781 = n9440 ;
  assign y3782 = ~n9442 ;
  assign y3783 = n9444 ;
  assign y3784 = ~n9445 ;
  assign y3785 = n9447 ;
  assign y3786 = ~1'b0 ;
  assign y3787 = n9448 ;
  assign y3788 = ~n9450 ;
  assign y3789 = ~n9455 ;
  assign y3790 = ~1'b0 ;
  assign y3791 = n9456 ;
  assign y3792 = ~1'b0 ;
  assign y3793 = ~n9465 ;
  assign y3794 = 1'b0 ;
  assign y3795 = ~1'b0 ;
  assign y3796 = n9471 ;
  assign y3797 = ~n9476 ;
  assign y3798 = n9488 ;
  assign y3799 = ~1'b0 ;
  assign y3800 = n9496 ;
  assign y3801 = n9497 ;
  assign y3802 = ~n9504 ;
  assign y3803 = ~n9510 ;
  assign y3804 = ~1'b0 ;
  assign y3805 = ~n9514 ;
  assign y3806 = n9515 ;
  assign y3807 = ~1'b0 ;
  assign y3808 = n9517 ;
  assign y3809 = ~1'b0 ;
  assign y3810 = ~1'b0 ;
  assign y3811 = n9524 ;
  assign y3812 = n1961 ;
  assign y3813 = ~1'b0 ;
  assign y3814 = ~1'b0 ;
  assign y3815 = n9527 ;
  assign y3816 = n9528 ;
  assign y3817 = n9529 ;
  assign y3818 = ~n9532 ;
  assign y3819 = ~1'b0 ;
  assign y3820 = ~1'b0 ;
  assign y3821 = n9535 ;
  assign y3822 = ~n9538 ;
  assign y3823 = n9541 ;
  assign y3824 = n9546 ;
  assign y3825 = ~1'b0 ;
  assign y3826 = n9550 ;
  assign y3827 = ~n9553 ;
  assign y3828 = n9555 ;
  assign y3829 = n9559 ;
  assign y3830 = ~n9564 ;
  assign y3831 = ~1'b0 ;
  assign y3832 = n9567 ;
  assign y3833 = n9568 ;
  assign y3834 = n9569 ;
  assign y3835 = ~1'b0 ;
  assign y3836 = n9575 ;
  assign y3837 = n9577 ;
  assign y3838 = ~1'b0 ;
  assign y3839 = ~n9581 ;
  assign y3840 = n9583 ;
  assign y3841 = n9585 ;
  assign y3842 = ~n9588 ;
  assign y3843 = n9592 ;
  assign y3844 = n9595 ;
  assign y3845 = ~1'b0 ;
  assign y3846 = ~n9599 ;
  assign y3847 = n9601 ;
  assign y3848 = ~n9603 ;
  assign y3849 = ~1'b0 ;
  assign y3850 = ~1'b0 ;
  assign y3851 = n9605 ;
  assign y3852 = n9610 ;
  assign y3853 = ~1'b0 ;
  assign y3854 = ~n9611 ;
  assign y3855 = ~n9613 ;
  assign y3856 = ~1'b0 ;
  assign y3857 = ~1'b0 ;
  assign y3858 = n9616 ;
  assign y3859 = ~1'b0 ;
  assign y3860 = ~n9619 ;
  assign y3861 = ~n9622 ;
  assign y3862 = ~1'b0 ;
  assign y3863 = ~1'b0 ;
  assign y3864 = ~n9623 ;
  assign y3865 = ~n9629 ;
  assign y3866 = ~1'b0 ;
  assign y3867 = ~1'b0 ;
  assign y3868 = ~n9634 ;
  assign y3869 = ~n9636 ;
  assign y3870 = n9645 ;
  assign y3871 = ~n9646 ;
  assign y3872 = ~1'b0 ;
  assign y3873 = n9655 ;
  assign y3874 = n9661 ;
  assign y3875 = ~n9663 ;
  assign y3876 = n9665 ;
  assign y3877 = ~1'b0 ;
  assign y3878 = n9670 ;
  assign y3879 = ~n9674 ;
  assign y3880 = ~1'b0 ;
  assign y3881 = ~n9675 ;
  assign y3882 = ~n9686 ;
  assign y3883 = ~n8411 ;
  assign y3884 = ~n9689 ;
  assign y3885 = ~1'b0 ;
  assign y3886 = n9692 ;
  assign y3887 = n9694 ;
  assign y3888 = n9700 ;
  assign y3889 = ~1'b0 ;
  assign y3890 = ~1'b0 ;
  assign y3891 = n9701 ;
  assign y3892 = n9704 ;
  assign y3893 = n9708 ;
  assign y3894 = ~1'b0 ;
  assign y3895 = ~n9714 ;
  assign y3896 = n9581 ;
  assign y3897 = ~n9715 ;
  assign y3898 = n9726 ;
  assign y3899 = n9727 ;
  assign y3900 = ~n9737 ;
  assign y3901 = n9738 ;
  assign y3902 = ~n9742 ;
  assign y3903 = n9745 ;
  assign y3904 = ~n9747 ;
  assign y3905 = ~1'b0 ;
  assign y3906 = ~1'b0 ;
  assign y3907 = ~n9748 ;
  assign y3908 = ~n6373 ;
  assign y3909 = ~n9751 ;
  assign y3910 = ~n9752 ;
  assign y3911 = ~n9755 ;
  assign y3912 = ~n9761 ;
  assign y3913 = n9763 ;
  assign y3914 = n9765 ;
  assign y3915 = ~n9768 ;
  assign y3916 = ~n9772 ;
  assign y3917 = ~1'b0 ;
  assign y3918 = ~n9774 ;
  assign y3919 = n5099 ;
  assign y3920 = x98 ;
  assign y3921 = ~n9779 ;
  assign y3922 = 1'b0 ;
  assign y3923 = ~1'b0 ;
  assign y3924 = n9782 ;
  assign y3925 = ~1'b0 ;
  assign y3926 = n9783 ;
  assign y3927 = ~n9785 ;
  assign y3928 = n9788 ;
  assign y3929 = ~1'b0 ;
  assign y3930 = ~n9792 ;
  assign y3931 = n9793 ;
  assign y3932 = ~n9795 ;
  assign y3933 = ~n9797 ;
  assign y3934 = n9804 ;
  assign y3935 = n9807 ;
  assign y3936 = ~n9811 ;
  assign y3937 = ~1'b0 ;
  assign y3938 = ~1'b0 ;
  assign y3939 = n9817 ;
  assign y3940 = n9820 ;
  assign y3941 = ~n9831 ;
  assign y3942 = ~n9835 ;
  assign y3943 = ~n9836 ;
  assign y3944 = ~n9842 ;
  assign y3945 = n9843 ;
  assign y3946 = ~1'b0 ;
  assign y3947 = ~n9846 ;
  assign y3948 = ~n9847 ;
  assign y3949 = ~n9848 ;
  assign y3950 = ~n9849 ;
  assign y3951 = n9853 ;
  assign y3952 = ~n9863 ;
  assign y3953 = ~1'b0 ;
  assign y3954 = n9869 ;
  assign y3955 = n9871 ;
  assign y3956 = ~n9877 ;
  assign y3957 = ~n9879 ;
  assign y3958 = n9880 ;
  assign y3959 = n9881 ;
  assign y3960 = ~1'b0 ;
  assign y3961 = ~1'b0 ;
  assign y3962 = n9882 ;
  assign y3963 = ~n9884 ;
  assign y3964 = ~n3641 ;
  assign y3965 = n9894 ;
  assign y3966 = ~1'b0 ;
  assign y3967 = n9895 ;
  assign y3968 = ~n9900 ;
  assign y3969 = ~n9901 ;
  assign y3970 = ~n9903 ;
  assign y3971 = ~n9529 ;
  assign y3972 = ~n9904 ;
  assign y3973 = ~1'b0 ;
  assign y3974 = n9908 ;
  assign y3975 = n9909 ;
  assign y3976 = ~1'b0 ;
  assign y3977 = n5550 ;
  assign y3978 = ~n9917 ;
  assign y3979 = ~n9919 ;
  assign y3980 = ~n9920 ;
  assign y3981 = ~n9923 ;
  assign y3982 = ~n9932 ;
  assign y3983 = ~1'b0 ;
  assign y3984 = ~n9934 ;
  assign y3985 = ~n9937 ;
  assign y3986 = ~1'b0 ;
  assign y3987 = ~1'b0 ;
  assign y3988 = ~n9938 ;
  assign y3989 = ~n9939 ;
  assign y3990 = n9944 ;
  assign y3991 = ~n9946 ;
  assign y3992 = ~n9948 ;
  assign y3993 = ~1'b0 ;
  assign y3994 = n9949 ;
  assign y3995 = n9953 ;
  assign y3996 = ~n9956 ;
  assign y3997 = ~n9960 ;
  assign y3998 = n9966 ;
  assign y3999 = ~n9971 ;
  assign y4000 = ~n9981 ;
  assign y4001 = ~1'b0 ;
  assign y4002 = ~n9983 ;
  assign y4003 = ~n9985 ;
  assign y4004 = ~1'b0 ;
  assign y4005 = n9989 ;
  assign y4006 = n9991 ;
  assign y4007 = ~1'b0 ;
  assign y4008 = ~n9995 ;
  assign y4009 = ~1'b0 ;
  assign y4010 = ~n9999 ;
  assign y4011 = ~n10001 ;
  assign y4012 = ~n10002 ;
  assign y4013 = 1'b0 ;
  assign y4014 = ~n10006 ;
  assign y4015 = ~n10013 ;
  assign y4016 = n10016 ;
  assign y4017 = ~1'b0 ;
  assign y4018 = ~x138 ;
  assign y4019 = ~1'b0 ;
  assign y4020 = ~1'b0 ;
  assign y4021 = n10017 ;
  assign y4022 = ~1'b0 ;
  assign y4023 = ~n10023 ;
  assign y4024 = n10026 ;
  assign y4025 = ~n10027 ;
  assign y4026 = 1'b0 ;
  assign y4027 = n10028 ;
  assign y4028 = n10030 ;
  assign y4029 = ~1'b0 ;
  assign y4030 = n10033 ;
  assign y4031 = ~n10040 ;
  assign y4032 = n10043 ;
  assign y4033 = n10051 ;
  assign y4034 = n10057 ;
  assign y4035 = ~n8824 ;
  assign y4036 = ~n10059 ;
  assign y4037 = n10064 ;
  assign y4038 = ~1'b0 ;
  assign y4039 = ~n10066 ;
  assign y4040 = n10072 ;
  assign y4041 = n10078 ;
  assign y4042 = ~1'b0 ;
  assign y4043 = n10085 ;
  assign y4044 = ~n10088 ;
  assign y4045 = ~1'b0 ;
  assign y4046 = n10091 ;
  assign y4047 = ~n10094 ;
  assign y4048 = ~n8163 ;
  assign y4049 = ~1'b0 ;
  assign y4050 = ~n10095 ;
  assign y4051 = n10106 ;
  assign y4052 = ~n10108 ;
  assign y4053 = ~n10112 ;
  assign y4054 = n10123 ;
  assign y4055 = ~n10127 ;
  assign y4056 = ~1'b0 ;
  assign y4057 = ~1'b0 ;
  assign y4058 = n10132 ;
  assign y4059 = ~n10133 ;
  assign y4060 = ~1'b0 ;
  assign y4061 = n10135 ;
  assign y4062 = ~n10138 ;
  assign y4063 = 1'b0 ;
  assign y4064 = n10140 ;
  assign y4065 = n10142 ;
  assign y4066 = n10145 ;
  assign y4067 = ~1'b0 ;
  assign y4068 = ~1'b0 ;
  assign y4069 = n10148 ;
  assign y4070 = ~1'b0 ;
  assign y4071 = n10158 ;
  assign y4072 = ~n10167 ;
  assign y4073 = ~1'b0 ;
  assign y4074 = ~n10169 ;
  assign y4075 = n10170 ;
  assign y4076 = n10172 ;
  assign y4077 = n10174 ;
  assign y4078 = ~n10175 ;
  assign y4079 = n10178 ;
  assign y4080 = ~1'b0 ;
  assign y4081 = ~n10179 ;
  assign y4082 = n10185 ;
  assign y4083 = ~n10192 ;
  assign y4084 = ~n10193 ;
  assign y4085 = 1'b0 ;
  assign y4086 = ~1'b0 ;
  assign y4087 = ~1'b0 ;
  assign y4088 = n10196 ;
  assign y4089 = ~n10200 ;
  assign y4090 = ~n10207 ;
  assign y4091 = n8894 ;
  assign y4092 = ~n10209 ;
  assign y4093 = ~n10212 ;
  assign y4094 = n10213 ;
  assign y4095 = ~1'b0 ;
  assign y4096 = n10214 ;
  assign y4097 = ~n10215 ;
  assign y4098 = ~1'b0 ;
  assign y4099 = ~1'b0 ;
  assign y4100 = ~1'b0 ;
  assign y4101 = n10217 ;
  assign y4102 = ~n10228 ;
  assign y4103 = ~1'b0 ;
  assign y4104 = ~n10231 ;
  assign y4105 = n10232 ;
  assign y4106 = n10234 ;
  assign y4107 = n10239 ;
  assign y4108 = ~1'b0 ;
  assign y4109 = ~n6198 ;
  assign y4110 = 1'b0 ;
  assign y4111 = ~1'b0 ;
  assign y4112 = ~n10241 ;
  assign y4113 = ~n10243 ;
  assign y4114 = ~1'b0 ;
  assign y4115 = ~n10244 ;
  assign y4116 = n10245 ;
  assign y4117 = ~1'b0 ;
  assign y4118 = ~n10248 ;
  assign y4119 = ~1'b0 ;
  assign y4120 = ~n10252 ;
  assign y4121 = n10253 ;
  assign y4122 = n10255 ;
  assign y4123 = n10258 ;
  assign y4124 = ~1'b0 ;
  assign y4125 = ~n10261 ;
  assign y4126 = n10262 ;
  assign y4127 = ~1'b0 ;
  assign y4128 = ~n10270 ;
  assign y4129 = ~n10273 ;
  assign y4130 = ~n10277 ;
  assign y4131 = ~n10279 ;
  assign y4132 = n10282 ;
  assign y4133 = n10285 ;
  assign y4134 = ~n4953 ;
  assign y4135 = ~1'b0 ;
  assign y4136 = ~1'b0 ;
  assign y4137 = ~n10288 ;
  assign y4138 = ~n10291 ;
  assign y4139 = n10293 ;
  assign y4140 = n6312 ;
  assign y4141 = ~1'b0 ;
  assign y4142 = ~1'b0 ;
  assign y4143 = n10298 ;
  assign y4144 = ~n10303 ;
  assign y4145 = ~n10306 ;
  assign y4146 = n10315 ;
  assign y4147 = n10321 ;
  assign y4148 = n10322 ;
  assign y4149 = n10323 ;
  assign y4150 = n10327 ;
  assign y4151 = ~n10331 ;
  assign y4152 = ~1'b0 ;
  assign y4153 = ~1'b0 ;
  assign y4154 = n10333 ;
  assign y4155 = n10341 ;
  assign y4156 = n10343 ;
  assign y4157 = ~n7714 ;
  assign y4158 = n10344 ;
  assign y4159 = n10349 ;
  assign y4160 = ~n10354 ;
  assign y4161 = n10356 ;
  assign y4162 = ~n10359 ;
  assign y4163 = ~1'b0 ;
  assign y4164 = ~n10361 ;
  assign y4165 = n10365 ;
  assign y4166 = n10366 ;
  assign y4167 = ~n10374 ;
  assign y4168 = n10375 ;
  assign y4169 = ~1'b0 ;
  assign y4170 = ~1'b0 ;
  assign y4171 = n10379 ;
  assign y4172 = ~n10380 ;
  assign y4173 = ~n10383 ;
  assign y4174 = n10386 ;
  assign y4175 = n10387 ;
  assign y4176 = ~1'b0 ;
  assign y4177 = n10389 ;
  assign y4178 = ~n10391 ;
  assign y4179 = n10393 ;
  assign y4180 = n8790 ;
  assign y4181 = ~1'b0 ;
  assign y4182 = n10394 ;
  assign y4183 = n1826 ;
  assign y4184 = n10395 ;
  assign y4185 = n10396 ;
  assign y4186 = ~n10397 ;
  assign y4187 = ~n10398 ;
  assign y4188 = n10402 ;
  assign y4189 = ~n10404 ;
  assign y4190 = n10408 ;
  assign y4191 = n9531 ;
  assign y4192 = n10413 ;
  assign y4193 = ~n10414 ;
  assign y4194 = ~n10416 ;
  assign y4195 = ~n10417 ;
  assign y4196 = n10420 ;
  assign y4197 = 1'b0 ;
  assign y4198 = ~n10422 ;
  assign y4199 = n10425 ;
  assign y4200 = n10431 ;
  assign y4201 = ~n10436 ;
  assign y4202 = ~n10439 ;
  assign y4203 = 1'b0 ;
  assign y4204 = ~n10440 ;
  assign y4205 = ~1'b0 ;
  assign y4206 = ~1'b0 ;
  assign y4207 = ~1'b0 ;
  assign y4208 = n10453 ;
  assign y4209 = ~1'b0 ;
  assign y4210 = ~n10457 ;
  assign y4211 = ~n10462 ;
  assign y4212 = ~n10466 ;
  assign y4213 = n10468 ;
  assign y4214 = ~n10473 ;
  assign y4215 = n10474 ;
  assign y4216 = ~n10479 ;
  assign y4217 = ~n10483 ;
  assign y4218 = ~n10486 ;
  assign y4219 = ~n10488 ;
  assign y4220 = n10491 ;
  assign y4221 = ~1'b0 ;
  assign y4222 = n10492 ;
  assign y4223 = n10494 ;
  assign y4224 = ~1'b0 ;
  assign y4225 = ~n10497 ;
  assign y4226 = n10499 ;
  assign y4227 = n10502 ;
  assign y4228 = n10508 ;
  assign y4229 = ~n10514 ;
  assign y4230 = n10515 ;
  assign y4231 = ~n10516 ;
  assign y4232 = n10518 ;
  assign y4233 = n10521 ;
  assign y4234 = ~n10529 ;
  assign y4235 = ~n10545 ;
  assign y4236 = ~n10547 ;
  assign y4237 = ~n10548 ;
  assign y4238 = ~n10550 ;
  assign y4239 = ~n10552 ;
  assign y4240 = ~n10553 ;
  assign y4241 = n10555 ;
  assign y4242 = ~n10558 ;
  assign y4243 = ~1'b0 ;
  assign y4244 = n10560 ;
  assign y4245 = ~n10562 ;
  assign y4246 = n10568 ;
  assign y4247 = ~1'b0 ;
  assign y4248 = ~1'b0 ;
  assign y4249 = n10573 ;
  assign y4250 = n10575 ;
  assign y4251 = n10578 ;
  assign y4252 = n10580 ;
  assign y4253 = ~1'b0 ;
  assign y4254 = ~n10582 ;
  assign y4255 = ~n10584 ;
  assign y4256 = ~n6313 ;
  assign y4257 = n10589 ;
  assign y4258 = ~1'b0 ;
  assign y4259 = n10592 ;
  assign y4260 = n10593 ;
  assign y4261 = n10595 ;
  assign y4262 = n10603 ;
  assign y4263 = ~1'b0 ;
  assign y4264 = ~n10606 ;
  assign y4265 = n10607 ;
  assign y4266 = ~n10609 ;
  assign y4267 = n10611 ;
  assign y4268 = ~1'b0 ;
  assign y4269 = n10617 ;
  assign y4270 = ~x131 ;
  assign y4271 = ~n10620 ;
  assign y4272 = n10621 ;
  assign y4273 = n10623 ;
  assign y4274 = n10627 ;
  assign y4275 = 1'b0 ;
  assign y4276 = n10632 ;
  assign y4277 = ~n10634 ;
  assign y4278 = n10637 ;
  assign y4279 = ~n10644 ;
  assign y4280 = n10646 ;
  assign y4281 = ~n10647 ;
  assign y4282 = n10649 ;
  assign y4283 = ~1'b0 ;
  assign y4284 = ~n9403 ;
  assign y4285 = n10651 ;
  assign y4286 = ~n10660 ;
  assign y4287 = ~1'b0 ;
  assign y4288 = ~n10664 ;
  assign y4289 = n9112 ;
  assign y4290 = n10667 ;
  assign y4291 = ~1'b0 ;
  assign y4292 = n10669 ;
  assign y4293 = ~1'b0 ;
  assign y4294 = ~n10677 ;
  assign y4295 = ~1'b0 ;
  assign y4296 = ~n10679 ;
  assign y4297 = ~1'b0 ;
  assign y4298 = ~n10680 ;
  assign y4299 = n10683 ;
  assign y4300 = n2930 ;
  assign y4301 = ~1'b0 ;
  assign y4302 = ~n10684 ;
  assign y4303 = n10685 ;
  assign y4304 = ~n10686 ;
  assign y4305 = ~1'b0 ;
  assign y4306 = ~n10692 ;
  assign y4307 = n10696 ;
  assign y4308 = n10697 ;
  assign y4309 = n10702 ;
  assign y4310 = ~n10706 ;
  assign y4311 = ~1'b0 ;
  assign y4312 = ~n10711 ;
  assign y4313 = ~n7928 ;
  assign y4314 = ~1'b0 ;
  assign y4315 = ~n5720 ;
  assign y4316 = ~1'b0 ;
  assign y4317 = ~1'b0 ;
  assign y4318 = ~n10715 ;
  assign y4319 = ~n10718 ;
  assign y4320 = ~1'b0 ;
  assign y4321 = ~n10721 ;
  assign y4322 = ~1'b0 ;
  assign y4323 = ~n10732 ;
  assign y4324 = ~n10733 ;
  assign y4325 = n10737 ;
  assign y4326 = n10743 ;
  assign y4327 = n10744 ;
  assign y4328 = ~n10745 ;
  assign y4329 = ~1'b0 ;
  assign y4330 = n10746 ;
  assign y4331 = 1'b0 ;
  assign y4332 = ~n10747 ;
  assign y4333 = n10750 ;
  assign y4334 = ~n10753 ;
  assign y4335 = n10755 ;
  assign y4336 = ~n10759 ;
  assign y4337 = n10761 ;
  assign y4338 = ~n10763 ;
  assign y4339 = ~n10774 ;
  assign y4340 = ~1'b0 ;
  assign y4341 = ~n10776 ;
  assign y4342 = ~1'b0 ;
  assign y4343 = n10778 ;
  assign y4344 = n10783 ;
  assign y4345 = ~n1285 ;
  assign y4346 = ~1'b0 ;
  assign y4347 = n10786 ;
  assign y4348 = n10787 ;
  assign y4349 = n10793 ;
  assign y4350 = ~1'b0 ;
  assign y4351 = ~n10806 ;
  assign y4352 = n10808 ;
  assign y4353 = n10812 ;
  assign y4354 = n10815 ;
  assign y4355 = ~1'b0 ;
  assign y4356 = n10820 ;
  assign y4357 = ~n10827 ;
  assign y4358 = ~1'b0 ;
  assign y4359 = ~1'b0 ;
  assign y4360 = ~1'b0 ;
  assign y4361 = ~1'b0 ;
  assign y4362 = n10828 ;
  assign y4363 = ~n10833 ;
  assign y4364 = n10839 ;
  assign y4365 = ~1'b0 ;
  assign y4366 = ~n10842 ;
  assign y4367 = ~n10844 ;
  assign y4368 = ~1'b0 ;
  assign y4369 = n10845 ;
  assign y4370 = n10846 ;
  assign y4371 = ~n1187 ;
  assign y4372 = n10848 ;
  assign y4373 = ~n10850 ;
  assign y4374 = ~n10853 ;
  assign y4375 = n8648 ;
  assign y4376 = n10855 ;
  assign y4377 = ~1'b0 ;
  assign y4378 = ~1'b0 ;
  assign y4379 = ~n10856 ;
  assign y4380 = ~n10864 ;
  assign y4381 = ~1'b0 ;
  assign y4382 = n10865 ;
  assign y4383 = ~n10870 ;
  assign y4384 = ~n10873 ;
  assign y4385 = ~1'b0 ;
  assign y4386 = n10874 ;
  assign y4387 = n10891 ;
  assign y4388 = n10895 ;
  assign y4389 = ~n10896 ;
  assign y4390 = ~1'b0 ;
  assign y4391 = n10898 ;
  assign y4392 = n10900 ;
  assign y4393 = ~x17 ;
  assign y4394 = ~n10901 ;
  assign y4395 = n10908 ;
  assign y4396 = ~n10909 ;
  assign y4397 = ~n10917 ;
  assign y4398 = ~n10920 ;
  assign y4399 = n10921 ;
  assign y4400 = n10930 ;
  assign y4401 = n10934 ;
  assign y4402 = ~n10939 ;
  assign y4403 = ~n10943 ;
  assign y4404 = ~1'b0 ;
  assign y4405 = n10944 ;
  assign y4406 = n10946 ;
  assign y4407 = n9544 ;
  assign y4408 = ~n10949 ;
  assign y4409 = ~1'b0 ;
  assign y4410 = n10787 ;
  assign y4411 = n10951 ;
  assign y4412 = ~n10958 ;
  assign y4413 = ~1'b0 ;
  assign y4414 = ~n10960 ;
  assign y4415 = ~1'b0 ;
  assign y4416 = ~1'b0 ;
  assign y4417 = ~n10962 ;
  assign y4418 = ~1'b0 ;
  assign y4419 = ~n10968 ;
  assign y4420 = ~n10970 ;
  assign y4421 = ~n10971 ;
  assign y4422 = ~n10975 ;
  assign y4423 = n10976 ;
  assign y4424 = ~n10978 ;
  assign y4425 = ~1'b0 ;
  assign y4426 = ~1'b0 ;
  assign y4427 = ~1'b0 ;
  assign y4428 = ~n10979 ;
  assign y4429 = ~n10984 ;
  assign y4430 = n10985 ;
  assign y4431 = 1'b0 ;
  assign y4432 = ~1'b0 ;
  assign y4433 = ~n10991 ;
  assign y4434 = n10995 ;
  assign y4435 = ~1'b0 ;
  assign y4436 = ~n10999 ;
  assign y4437 = n10973 ;
  assign y4438 = ~n4931 ;
  assign y4439 = ~n11006 ;
  assign y4440 = ~n11008 ;
  assign y4441 = ~n11010 ;
  assign y4442 = 1'b0 ;
  assign y4443 = n11011 ;
  assign y4444 = ~n11012 ;
  assign y4445 = n11013 ;
  assign y4446 = ~1'b0 ;
  assign y4447 = n11015 ;
  assign y4448 = n11017 ;
  assign y4449 = ~n11022 ;
  assign y4450 = n11026 ;
  assign y4451 = ~1'b0 ;
  assign y4452 = ~1'b0 ;
  assign y4453 = ~n11028 ;
  assign y4454 = n2026 ;
  assign y4455 = ~1'b0 ;
  assign y4456 = ~n11032 ;
  assign y4457 = ~1'b0 ;
  assign y4458 = ~n11037 ;
  assign y4459 = n11042 ;
  assign y4460 = ~n11045 ;
  assign y4461 = ~1'b0 ;
  assign y4462 = ~n11047 ;
  assign y4463 = n11053 ;
  assign y4464 = ~1'b0 ;
  assign y4465 = n11058 ;
  assign y4466 = ~1'b0 ;
  assign y4467 = ~n11061 ;
  assign y4468 = ~n11063 ;
  assign y4469 = n11065 ;
  assign y4470 = 1'b0 ;
  assign y4471 = n11066 ;
  assign y4472 = ~n11069 ;
  assign y4473 = ~1'b0 ;
  assign y4474 = 1'b0 ;
  assign y4475 = ~n11070 ;
  assign y4476 = ~1'b0 ;
  assign y4477 = n11074 ;
  assign y4478 = ~n11076 ;
  assign y4479 = n11077 ;
  assign y4480 = n11082 ;
  assign y4481 = ~n11083 ;
  assign y4482 = ~n11085 ;
  assign y4483 = ~n11086 ;
  assign y4484 = ~n11087 ;
  assign y4485 = n8632 ;
  assign y4486 = ~1'b0 ;
  assign y4487 = n11088 ;
  assign y4488 = ~n11090 ;
  assign y4489 = ~1'b0 ;
  assign y4490 = n11091 ;
  assign y4491 = ~n11097 ;
  assign y4492 = ~n11098 ;
  assign y4493 = ~n11101 ;
  assign y4494 = n11108 ;
  assign y4495 = ~1'b0 ;
  assign y4496 = ~n11113 ;
  assign y4497 = n1350 ;
  assign y4498 = n11115 ;
  assign y4499 = ~1'b0 ;
  assign y4500 = ~1'b0 ;
  assign y4501 = n11121 ;
  assign y4502 = n11122 ;
  assign y4503 = n11123 ;
  assign y4504 = ~n11127 ;
  assign y4505 = ~n11129 ;
  assign y4506 = ~1'b0 ;
  assign y4507 = n11133 ;
  assign y4508 = n11135 ;
  assign y4509 = ~1'b0 ;
  assign y4510 = n11136 ;
  assign y4511 = ~1'b0 ;
  assign y4512 = ~n11141 ;
  assign y4513 = n11147 ;
  assign y4514 = ~n11151 ;
  assign y4515 = ~1'b0 ;
  assign y4516 = ~n11152 ;
  assign y4517 = ~n11153 ;
  assign y4518 = ~n11161 ;
  assign y4519 = n11163 ;
  assign y4520 = ~1'b0 ;
  assign y4521 = ~1'b0 ;
  assign y4522 = ~1'b0 ;
  assign y4523 = n271 ;
  assign y4524 = ~n11164 ;
  assign y4525 = ~1'b0 ;
  assign y4526 = ~n11165 ;
  assign y4527 = ~n11168 ;
  assign y4528 = ~n11169 ;
  assign y4529 = ~1'b0 ;
  assign y4530 = n11171 ;
  assign y4531 = n11174 ;
  assign y4532 = ~n11175 ;
  assign y4533 = ~n11187 ;
  assign y4534 = n11190 ;
  assign y4535 = n11194 ;
  assign y4536 = ~1'b0 ;
  assign y4537 = ~n11196 ;
  assign y4538 = ~n11198 ;
  assign y4539 = n11200 ;
  assign y4540 = n11202 ;
  assign y4541 = n11204 ;
  assign y4542 = ~n11208 ;
  assign y4543 = ~1'b0 ;
  assign y4544 = ~1'b0 ;
  assign y4545 = ~n11213 ;
  assign y4546 = ~n11215 ;
  assign y4547 = n11221 ;
  assign y4548 = n11231 ;
  assign y4549 = ~n706 ;
  assign y4550 = ~n11235 ;
  assign y4551 = n11236 ;
  assign y4552 = ~n11246 ;
  assign y4553 = ~n11249 ;
  assign y4554 = n11252 ;
  assign y4555 = ~1'b0 ;
  assign y4556 = ~1'b0 ;
  assign y4557 = ~1'b0 ;
  assign y4558 = n11256 ;
  assign y4559 = n6683 ;
  assign y4560 = n11266 ;
  assign y4561 = ~n11267 ;
  assign y4562 = ~1'b0 ;
  assign y4563 = ~1'b0 ;
  assign y4564 = n11268 ;
  assign y4565 = n11269 ;
  assign y4566 = ~n11271 ;
  assign y4567 = ~n11272 ;
  assign y4568 = ~n11275 ;
  assign y4569 = n11276 ;
  assign y4570 = ~n11280 ;
  assign y4571 = ~1'b0 ;
  assign y4572 = ~1'b0 ;
  assign y4573 = n11284 ;
  assign y4574 = 1'b0 ;
  assign y4575 = n11286 ;
  assign y4576 = ~n11289 ;
  assign y4577 = ~n279 ;
  assign y4578 = ~n11290 ;
  assign y4579 = ~1'b0 ;
  assign y4580 = n11292 ;
  assign y4581 = n11295 ;
  assign y4582 = n11300 ;
  assign y4583 = ~1'b0 ;
  assign y4584 = ~n11302 ;
  assign y4585 = ~1'b0 ;
  assign y4586 = ~n11303 ;
  assign y4587 = ~n11304 ;
  assign y4588 = ~1'b0 ;
  assign y4589 = ~1'b0 ;
  assign y4590 = ~n11306 ;
  assign y4591 = ~n7490 ;
  assign y4592 = ~n11308 ;
  assign y4593 = ~1'b0 ;
  assign y4594 = n11313 ;
  assign y4595 = ~n11324 ;
  assign y4596 = ~1'b0 ;
  assign y4597 = ~1'b0 ;
  assign y4598 = ~1'b0 ;
  assign y4599 = ~n11330 ;
  assign y4600 = n11332 ;
  assign y4601 = ~1'b0 ;
  assign y4602 = n11335 ;
  assign y4603 = ~n11336 ;
  assign y4604 = n11338 ;
  assign y4605 = n11339 ;
  assign y4606 = ~n11341 ;
  assign y4607 = n11346 ;
  assign y4608 = ~1'b0 ;
  assign y4609 = n10803 ;
  assign y4610 = ~n11348 ;
  assign y4611 = ~1'b0 ;
  assign y4612 = ~n11350 ;
  assign y4613 = n11351 ;
  assign y4614 = n11355 ;
  assign y4615 = ~1'b0 ;
  assign y4616 = ~n11359 ;
  assign y4617 = ~1'b0 ;
  assign y4618 = n11360 ;
  assign y4619 = ~n1801 ;
  assign y4620 = n11365 ;
  assign y4621 = ~n11367 ;
  assign y4622 = n11368 ;
  assign y4623 = ~n11370 ;
  assign y4624 = n11372 ;
  assign y4625 = ~n11380 ;
  assign y4626 = ~n11385 ;
  assign y4627 = ~n11394 ;
  assign y4628 = ~n11402 ;
  assign y4629 = ~n11404 ;
  assign y4630 = ~n11405 ;
  assign y4631 = n11406 ;
  assign y4632 = n11410 ;
  assign y4633 = ~n11413 ;
  assign y4634 = ~1'b0 ;
  assign y4635 = n11415 ;
  assign y4636 = ~n11419 ;
  assign y4637 = n11422 ;
  assign y4638 = n11428 ;
  assign y4639 = ~n11429 ;
  assign y4640 = ~n11438 ;
  assign y4641 = ~1'b0 ;
  assign y4642 = ~1'b0 ;
  assign y4643 = ~1'b0 ;
  assign y4644 = n11440 ;
  assign y4645 = ~1'b0 ;
  assign y4646 = ~1'b0 ;
  assign y4647 = ~1'b0 ;
  assign y4648 = ~n11444 ;
  assign y4649 = n11446 ;
  assign y4650 = ~n11448 ;
  assign y4651 = n11454 ;
  assign y4652 = ~1'b0 ;
  assign y4653 = n11455 ;
  assign y4654 = n11459 ;
  assign y4655 = n2725 ;
  assign y4656 = ~1'b0 ;
  assign y4657 = n11464 ;
  assign y4658 = ~1'b0 ;
  assign y4659 = n11465 ;
  assign y4660 = ~1'b0 ;
  assign y4661 = ~n7915 ;
  assign y4662 = ~1'b0 ;
  assign y4663 = n11467 ;
  assign y4664 = ~n11468 ;
  assign y4665 = ~n11471 ;
  assign y4666 = n11477 ;
  assign y4667 = n11478 ;
  assign y4668 = ~1'b0 ;
  assign y4669 = n11482 ;
  assign y4670 = ~1'b0 ;
  assign y4671 = n11483 ;
  assign y4672 = n11484 ;
  assign y4673 = ~n11488 ;
  assign y4674 = n11490 ;
  assign y4675 = n11496 ;
  assign y4676 = n11499 ;
  assign y4677 = ~n11501 ;
  assign y4678 = ~n11503 ;
  assign y4679 = ~n11505 ;
  assign y4680 = ~n11508 ;
  assign y4681 = ~1'b0 ;
  assign y4682 = ~n11515 ;
  assign y4683 = ~1'b0 ;
  assign y4684 = n11518 ;
  assign y4685 = n11519 ;
  assign y4686 = ~n11522 ;
  assign y4687 = n11528 ;
  assign y4688 = n11530 ;
  assign y4689 = ~n11534 ;
  assign y4690 = ~1'b0 ;
  assign y4691 = 1'b0 ;
  assign y4692 = n11541 ;
  assign y4693 = ~1'b0 ;
  assign y4694 = ~n7399 ;
  assign y4695 = ~n11545 ;
  assign y4696 = n11552 ;
  assign y4697 = n11553 ;
  assign y4698 = ~n11554 ;
  assign y4699 = ~n11558 ;
  assign y4700 = ~1'b0 ;
  assign y4701 = n11560 ;
  assign y4702 = ~n11561 ;
  assign y4703 = ~n11564 ;
  assign y4704 = n11565 ;
  assign y4705 = ~1'b0 ;
  assign y4706 = n11566 ;
  assign y4707 = ~n11567 ;
  assign y4708 = ~1'b0 ;
  assign y4709 = n11569 ;
  assign y4710 = ~1'b0 ;
  assign y4711 = ~1'b0 ;
  assign y4712 = ~n11570 ;
  assign y4713 = n11571 ;
  assign y4714 = ~1'b0 ;
  assign y4715 = ~n11574 ;
  assign y4716 = ~n11579 ;
  assign y4717 = ~n11583 ;
  assign y4718 = ~n11585 ;
  assign y4719 = n11588 ;
  assign y4720 = n11591 ;
  assign y4721 = ~1'b0 ;
  assign y4722 = ~n11594 ;
  assign y4723 = n2226 ;
  assign y4724 = 1'b0 ;
  assign y4725 = ~n11597 ;
  assign y4726 = ~1'b0 ;
  assign y4727 = ~1'b0 ;
  assign y4728 = ~n11604 ;
  assign y4729 = ~n11607 ;
  assign y4730 = n11616 ;
  assign y4731 = n11618 ;
  assign y4732 = n11624 ;
  assign y4733 = ~n11626 ;
  assign y4734 = n11628 ;
  assign y4735 = ~1'b0 ;
  assign y4736 = ~1'b0 ;
  assign y4737 = ~1'b0 ;
  assign y4738 = ~n3053 ;
  assign y4739 = ~n11633 ;
  assign y4740 = ~n11635 ;
  assign y4741 = n11636 ;
  assign y4742 = ~1'b0 ;
  assign y4743 = ~n11645 ;
  assign y4744 = ~1'b0 ;
  assign y4745 = ~n11647 ;
  assign y4746 = n11655 ;
  assign y4747 = ~n11657 ;
  assign y4748 = ~n11660 ;
  assign y4749 = ~n11665 ;
  assign y4750 = ~n11668 ;
  assign y4751 = ~n11674 ;
  assign y4752 = ~n11678 ;
  assign y4753 = n11679 ;
  assign y4754 = n11683 ;
  assign y4755 = ~n11690 ;
  assign y4756 = ~1'b0 ;
  assign y4757 = n11698 ;
  assign y4758 = n11699 ;
  assign y4759 = ~1'b0 ;
  assign y4760 = ~1'b0 ;
  assign y4761 = n11713 ;
  assign y4762 = n11716 ;
  assign y4763 = ~1'b0 ;
  assign y4764 = ~n11717 ;
  assign y4765 = n11721 ;
  assign y4766 = 1'b0 ;
  assign y4767 = ~n11724 ;
  assign y4768 = ~1'b0 ;
  assign y4769 = n11725 ;
  assign y4770 = ~1'b0 ;
  assign y4771 = ~n11730 ;
  assign y4772 = ~n11737 ;
  assign y4773 = ~1'b0 ;
  assign y4774 = n11741 ;
  assign y4775 = ~n11746 ;
  assign y4776 = 1'b0 ;
  assign y4777 = ~n11747 ;
  assign y4778 = ~n11750 ;
  assign y4779 = ~n11751 ;
  assign y4780 = ~1'b0 ;
  assign y4781 = ~n11752 ;
  assign y4782 = n7603 ;
  assign y4783 = n11753 ;
  assign y4784 = ~1'b0 ;
  assign y4785 = ~n11754 ;
  assign y4786 = n11764 ;
  assign y4787 = n11770 ;
  assign y4788 = ~n11771 ;
  assign y4789 = ~n11776 ;
  assign y4790 = n11777 ;
  assign y4791 = n11778 ;
  assign y4792 = n11780 ;
  assign y4793 = n11781 ;
  assign y4794 = n11796 ;
  assign y4795 = ~n11799 ;
  assign y4796 = ~n11804 ;
  assign y4797 = ~n11809 ;
  assign y4798 = ~n11812 ;
  assign y4799 = ~n11813 ;
  assign y4800 = ~1'b0 ;
  assign y4801 = n11815 ;
  assign y4802 = n11817 ;
  assign y4803 = n11819 ;
  assign y4804 = ~1'b0 ;
  assign y4805 = ~n11821 ;
  assign y4806 = ~1'b0 ;
  assign y4807 = ~n11823 ;
  assign y4808 = ~n11827 ;
  assign y4809 = ~1'b0 ;
  assign y4810 = ~n11829 ;
  assign y4811 = ~n11830 ;
  assign y4812 = ~n11834 ;
  assign y4813 = ~n11841 ;
  assign y4814 = n11844 ;
  assign y4815 = n11845 ;
  assign y4816 = n11846 ;
  assign y4817 = n11848 ;
  assign y4818 = ~n11853 ;
  assign y4819 = n11854 ;
  assign y4820 = ~n11855 ;
  assign y4821 = ~n11858 ;
  assign y4822 = ~1'b0 ;
  assign y4823 = n11863 ;
  assign y4824 = ~n11870 ;
  assign y4825 = ~n11876 ;
  assign y4826 = ~1'b0 ;
  assign y4827 = ~n11879 ;
  assign y4828 = n11888 ;
  assign y4829 = ~n11889 ;
  assign y4830 = ~n11893 ;
  assign y4831 = n11898 ;
  assign y4832 = ~1'b0 ;
  assign y4833 = n11900 ;
  assign y4834 = ~1'b0 ;
  assign y4835 = n11901 ;
  assign y4836 = ~n11902 ;
  assign y4837 = ~n11905 ;
  assign y4838 = ~n11908 ;
  assign y4839 = n11917 ;
  assign y4840 = ~1'b0 ;
  assign y4841 = ~n11918 ;
  assign y4842 = ~n11921 ;
  assign y4843 = n11924 ;
  assign y4844 = ~n11928 ;
  assign y4845 = n11929 ;
  assign y4846 = ~n11933 ;
  assign y4847 = n11934 ;
  assign y4848 = n11937 ;
  assign y4849 = ~1'b0 ;
  assign y4850 = ~1'b0 ;
  assign y4851 = n11939 ;
  assign y4852 = ~n11942 ;
  assign y4853 = ~n11948 ;
  assign y4854 = n11949 ;
  assign y4855 = n11953 ;
  assign y4856 = n11955 ;
  assign y4857 = ~n11956 ;
  assign y4858 = ~n4148 ;
  assign y4859 = ~n11959 ;
  assign y4860 = n11960 ;
  assign y4861 = ~n11963 ;
  assign y4862 = ~1'b0 ;
  assign y4863 = ~n4953 ;
  assign y4864 = ~1'b0 ;
  assign y4865 = ~n11968 ;
  assign y4866 = ~n11972 ;
  assign y4867 = ~1'b0 ;
  assign y4868 = ~1'b0 ;
  assign y4869 = n11973 ;
  assign y4870 = ~n11974 ;
  assign y4871 = ~n11977 ;
  assign y4872 = ~n11981 ;
  assign y4873 = ~1'b0 ;
  assign y4874 = ~n11983 ;
  assign y4875 = n11988 ;
  assign y4876 = ~n11989 ;
  assign y4877 = ~1'b0 ;
  assign y4878 = ~n11990 ;
  assign y4879 = n11991 ;
  assign y4880 = n11997 ;
  assign y4881 = n11998 ;
  assign y4882 = n11999 ;
  assign y4883 = ~n12007 ;
  assign y4884 = n12008 ;
  assign y4885 = ~n12013 ;
  assign y4886 = ~n12018 ;
  assign y4887 = ~1'b0 ;
  assign y4888 = ~n12019 ;
  assign y4889 = ~n12025 ;
  assign y4890 = ~n12027 ;
  assign y4891 = ~1'b0 ;
  assign y4892 = ~1'b0 ;
  assign y4893 = n12029 ;
  assign y4894 = ~n12033 ;
  assign y4895 = ~n12035 ;
  assign y4896 = n12037 ;
  assign y4897 = ~n12039 ;
  assign y4898 = ~n12044 ;
  assign y4899 = ~n4016 ;
  assign y4900 = ~n12045 ;
  assign y4901 = ~1'b0 ;
  assign y4902 = ~n12048 ;
  assign y4903 = ~n12051 ;
  assign y4904 = ~n12053 ;
  assign y4905 = n5740 ;
  assign y4906 = ~n5788 ;
  assign y4907 = ~1'b0 ;
  assign y4908 = ~n12058 ;
  assign y4909 = n12060 ;
  assign y4910 = ~1'b0 ;
  assign y4911 = ~n12061 ;
  assign y4912 = ~n12065 ;
  assign y4913 = ~1'b0 ;
  assign y4914 = n12070 ;
  assign y4915 = ~1'b0 ;
  assign y4916 = ~n12071 ;
  assign y4917 = ~1'b0 ;
  assign y4918 = n12072 ;
  assign y4919 = ~1'b0 ;
  assign y4920 = ~n12075 ;
  assign y4921 = ~n12078 ;
  assign y4922 = n12083 ;
  assign y4923 = ~n12085 ;
  assign y4924 = ~n12090 ;
  assign y4925 = ~n12097 ;
  assign y4926 = n12099 ;
  assign y4927 = n12103 ;
  assign y4928 = n12106 ;
  assign y4929 = n12112 ;
  assign y4930 = ~1'b0 ;
  assign y4931 = n12114 ;
  assign y4932 = ~n6844 ;
  assign y4933 = ~1'b0 ;
  assign y4934 = n12115 ;
  assign y4935 = n12117 ;
  assign y4936 = ~n6683 ;
  assign y4937 = ~1'b0 ;
  assign y4938 = ~1'b0 ;
  assign y4939 = ~1'b0 ;
  assign y4940 = n12124 ;
  assign y4941 = ~n12125 ;
  assign y4942 = n12131 ;
  assign y4943 = ~n12132 ;
  assign y4944 = ~n12136 ;
  assign y4945 = n12140 ;
  assign y4946 = ~n12150 ;
  assign y4947 = ~1'b0 ;
  assign y4948 = ~1'b0 ;
  assign y4949 = ~1'b0 ;
  assign y4950 = ~n12151 ;
  assign y4951 = ~n12155 ;
  assign y4952 = ~n12157 ;
  assign y4953 = ~n12158 ;
  assign y4954 = ~1'b0 ;
  assign y4955 = ~n12160 ;
  assign y4956 = ~1'b0 ;
  assign y4957 = n12165 ;
  assign y4958 = n12168 ;
  assign y4959 = ~n12172 ;
  assign y4960 = ~1'b0 ;
  assign y4961 = ~n12176 ;
  assign y4962 = ~n12178 ;
  assign y4963 = ~1'b0 ;
  assign y4964 = ~n12180 ;
  assign y4965 = ~n12186 ;
  assign y4966 = n12187 ;
  assign y4967 = ~1'b0 ;
  assign y4968 = ~n12190 ;
  assign y4969 = ~n9002 ;
  assign y4970 = n12195 ;
  assign y4971 = n12197 ;
  assign y4972 = n12198 ;
  assign y4973 = n12202 ;
  assign y4974 = ~1'b0 ;
  assign y4975 = n12204 ;
  assign y4976 = ~n12205 ;
  assign y4977 = n12208 ;
  assign y4978 = n12213 ;
  assign y4979 = n10455 ;
  assign y4980 = n12219 ;
  assign y4981 = n12223 ;
  assign y4982 = ~n12231 ;
  assign y4983 = ~n12233 ;
  assign y4984 = ~1'b0 ;
  assign y4985 = ~n12235 ;
  assign y4986 = ~n12236 ;
  assign y4987 = n12237 ;
  assign y4988 = ~n12242 ;
  assign y4989 = n12243 ;
  assign y4990 = ~1'b0 ;
  assign y4991 = n12245 ;
  assign y4992 = ~n9539 ;
  assign y4993 = ~n12247 ;
  assign y4994 = ~1'b0 ;
  assign y4995 = ~1'b0 ;
  assign y4996 = ~n12248 ;
  assign y4997 = ~1'b0 ;
  assign y4998 = n12258 ;
  assign y4999 = n12265 ;
  assign y5000 = ~n12273 ;
  assign y5001 = ~n12275 ;
  assign y5002 = ~n12278 ;
  assign y5003 = ~n12279 ;
  assign y5004 = n5695 ;
  assign y5005 = ~n7349 ;
  assign y5006 = ~1'b0 ;
  assign y5007 = n12281 ;
  assign y5008 = n12286 ;
  assign y5009 = ~1'b0 ;
  assign y5010 = ~1'b0 ;
  assign y5011 = ~n12297 ;
  assign y5012 = ~n12300 ;
  assign y5013 = ~n12302 ;
  assign y5014 = 1'b0 ;
  assign y5015 = ~1'b0 ;
  assign y5016 = n12304 ;
  assign y5017 = n12305 ;
  assign y5018 = ~1'b0 ;
  assign y5019 = n12322 ;
  assign y5020 = ~n12324 ;
  assign y5021 = ~n12329 ;
  assign y5022 = n12334 ;
  assign y5023 = ~n12337 ;
  assign y5024 = ~1'b0 ;
  assign y5025 = n12339 ;
  assign y5026 = ~n12341 ;
  assign y5027 = n12342 ;
  assign y5028 = ~1'b0 ;
  assign y5029 = ~n12343 ;
  assign y5030 = ~1'b0 ;
  assign y5031 = ~n12344 ;
  assign y5032 = n12346 ;
  assign y5033 = n12356 ;
  assign y5034 = ~n12360 ;
  assign y5035 = n12362 ;
  assign y5036 = n12368 ;
  assign y5037 = ~n12370 ;
  assign y5038 = n12375 ;
  assign y5039 = n12376 ;
  assign y5040 = ~1'b0 ;
  assign y5041 = n12385 ;
  assign y5042 = ~n12394 ;
  assign y5043 = n12396 ;
  assign y5044 = ~n12399 ;
  assign y5045 = n12402 ;
  assign y5046 = n12403 ;
  assign y5047 = n12405 ;
  assign y5048 = n12408 ;
  assign y5049 = ~1'b0 ;
  assign y5050 = n12417 ;
  assign y5051 = n12420 ;
  assign y5052 = ~1'b0 ;
  assign y5053 = ~n12421 ;
  assign y5054 = ~1'b0 ;
  assign y5055 = ~1'b0 ;
  assign y5056 = ~n12426 ;
  assign y5057 = n12432 ;
  assign y5058 = n6569 ;
  assign y5059 = ~n12436 ;
  assign y5060 = ~n12437 ;
  assign y5061 = ~n9733 ;
  assign y5062 = 1'b0 ;
  assign y5063 = ~n12445 ;
  assign y5064 = n12448 ;
  assign y5065 = n12449 ;
  assign y5066 = n12453 ;
  assign y5067 = ~1'b0 ;
  assign y5068 = ~n12454 ;
  assign y5069 = 1'b0 ;
  assign y5070 = ~n12456 ;
  assign y5071 = n12466 ;
  assign y5072 = ~n12469 ;
  assign y5073 = n12470 ;
  assign y5074 = n12471 ;
  assign y5075 = ~n12474 ;
  assign y5076 = ~1'b0 ;
  assign y5077 = ~n12481 ;
  assign y5078 = ~1'b0 ;
  assign y5079 = ~n12484 ;
  assign y5080 = ~1'b0 ;
  assign y5081 = n12488 ;
  assign y5082 = ~n12490 ;
  assign y5083 = ~n12493 ;
  assign y5084 = n12497 ;
  assign y5085 = n12502 ;
  assign y5086 = n12503 ;
  assign y5087 = ~n12512 ;
  assign y5088 = ~n12518 ;
  assign y5089 = n12522 ;
  assign y5090 = n12523 ;
  assign y5091 = ~1'b0 ;
  assign y5092 = ~1'b0 ;
  assign y5093 = ~1'b0 ;
  assign y5094 = n3365 ;
  assign y5095 = ~n12527 ;
  assign y5096 = ~n8340 ;
  assign y5097 = n12529 ;
  assign y5098 = ~n12533 ;
  assign y5099 = ~n12534 ;
  assign y5100 = ~n12538 ;
  assign y5101 = n12540 ;
  assign y5102 = n12547 ;
  assign y5103 = ~1'b0 ;
  assign y5104 = n12548 ;
  assign y5105 = n12552 ;
  assign y5106 = n12555 ;
  assign y5107 = ~1'b0 ;
  assign y5108 = ~1'b0 ;
  assign y5109 = n12563 ;
  assign y5110 = n12567 ;
  assign y5111 = ~n12568 ;
  assign y5112 = ~1'b0 ;
  assign y5113 = n12575 ;
  assign y5114 = ~n12579 ;
  assign y5115 = ~n12580 ;
  assign y5116 = n12582 ;
  assign y5117 = ~1'b0 ;
  assign y5118 = n12588 ;
  assign y5119 = ~1'b0 ;
  assign y5120 = ~1'b0 ;
  assign y5121 = n12594 ;
  assign y5122 = ~1'b0 ;
  assign y5123 = n12598 ;
  assign y5124 = n12604 ;
  assign y5125 = n12608 ;
  assign y5126 = ~n12609 ;
  assign y5127 = ~1'b0 ;
  assign y5128 = ~n12611 ;
  assign y5129 = ~n12614 ;
  assign y5130 = n12617 ;
  assign y5131 = n12620 ;
  assign y5132 = ~n12622 ;
  assign y5133 = n12629 ;
  assign y5134 = ~n10973 ;
  assign y5135 = n12638 ;
  assign y5136 = n12648 ;
  assign y5137 = ~n12653 ;
  assign y5138 = n12655 ;
  assign y5139 = ~n12656 ;
  assign y5140 = ~n12657 ;
  assign y5141 = ~n12659 ;
  assign y5142 = ~n12660 ;
  assign y5143 = ~1'b0 ;
  assign y5144 = ~n12661 ;
  assign y5145 = ~n12662 ;
  assign y5146 = ~1'b0 ;
  assign y5147 = n12665 ;
  assign y5148 = n12668 ;
  assign y5149 = ~1'b0 ;
  assign y5150 = ~1'b0 ;
  assign y5151 = ~n12672 ;
  assign y5152 = n12676 ;
  assign y5153 = ~1'b0 ;
  assign y5154 = ~1'b0 ;
  assign y5155 = n12677 ;
  assign y5156 = ~n12678 ;
  assign y5157 = n12680 ;
  assign y5158 = n12683 ;
  assign y5159 = ~n12687 ;
  assign y5160 = n12688 ;
  assign y5161 = ~1'b0 ;
  assign y5162 = n12689 ;
  assign y5163 = n12690 ;
  assign y5164 = ~1'b0 ;
  assign y5165 = ~n12691 ;
  assign y5166 = ~n12693 ;
  assign y5167 = ~n12694 ;
  assign y5168 = ~n12696 ;
  assign y5169 = ~1'b0 ;
  assign y5170 = ~n12698 ;
  assign y5171 = ~n12700 ;
  assign y5172 = ~n12701 ;
  assign y5173 = ~1'b0 ;
  assign y5174 = ~n12703 ;
  assign y5175 = ~1'b0 ;
  assign y5176 = n12709 ;
  assign y5177 = n12710 ;
  assign y5178 = ~1'b0 ;
  assign y5179 = ~1'b0 ;
  assign y5180 = n12711 ;
  assign y5181 = n12712 ;
  assign y5182 = n12713 ;
  assign y5183 = n12715 ;
  assign y5184 = n12717 ;
  assign y5185 = n12720 ;
  assign y5186 = n12721 ;
  assign y5187 = n12724 ;
  assign y5188 = ~1'b0 ;
  assign y5189 = ~n12731 ;
  assign y5190 = n12733 ;
  assign y5191 = ~1'b0 ;
  assign y5192 = n12741 ;
  assign y5193 = ~n12743 ;
  assign y5194 = ~n12745 ;
  assign y5195 = ~n12746 ;
  assign y5196 = ~n12748 ;
  assign y5197 = ~1'b0 ;
  assign y5198 = ~n12752 ;
  assign y5199 = ~n12754 ;
  assign y5200 = n12763 ;
  assign y5201 = ~1'b0 ;
  assign y5202 = n10121 ;
  assign y5203 = n12769 ;
  assign y5204 = n12772 ;
  assign y5205 = n12773 ;
  assign y5206 = ~n12775 ;
  assign y5207 = ~1'b0 ;
  assign y5208 = ~1'b0 ;
  assign y5209 = n12780 ;
  assign y5210 = ~n12786 ;
  assign y5211 = ~n3480 ;
  assign y5212 = n12798 ;
  assign y5213 = ~1'b0 ;
  assign y5214 = ~n12799 ;
  assign y5215 = n12802 ;
  assign y5216 = n12804 ;
  assign y5217 = 1'b0 ;
  assign y5218 = ~1'b0 ;
  assign y5219 = n12806 ;
  assign y5220 = ~n12808 ;
  assign y5221 = ~n12809 ;
  assign y5222 = ~n12812 ;
  assign y5223 = n12815 ;
  assign y5224 = n12816 ;
  assign y5225 = ~n12820 ;
  assign y5226 = ~n12828 ;
  assign y5227 = ~1'b0 ;
  assign y5228 = n12830 ;
  assign y5229 = n12832 ;
  assign y5230 = ~n12835 ;
  assign y5231 = 1'b0 ;
  assign y5232 = ~n3490 ;
  assign y5233 = ~n12841 ;
  assign y5234 = n12843 ;
  assign y5235 = n12846 ;
  assign y5236 = n12851 ;
  assign y5237 = ~n12855 ;
  assign y5238 = n12860 ;
  assign y5239 = ~1'b0 ;
  assign y5240 = ~n12862 ;
  assign y5241 = ~n12863 ;
  assign y5242 = ~n12865 ;
  assign y5243 = ~1'b0 ;
  assign y5244 = n12866 ;
  assign y5245 = n12874 ;
  assign y5246 = ~n12879 ;
  assign y5247 = ~1'b0 ;
  assign y5248 = n1291 ;
  assign y5249 = ~n12884 ;
  assign y5250 = ~n12887 ;
  assign y5251 = ~n12888 ;
  assign y5252 = n12892 ;
  assign y5253 = ~n12895 ;
  assign y5254 = n12902 ;
  assign y5255 = n12905 ;
  assign y5256 = ~1'b0 ;
  assign y5257 = n12660 ;
  assign y5258 = ~n12910 ;
  assign y5259 = ~1'b0 ;
  assign y5260 = ~1'b0 ;
  assign y5261 = ~1'b0 ;
  assign y5262 = ~n12916 ;
  assign y5263 = ~n12918 ;
  assign y5264 = n12927 ;
  assign y5265 = ~n12933 ;
  assign y5266 = n12934 ;
  assign y5267 = ~n12936 ;
  assign y5268 = ~1'b0 ;
  assign y5269 = n12940 ;
  assign y5270 = ~n9317 ;
  assign y5271 = ~n12944 ;
  assign y5272 = n12946 ;
  assign y5273 = ~n12950 ;
  assign y5274 = ~n12952 ;
  assign y5275 = ~n12955 ;
  assign y5276 = n12958 ;
  assign y5277 = ~n12959 ;
  assign y5278 = n12961 ;
  assign y5279 = ~n12963 ;
  assign y5280 = ~n12970 ;
  assign y5281 = n12971 ;
  assign y5282 = n12973 ;
  assign y5283 = ~n12976 ;
  assign y5284 = n12908 ;
  assign y5285 = ~n12977 ;
  assign y5286 = ~1'b0 ;
  assign y5287 = ~n2495 ;
  assign y5288 = n12983 ;
  assign y5289 = ~n12990 ;
  assign y5290 = ~n12991 ;
  assign y5291 = ~1'b0 ;
  assign y5292 = ~1'b0 ;
  assign y5293 = ~n12993 ;
  assign y5294 = n12994 ;
  assign y5295 = n12998 ;
  assign y5296 = ~1'b0 ;
  assign y5297 = ~1'b0 ;
  assign y5298 = 1'b0 ;
  assign y5299 = ~1'b0 ;
  assign y5300 = ~n13004 ;
  assign y5301 = n13007 ;
  assign y5302 = ~n13011 ;
  assign y5303 = ~n13012 ;
  assign y5304 = ~1'b0 ;
  assign y5305 = n13015 ;
  assign y5306 = ~n13026 ;
  assign y5307 = ~1'b0 ;
  assign y5308 = ~n13028 ;
  assign y5309 = ~1'b0 ;
  assign y5310 = ~n13033 ;
  assign y5311 = ~n13037 ;
  assign y5312 = ~n13044 ;
  assign y5313 = n13050 ;
  assign y5314 = n13053 ;
  assign y5315 = ~n13055 ;
  assign y5316 = n13056 ;
  assign y5317 = n13057 ;
  assign y5318 = ~n13061 ;
  assign y5319 = ~n13064 ;
  assign y5320 = n13075 ;
  assign y5321 = n13079 ;
  assign y5322 = n13080 ;
  assign y5323 = ~1'b0 ;
  assign y5324 = ~1'b0 ;
  assign y5325 = n13090 ;
  assign y5326 = ~n5997 ;
  assign y5327 = ~1'b0 ;
  assign y5328 = n13094 ;
  assign y5329 = ~n13095 ;
  assign y5330 = n13096 ;
  assign y5331 = n13113 ;
  assign y5332 = ~n13114 ;
  assign y5333 = ~n13116 ;
  assign y5334 = ~n13117 ;
  assign y5335 = ~n13119 ;
  assign y5336 = ~n13121 ;
  assign y5337 = ~n13123 ;
  assign y5338 = n13125 ;
  assign y5339 = ~n13128 ;
  assign y5340 = 1'b0 ;
  assign y5341 = ~1'b0 ;
  assign y5342 = ~n13134 ;
  assign y5343 = ~n13135 ;
  assign y5344 = ~n13139 ;
  assign y5345 = ~n13144 ;
  assign y5346 = n13146 ;
  assign y5347 = ~n13151 ;
  assign y5348 = ~1'b0 ;
  assign y5349 = ~n7796 ;
  assign y5350 = n13155 ;
  assign y5351 = ~1'b0 ;
  assign y5352 = ~1'b0 ;
  assign y5353 = ~n13160 ;
  assign y5354 = ~n13169 ;
  assign y5355 = ~n13172 ;
  assign y5356 = ~n13174 ;
  assign y5357 = ~n4060 ;
  assign y5358 = n13175 ;
  assign y5359 = n13176 ;
  assign y5360 = ~1'b0 ;
  assign y5361 = ~1'b0 ;
  assign y5362 = n13181 ;
  assign y5363 = ~1'b0 ;
  assign y5364 = n13182 ;
  assign y5365 = ~1'b0 ;
  assign y5366 = ~n13185 ;
  assign y5367 = n13188 ;
  assign y5368 = ~n13191 ;
  assign y5369 = ~n10032 ;
  assign y5370 = n13192 ;
  assign y5371 = ~1'b0 ;
  assign y5372 = n8627 ;
  assign y5373 = ~n13198 ;
  assign y5374 = n13199 ;
  assign y5375 = n13202 ;
  assign y5376 = ~n13203 ;
  assign y5377 = n13204 ;
  assign y5378 = n13206 ;
  assign y5379 = n13207 ;
  assign y5380 = ~n13211 ;
  assign y5381 = ~1'b0 ;
  assign y5382 = ~n13214 ;
  assign y5383 = ~n13215 ;
  assign y5384 = n13217 ;
  assign y5385 = ~n13218 ;
  assign y5386 = n13221 ;
  assign y5387 = ~n13225 ;
  assign y5388 = ~n13227 ;
  assign y5389 = ~n13234 ;
  assign y5390 = ~n13235 ;
  assign y5391 = ~n13236 ;
  assign y5392 = n13237 ;
  assign y5393 = ~1'b0 ;
  assign y5394 = ~n13238 ;
  assign y5395 = ~n13244 ;
  assign y5396 = ~n13249 ;
  assign y5397 = ~n13253 ;
  assign y5398 = ~1'b0 ;
  assign y5399 = ~n13254 ;
  assign y5400 = n13255 ;
  assign y5401 = n13257 ;
  assign y5402 = ~1'b0 ;
  assign y5403 = n13262 ;
  assign y5404 = n13264 ;
  assign y5405 = ~1'b0 ;
  assign y5406 = n13265 ;
  assign y5407 = ~n13268 ;
  assign y5408 = ~1'b0 ;
  assign y5409 = ~n13271 ;
  assign y5410 = n13274 ;
  assign y5411 = n13276 ;
  assign y5412 = n6895 ;
  assign y5413 = ~n13278 ;
  assign y5414 = ~n13282 ;
  assign y5415 = ~n13286 ;
  assign y5416 = ~n13289 ;
  assign y5417 = ~1'b0 ;
  assign y5418 = ~n13291 ;
  assign y5419 = ~n13292 ;
  assign y5420 = n13296 ;
  assign y5421 = ~n13299 ;
  assign y5422 = ~n13307 ;
  assign y5423 = n13313 ;
  assign y5424 = ~1'b0 ;
  assign y5425 = ~n13314 ;
  assign y5426 = ~n13319 ;
  assign y5427 = n13320 ;
  assign y5428 = n13325 ;
  assign y5429 = ~n13327 ;
  assign y5430 = 1'b0 ;
  assign y5431 = ~n13332 ;
  assign y5432 = ~1'b0 ;
  assign y5433 = n13339 ;
  assign y5434 = ~1'b0 ;
  assign y5435 = ~n13340 ;
  assign y5436 = ~1'b0 ;
  assign y5437 = n13342 ;
  assign y5438 = ~n12947 ;
  assign y5439 = ~n13344 ;
  assign y5440 = ~1'b0 ;
  assign y5441 = n13351 ;
  assign y5442 = ~1'b0 ;
  assign y5443 = n13353 ;
  assign y5444 = ~1'b0 ;
  assign y5445 = ~1'b0 ;
  assign y5446 = ~1'b0 ;
  assign y5447 = ~1'b0 ;
  assign y5448 = n13354 ;
  assign y5449 = n13359 ;
  assign y5450 = ~n13367 ;
  assign y5451 = n13371 ;
  assign y5452 = ~n13372 ;
  assign y5453 = ~1'b0 ;
  assign y5454 = ~1'b0 ;
  assign y5455 = ~n13375 ;
  assign y5456 = n13378 ;
  assign y5457 = ~1'b0 ;
  assign y5458 = ~n13381 ;
  assign y5459 = ~1'b0 ;
  assign y5460 = ~1'b0 ;
  assign y5461 = ~n13390 ;
  assign y5462 = n13394 ;
  assign y5463 = ~n13396 ;
  assign y5464 = n13397 ;
  assign y5465 = ~1'b0 ;
  assign y5466 = ~n13402 ;
  assign y5467 = n13407 ;
  assign y5468 = ~n13408 ;
  assign y5469 = ~n13409 ;
  assign y5470 = ~n13411 ;
  assign y5471 = ~n13413 ;
  assign y5472 = ~n13415 ;
  assign y5473 = n261 ;
  assign y5474 = ~1'b0 ;
  assign y5475 = ~n13418 ;
  assign y5476 = ~1'b0 ;
  assign y5477 = ~1'b0 ;
  assign y5478 = n13421 ;
  assign y5479 = 1'b0 ;
  assign y5480 = ~n13433 ;
  assign y5481 = ~n13439 ;
  assign y5482 = n13445 ;
  assign y5483 = ~n13447 ;
  assign y5484 = ~1'b0 ;
  assign y5485 = ~1'b0 ;
  assign y5486 = n13454 ;
  assign y5487 = n13462 ;
  assign y5488 = ~n13466 ;
  assign y5489 = n13471 ;
  assign y5490 = ~n4136 ;
  assign y5491 = n13474 ;
  assign y5492 = ~n13477 ;
  assign y5493 = ~1'b0 ;
  assign y5494 = ~n13479 ;
  assign y5495 = ~1'b0 ;
  assign y5496 = ~n4150 ;
  assign y5497 = n13482 ;
  assign y5498 = ~n13484 ;
  assign y5499 = ~1'b0 ;
  assign y5500 = ~1'b0 ;
  assign y5501 = ~n3480 ;
  assign y5502 = ~n13488 ;
  assign y5503 = n13491 ;
  assign y5504 = n13494 ;
  assign y5505 = ~n13497 ;
  assign y5506 = ~n13508 ;
  assign y5507 = n13509 ;
  assign y5508 = ~n13515 ;
  assign y5509 = ~n13528 ;
  assign y5510 = ~1'b0 ;
  assign y5511 = ~n8102 ;
  assign y5512 = n13531 ;
  assign y5513 = ~1'b0 ;
  assign y5514 = n13535 ;
  assign y5515 = ~1'b0 ;
  assign y5516 = n13536 ;
  assign y5517 = ~n13537 ;
  assign y5518 = n13540 ;
  assign y5519 = ~n13542 ;
  assign y5520 = n13546 ;
  assign y5521 = n13550 ;
  assign y5522 = n13551 ;
  assign y5523 = ~n13558 ;
  assign y5524 = ~n13559 ;
  assign y5525 = ~n13560 ;
  assign y5526 = ~n13563 ;
  assign y5527 = ~n13564 ;
  assign y5528 = ~1'b0 ;
  assign y5529 = ~1'b0 ;
  assign y5530 = n13565 ;
  assign y5531 = ~n13568 ;
  assign y5532 = ~n13571 ;
  assign y5533 = n13572 ;
  assign y5534 = ~n13575 ;
  assign y5535 = n13578 ;
  assign y5536 = n13579 ;
  assign y5537 = ~n13581 ;
  assign y5538 = ~n13588 ;
  assign y5539 = n2816 ;
  assign y5540 = ~n13598 ;
  assign y5541 = ~n13601 ;
  assign y5542 = ~1'b0 ;
  assign y5543 = ~n13604 ;
  assign y5544 = n11573 ;
  assign y5545 = ~1'b0 ;
  assign y5546 = ~1'b0 ;
  assign y5547 = 1'b0 ;
  assign y5548 = ~n13605 ;
  assign y5549 = ~1'b0 ;
  assign y5550 = ~n13606 ;
  assign y5551 = n13607 ;
  assign y5552 = n13613 ;
  assign y5553 = ~n13631 ;
  assign y5554 = ~n13632 ;
  assign y5555 = n13634 ;
  assign y5556 = ~n13635 ;
  assign y5557 = n13639 ;
  assign y5558 = n13649 ;
  assign y5559 = ~1'b0 ;
  assign y5560 = ~1'b0 ;
  assign y5561 = ~n13650 ;
  assign y5562 = ~n13662 ;
  assign y5563 = ~n13663 ;
  assign y5564 = n13664 ;
  assign y5565 = ~n13670 ;
  assign y5566 = ~1'b0 ;
  assign y5567 = n13671 ;
  assign y5568 = n13673 ;
  assign y5569 = n13674 ;
  assign y5570 = n13676 ;
  assign y5571 = ~n13677 ;
  assign y5572 = 1'b0 ;
  assign y5573 = ~n13682 ;
  assign y5574 = ~n13683 ;
  assign y5575 = ~n13684 ;
  assign y5576 = ~1'b0 ;
  assign y5577 = ~1'b0 ;
  assign y5578 = n13685 ;
  assign y5579 = ~1'b0 ;
  assign y5580 = ~1'b0 ;
  assign y5581 = ~n13693 ;
  assign y5582 = ~1'b0 ;
  assign y5583 = n13698 ;
  assign y5584 = n13700 ;
  assign y5585 = ~n13703 ;
  assign y5586 = ~1'b0 ;
  assign y5587 = ~1'b0 ;
  assign y5588 = ~n10850 ;
  assign y5589 = ~n12360 ;
  assign y5590 = ~1'b0 ;
  assign y5591 = n13704 ;
  assign y5592 = ~n13707 ;
  assign y5593 = ~n13708 ;
  assign y5594 = n13709 ;
  assign y5595 = ~n13713 ;
  assign y5596 = x158 ;
  assign y5597 = n13718 ;
  assign y5598 = ~1'b0 ;
  assign y5599 = ~n13720 ;
  assign y5600 = ~n13722 ;
  assign y5601 = ~n13723 ;
  assign y5602 = ~n13726 ;
  assign y5603 = n5369 ;
  assign y5604 = n13729 ;
  assign y5605 = ~1'b0 ;
  assign y5606 = ~n13730 ;
  assign y5607 = ~n13737 ;
  assign y5608 = n13739 ;
  assign y5609 = ~n13741 ;
  assign y5610 = ~1'b0 ;
  assign y5611 = n8888 ;
  assign y5612 = n13747 ;
  assign y5613 = ~n13752 ;
  assign y5614 = n13754 ;
  assign y5615 = n13758 ;
  assign y5616 = ~1'b0 ;
  assign y5617 = ~1'b0 ;
  assign y5618 = n13762 ;
  assign y5619 = n13765 ;
  assign y5620 = n13766 ;
  assign y5621 = n13768 ;
  assign y5622 = ~n13769 ;
  assign y5623 = ~1'b0 ;
  assign y5624 = n13772 ;
  assign y5625 = n13777 ;
  assign y5626 = n13778 ;
  assign y5627 = n13780 ;
  assign y5628 = ~n13783 ;
  assign y5629 = ~n13789 ;
  assign y5630 = ~n13790 ;
  assign y5631 = n13791 ;
  assign y5632 = ~n13795 ;
  assign y5633 = ~1'b0 ;
  assign y5634 = ~n13796 ;
  assign y5635 = ~1'b0 ;
  assign y5636 = n13797 ;
  assign y5637 = n13803 ;
  assign y5638 = ~1'b0 ;
  assign y5639 = n13806 ;
  assign y5640 = ~1'b0 ;
  assign y5641 = ~1'b0 ;
  assign y5642 = ~1'b0 ;
  assign y5643 = ~1'b0 ;
  assign y5644 = n13807 ;
  assign y5645 = ~1'b0 ;
  assign y5646 = ~1'b0 ;
  assign y5647 = ~n13809 ;
  assign y5648 = n13812 ;
  assign y5649 = ~1'b0 ;
  assign y5650 = ~n5013 ;
  assign y5651 = n13818 ;
  assign y5652 = ~n13819 ;
  assign y5653 = ~n13821 ;
  assign y5654 = n13824 ;
  assign y5655 = ~n13827 ;
  assign y5656 = n13830 ;
  assign y5657 = ~n13834 ;
  assign y5658 = n13835 ;
  assign y5659 = ~n13841 ;
  assign y5660 = 1'b0 ;
  assign y5661 = n5028 ;
  assign y5662 = ~1'b0 ;
  assign y5663 = n13842 ;
  assign y5664 = ~n13844 ;
  assign y5665 = ~1'b0 ;
  assign y5666 = n13846 ;
  assign y5667 = n13847 ;
  assign y5668 = ~n13850 ;
  assign y5669 = n13852 ;
  assign y5670 = n13853 ;
  assign y5671 = ~n13854 ;
  assign y5672 = ~n13859 ;
  assign y5673 = n13861 ;
  assign y5674 = 1'b0 ;
  assign y5675 = ~1'b0 ;
  assign y5676 = ~n13863 ;
  assign y5677 = ~n13867 ;
  assign y5678 = ~n13878 ;
  assign y5679 = n13879 ;
  assign y5680 = ~1'b0 ;
  assign y5681 = ~1'b0 ;
  assign y5682 = ~1'b0 ;
  assign y5683 = ~n13883 ;
  assign y5684 = ~1'b0 ;
  assign y5685 = ~1'b0 ;
  assign y5686 = ~n13890 ;
  assign y5687 = ~n13893 ;
  assign y5688 = ~n13903 ;
  assign y5689 = 1'b0 ;
  assign y5690 = ~1'b0 ;
  assign y5691 = ~1'b0 ;
  assign y5692 = ~n13904 ;
  assign y5693 = ~1'b0 ;
  assign y5694 = ~n13906 ;
  assign y5695 = n13909 ;
  assign y5696 = n13919 ;
  assign y5697 = n13921 ;
  assign y5698 = n13923 ;
  assign y5699 = ~n13931 ;
  assign y5700 = ~n13932 ;
  assign y5701 = ~n13934 ;
  assign y5702 = ~1'b0 ;
  assign y5703 = ~n13937 ;
  assign y5704 = 1'b0 ;
  assign y5705 = ~n13938 ;
  assign y5706 = n7270 ;
  assign y5707 = n13947 ;
  assign y5708 = n13948 ;
  assign y5709 = n13949 ;
  assign y5710 = ~1'b0 ;
  assign y5711 = ~n13955 ;
  assign y5712 = n13956 ;
  assign y5713 = ~n13957 ;
  assign y5714 = ~1'b0 ;
  assign y5715 = n13964 ;
  assign y5716 = ~n7380 ;
  assign y5717 = ~1'b0 ;
  assign y5718 = ~n13968 ;
  assign y5719 = ~1'b0 ;
  assign y5720 = n13972 ;
  assign y5721 = n13973 ;
  assign y5722 = ~n13976 ;
  assign y5723 = ~1'b0 ;
  assign y5724 = n13980 ;
  assign y5725 = n13992 ;
  assign y5726 = n13994 ;
  assign y5727 = ~n14002 ;
  assign y5728 = ~n14009 ;
  assign y5729 = n14014 ;
  assign y5730 = ~n14015 ;
  assign y5731 = n6188 ;
  assign y5732 = ~1'b0 ;
  assign y5733 = ~n14027 ;
  assign y5734 = ~1'b0 ;
  assign y5735 = n14032 ;
  assign y5736 = n14034 ;
  assign y5737 = n14040 ;
  assign y5738 = n14041 ;
  assign y5739 = ~1'b0 ;
  assign y5740 = n14045 ;
  assign y5741 = ~n14048 ;
  assign y5742 = n14052 ;
  assign y5743 = n14054 ;
  assign y5744 = ~n14055 ;
  assign y5745 = n14058 ;
  assign y5746 = ~n14061 ;
  assign y5747 = n14065 ;
  assign y5748 = ~1'b0 ;
  assign y5749 = n14068 ;
  assign y5750 = n9302 ;
  assign y5751 = ~1'b0 ;
  assign y5752 = ~1'b0 ;
  assign y5753 = n14070 ;
  assign y5754 = ~n14075 ;
  assign y5755 = n14076 ;
  assign y5756 = n14081 ;
  assign y5757 = ~1'b0 ;
  assign y5758 = n14088 ;
  assign y5759 = ~1'b0 ;
  assign y5760 = ~1'b0 ;
  assign y5761 = n14092 ;
  assign y5762 = ~n14098 ;
  assign y5763 = n14102 ;
  assign y5764 = n14104 ;
  assign y5765 = ~1'b0 ;
  assign y5766 = n5404 ;
  assign y5767 = n14111 ;
  assign y5768 = n14112 ;
  assign y5769 = ~1'b0 ;
  assign y5770 = ~1'b0 ;
  assign y5771 = n14113 ;
  assign y5772 = ~1'b0 ;
  assign y5773 = n14115 ;
  assign y5774 = ~n14117 ;
  assign y5775 = ~n14119 ;
  assign y5776 = n14120 ;
  assign y5777 = n14125 ;
  assign y5778 = ~1'b0 ;
  assign y5779 = n14129 ;
  assign y5780 = ~1'b0 ;
  assign y5781 = ~1'b0 ;
  assign y5782 = ~n14136 ;
  assign y5783 = ~n14137 ;
  assign y5784 = ~n14138 ;
  assign y5785 = ~1'b0 ;
  assign y5786 = ~1'b0 ;
  assign y5787 = n14140 ;
  assign y5788 = ~n14141 ;
  assign y5789 = n7718 ;
  assign y5790 = ~n14147 ;
  assign y5791 = ~1'b0 ;
  assign y5792 = n9688 ;
  assign y5793 = ~1'b0 ;
  assign y5794 = ~n14149 ;
  assign y5795 = n14155 ;
  assign y5796 = ~1'b0 ;
  assign y5797 = ~n14157 ;
  assign y5798 = ~1'b0 ;
  assign y5799 = n14161 ;
  assign y5800 = ~n14165 ;
  assign y5801 = ~1'b0 ;
  assign y5802 = n14166 ;
  assign y5803 = ~n14170 ;
  assign y5804 = ~n14173 ;
  assign y5805 = n14176 ;
  assign y5806 = ~n14177 ;
  assign y5807 = ~n14183 ;
  assign y5808 = n14185 ;
  assign y5809 = ~n14188 ;
  assign y5810 = 1'b0 ;
  assign y5811 = n14190 ;
  assign y5812 = ~n14192 ;
  assign y5813 = ~n14196 ;
  assign y5814 = ~n14197 ;
  assign y5815 = n2120 ;
  assign y5816 = n14198 ;
  assign y5817 = ~n14200 ;
  assign y5818 = n14206 ;
  assign y5819 = ~1'b0 ;
  assign y5820 = n14207 ;
  assign y5821 = n14210 ;
  assign y5822 = ~n14216 ;
  assign y5823 = n14217 ;
  assign y5824 = ~n14218 ;
  assign y5825 = ~1'b0 ;
  assign y5826 = n14219 ;
  assign y5827 = n14224 ;
  assign y5828 = n14226 ;
  assign y5829 = n14228 ;
  assign y5830 = n14237 ;
  assign y5831 = ~n14242 ;
  assign y5832 = x70 ;
  assign y5833 = n14244 ;
  assign y5834 = n14246 ;
  assign y5835 = ~1'b0 ;
  assign y5836 = ~1'b0 ;
  assign y5837 = ~n14247 ;
  assign y5838 = ~n14250 ;
  assign y5839 = ~n14253 ;
  assign y5840 = n14255 ;
  assign y5841 = 1'b0 ;
  assign y5842 = ~n14257 ;
  assign y5843 = n14259 ;
  assign y5844 = n14267 ;
  assign y5845 = ~1'b0 ;
  assign y5846 = ~n14269 ;
  assign y5847 = ~1'b0 ;
  assign y5848 = ~n14270 ;
  assign y5849 = n12802 ;
  assign y5850 = ~1'b0 ;
  assign y5851 = ~1'b0 ;
  assign y5852 = n14273 ;
  assign y5853 = ~1'b0 ;
  assign y5854 = n14278 ;
  assign y5855 = ~n14281 ;
  assign y5856 = n14284 ;
  assign y5857 = ~1'b0 ;
  assign y5858 = ~n14293 ;
  assign y5859 = ~1'b0 ;
  assign y5860 = n14294 ;
  assign y5861 = ~1'b0 ;
  assign y5862 = ~1'b0 ;
  assign y5863 = ~1'b0 ;
  assign y5864 = ~1'b0 ;
  assign y5865 = ~1'b0 ;
  assign y5866 = ~1'b0 ;
  assign y5867 = ~n14296 ;
  assign y5868 = n13982 ;
  assign y5869 = n9900 ;
  assign y5870 = ~1'b0 ;
  assign y5871 = n14300 ;
  assign y5872 = ~n14308 ;
  assign y5873 = ~n14312 ;
  assign y5874 = ~n14313 ;
  assign y5875 = ~n14318 ;
  assign y5876 = ~1'b0 ;
  assign y5877 = n14319 ;
  assign y5878 = n14320 ;
  assign y5879 = n14324 ;
  assign y5880 = n14326 ;
  assign y5881 = n14328 ;
  assign y5882 = ~n14332 ;
  assign y5883 = n14334 ;
  assign y5884 = ~1'b0 ;
  assign y5885 = ~n14335 ;
  assign y5886 = n14338 ;
  assign y5887 = ~n14342 ;
  assign y5888 = ~n14346 ;
  assign y5889 = ~n14347 ;
  assign y5890 = n14350 ;
  assign y5891 = ~1'b0 ;
  assign y5892 = ~n14352 ;
  assign y5893 = ~n14354 ;
  assign y5894 = ~n14356 ;
  assign y5895 = ~n14357 ;
  assign y5896 = ~n14362 ;
  assign y5897 = ~1'b0 ;
  assign y5898 = ~1'b0 ;
  assign y5899 = ~n14364 ;
  assign y5900 = n14367 ;
  assign y5901 = ~1'b0 ;
  assign y5902 = ~1'b0 ;
  assign y5903 = n14370 ;
  assign y5904 = ~n14372 ;
  assign y5905 = ~1'b0 ;
  assign y5906 = ~1'b0 ;
  assign y5907 = 1'b0 ;
  assign y5908 = ~1'b0 ;
  assign y5909 = n14373 ;
  assign y5910 = ~n4468 ;
  assign y5911 = n14375 ;
  assign y5912 = n14379 ;
  assign y5913 = n14380 ;
  assign y5914 = n14383 ;
  assign y5915 = ~n14392 ;
  assign y5916 = n14394 ;
  assign y5917 = ~n802 ;
  assign y5918 = ~1'b0 ;
  assign y5919 = n14401 ;
  assign y5920 = ~n14406 ;
  assign y5921 = ~1'b0 ;
  assign y5922 = n14408 ;
  assign y5923 = ~n14412 ;
  assign y5924 = ~n14417 ;
  assign y5925 = ~n14419 ;
  assign y5926 = ~n14422 ;
  assign y5927 = ~1'b0 ;
  assign y5928 = ~1'b0 ;
  assign y5929 = ~1'b0 ;
  assign y5930 = ~1'b0 ;
  assign y5931 = n14424 ;
  assign y5932 = ~n14425 ;
  assign y5933 = ~n14429 ;
  assign y5934 = n14430 ;
  assign y5935 = ~1'b0 ;
  assign y5936 = ~1'b0 ;
  assign y5937 = ~n14435 ;
  assign y5938 = ~n14439 ;
  assign y5939 = ~1'b0 ;
  assign y5940 = ~n14443 ;
  assign y5941 = n14449 ;
  assign y5942 = ~n14460 ;
  assign y5943 = n14467 ;
  assign y5944 = n14468 ;
  assign y5945 = ~n14470 ;
  assign y5946 = ~1'b0 ;
  assign y5947 = ~n14471 ;
  assign y5948 = ~1'b0 ;
  assign y5949 = ~1'b0 ;
  assign y5950 = n14473 ;
  assign y5951 = ~1'b0 ;
  assign y5952 = n14477 ;
  assign y5953 = n14481 ;
  assign y5954 = n14490 ;
  assign y5955 = n14493 ;
  assign y5956 = n14495 ;
  assign y5957 = ~n14500 ;
  assign y5958 = ~n14505 ;
  assign y5959 = ~1'b0 ;
  assign y5960 = ~1'b0 ;
  assign y5961 = n14509 ;
  assign y5962 = ~n14515 ;
  assign y5963 = ~1'b0 ;
  assign y5964 = ~n14518 ;
  assign y5965 = n14521 ;
  assign y5966 = ~1'b0 ;
  assign y5967 = ~1'b0 ;
  assign y5968 = ~n14525 ;
  assign y5969 = ~n14527 ;
  assign y5970 = ~n14533 ;
  assign y5971 = n14534 ;
  assign y5972 = ~n14539 ;
  assign y5973 = ~n14540 ;
  assign y5974 = n13685 ;
  assign y5975 = n14547 ;
  assign y5976 = n14548 ;
  assign y5977 = n14550 ;
  assign y5978 = n14553 ;
  assign y5979 = ~1'b0 ;
  assign y5980 = ~1'b0 ;
  assign y5981 = ~1'b0 ;
  assign y5982 = ~n14556 ;
  assign y5983 = ~n14560 ;
  assign y5984 = n14567 ;
  assign y5985 = ~1'b0 ;
  assign y5986 = n14569 ;
  assign y5987 = ~n14578 ;
  assign y5988 = n14581 ;
  assign y5989 = ~1'b0 ;
  assign y5990 = ~n14586 ;
  assign y5991 = 1'b0 ;
  assign y5992 = ~n14592 ;
  assign y5993 = ~n14593 ;
  assign y5994 = ~n14594 ;
  assign y5995 = n14596 ;
  assign y5996 = n14598 ;
  assign y5997 = n14605 ;
  assign y5998 = ~n14607 ;
  assign y5999 = n14612 ;
  assign y6000 = ~1'b0 ;
  assign y6001 = ~n14613 ;
  assign y6002 = n14621 ;
  assign y6003 = ~1'b0 ;
  assign y6004 = ~1'b0 ;
  assign y6005 = ~n14624 ;
  assign y6006 = ~n14627 ;
  assign y6007 = n14629 ;
  assign y6008 = n14630 ;
  assign y6009 = ~1'b0 ;
  assign y6010 = ~1'b0 ;
  assign y6011 = ~n14632 ;
  assign y6012 = n14635 ;
  assign y6013 = ~1'b0 ;
  assign y6014 = ~1'b0 ;
  assign y6015 = n14642 ;
  assign y6016 = ~n14645 ;
  assign y6017 = ~1'b0 ;
  assign y6018 = n14650 ;
  assign y6019 = n14660 ;
  assign y6020 = n14662 ;
  assign y6021 = n14665 ;
  assign y6022 = ~1'b0 ;
  assign y6023 = n14666 ;
  assign y6024 = ~n14669 ;
  assign y6025 = ~1'b0 ;
  assign y6026 = ~n14672 ;
  assign y6027 = ~n11532 ;
  assign y6028 = n14673 ;
  assign y6029 = n14677 ;
  assign y6030 = ~1'b0 ;
  assign y6031 = ~1'b0 ;
  assign y6032 = ~n14679 ;
  assign y6033 = n14681 ;
  assign y6034 = n14689 ;
  assign y6035 = ~1'b0 ;
  assign y6036 = ~n14694 ;
  assign y6037 = n14706 ;
  assign y6038 = n14709 ;
  assign y6039 = 1'b0 ;
  assign y6040 = ~1'b0 ;
  assign y6041 = ~n9577 ;
  assign y6042 = ~n14710 ;
  assign y6043 = ~1'b0 ;
  assign y6044 = ~1'b0 ;
  assign y6045 = n14716 ;
  assign y6046 = ~1'b0 ;
  assign y6047 = ~1'b0 ;
  assign y6048 = ~1'b0 ;
  assign y6049 = n14720 ;
  assign y6050 = n14723 ;
  assign y6051 = n14724 ;
  assign y6052 = ~n14726 ;
  assign y6053 = n14731 ;
  assign y6054 = ~n14733 ;
  assign y6055 = n14735 ;
  assign y6056 = ~1'b0 ;
  assign y6057 = ~n14739 ;
  assign y6058 = ~n14742 ;
  assign y6059 = ~1'b0 ;
  assign y6060 = ~n14744 ;
  assign y6061 = ~n14746 ;
  assign y6062 = ~1'b0 ;
  assign y6063 = ~n14749 ;
  assign y6064 = ~1'b0 ;
  assign y6065 = ~n14751 ;
  assign y6066 = ~n14752 ;
  assign y6067 = n3422 ;
  assign y6068 = ~n6950 ;
  assign y6069 = ~n14753 ;
  assign y6070 = n14754 ;
  assign y6071 = ~n14765 ;
  assign y6072 = ~n14766 ;
  assign y6073 = ~1'b0 ;
  assign y6074 = ~n14768 ;
  assign y6075 = ~n14772 ;
  assign y6076 = ~n8129 ;
  assign y6077 = ~n14773 ;
  assign y6078 = n14775 ;
  assign y6079 = ~n14776 ;
  assign y6080 = ~n14778 ;
  assign y6081 = ~1'b0 ;
  assign y6082 = n14782 ;
  assign y6083 = ~n14789 ;
  assign y6084 = n14795 ;
  assign y6085 = ~n14796 ;
  assign y6086 = n14798 ;
  assign y6087 = ~n3490 ;
  assign y6088 = n14799 ;
  assign y6089 = n14801 ;
  assign y6090 = n14803 ;
  assign y6091 = ~x158 ;
  assign y6092 = n14804 ;
  assign y6093 = ~1'b0 ;
  assign y6094 = ~n14811 ;
  assign y6095 = n14813 ;
  assign y6096 = n14814 ;
  assign y6097 = n14815 ;
  assign y6098 = ~n14821 ;
  assign y6099 = ~n1801 ;
  assign y6100 = ~n14829 ;
  assign y6101 = ~1'b0 ;
  assign y6102 = ~n14830 ;
  assign y6103 = n14831 ;
  assign y6104 = ~1'b0 ;
  assign y6105 = ~n14835 ;
  assign y6106 = ~n14837 ;
  assign y6107 = ~n14838 ;
  assign y6108 = ~n14839 ;
  assign y6109 = n14841 ;
  assign y6110 = ~n14842 ;
  assign y6111 = ~n7700 ;
  assign y6112 = n14844 ;
  assign y6113 = ~1'b0 ;
  assign y6114 = ~n14845 ;
  assign y6115 = n14851 ;
  assign y6116 = n14854 ;
  assign y6117 = n14859 ;
  assign y6118 = ~1'b0 ;
  assign y6119 = ~1'b0 ;
  assign y6120 = ~1'b0 ;
  assign y6121 = n14860 ;
  assign y6122 = n12277 ;
  assign y6123 = n14863 ;
  assign y6124 = ~1'b0 ;
  assign y6125 = ~1'b0 ;
  assign y6126 = n14867 ;
  assign y6127 = ~1'b0 ;
  assign y6128 = n14870 ;
  assign y6129 = n14872 ;
  assign y6130 = n14875 ;
  assign y6131 = n14877 ;
  assign y6132 = ~1'b0 ;
  assign y6133 = n14879 ;
  assign y6134 = n14881 ;
  assign y6135 = 1'b0 ;
  assign y6136 = ~n14883 ;
  assign y6137 = ~1'b0 ;
  assign y6138 = n14886 ;
  assign y6139 = ~n14895 ;
  assign y6140 = n14898 ;
  assign y6141 = ~n14900 ;
  assign y6142 = ~n14901 ;
  assign y6143 = n14904 ;
  assign y6144 = n14907 ;
  assign y6145 = ~n14908 ;
  assign y6146 = ~1'b0 ;
  assign y6147 = ~n14915 ;
  assign y6148 = ~1'b0 ;
  assign y6149 = n4950 ;
  assign y6150 = n14920 ;
  assign y6151 = n14922 ;
  assign y6152 = ~1'b0 ;
  assign y6153 = ~n14923 ;
  assign y6154 = ~n661 ;
  assign y6155 = ~n14930 ;
  assign y6156 = ~1'b0 ;
  assign y6157 = ~n14933 ;
  assign y6158 = n14936 ;
  assign y6159 = ~n14945 ;
  assign y6160 = n14948 ;
  assign y6161 = ~n11117 ;
  assign y6162 = 1'b0 ;
  assign y6163 = ~n14949 ;
  assign y6164 = n14955 ;
  assign y6165 = ~1'b0 ;
  assign y6166 = ~1'b0 ;
  assign y6167 = ~1'b0 ;
  assign y6168 = ~n14961 ;
  assign y6169 = n14963 ;
  assign y6170 = ~n14966 ;
  assign y6171 = ~n14967 ;
  assign y6172 = ~1'b0 ;
  assign y6173 = n14968 ;
  assign y6174 = ~1'b0 ;
  assign y6175 = ~1'b0 ;
  assign y6176 = ~n14970 ;
  assign y6177 = ~n14972 ;
  assign y6178 = ~n14976 ;
  assign y6179 = n14979 ;
  assign y6180 = ~n14982 ;
  assign y6181 = n14988 ;
  assign y6182 = ~1'b0 ;
  assign y6183 = n14989 ;
  assign y6184 = ~n14990 ;
  assign y6185 = ~n14991 ;
  assign y6186 = n14993 ;
  assign y6187 = ~n14996 ;
  assign y6188 = ~1'b0 ;
  assign y6189 = ~n14998 ;
  assign y6190 = 1'b0 ;
  assign y6191 = n14999 ;
  assign y6192 = n15001 ;
  assign y6193 = n15004 ;
  assign y6194 = n15006 ;
  assign y6195 = n15011 ;
  assign y6196 = ~n9491 ;
  assign y6197 = ~n15014 ;
  assign y6198 = ~n15016 ;
  assign y6199 = ~n15018 ;
  assign y6200 = ~n15019 ;
  assign y6201 = n15031 ;
  assign y6202 = ~1'b0 ;
  assign y6203 = n15032 ;
  assign y6204 = ~1'b0 ;
  assign y6205 = ~n15033 ;
  assign y6206 = ~n15040 ;
  assign y6207 = ~1'b0 ;
  assign y6208 = n15043 ;
  assign y6209 = ~n15044 ;
  assign y6210 = n15047 ;
  assign y6211 = 1'b0 ;
  assign y6212 = ~n15051 ;
  assign y6213 = ~n15055 ;
  assign y6214 = n15056 ;
  assign y6215 = n15058 ;
  assign y6216 = ~1'b0 ;
  assign y6217 = ~1'b0 ;
  assign y6218 = n15060 ;
  assign y6219 = ~1'b0 ;
  assign y6220 = ~1'b0 ;
  assign y6221 = ~n15062 ;
  assign y6222 = ~1'b0 ;
  assign y6223 = 1'b0 ;
  assign y6224 = ~n15064 ;
  assign y6225 = ~n15065 ;
  assign y6226 = n15067 ;
  assign y6227 = n15068 ;
  assign y6228 = n15072 ;
  assign y6229 = ~1'b0 ;
  assign y6230 = ~n15073 ;
  assign y6231 = ~n15077 ;
  assign y6232 = ~n15079 ;
  assign y6233 = n15083 ;
  assign y6234 = ~1'b0 ;
  assign y6235 = ~1'b0 ;
  assign y6236 = ~1'b0 ;
  assign y6237 = ~n15084 ;
  assign y6238 = ~1'b0 ;
  assign y6239 = n5914 ;
  assign y6240 = ~1'b0 ;
  assign y6241 = n15086 ;
  assign y6242 = ~n15087 ;
  assign y6243 = n15089 ;
  assign y6244 = ~n15091 ;
  assign y6245 = ~n15093 ;
  assign y6246 = n15113 ;
  assign y6247 = ~1'b0 ;
  assign y6248 = ~1'b0 ;
  assign y6249 = ~n15114 ;
  assign y6250 = n15117 ;
  assign y6251 = ~n11490 ;
  assign y6252 = n15119 ;
  assign y6253 = ~1'b0 ;
  assign y6254 = n15124 ;
  assign y6255 = ~n15130 ;
  assign y6256 = ~n15131 ;
  assign y6257 = ~n15132 ;
  assign y6258 = ~n15133 ;
  assign y6259 = n15134 ;
  assign y6260 = ~n15137 ;
  assign y6261 = ~1'b0 ;
  assign y6262 = ~n15138 ;
  assign y6263 = n15140 ;
  assign y6264 = ~1'b0 ;
  assign y6265 = ~n15144 ;
  assign y6266 = ~1'b0 ;
  assign y6267 = ~n15147 ;
  assign y6268 = ~1'b0 ;
  assign y6269 = n15149 ;
  assign y6270 = n15152 ;
  assign y6271 = ~1'b0 ;
  assign y6272 = ~1'b0 ;
  assign y6273 = ~1'b0 ;
  assign y6274 = ~n15162 ;
  assign y6275 = n15166 ;
  assign y6276 = ~n15169 ;
  assign y6277 = n15174 ;
  assign y6278 = n15175 ;
  assign y6279 = ~1'b0 ;
  assign y6280 = ~n15176 ;
  assign y6281 = ~n10856 ;
  assign y6282 = ~1'b0 ;
  assign y6283 = 1'b0 ;
  assign y6284 = n15178 ;
  assign y6285 = ~1'b0 ;
  assign y6286 = n15184 ;
  assign y6287 = ~1'b0 ;
  assign y6288 = ~1'b0 ;
  assign y6289 = ~1'b0 ;
  assign y6290 = ~n2253 ;
  assign y6291 = n15190 ;
  assign y6292 = ~1'b0 ;
  assign y6293 = ~1'b0 ;
  assign y6294 = ~n15191 ;
  assign y6295 = n7573 ;
  assign y6296 = ~n15198 ;
  assign y6297 = ~n15199 ;
  assign y6298 = n15202 ;
  assign y6299 = n15217 ;
  assign y6300 = ~n15218 ;
  assign y6301 = n15221 ;
  assign y6302 = n15222 ;
  assign y6303 = n15223 ;
  assign y6304 = ~n15225 ;
  assign y6305 = ~1'b0 ;
  assign y6306 = n15226 ;
  assign y6307 = ~n15229 ;
  assign y6308 = n15236 ;
  assign y6309 = ~1'b0 ;
  assign y6310 = n15237 ;
  assign y6311 = ~n15238 ;
  assign y6312 = ~n15244 ;
  assign y6313 = ~n15247 ;
  assign y6314 = n15248 ;
  assign y6315 = ~1'b0 ;
  assign y6316 = ~1'b0 ;
  assign y6317 = ~1'b0 ;
  assign y6318 = ~n15249 ;
  assign y6319 = n15250 ;
  assign y6320 = n15253 ;
  assign y6321 = n15256 ;
  assign y6322 = ~n15259 ;
  assign y6323 = ~n15260 ;
  assign y6324 = ~1'b0 ;
  assign y6325 = n15272 ;
  assign y6326 = ~1'b0 ;
  assign y6327 = ~1'b0 ;
  assign y6328 = ~n15279 ;
  assign y6329 = ~1'b0 ;
  assign y6330 = ~n15280 ;
  assign y6331 = n15286 ;
  assign y6332 = ~1'b0 ;
  assign y6333 = ~n15287 ;
  assign y6334 = n15290 ;
  assign y6335 = n15292 ;
  assign y6336 = ~n15296 ;
  assign y6337 = ~n15298 ;
  assign y6338 = n15301 ;
  assign y6339 = n15306 ;
  assign y6340 = ~1'b0 ;
  assign y6341 = n15307 ;
  assign y6342 = ~1'b0 ;
  assign y6343 = ~n15309 ;
  assign y6344 = ~1'b0 ;
  assign y6345 = ~n15310 ;
  assign y6346 = ~n15314 ;
  assign y6347 = ~1'b0 ;
  assign y6348 = ~1'b0 ;
  assign y6349 = ~n15319 ;
  assign y6350 = ~n15321 ;
  assign y6351 = ~1'b0 ;
  assign y6352 = ~n15324 ;
  assign y6353 = ~1'b0 ;
  assign y6354 = ~n15332 ;
  assign y6355 = ~n15333 ;
  assign y6356 = 1'b0 ;
  assign y6357 = ~1'b0 ;
  assign y6358 = n15338 ;
  assign y6359 = n15339 ;
  assign y6360 = ~1'b0 ;
  assign y6361 = ~n15343 ;
  assign y6362 = n15345 ;
  assign y6363 = ~n15348 ;
  assign y6364 = ~n15353 ;
  assign y6365 = ~n15363 ;
  assign y6366 = n15365 ;
  assign y6367 = n15368 ;
  assign y6368 = ~n15376 ;
  assign y6369 = ~n15379 ;
  assign y6370 = n15381 ;
  assign y6371 = ~1'b0 ;
  assign y6372 = n15385 ;
  assign y6373 = n15388 ;
  assign y6374 = n15389 ;
  assign y6375 = n15390 ;
  assign y6376 = ~1'b0 ;
  assign y6377 = ~1'b0 ;
  assign y6378 = ~n15394 ;
  assign y6379 = n15400 ;
  assign y6380 = ~n15401 ;
  assign y6381 = n15404 ;
  assign y6382 = ~n15408 ;
  assign y6383 = ~n15409 ;
  assign y6384 = n15411 ;
  assign y6385 = ~1'b0 ;
  assign y6386 = ~n15412 ;
  assign y6387 = ~n15416 ;
  assign y6388 = ~1'b0 ;
  assign y6389 = ~1'b0 ;
  assign y6390 = ~n15420 ;
  assign y6391 = ~n15421 ;
  assign y6392 = ~1'b0 ;
  assign y6393 = n15422 ;
  assign y6394 = n15427 ;
  assign y6395 = ~1'b0 ;
  assign y6396 = n15430 ;
  assign y6397 = ~n15432 ;
  assign y6398 = ~1'b0 ;
  assign y6399 = ~1'b0 ;
  assign y6400 = ~n15433 ;
  assign y6401 = n15436 ;
  assign y6402 = ~1'b0 ;
  assign y6403 = ~1'b0 ;
  assign y6404 = n15437 ;
  assign y6405 = ~n15438 ;
  assign y6406 = n15441 ;
  assign y6407 = ~n15442 ;
  assign y6408 = ~1'b0 ;
  assign y6409 = ~1'b0 ;
  assign y6410 = ~1'b0 ;
  assign y6411 = ~1'b0 ;
  assign y6412 = n15447 ;
  assign y6413 = ~n15449 ;
  assign y6414 = ~n15451 ;
  assign y6415 = ~n15452 ;
  assign y6416 = n15453 ;
  assign y6417 = ~n15454 ;
  assign y6418 = ~1'b0 ;
  assign y6419 = ~n15456 ;
  assign y6420 = ~n9170 ;
  assign y6421 = n15458 ;
  assign y6422 = ~n15459 ;
  assign y6423 = 1'b0 ;
  assign y6424 = ~1'b0 ;
  assign y6425 = ~n15460 ;
  assign y6426 = ~n15464 ;
  assign y6427 = ~1'b0 ;
  assign y6428 = ~n15468 ;
  assign y6429 = n15469 ;
  assign y6430 = ~n11878 ;
  assign y6431 = ~n15474 ;
  assign y6432 = ~n15485 ;
  assign y6433 = n15491 ;
  assign y6434 = n15493 ;
  assign y6435 = ~n15494 ;
  assign y6436 = ~n15495 ;
  assign y6437 = ~1'b0 ;
  assign y6438 = ~n15496 ;
  assign y6439 = n15497 ;
  assign y6440 = ~n15498 ;
  assign y6441 = ~n15507 ;
  assign y6442 = ~1'b0 ;
  assign y6443 = n15509 ;
  assign y6444 = ~n15511 ;
  assign y6445 = n15527 ;
  assign y6446 = ~1'b0 ;
  assign y6447 = ~n15529 ;
  assign y6448 = ~n15530 ;
  assign y6449 = n15532 ;
  assign y6450 = n15534 ;
  assign y6451 = n15538 ;
  assign y6452 = ~n15541 ;
  assign y6453 = n15542 ;
  assign y6454 = 1'b0 ;
  assign y6455 = ~n15544 ;
  assign y6456 = ~1'b0 ;
  assign y6457 = ~1'b0 ;
  assign y6458 = ~n15552 ;
  assign y6459 = n15554 ;
  assign y6460 = n15555 ;
  assign y6461 = ~n15560 ;
  assign y6462 = ~1'b0 ;
  assign y6463 = n15562 ;
  assign y6464 = ~n15564 ;
  assign y6465 = ~1'b0 ;
  assign y6466 = ~n15566 ;
  assign y6467 = ~n15567 ;
  assign y6468 = n15574 ;
  assign y6469 = n15577 ;
  assign y6470 = n13122 ;
  assign y6471 = n15578 ;
  assign y6472 = n15584 ;
  assign y6473 = ~n15586 ;
  assign y6474 = ~1'b0 ;
  assign y6475 = ~1'b0 ;
  assign y6476 = n15588 ;
  assign y6477 = n15589 ;
  assign y6478 = n15594 ;
  assign y6479 = ~1'b0 ;
  assign y6480 = ~n15605 ;
  assign y6481 = ~1'b0 ;
  assign y6482 = ~n15608 ;
  assign y6483 = ~n15609 ;
  assign y6484 = ~n15614 ;
  assign y6485 = n15620 ;
  assign y6486 = n15623 ;
  assign y6487 = 1'b0 ;
  assign y6488 = ~1'b0 ;
  assign y6489 = n8645 ;
  assign y6490 = ~n15624 ;
  assign y6491 = n15625 ;
  assign y6492 = ~1'b0 ;
  assign y6493 = ~1'b0 ;
  assign y6494 = n15627 ;
  assign y6495 = n15631 ;
  assign y6496 = n15632 ;
  assign y6497 = ~n15634 ;
  assign y6498 = n15636 ;
  assign y6499 = ~n15640 ;
  assign y6500 = ~1'b0 ;
  assign y6501 = ~1'b0 ;
  assign y6502 = n15645 ;
  assign y6503 = ~n15650 ;
  assign y6504 = ~n15655 ;
  assign y6505 = n15657 ;
  assign y6506 = n15659 ;
  assign y6507 = ~n15661 ;
  assign y6508 = ~1'b0 ;
  assign y6509 = ~x94 ;
  assign y6510 = ~n15663 ;
  assign y6511 = ~n15669 ;
  assign y6512 = n15671 ;
  assign y6513 = ~n8146 ;
  assign y6514 = ~1'b0 ;
  assign y6515 = n15672 ;
  assign y6516 = n12918 ;
  assign y6517 = ~1'b0 ;
  assign y6518 = n15676 ;
  assign y6519 = ~n15677 ;
  assign y6520 = n15682 ;
  assign y6521 = ~1'b0 ;
  assign y6522 = n15683 ;
  assign y6523 = ~n15688 ;
  assign y6524 = ~1'b0 ;
  assign y6525 = ~1'b0 ;
  assign y6526 = n15689 ;
  assign y6527 = ~1'b0 ;
  assign y6528 = ~1'b0 ;
  assign y6529 = ~n15692 ;
  assign y6530 = ~n15695 ;
  assign y6531 = ~n15699 ;
  assign y6532 = ~n15704 ;
  assign y6533 = ~n15706 ;
  assign y6534 = ~n15707 ;
  assign y6535 = ~n15708 ;
  assign y6536 = ~n15726 ;
  assign y6537 = n15728 ;
  assign y6538 = n15729 ;
  assign y6539 = ~n3737 ;
  assign y6540 = ~1'b0 ;
  assign y6541 = n15730 ;
  assign y6542 = ~1'b0 ;
  assign y6543 = n15733 ;
  assign y6544 = ~n15736 ;
  assign y6545 = n15741 ;
  assign y6546 = n15743 ;
  assign y6547 = n15744 ;
  assign y6548 = ~n15746 ;
  assign y6549 = ~1'b0 ;
  assign y6550 = n15750 ;
  assign y6551 = ~1'b0 ;
  assign y6552 = ~n15751 ;
  assign y6553 = ~n15754 ;
  assign y6554 = ~1'b0 ;
  assign y6555 = n15755 ;
  assign y6556 = n15757 ;
  assign y6557 = ~1'b0 ;
  assign y6558 = ~1'b0 ;
  assign y6559 = ~1'b0 ;
  assign y6560 = n10127 ;
  assign y6561 = n8029 ;
  assign y6562 = n15760 ;
  assign y6563 = n15761 ;
  assign y6564 = n15762 ;
  assign y6565 = ~n15765 ;
  assign y6566 = n15767 ;
  assign y6567 = ~n15768 ;
  assign y6568 = n15772 ;
  assign y6569 = ~n15774 ;
  assign y6570 = ~n15778 ;
  assign y6571 = n15781 ;
  assign y6572 = ~n15787 ;
  assign y6573 = ~n15791 ;
  assign y6574 = ~n15792 ;
  assign y6575 = n15795 ;
  assign y6576 = ~n3147 ;
  assign y6577 = ~n15799 ;
  assign y6578 = ~n15800 ;
  assign y6579 = n15802 ;
  assign y6580 = n15803 ;
  assign y6581 = ~1'b0 ;
  assign y6582 = ~1'b0 ;
  assign y6583 = ~1'b0 ;
  assign y6584 = n15805 ;
  assign y6585 = ~1'b0 ;
  assign y6586 = n15811 ;
  assign y6587 = ~n15815 ;
  assign y6588 = ~n15816 ;
  assign y6589 = ~1'b0 ;
  assign y6590 = n15828 ;
  assign y6591 = ~n15829 ;
  assign y6592 = ~1'b0 ;
  assign y6593 = ~1'b0 ;
  assign y6594 = n15831 ;
  assign y6595 = ~1'b0 ;
  assign y6596 = ~n15833 ;
  assign y6597 = ~1'b0 ;
  assign y6598 = n10569 ;
  assign y6599 = ~1'b0 ;
  assign y6600 = n15838 ;
  assign y6601 = ~1'b0 ;
  assign y6602 = n15840 ;
  assign y6603 = ~1'b0 ;
  assign y6604 = n15841 ;
  assign y6605 = n15842 ;
  assign y6606 = ~1'b0 ;
  assign y6607 = ~n15845 ;
  assign y6608 = n15849 ;
  assign y6609 = ~1'b0 ;
  assign y6610 = n15852 ;
  assign y6611 = n15859 ;
  assign y6612 = n15861 ;
  assign y6613 = n15862 ;
  assign y6614 = ~n15865 ;
  assign y6615 = n15870 ;
  assign y6616 = n15871 ;
  assign y6617 = n15874 ;
  assign y6618 = n15878 ;
  assign y6619 = n15880 ;
  assign y6620 = ~n15887 ;
  assign y6621 = ~n15898 ;
  assign y6622 = ~1'b0 ;
  assign y6623 = ~1'b0 ;
  assign y6624 = ~n15901 ;
  assign y6625 = ~1'b0 ;
  assign y6626 = ~1'b0 ;
  assign y6627 = ~n15904 ;
  assign y6628 = n13829 ;
  assign y6629 = ~1'b0 ;
  assign y6630 = ~n15905 ;
  assign y6631 = n15910 ;
  assign y6632 = ~n15912 ;
  assign y6633 = ~n15913 ;
  assign y6634 = n15917 ;
  assign y6635 = ~n15919 ;
  assign y6636 = n15927 ;
  assign y6637 = ~1'b0 ;
  assign y6638 = ~n15928 ;
  assign y6639 = ~n15932 ;
  assign y6640 = n15935 ;
  assign y6641 = ~1'b0 ;
  assign y6642 = ~1'b0 ;
  assign y6643 = ~1'b0 ;
  assign y6644 = ~n15944 ;
  assign y6645 = n15945 ;
  assign y6646 = ~n15946 ;
  assign y6647 = ~n15947 ;
  assign y6648 = ~n15952 ;
  assign y6649 = ~1'b0 ;
  assign y6650 = n15953 ;
  assign y6651 = ~1'b0 ;
  assign y6652 = n15957 ;
  assign y6653 = n15962 ;
  assign y6654 = 1'b0 ;
  assign y6655 = n15973 ;
  assign y6656 = n15976 ;
  assign y6657 = ~n15979 ;
  assign y6658 = ~n15980 ;
  assign y6659 = ~1'b0 ;
  assign y6660 = ~n12601 ;
  assign y6661 = n15984 ;
  assign y6662 = n15985 ;
  assign y6663 = n15991 ;
  assign y6664 = ~n15993 ;
  assign y6665 = n16001 ;
  assign y6666 = n16006 ;
  assign y6667 = n16008 ;
  assign y6668 = ~n4895 ;
  assign y6669 = ~1'b0 ;
  assign y6670 = ~n16009 ;
  assign y6671 = n16010 ;
  assign y6672 = ~n16015 ;
  assign y6673 = ~1'b0 ;
  assign y6674 = ~n16016 ;
  assign y6675 = ~n16021 ;
  assign y6676 = ~1'b0 ;
  assign y6677 = ~n16022 ;
  assign y6678 = n16023 ;
  assign y6679 = ~n16026 ;
  assign y6680 = n16037 ;
  assign y6681 = n16039 ;
  assign y6682 = ~n16040 ;
  assign y6683 = ~n16041 ;
  assign y6684 = ~n4045 ;
  assign y6685 = ~n16042 ;
  assign y6686 = ~n16043 ;
  assign y6687 = ~n16046 ;
  assign y6688 = n16049 ;
  assign y6689 = n16051 ;
  assign y6690 = ~n16055 ;
  assign y6691 = ~n9835 ;
  assign y6692 = ~n16062 ;
  assign y6693 = n16064 ;
  assign y6694 = n16066 ;
  assign y6695 = n16068 ;
  assign y6696 = ~n16080 ;
  assign y6697 = ~1'b0 ;
  assign y6698 = ~n16083 ;
  assign y6699 = ~n16095 ;
  assign y6700 = ~1'b0 ;
  assign y6701 = n16097 ;
  assign y6702 = n16099 ;
  assign y6703 = ~1'b0 ;
  assign y6704 = ~1'b0 ;
  assign y6705 = n16104 ;
  assign y6706 = n16105 ;
  assign y6707 = n16107 ;
  assign y6708 = ~1'b0 ;
  assign y6709 = n16111 ;
  assign y6710 = n16112 ;
  assign y6711 = n16113 ;
  assign y6712 = 1'b0 ;
  assign y6713 = ~1'b0 ;
  assign y6714 = ~n16115 ;
  assign y6715 = ~1'b0 ;
  assign y6716 = ~n16116 ;
  assign y6717 = n16131 ;
  assign y6718 = n16134 ;
  assign y6719 = n16136 ;
  assign y6720 = n16137 ;
  assign y6721 = n16144 ;
  assign y6722 = ~n16146 ;
  assign y6723 = ~n16151 ;
  assign y6724 = n16153 ;
  assign y6725 = ~1'b0 ;
  assign y6726 = n16156 ;
  assign y6727 = n16157 ;
  assign y6728 = ~n16161 ;
  assign y6729 = ~n16163 ;
  assign y6730 = ~1'b0 ;
  assign y6731 = n16165 ;
  assign y6732 = ~1'b0 ;
  assign y6733 = 1'b0 ;
  assign y6734 = ~1'b0 ;
  assign y6735 = n16169 ;
  assign y6736 = ~1'b0 ;
  assign y6737 = n16172 ;
  assign y6738 = n3659 ;
  assign y6739 = ~n16173 ;
  assign y6740 = ~n16174 ;
  assign y6741 = ~n16177 ;
  assign y6742 = ~n16181 ;
  assign y6743 = ~n16183 ;
  assign y6744 = ~1'b0 ;
  assign y6745 = n16187 ;
  assign y6746 = ~1'b0 ;
  assign y6747 = ~1'b0 ;
  assign y6748 = ~1'b0 ;
  assign y6749 = ~n16188 ;
  assign y6750 = n16190 ;
  assign y6751 = ~n16201 ;
  assign y6752 = ~n16215 ;
  assign y6753 = n16218 ;
  assign y6754 = ~1'b0 ;
  assign y6755 = ~n16220 ;
  assign y6756 = n16222 ;
  assign y6757 = ~1'b0 ;
  assign y6758 = ~n16223 ;
  assign y6759 = n16225 ;
  assign y6760 = ~1'b0 ;
  assign y6761 = ~1'b0 ;
  assign y6762 = ~n16226 ;
  assign y6763 = ~n16227 ;
  assign y6764 = n16228 ;
  assign y6765 = ~n16229 ;
  assign y6766 = ~1'b0 ;
  assign y6767 = ~1'b0 ;
  assign y6768 = n16230 ;
  assign y6769 = ~n16231 ;
  assign y6770 = n16234 ;
  assign y6771 = n16240 ;
  assign y6772 = n16242 ;
  assign y6773 = n16244 ;
  assign y6774 = ~n11524 ;
  assign y6775 = ~1'b0 ;
  assign y6776 = ~n16251 ;
  assign y6777 = n16252 ;
  assign y6778 = ~n16255 ;
  assign y6779 = n16265 ;
  assign y6780 = ~n16266 ;
  assign y6781 = ~n16271 ;
  assign y6782 = n16276 ;
  assign y6783 = ~n16278 ;
  assign y6784 = ~1'b0 ;
  assign y6785 = n16280 ;
  assign y6786 = n16290 ;
  assign y6787 = ~n16294 ;
  assign y6788 = ~n16297 ;
  assign y6789 = n16298 ;
  assign y6790 = ~1'b0 ;
  assign y6791 = n16301 ;
  assign y6792 = ~1'b0 ;
  assign y6793 = ~n14341 ;
  assign y6794 = n16302 ;
  assign y6795 = ~n16303 ;
  assign y6796 = n16309 ;
  assign y6797 = 1'b0 ;
  assign y6798 = ~n16311 ;
  assign y6799 = ~1'b0 ;
  assign y6800 = ~1'b0 ;
  assign y6801 = ~1'b0 ;
  assign y6802 = ~n16313 ;
  assign y6803 = ~n3313 ;
  assign y6804 = ~n16314 ;
  assign y6805 = n16315 ;
  assign y6806 = n16318 ;
  assign y6807 = n418 ;
  assign y6808 = ~n16320 ;
  assign y6809 = ~n16322 ;
  assign y6810 = ~n16324 ;
  assign y6811 = ~1'b0 ;
  assign y6812 = ~n16331 ;
  assign y6813 = ~1'b0 ;
  assign y6814 = n16337 ;
  assign y6815 = ~n16339 ;
  assign y6816 = ~n16341 ;
  assign y6817 = n16344 ;
  assign y6818 = n16346 ;
  assign y6819 = ~n16349 ;
  assign y6820 = ~n16356 ;
  assign y6821 = n16357 ;
  assign y6822 = ~1'b0 ;
  assign y6823 = ~n9421 ;
  assign y6824 = ~1'b0 ;
  assign y6825 = ~n16361 ;
  assign y6826 = ~1'b0 ;
  assign y6827 = ~1'b0 ;
  assign y6828 = ~n16363 ;
  assign y6829 = ~n16365 ;
  assign y6830 = ~1'b0 ;
  assign y6831 = n16366 ;
  assign y6832 = ~1'b0 ;
  assign y6833 = ~1'b0 ;
  assign y6834 = ~n16367 ;
  assign y6835 = ~n16370 ;
  assign y6836 = n16375 ;
  assign y6837 = n16378 ;
  assign y6838 = ~n16382 ;
  assign y6839 = ~n16387 ;
  assign y6840 = ~1'b0 ;
  assign y6841 = n16389 ;
  assign y6842 = 1'b0 ;
  assign y6843 = n16392 ;
  assign y6844 = n16394 ;
  assign y6845 = ~1'b0 ;
  assign y6846 = n16395 ;
  assign y6847 = ~n16408 ;
  assign y6848 = n16411 ;
  assign y6849 = n16420 ;
  assign y6850 = n16422 ;
  assign y6851 = n16424 ;
  assign y6852 = n16427 ;
  assign y6853 = n16431 ;
  assign y6854 = ~1'b0 ;
  assign y6855 = n4215 ;
  assign y6856 = ~1'b0 ;
  assign y6857 = n16432 ;
  assign y6858 = 1'b0 ;
  assign y6859 = ~n16433 ;
  assign y6860 = n16435 ;
  assign y6861 = ~1'b0 ;
  assign y6862 = ~n16437 ;
  assign y6863 = ~1'b0 ;
  assign y6864 = ~1'b0 ;
  assign y6865 = ~n16438 ;
  assign y6866 = ~1'b0 ;
  assign y6867 = ~1'b0 ;
  assign y6868 = ~n16440 ;
  assign y6869 = n16443 ;
  assign y6870 = ~n16446 ;
  assign y6871 = ~1'b0 ;
  assign y6872 = ~n16448 ;
  assign y6873 = ~n16449 ;
  assign y6874 = ~n16451 ;
  assign y6875 = n16455 ;
  assign y6876 = ~n16459 ;
  assign y6877 = n16460 ;
  assign y6878 = n16462 ;
  assign y6879 = ~1'b0 ;
  assign y6880 = ~n16467 ;
  assign y6881 = ~n16470 ;
  assign y6882 = n16476 ;
  assign y6883 = n16479 ;
  assign y6884 = ~n16481 ;
  assign y6885 = ~n16484 ;
  assign y6886 = ~n16486 ;
  assign y6887 = n16488 ;
  assign y6888 = ~1'b0 ;
  assign y6889 = ~1'b0 ;
  assign y6890 = ~n16490 ;
  assign y6891 = ~1'b0 ;
  assign y6892 = n16493 ;
  assign y6893 = ~1'b0 ;
  assign y6894 = ~n16498 ;
  assign y6895 = ~n16499 ;
  assign y6896 = ~n16501 ;
  assign y6897 = ~n16502 ;
  assign y6898 = ~n16506 ;
  assign y6899 = ~n16507 ;
  assign y6900 = n16509 ;
  assign y6901 = n16510 ;
  assign y6902 = n16511 ;
  assign y6903 = n16516 ;
  assign y6904 = n16525 ;
  assign y6905 = n14112 ;
  assign y6906 = n16527 ;
  assign y6907 = 1'b0 ;
  assign y6908 = ~n16528 ;
  assign y6909 = ~n16530 ;
  assign y6910 = ~1'b0 ;
  assign y6911 = ~n16542 ;
  assign y6912 = ~1'b0 ;
  assign y6913 = n327 ;
  assign y6914 = ~n1264 ;
  assign y6915 = ~1'b0 ;
  assign y6916 = ~n16545 ;
  assign y6917 = n16547 ;
  assign y6918 = n16549 ;
  assign y6919 = n16552 ;
  assign y6920 = n16553 ;
  assign y6921 = ~n16560 ;
  assign y6922 = n16561 ;
  assign y6923 = ~n16566 ;
  assign y6924 = n16572 ;
  assign y6925 = ~1'b0 ;
  assign y6926 = n10396 ;
  assign y6927 = ~n16575 ;
  assign y6928 = ~n16576 ;
  assign y6929 = ~1'b0 ;
  assign y6930 = ~1'b0 ;
  assign y6931 = ~1'b0 ;
  assign y6932 = ~n16577 ;
  assign y6933 = ~n16579 ;
  assign y6934 = ~n16580 ;
  assign y6935 = n16581 ;
  assign y6936 = n16584 ;
  assign y6937 = ~1'b0 ;
  assign y6938 = ~n16585 ;
  assign y6939 = ~n16589 ;
  assign y6940 = ~1'b0 ;
  assign y6941 = ~n16591 ;
  assign y6942 = n16598 ;
  assign y6943 = ~1'b0 ;
  assign y6944 = ~n16606 ;
  assign y6945 = ~1'b0 ;
  assign y6946 = n7590 ;
  assign y6947 = ~1'b0 ;
  assign y6948 = ~1'b0 ;
  assign y6949 = ~1'b0 ;
  assign y6950 = ~1'b0 ;
  assign y6951 = ~n16607 ;
  assign y6952 = 1'b0 ;
  assign y6953 = n16612 ;
  assign y6954 = ~n16614 ;
  assign y6955 = ~1'b0 ;
  assign y6956 = n16616 ;
  assign y6957 = n16622 ;
  assign y6958 = ~n16630 ;
  assign y6959 = ~n16631 ;
  assign y6960 = n16638 ;
  assign y6961 = n16641 ;
  assign y6962 = 1'b0 ;
  assign y6963 = ~n16642 ;
  assign y6964 = ~n16644 ;
  assign y6965 = ~1'b0 ;
  assign y6966 = ~n16646 ;
  assign y6967 = n16648 ;
  assign y6968 = ~n16654 ;
  assign y6969 = n16657 ;
  assign y6970 = ~n16662 ;
  assign y6971 = n16669 ;
  assign y6972 = ~n16680 ;
  assign y6973 = ~1'b0 ;
  assign y6974 = ~n16681 ;
  assign y6975 = n16682 ;
  assign y6976 = ~n16686 ;
  assign y6977 = ~n16687 ;
  assign y6978 = ~1'b0 ;
  assign y6979 = ~1'b0 ;
  assign y6980 = ~1'b0 ;
  assign y6981 = n16690 ;
  assign y6982 = n16693 ;
  assign y6983 = 1'b0 ;
  assign y6984 = ~n16694 ;
  assign y6985 = ~1'b0 ;
  assign y6986 = n16695 ;
  assign y6987 = ~n16697 ;
  assign y6988 = n16698 ;
  assign y6989 = ~n16700 ;
  assign y6990 = ~n16701 ;
  assign y6991 = ~1'b0 ;
  assign y6992 = ~n16703 ;
  assign y6993 = ~1'b0 ;
  assign y6994 = ~n16708 ;
  assign y6995 = ~n16709 ;
  assign y6996 = ~n16710 ;
  assign y6997 = ~n16713 ;
  assign y6998 = n16714 ;
  assign y6999 = n16715 ;
  assign y7000 = ~1'b0 ;
  assign y7001 = ~n16722 ;
  assign y7002 = ~n16727 ;
  assign y7003 = ~1'b0 ;
  assign y7004 = ~1'b0 ;
  assign y7005 = n16730 ;
  assign y7006 = n12907 ;
  assign y7007 = ~1'b0 ;
  assign y7008 = ~n16731 ;
  assign y7009 = n16732 ;
  assign y7010 = n16734 ;
  assign y7011 = ~1'b0 ;
  assign y7012 = n16736 ;
  assign y7013 = n16737 ;
  assign y7014 = n16739 ;
  assign y7015 = n13230 ;
  assign y7016 = ~1'b0 ;
  assign y7017 = n16741 ;
  assign y7018 = ~1'b0 ;
  assign y7019 = n6361 ;
  assign y7020 = n16743 ;
  assign y7021 = ~n16745 ;
  assign y7022 = n16747 ;
  assign y7023 = n16751 ;
  assign y7024 = n16752 ;
  assign y7025 = n16760 ;
  assign y7026 = ~1'b0 ;
  assign y7027 = ~1'b0 ;
  assign y7028 = n14662 ;
  assign y7029 = ~n16763 ;
  assign y7030 = n16764 ;
  assign y7031 = n16765 ;
  assign y7032 = ~1'b0 ;
  assign y7033 = n16766 ;
  assign y7034 = n16770 ;
  assign y7035 = ~1'b0 ;
  assign y7036 = ~n16773 ;
  assign y7037 = ~n16775 ;
  assign y7038 = n16777 ;
  assign y7039 = n16784 ;
  assign y7040 = ~n16785 ;
  assign y7041 = n16794 ;
  assign y7042 = ~n16805 ;
  assign y7043 = ~1'b0 ;
  assign y7044 = ~n16809 ;
  assign y7045 = n10950 ;
  assign y7046 = n16814 ;
  assign y7047 = ~n16818 ;
  assign y7048 = ~n16824 ;
  assign y7049 = ~1'b0 ;
  assign y7050 = ~n16826 ;
  assign y7051 = ~n16829 ;
  assign y7052 = n16833 ;
  assign y7053 = ~1'b0 ;
  assign y7054 = ~1'b0 ;
  assign y7055 = ~n16838 ;
  assign y7056 = n16839 ;
  assign y7057 = ~n16846 ;
  assign y7058 = ~1'b0 ;
  assign y7059 = ~1'b0 ;
  assign y7060 = ~n16847 ;
  assign y7061 = n16851 ;
  assign y7062 = n16855 ;
  assign y7063 = ~1'b0 ;
  assign y7064 = ~n16857 ;
  assign y7065 = n9356 ;
  assign y7066 = n16858 ;
  assign y7067 = n16864 ;
  assign y7068 = n4286 ;
  assign y7069 = ~n16867 ;
  assign y7070 = ~n16870 ;
  assign y7071 = ~n16871 ;
  assign y7072 = ~n16872 ;
  assign y7073 = n16878 ;
  assign y7074 = ~n16880 ;
  assign y7075 = n16887 ;
  assign y7076 = ~n16891 ;
  assign y7077 = ~n16896 ;
  assign y7078 = ~1'b0 ;
  assign y7079 = ~n16899 ;
  assign y7080 = n16901 ;
  assign y7081 = n16904 ;
  assign y7082 = n16907 ;
  assign y7083 = ~n16912 ;
  assign y7084 = ~n16913 ;
  assign y7085 = n16916 ;
  assign y7086 = ~n16917 ;
  assign y7087 = ~1'b0 ;
  assign y7088 = n16919 ;
  assign y7089 = n681 ;
  assign y7090 = n16920 ;
  assign y7091 = ~1'b0 ;
  assign y7092 = ~1'b0 ;
  assign y7093 = ~1'b0 ;
  assign y7094 = n16923 ;
  assign y7095 = ~n16924 ;
  assign y7096 = n16925 ;
  assign y7097 = n8531 ;
  assign y7098 = n16928 ;
  assign y7099 = n16929 ;
  assign y7100 = n16932 ;
  assign y7101 = ~n16934 ;
  assign y7102 = 1'b0 ;
  assign y7103 = n16935 ;
  assign y7104 = n16936 ;
  assign y7105 = n16937 ;
  assign y7106 = ~n16943 ;
  assign y7107 = ~1'b0 ;
  assign y7108 = ~n16944 ;
  assign y7109 = ~1'b0 ;
  assign y7110 = n16946 ;
  assign y7111 = ~n16947 ;
  assign y7112 = ~n16950 ;
  assign y7113 = n16953 ;
  assign y7114 = ~n16955 ;
  assign y7115 = ~1'b0 ;
  assign y7116 = n16957 ;
  assign y7117 = n6458 ;
  assign y7118 = ~1'b0 ;
  assign y7119 = ~n16959 ;
  assign y7120 = ~1'b0 ;
  assign y7121 = ~1'b0 ;
  assign y7122 = ~n16964 ;
  assign y7123 = ~n16965 ;
  assign y7124 = n16966 ;
  assign y7125 = ~n16974 ;
  assign y7126 = ~n16975 ;
  assign y7127 = n16980 ;
  assign y7128 = n16987 ;
  assign y7129 = ~1'b0 ;
  assign y7130 = ~n16989 ;
  assign y7131 = ~1'b0 ;
  assign y7132 = ~n16998 ;
  assign y7133 = n16999 ;
  assign y7134 = ~n17000 ;
  assign y7135 = ~1'b0 ;
  assign y7136 = n17001 ;
  assign y7137 = ~n17005 ;
  assign y7138 = n17006 ;
  assign y7139 = ~n17008 ;
  assign y7140 = ~n17013 ;
  assign y7141 = ~n17015 ;
  assign y7142 = n17016 ;
  assign y7143 = ~n17020 ;
  assign y7144 = ~1'b0 ;
  assign y7145 = ~n17021 ;
  assign y7146 = n17022 ;
  assign y7147 = ~1'b0 ;
  assign y7148 = ~1'b0 ;
  assign y7149 = ~n17023 ;
  assign y7150 = n17025 ;
  assign y7151 = ~n17031 ;
  assign y7152 = ~n17039 ;
  assign y7153 = ~1'b0 ;
  assign y7154 = ~n17040 ;
  assign y7155 = n17044 ;
  assign y7156 = ~1'b0 ;
  assign y7157 = ~1'b0 ;
  assign y7158 = ~1'b0 ;
  assign y7159 = ~n17045 ;
  assign y7160 = n17065 ;
  assign y7161 = ~n17068 ;
  assign y7162 = n17072 ;
  assign y7163 = n17073 ;
  assign y7164 = ~1'b0 ;
  assign y7165 = ~n17080 ;
  assign y7166 = ~n17081 ;
  assign y7167 = n17083 ;
  assign y7168 = n17089 ;
  assign y7169 = ~n17091 ;
  assign y7170 = n17107 ;
  assign y7171 = ~n17110 ;
  assign y7172 = ~1'b0 ;
  assign y7173 = ~1'b0 ;
  assign y7174 = n17112 ;
  assign y7175 = ~n17115 ;
  assign y7176 = ~n9356 ;
  assign y7177 = ~1'b0 ;
  assign y7178 = ~n7756 ;
  assign y7179 = ~n17117 ;
  assign y7180 = ~n17118 ;
  assign y7181 = ~n17132 ;
  assign y7182 = ~1'b0 ;
  assign y7183 = ~n17133 ;
  assign y7184 = ~n17135 ;
  assign y7185 = ~1'b0 ;
  assign y7186 = ~1'b0 ;
  assign y7187 = ~n17136 ;
  assign y7188 = ~n17137 ;
  assign y7189 = n17139 ;
  assign y7190 = ~1'b0 ;
  assign y7191 = n17144 ;
  assign y7192 = n17152 ;
  assign y7193 = n17153 ;
  assign y7194 = ~1'b0 ;
  assign y7195 = n17155 ;
  assign y7196 = ~1'b0 ;
  assign y7197 = n17156 ;
  assign y7198 = ~n17162 ;
  assign y7199 = n17166 ;
  assign y7200 = ~n17167 ;
  assign y7201 = ~n17168 ;
  assign y7202 = n17169 ;
  assign y7203 = n17175 ;
  assign y7204 = ~n17176 ;
  assign y7205 = ~n17178 ;
  assign y7206 = ~n17179 ;
  assign y7207 = n17181 ;
  assign y7208 = ~1'b0 ;
  assign y7209 = ~n17185 ;
  assign y7210 = ~n17186 ;
  assign y7211 = ~n17188 ;
  assign y7212 = ~1'b0 ;
  assign y7213 = n17190 ;
  assign y7214 = n17191 ;
  assign y7215 = ~n17196 ;
  assign y7216 = n17203 ;
  assign y7217 = ~n17206 ;
  assign y7218 = ~n17207 ;
  assign y7219 = 1'b0 ;
  assign y7220 = n17210 ;
  assign y7221 = n17211 ;
  assign y7222 = ~n17213 ;
  assign y7223 = n17214 ;
  assign y7224 = ~1'b0 ;
  assign y7225 = n17218 ;
  assign y7226 = ~1'b0 ;
  assign y7227 = ~n17221 ;
  assign y7228 = ~n17224 ;
  assign y7229 = ~n15985 ;
  assign y7230 = ~1'b0 ;
  assign y7231 = ~n17226 ;
  assign y7232 = ~n17228 ;
  assign y7233 = ~1'b0 ;
  assign y7234 = ~n17232 ;
  assign y7235 = ~1'b0 ;
  assign y7236 = ~1'b0 ;
  assign y7237 = ~n17237 ;
  assign y7238 = ~n17240 ;
  assign y7239 = ~n17242 ;
  assign y7240 = n17245 ;
  assign y7241 = n17252 ;
  assign y7242 = ~n3246 ;
  assign y7243 = n17254 ;
  assign y7244 = ~1'b0 ;
  assign y7245 = ~1'b0 ;
  assign y7246 = ~1'b0 ;
  assign y7247 = n17258 ;
  assign y7248 = ~n3318 ;
  assign y7249 = ~n17260 ;
  assign y7250 = ~n17261 ;
  assign y7251 = ~1'b0 ;
  assign y7252 = ~1'b0 ;
  assign y7253 = ~n17270 ;
  assign y7254 = ~1'b0 ;
  assign y7255 = ~1'b0 ;
  assign y7256 = ~1'b0 ;
  assign y7257 = ~n17272 ;
  assign y7258 = n17273 ;
  assign y7259 = n17275 ;
  assign y7260 = ~1'b0 ;
  assign y7261 = n17277 ;
  assign y7262 = ~n17279 ;
  assign y7263 = ~1'b0 ;
  assign y7264 = n17280 ;
  assign y7265 = ~n17287 ;
  assign y7266 = 1'b0 ;
  assign y7267 = n17298 ;
  assign y7268 = n17300 ;
  assign y7269 = ~1'b0 ;
  assign y7270 = ~n1500 ;
  assign y7271 = ~1'b0 ;
  assign y7272 = ~n17307 ;
  assign y7273 = n17311 ;
  assign y7274 = ~1'b0 ;
  assign y7275 = n17314 ;
  assign y7276 = n17316 ;
  assign y7277 = ~n17322 ;
  assign y7278 = ~1'b0 ;
  assign y7279 = n17324 ;
  assign y7280 = n17328 ;
  assign y7281 = n17333 ;
  assign y7282 = ~n3918 ;
  assign y7283 = ~1'b0 ;
  assign y7284 = ~n17337 ;
  assign y7285 = n17340 ;
  assign y7286 = n17342 ;
  assign y7287 = ~n17346 ;
  assign y7288 = ~n17348 ;
  assign y7289 = ~1'b0 ;
  assign y7290 = ~1'b0 ;
  assign y7291 = n17350 ;
  assign y7292 = n17353 ;
  assign y7293 = ~n8115 ;
  assign y7294 = ~n17354 ;
  assign y7295 = ~1'b0 ;
  assign y7296 = n17355 ;
  assign y7297 = ~n17357 ;
  assign y7298 = n17359 ;
  assign y7299 = ~1'b0 ;
  assign y7300 = ~1'b0 ;
  assign y7301 = ~n17362 ;
  assign y7302 = n17371 ;
  assign y7303 = n17373 ;
  assign y7304 = ~n17377 ;
  assign y7305 = ~n17381 ;
  assign y7306 = n17383 ;
  assign y7307 = ~1'b0 ;
  assign y7308 = ~n17385 ;
  assign y7309 = n17393 ;
  assign y7310 = ~n17403 ;
  assign y7311 = ~1'b0 ;
  assign y7312 = ~1'b0 ;
  assign y7313 = n17406 ;
  assign y7314 = ~1'b0 ;
  assign y7315 = n17409 ;
  assign y7316 = n17413 ;
  assign y7317 = ~n17414 ;
  assign y7318 = n17417 ;
  assign y7319 = n17418 ;
  assign y7320 = ~1'b0 ;
  assign y7321 = n17432 ;
  assign y7322 = 1'b0 ;
  assign y7323 = n17433 ;
  assign y7324 = n17439 ;
  assign y7325 = n17440 ;
  assign y7326 = n17443 ;
  assign y7327 = n17444 ;
  assign y7328 = ~1'b0 ;
  assign y7329 = ~n17445 ;
  assign y7330 = ~1'b0 ;
  assign y7331 = n17448 ;
  assign y7332 = ~n17453 ;
  assign y7333 = ~n17454 ;
  assign y7334 = n17456 ;
  assign y7335 = ~1'b0 ;
  assign y7336 = n627 ;
  assign y7337 = ~1'b0 ;
  assign y7338 = n17459 ;
  assign y7339 = ~n17464 ;
  assign y7340 = n17465 ;
  assign y7341 = n17469 ;
  assign y7342 = ~n17471 ;
  assign y7343 = ~n17473 ;
  assign y7344 = n17474 ;
  assign y7345 = n17479 ;
  assign y7346 = n17481 ;
  assign y7347 = n17489 ;
  assign y7348 = 1'b0 ;
  assign y7349 = 1'b0 ;
  assign y7350 = n17492 ;
  assign y7351 = ~n17493 ;
  assign y7352 = ~n17502 ;
  assign y7353 = ~n17507 ;
  assign y7354 = ~1'b0 ;
  assign y7355 = ~1'b0 ;
  assign y7356 = ~n17510 ;
  assign y7357 = ~n3016 ;
  assign y7358 = ~n17512 ;
  assign y7359 = ~1'b0 ;
  assign y7360 = ~1'b0 ;
  assign y7361 = n17515 ;
  assign y7362 = ~n17520 ;
  assign y7363 = ~1'b0 ;
  assign y7364 = ~1'b0 ;
  assign y7365 = ~1'b0 ;
  assign y7366 = ~n7871 ;
  assign y7367 = n17522 ;
  assign y7368 = ~1'b0 ;
  assign y7369 = ~n17525 ;
  assign y7370 = ~n17528 ;
  assign y7371 = n17530 ;
  assign y7372 = ~n17539 ;
  assign y7373 = ~1'b0 ;
  assign y7374 = n17540 ;
  assign y7375 = ~n17543 ;
  assign y7376 = ~n17546 ;
  assign y7377 = ~n17550 ;
  assign y7378 = n17555 ;
  assign y7379 = ~1'b0 ;
  assign y7380 = ~n17560 ;
  assign y7381 = ~n17561 ;
  assign y7382 = n17567 ;
  assign y7383 = n17568 ;
  assign y7384 = ~n17571 ;
  assign y7385 = n17576 ;
  assign y7386 = ~1'b0 ;
  assign y7387 = ~n1365 ;
  assign y7388 = ~n17578 ;
  assign y7389 = ~n17580 ;
  assign y7390 = ~n17584 ;
  assign y7391 = n17586 ;
  assign y7392 = n17590 ;
  assign y7393 = n17592 ;
  assign y7394 = ~1'b0 ;
  assign y7395 = ~1'b0 ;
  assign y7396 = ~n326 ;
  assign y7397 = ~n17593 ;
  assign y7398 = ~1'b0 ;
  assign y7399 = ~1'b0 ;
  assign y7400 = n17595 ;
  assign y7401 = ~n17596 ;
  assign y7402 = n17597 ;
  assign y7403 = ~n17601 ;
  assign y7404 = n17602 ;
  assign y7405 = ~n17605 ;
  assign y7406 = ~1'b0 ;
  assign y7407 = n17609 ;
  assign y7408 = ~n17616 ;
  assign y7409 = n17617 ;
  assign y7410 = n17619 ;
  assign y7411 = n17622 ;
  assign y7412 = ~n17624 ;
  assign y7413 = n17629 ;
  assign y7414 = n17635 ;
  assign y7415 = n17645 ;
  assign y7416 = n17646 ;
  assign y7417 = n17648 ;
  assign y7418 = n17653 ;
  assign y7419 = ~1'b0 ;
  assign y7420 = ~1'b0 ;
  assign y7421 = ~n17667 ;
  assign y7422 = n17672 ;
  assign y7423 = ~1'b0 ;
  assign y7424 = 1'b0 ;
  assign y7425 = n7324 ;
  assign y7426 = ~1'b0 ;
  assign y7427 = ~1'b0 ;
  assign y7428 = n17674 ;
  assign y7429 = ~n17676 ;
  assign y7430 = ~n17677 ;
  assign y7431 = ~n17680 ;
  assign y7432 = ~1'b0 ;
  assign y7433 = ~1'b0 ;
  assign y7434 = n17683 ;
  assign y7435 = n17685 ;
  assign y7436 = n17690 ;
  assign y7437 = ~1'b0 ;
  assign y7438 = ~1'b0 ;
  assign y7439 = ~1'b0 ;
  assign y7440 = ~1'b0 ;
  assign y7441 = n15604 ;
  assign y7442 = ~1'b0 ;
  assign y7443 = ~1'b0 ;
  assign y7444 = ~n17691 ;
  assign y7445 = n17695 ;
  assign y7446 = n17697 ;
  assign y7447 = ~n17700 ;
  assign y7448 = ~n17701 ;
  assign y7449 = n17702 ;
  assign y7450 = ~n17708 ;
  assign y7451 = ~1'b0 ;
  assign y7452 = ~n17712 ;
  assign y7453 = ~1'b0 ;
  assign y7454 = ~n17713 ;
  assign y7455 = ~1'b0 ;
  assign y7456 = n17714 ;
  assign y7457 = n17715 ;
  assign y7458 = ~n17719 ;
  assign y7459 = ~n8294 ;
  assign y7460 = ~n17723 ;
  assign y7461 = ~n17725 ;
  assign y7462 = n17727 ;
  assign y7463 = n17729 ;
  assign y7464 = ~1'b0 ;
  assign y7465 = n7204 ;
  assign y7466 = n17730 ;
  assign y7467 = ~1'b0 ;
  assign y7468 = ~n17737 ;
  assign y7469 = ~n17738 ;
  assign y7470 = n17742 ;
  assign y7471 = ~n17744 ;
  assign y7472 = n17749 ;
  assign y7473 = ~1'b0 ;
  assign y7474 = ~n17753 ;
  assign y7475 = ~1'b0 ;
  assign y7476 = ~n17755 ;
  assign y7477 = ~1'b0 ;
  assign y7478 = ~1'b0 ;
  assign y7479 = n17757 ;
  assign y7480 = ~n17760 ;
  assign y7481 = n17763 ;
  assign y7482 = ~1'b0 ;
  assign y7483 = n17768 ;
  assign y7484 = ~n17774 ;
  assign y7485 = n17778 ;
  assign y7486 = n16513 ;
  assign y7487 = ~n17783 ;
  assign y7488 = ~n17786 ;
  assign y7489 = ~n17791 ;
  assign y7490 = ~1'b0 ;
  assign y7491 = n17794 ;
  assign y7492 = ~1'b0 ;
  assign y7493 = n17802 ;
  assign y7494 = ~n17803 ;
  assign y7495 = ~n17804 ;
  assign y7496 = n17810 ;
  assign y7497 = n17812 ;
  assign y7498 = ~1'b0 ;
  assign y7499 = n17818 ;
  assign y7500 = ~n17825 ;
  assign y7501 = ~1'b0 ;
  assign y7502 = 1'b0 ;
  assign y7503 = n17828 ;
  assign y7504 = ~n17834 ;
  assign y7505 = n17835 ;
  assign y7506 = n17838 ;
  assign y7507 = ~n17839 ;
  assign y7508 = ~n17841 ;
  assign y7509 = ~n17843 ;
  assign y7510 = ~n17851 ;
  assign y7511 = ~1'b0 ;
  assign y7512 = n17853 ;
  assign y7513 = ~1'b0 ;
  assign y7514 = ~n17854 ;
  assign y7515 = n17855 ;
  assign y7516 = n17857 ;
  assign y7517 = ~1'b0 ;
  assign y7518 = ~1'b0 ;
  assign y7519 = ~n17864 ;
  assign y7520 = n17865 ;
  assign y7521 = ~n17874 ;
  assign y7522 = ~n17876 ;
  assign y7523 = n17878 ;
  assign y7524 = n17880 ;
  assign y7525 = n17882 ;
  assign y7526 = ~1'b0 ;
  assign y7527 = ~1'b0 ;
  assign y7528 = ~1'b0 ;
  assign y7529 = ~n17887 ;
  assign y7530 = n15276 ;
  assign y7531 = ~n17888 ;
  assign y7532 = n17891 ;
  assign y7533 = ~n17895 ;
  assign y7534 = n17896 ;
  assign y7535 = n17897 ;
  assign y7536 = ~n17899 ;
  assign y7537 = ~n17902 ;
  assign y7538 = ~n17909 ;
  assign y7539 = n17910 ;
  assign y7540 = n17912 ;
  assign y7541 = ~n17913 ;
  assign y7542 = n17914 ;
  assign y7543 = ~n3296 ;
  assign y7544 = n17916 ;
  assign y7545 = n17918 ;
  assign y7546 = ~1'b0 ;
  assign y7547 = n17921 ;
  assign y7548 = ~1'b0 ;
  assign y7549 = n15320 ;
  assign y7550 = n17923 ;
  assign y7551 = ~1'b0 ;
  assign y7552 = ~n17925 ;
  assign y7553 = ~1'b0 ;
  assign y7554 = n7567 ;
  assign y7555 = ~1'b0 ;
  assign y7556 = ~n17928 ;
  assign y7557 = ~n17929 ;
  assign y7558 = n17931 ;
  assign y7559 = ~n5314 ;
  assign y7560 = ~n17936 ;
  assign y7561 = n17939 ;
  assign y7562 = n8443 ;
  assign y7563 = ~n17941 ;
  assign y7564 = n13796 ;
  assign y7565 = ~1'b0 ;
  assign y7566 = 1'b0 ;
  assign y7567 = ~n17943 ;
  assign y7568 = 1'b0 ;
  assign y7569 = n3738 ;
  assign y7570 = ~1'b0 ;
  assign y7571 = ~n17945 ;
  assign y7572 = ~1'b0 ;
  assign y7573 = ~n17946 ;
  assign y7574 = ~n6174 ;
  assign y7575 = ~n17951 ;
  assign y7576 = n17956 ;
  assign y7577 = n17960 ;
  assign y7578 = n17964 ;
  assign y7579 = n17965 ;
  assign y7580 = ~n17967 ;
  assign y7581 = ~n17969 ;
  assign y7582 = n17973 ;
  assign y7583 = n17976 ;
  assign y7584 = n17983 ;
  assign y7585 = ~n17986 ;
  assign y7586 = n17991 ;
  assign y7587 = ~n17996 ;
  assign y7588 = ~1'b0 ;
  assign y7589 = n17998 ;
  assign y7590 = n8262 ;
  assign y7591 = ~n18000 ;
  assign y7592 = ~1'b0 ;
  assign y7593 = 1'b0 ;
  assign y7594 = ~1'b0 ;
  assign y7595 = n18007 ;
  assign y7596 = ~n18008 ;
  assign y7597 = ~n18011 ;
  assign y7598 = ~n18022 ;
  assign y7599 = n18027 ;
  assign y7600 = n18029 ;
  assign y7601 = ~n18031 ;
  assign y7602 = n18035 ;
  assign y7603 = n18039 ;
  assign y7604 = ~n18046 ;
  assign y7605 = ~1'b0 ;
  assign y7606 = ~1'b0 ;
  assign y7607 = 1'b0 ;
  assign y7608 = n18049 ;
  assign y7609 = ~n18051 ;
  assign y7610 = n18052 ;
  assign y7611 = n18054 ;
  assign y7612 = ~n18062 ;
  assign y7613 = ~n18068 ;
  assign y7614 = ~n18075 ;
  assign y7615 = ~n18078 ;
  assign y7616 = n18083 ;
  assign y7617 = n18090 ;
  assign y7618 = ~1'b0 ;
  assign y7619 = ~1'b0 ;
  assign y7620 = n18092 ;
  assign y7621 = n18095 ;
  assign y7622 = ~n18098 ;
  assign y7623 = ~n18099 ;
  assign y7624 = n5384 ;
  assign y7625 = ~n18100 ;
  assign y7626 = n18103 ;
  assign y7627 = n18105 ;
  assign y7628 = ~n18107 ;
  assign y7629 = ~1'b0 ;
  assign y7630 = ~1'b0 ;
  assign y7631 = ~n18108 ;
  assign y7632 = ~1'b0 ;
  assign y7633 = ~n18109 ;
  assign y7634 = ~n18110 ;
  assign y7635 = ~1'b0 ;
  assign y7636 = ~1'b0 ;
  assign y7637 = ~n18113 ;
  assign y7638 = ~n18115 ;
  assign y7639 = ~n18118 ;
  assign y7640 = n1488 ;
  assign y7641 = ~1'b0 ;
  assign y7642 = ~1'b0 ;
  assign y7643 = ~n18120 ;
  assign y7644 = n18122 ;
  assign y7645 = n1166 ;
  assign y7646 = ~n10879 ;
  assign y7647 = n18124 ;
  assign y7648 = ~n4134 ;
  assign y7649 = ~n8194 ;
  assign y7650 = ~n18125 ;
  assign y7651 = ~n18126 ;
  assign y7652 = n9949 ;
  assign y7653 = ~n18127 ;
  assign y7654 = ~1'b0 ;
  assign y7655 = ~n18129 ;
  assign y7656 = n18130 ;
  assign y7657 = n9513 ;
  assign y7658 = n18136 ;
  assign y7659 = n18139 ;
  assign y7660 = n18140 ;
  assign y7661 = n18147 ;
  assign y7662 = ~1'b0 ;
  assign y7663 = ~1'b0 ;
  assign y7664 = ~n18149 ;
  assign y7665 = ~1'b0 ;
  assign y7666 = ~n18155 ;
  assign y7667 = ~n18156 ;
  assign y7668 = ~n18166 ;
  assign y7669 = n18168 ;
  assign y7670 = n18175 ;
  assign y7671 = n2428 ;
  assign y7672 = ~n18179 ;
  assign y7673 = n18181 ;
  assign y7674 = n18183 ;
  assign y7675 = ~n18184 ;
  assign y7676 = 1'b0 ;
  assign y7677 = ~n18185 ;
  assign y7678 = n18194 ;
  assign y7679 = n18197 ;
  assign y7680 = ~n18201 ;
  assign y7681 = n18208 ;
  assign y7682 = n18211 ;
  assign y7683 = ~n18214 ;
  assign y7684 = ~n18220 ;
  assign y7685 = ~1'b0 ;
  assign y7686 = ~n5922 ;
  assign y7687 = ~n18224 ;
  assign y7688 = n18227 ;
  assign y7689 = n18229 ;
  assign y7690 = n18231 ;
  assign y7691 = ~1'b0 ;
  assign y7692 = n18233 ;
  assign y7693 = n18234 ;
  assign y7694 = n18240 ;
  assign y7695 = ~n18245 ;
  assign y7696 = ~n18250 ;
  assign y7697 = ~1'b0 ;
  assign y7698 = ~n18252 ;
  assign y7699 = ~n18256 ;
  assign y7700 = ~1'b0 ;
  assign y7701 = ~n18261 ;
  assign y7702 = n18262 ;
  assign y7703 = ~n18264 ;
  assign y7704 = ~n18265 ;
  assign y7705 = ~n18268 ;
  assign y7706 = n18275 ;
  assign y7707 = ~1'b0 ;
  assign y7708 = n18276 ;
  assign y7709 = n18289 ;
  assign y7710 = n18290 ;
  assign y7711 = ~1'b0 ;
  assign y7712 = n18292 ;
  assign y7713 = ~1'b0 ;
  assign y7714 = ~n18296 ;
  assign y7715 = ~1'b0 ;
  assign y7716 = ~n18297 ;
  assign y7717 = ~1'b0 ;
  assign y7718 = ~n18300 ;
  assign y7719 = ~n2941 ;
  assign y7720 = n18302 ;
  assign y7721 = ~n18303 ;
  assign y7722 = n18304 ;
  assign y7723 = n18305 ;
  assign y7724 = ~1'b0 ;
  assign y7725 = ~1'b0 ;
  assign y7726 = n11849 ;
  assign y7727 = ~n18307 ;
  assign y7728 = ~n18308 ;
  assign y7729 = ~1'b0 ;
  assign y7730 = ~n18312 ;
  assign y7731 = n18316 ;
  assign y7732 = ~n18317 ;
  assign y7733 = n18318 ;
  assign y7734 = n6298 ;
  assign y7735 = ~n18319 ;
  assign y7736 = ~n18322 ;
  assign y7737 = ~n18326 ;
  assign y7738 = ~n18332 ;
  assign y7739 = ~n18335 ;
  assign y7740 = n18342 ;
  assign y7741 = ~n18348 ;
  assign y7742 = ~1'b0 ;
  assign y7743 = n18349 ;
  assign y7744 = n18350 ;
  assign y7745 = n5043 ;
  assign y7746 = ~1'b0 ;
  assign y7747 = n18353 ;
  assign y7748 = n18358 ;
  assign y7749 = ~n18360 ;
  assign y7750 = ~n18361 ;
  assign y7751 = n1239 ;
  assign y7752 = 1'b0 ;
  assign y7753 = ~n18362 ;
  assign y7754 = n18364 ;
  assign y7755 = n18369 ;
  assign y7756 = n18370 ;
  assign y7757 = n18379 ;
  assign y7758 = ~1'b0 ;
  assign y7759 = ~1'b0 ;
  assign y7760 = ~n18382 ;
  assign y7761 = ~n18384 ;
  assign y7762 = n18386 ;
  assign y7763 = n18394 ;
  assign y7764 = ~1'b0 ;
  assign y7765 = n18400 ;
  assign y7766 = ~1'b0 ;
  assign y7767 = n18401 ;
  assign y7768 = ~1'b0 ;
  assign y7769 = n18403 ;
  assign y7770 = n18405 ;
  assign y7771 = n18409 ;
  assign y7772 = ~n18413 ;
  assign y7773 = ~1'b0 ;
  assign y7774 = 1'b0 ;
  assign y7775 = ~1'b0 ;
  assign y7776 = n18414 ;
  assign y7777 = ~1'b0 ;
  assign y7778 = n18416 ;
  assign y7779 = ~1'b0 ;
  assign y7780 = 1'b0 ;
  assign y7781 = ~1'b0 ;
  assign y7782 = n18417 ;
  assign y7783 = n18423 ;
  assign y7784 = ~1'b0 ;
  assign y7785 = n18426 ;
  assign y7786 = n18430 ;
  assign y7787 = ~n18435 ;
  assign y7788 = ~n18436 ;
  assign y7789 = n18437 ;
  assign y7790 = ~n18438 ;
  assign y7791 = n18439 ;
  assign y7792 = n18441 ;
  assign y7793 = n18444 ;
  assign y7794 = ~n18445 ;
  assign y7795 = n18447 ;
  assign y7796 = n18457 ;
  assign y7797 = n18460 ;
  assign y7798 = n18463 ;
  assign y7799 = ~n18464 ;
  assign y7800 = ~n18467 ;
  assign y7801 = ~1'b0 ;
  assign y7802 = n18470 ;
  assign y7803 = n18476 ;
  assign y7804 = n18486 ;
  assign y7805 = n18487 ;
  assign y7806 = ~n18489 ;
  assign y7807 = ~n18490 ;
  assign y7808 = ~n18494 ;
  assign y7809 = ~n18496 ;
  assign y7810 = ~n18499 ;
  assign y7811 = ~n18501 ;
  assign y7812 = ~n18504 ;
  assign y7813 = ~n18505 ;
  assign y7814 = n18506 ;
  assign y7815 = ~1'b0 ;
  assign y7816 = n18511 ;
  assign y7817 = n18512 ;
  assign y7818 = n18515 ;
  assign y7819 = ~n18517 ;
  assign y7820 = 1'b0 ;
  assign y7821 = ~1'b0 ;
  assign y7822 = n18525 ;
  assign y7823 = ~1'b0 ;
  assign y7824 = ~n18526 ;
  assign y7825 = n18528 ;
  assign y7826 = ~1'b0 ;
  assign y7827 = ~n18533 ;
  assign y7828 = ~n18534 ;
  assign y7829 = n18536 ;
  assign y7830 = n5915 ;
  assign y7831 = ~n18538 ;
  assign y7832 = n18539 ;
  assign y7833 = ~n14409 ;
  assign y7834 = ~n18542 ;
  assign y7835 = n18555 ;
  assign y7836 = n18557 ;
  assign y7837 = n18563 ;
  assign y7838 = ~1'b0 ;
  assign y7839 = ~n967 ;
  assign y7840 = ~n18568 ;
  assign y7841 = n18569 ;
  assign y7842 = n18570 ;
  assign y7843 = n18572 ;
  assign y7844 = n18577 ;
  assign y7845 = n18581 ;
  assign y7846 = ~n546 ;
  assign y7847 = n18586 ;
  assign y7848 = n18590 ;
  assign y7849 = n18591 ;
  assign y7850 = ~n18593 ;
  assign y7851 = n18594 ;
  assign y7852 = ~n18599 ;
  assign y7853 = ~n18605 ;
  assign y7854 = n18608 ;
  assign y7855 = n18612 ;
  assign y7856 = ~n18613 ;
  assign y7857 = ~n18619 ;
  assign y7858 = n18621 ;
  assign y7859 = ~1'b0 ;
  assign y7860 = n18626 ;
  assign y7861 = ~n18627 ;
  assign y7862 = n18628 ;
  assign y7863 = n18631 ;
  assign y7864 = ~n18632 ;
  assign y7865 = n18639 ;
  assign y7866 = ~1'b0 ;
  assign y7867 = n18643 ;
  assign y7868 = n18644 ;
  assign y7869 = n18648 ;
  assign y7870 = ~n18649 ;
  assign y7871 = n18650 ;
  assign y7872 = ~n18652 ;
  assign y7873 = ~n18655 ;
  assign y7874 = n18656 ;
  assign y7875 = ~n18658 ;
  assign y7876 = ~n18660 ;
  assign y7877 = n18666 ;
  assign y7878 = n18671 ;
  assign y7879 = ~n18674 ;
  assign y7880 = ~n18678 ;
  assign y7881 = n18679 ;
  assign y7882 = n18680 ;
  assign y7883 = ~1'b0 ;
  assign y7884 = n18682 ;
  assign y7885 = n18691 ;
  assign y7886 = n18693 ;
  assign y7887 = ~n18694 ;
  assign y7888 = ~n18695 ;
  assign y7889 = ~1'b0 ;
  assign y7890 = ~n18696 ;
  assign y7891 = n18699 ;
  assign y7892 = n18705 ;
  assign y7893 = ~1'b0 ;
  assign y7894 = ~1'b0 ;
  assign y7895 = ~1'b0 ;
  assign y7896 = n18706 ;
  assign y7897 = ~1'b0 ;
  assign y7898 = ~n18707 ;
  assign y7899 = n18708 ;
  assign y7900 = n18710 ;
  assign y7901 = n18712 ;
  assign y7902 = ~n18714 ;
  assign y7903 = ~1'b0 ;
  assign y7904 = ~n4802 ;
  assign y7905 = ~1'b0 ;
  assign y7906 = n18716 ;
  assign y7907 = n18721 ;
  assign y7908 = ~n18722 ;
  assign y7909 = ~n18723 ;
  assign y7910 = n2675 ;
  assign y7911 = ~1'b0 ;
  assign y7912 = ~1'b0 ;
  assign y7913 = n18726 ;
  assign y7914 = ~1'b0 ;
  assign y7915 = ~1'b0 ;
  assign y7916 = n18733 ;
  assign y7917 = ~n18734 ;
  assign y7918 = n18735 ;
  assign y7919 = n18739 ;
  assign y7920 = n18741 ;
  assign y7921 = n18746 ;
  assign y7922 = ~n18750 ;
  assign y7923 = n18752 ;
  assign y7924 = ~n18753 ;
  assign y7925 = n18754 ;
  assign y7926 = ~1'b0 ;
  assign y7927 = ~n18755 ;
  assign y7928 = n18759 ;
  assign y7929 = n18764 ;
  assign y7930 = ~n15275 ;
  assign y7931 = ~n18768 ;
  assign y7932 = ~n18769 ;
  assign y7933 = n18770 ;
  assign y7934 = ~1'b0 ;
  assign y7935 = ~n18772 ;
  assign y7936 = n18774 ;
  assign y7937 = ~n18777 ;
  assign y7938 = ~n18778 ;
  assign y7939 = ~1'b0 ;
  assign y7940 = n18779 ;
  assign y7941 = ~1'b0 ;
  assign y7942 = ~1'b0 ;
  assign y7943 = ~1'b0 ;
  assign y7944 = n18790 ;
  assign y7945 = n18795 ;
  assign y7946 = ~n18800 ;
  assign y7947 = ~n18801 ;
  assign y7948 = ~1'b0 ;
  assign y7949 = n18808 ;
  assign y7950 = n18810 ;
  assign y7951 = ~1'b0 ;
  assign y7952 = ~n18818 ;
  assign y7953 = ~n18820 ;
  assign y7954 = ~n18824 ;
  assign y7955 = ~n18825 ;
  assign y7956 = ~1'b0 ;
  assign y7957 = n18828 ;
  assign y7958 = n18833 ;
  assign y7959 = ~n18834 ;
  assign y7960 = n18842 ;
  assign y7961 = n18848 ;
  assign y7962 = n18850 ;
  assign y7963 = ~n18853 ;
  assign y7964 = n18857 ;
  assign y7965 = ~n18858 ;
  assign y7966 = ~1'b0 ;
  assign y7967 = n18860 ;
  assign y7968 = ~1'b0 ;
  assign y7969 = ~1'b0 ;
  assign y7970 = ~1'b0 ;
  assign y7971 = ~n18861 ;
  assign y7972 = n18862 ;
  assign y7973 = ~n16827 ;
  assign y7974 = n18863 ;
  assign y7975 = n18864 ;
  assign y7976 = n18865 ;
  assign y7977 = n18866 ;
  assign y7978 = ~n18869 ;
  assign y7979 = n18871 ;
  assign y7980 = ~1'b0 ;
  assign y7981 = n18876 ;
  assign y7982 = n18878 ;
  assign y7983 = n18882 ;
  assign y7984 = ~n18883 ;
  assign y7985 = n18886 ;
  assign y7986 = ~n18888 ;
  assign y7987 = n18896 ;
  assign y7988 = n18899 ;
  assign y7989 = ~n18902 ;
  assign y7990 = n18905 ;
  assign y7991 = ~1'b0 ;
  assign y7992 = ~n18906 ;
  assign y7993 = ~n18908 ;
  assign y7994 = ~n18914 ;
  assign y7995 = n18921 ;
  assign y7996 = 1'b0 ;
  assign y7997 = n18923 ;
  assign y7998 = ~1'b0 ;
  assign y7999 = ~n18924 ;
  assign y8000 = ~n18925 ;
  assign y8001 = ~n18927 ;
  assign y8002 = n18932 ;
  assign y8003 = ~1'b0 ;
  assign y8004 = ~1'b0 ;
  assign y8005 = n18934 ;
  assign y8006 = 1'b0 ;
  assign y8007 = ~n18945 ;
  assign y8008 = ~1'b0 ;
  assign y8009 = ~1'b0 ;
  assign y8010 = ~n18948 ;
  assign y8011 = n18951 ;
  assign y8012 = n18953 ;
  assign y8013 = ~n18955 ;
  assign y8014 = ~1'b0 ;
  assign y8015 = 1'b0 ;
  assign y8016 = ~n18957 ;
  assign y8017 = n18958 ;
  assign y8018 = ~n18959 ;
  assign y8019 = n18961 ;
  assign y8020 = ~n18964 ;
  assign y8021 = ~n18966 ;
  assign y8022 = n18970 ;
  assign y8023 = ~n18972 ;
  assign y8024 = ~1'b0 ;
  assign y8025 = ~1'b0 ;
  assign y8026 = ~1'b0 ;
  assign y8027 = ~n10745 ;
  assign y8028 = ~n18975 ;
  assign y8029 = ~n18977 ;
  assign y8030 = n18980 ;
  assign y8031 = n18984 ;
  assign y8032 = ~n18988 ;
  assign y8033 = ~1'b0 ;
  assign y8034 = n18989 ;
  assign y8035 = ~n18992 ;
  assign y8036 = ~1'b0 ;
  assign y8037 = n18993 ;
  assign y8038 = n18996 ;
  assign y8039 = n18997 ;
  assign y8040 = ~n19002 ;
  assign y8041 = ~n19003 ;
  assign y8042 = ~1'b0 ;
  assign y8043 = ~1'b0 ;
  assign y8044 = n19005 ;
  assign y8045 = ~n19007 ;
  assign y8046 = n19010 ;
  assign y8047 = 1'b0 ;
  assign y8048 = n19011 ;
  assign y8049 = ~1'b0 ;
  assign y8050 = ~1'b0 ;
  assign y8051 = ~1'b0 ;
  assign y8052 = n19012 ;
  assign y8053 = ~1'b0 ;
  assign y8054 = n19014 ;
  assign y8055 = n14138 ;
  assign y8056 = ~1'b0 ;
  assign y8057 = ~1'b0 ;
  assign y8058 = ~n19015 ;
  assign y8059 = ~1'b0 ;
  assign y8060 = ~1'b0 ;
  assign y8061 = ~n19018 ;
  assign y8062 = ~n2440 ;
  assign y8063 = ~n2130 ;
  assign y8064 = ~n9035 ;
  assign y8065 = n19020 ;
  assign y8066 = ~n19021 ;
  assign y8067 = n19023 ;
  assign y8068 = ~n19029 ;
  assign y8069 = n12154 ;
  assign y8070 = ~1'b0 ;
  assign y8071 = ~n19036 ;
  assign y8072 = n19037 ;
  assign y8073 = n19041 ;
  assign y8074 = ~n19047 ;
  assign y8075 = ~n19048 ;
  assign y8076 = n19049 ;
  assign y8077 = ~n19052 ;
  assign y8078 = n19054 ;
  assign y8079 = ~n19061 ;
  assign y8080 = n19062 ;
  assign y8081 = ~n19072 ;
  assign y8082 = ~n19078 ;
  assign y8083 = n19083 ;
  assign y8084 = ~1'b0 ;
  assign y8085 = ~1'b0 ;
  assign y8086 = n19088 ;
  assign y8087 = ~1'b0 ;
  assign y8088 = ~n19089 ;
  assign y8089 = ~1'b0 ;
  assign y8090 = ~n19092 ;
  assign y8091 = n19093 ;
  assign y8092 = ~n1851 ;
  assign y8093 = ~1'b0 ;
  assign y8094 = ~n19097 ;
  assign y8095 = n19106 ;
  assign y8096 = n19115 ;
  assign y8097 = ~1'b0 ;
  assign y8098 = ~1'b0 ;
  assign y8099 = n19117 ;
  assign y8100 = n19118 ;
  assign y8101 = ~n19123 ;
  assign y8102 = n19124 ;
  assign y8103 = n19125 ;
  assign y8104 = ~1'b0 ;
  assign y8105 = ~1'b0 ;
  assign y8106 = ~n19127 ;
  assign y8107 = ~n19132 ;
  assign y8108 = n19134 ;
  assign y8109 = n19135 ;
  assign y8110 = n19139 ;
  assign y8111 = ~n19144 ;
  assign y8112 = ~n19145 ;
  assign y8113 = n19149 ;
  assign y8114 = ~1'b0 ;
  assign y8115 = ~1'b0 ;
  assign y8116 = n19153 ;
  assign y8117 = ~n19157 ;
  assign y8118 = ~n19158 ;
  assign y8119 = ~1'b0 ;
  assign y8120 = ~n19159 ;
  assign y8121 = n19162 ;
  assign y8122 = ~1'b0 ;
  assign y8123 = ~1'b0 ;
  assign y8124 = ~1'b0 ;
  assign y8125 = ~1'b0 ;
  assign y8126 = n19164 ;
  assign y8127 = ~n19167 ;
  assign y8128 = ~n19168 ;
  assign y8129 = ~1'b0 ;
  assign y8130 = ~n19170 ;
  assign y8131 = n19173 ;
  assign y8132 = n19175 ;
  assign y8133 = ~n10289 ;
  assign y8134 = n19183 ;
  assign y8135 = n19189 ;
  assign y8136 = ~n19190 ;
  assign y8137 = ~n19193 ;
  assign y8138 = ~n19194 ;
  assign y8139 = ~n19214 ;
  assign y8140 = ~1'b0 ;
  assign y8141 = ~n19215 ;
  assign y8142 = n19228 ;
  assign y8143 = ~n19233 ;
  assign y8144 = ~1'b0 ;
  assign y8145 = ~1'b0 ;
  assign y8146 = n19234 ;
  assign y8147 = ~n19236 ;
  assign y8148 = ~n19238 ;
  assign y8149 = ~n19240 ;
  assign y8150 = ~n19242 ;
  assign y8151 = n19245 ;
  assign y8152 = ~1'b0 ;
  assign y8153 = ~1'b0 ;
  assign y8154 = n19248 ;
  assign y8155 = n19249 ;
  assign y8156 = ~1'b0 ;
  assign y8157 = ~n19251 ;
  assign y8158 = n19255 ;
  assign y8159 = ~n19257 ;
  assign y8160 = ~n19259 ;
  assign y8161 = n1314 ;
  assign y8162 = n19263 ;
  assign y8163 = ~n19264 ;
  assign y8164 = n19265 ;
  assign y8165 = n19274 ;
  assign y8166 = ~n19277 ;
  assign y8167 = n19289 ;
  assign y8168 = ~1'b0 ;
  assign y8169 = ~n19290 ;
  assign y8170 = ~n19293 ;
  assign y8171 = ~n19302 ;
  assign y8172 = ~n19313 ;
  assign y8173 = ~1'b0 ;
  assign y8174 = n19317 ;
  assign y8175 = n19318 ;
  assign y8176 = ~1'b0 ;
  assign y8177 = n19319 ;
  assign y8178 = ~1'b0 ;
  assign y8179 = ~n19320 ;
  assign y8180 = ~n19321 ;
  assign y8181 = ~n19328 ;
  assign y8182 = ~n19361 ;
  assign y8183 = ~1'b0 ;
  assign y8184 = 1'b0 ;
  assign y8185 = ~n19364 ;
  assign y8186 = n19365 ;
  assign y8187 = n19366 ;
  assign y8188 = ~1'b0 ;
  assign y8189 = n19367 ;
  assign y8190 = 1'b0 ;
  assign y8191 = ~n19369 ;
  assign y8192 = ~n19371 ;
  assign y8193 = n19374 ;
  assign y8194 = ~1'b0 ;
  assign y8195 = n19375 ;
  assign y8196 = ~n19378 ;
  assign y8197 = ~n19382 ;
  assign y8198 = n19384 ;
  assign y8199 = ~1'b0 ;
  assign y8200 = ~n19385 ;
  assign y8201 = ~n19387 ;
  assign y8202 = n19389 ;
  assign y8203 = ~1'b0 ;
  assign y8204 = ~n19393 ;
  assign y8205 = n19395 ;
  assign y8206 = ~1'b0 ;
  assign y8207 = ~n19398 ;
  assign y8208 = ~1'b0 ;
  assign y8209 = ~n19399 ;
  assign y8210 = ~n17178 ;
  assign y8211 = ~n19400 ;
  assign y8212 = ~n19402 ;
  assign y8213 = ~n19406 ;
  assign y8214 = n7376 ;
  assign y8215 = n19407 ;
  assign y8216 = ~n19410 ;
  assign y8217 = ~n19416 ;
  assign y8218 = ~1'b0 ;
  assign y8219 = 1'b0 ;
  assign y8220 = n19419 ;
  assign y8221 = ~n19421 ;
  assign y8222 = n19422 ;
  assign y8223 = n19427 ;
  assign y8224 = n19428 ;
  assign y8225 = n19430 ;
  assign y8226 = n19432 ;
  assign y8227 = ~1'b0 ;
  assign y8228 = ~n19435 ;
  assign y8229 = ~n19442 ;
  assign y8230 = ~n19445 ;
  assign y8231 = ~1'b0 ;
  assign y8232 = n19449 ;
  assign y8233 = n19450 ;
  assign y8234 = ~n19451 ;
  assign y8235 = n19453 ;
  assign y8236 = ~n19455 ;
  assign y8237 = n19459 ;
  assign y8238 = n19460 ;
  assign y8239 = n19461 ;
  assign y8240 = n19464 ;
  assign y8241 = ~n19465 ;
  assign y8242 = n2847 ;
  assign y8243 = n19467 ;
  assign y8244 = ~1'b0 ;
  assign y8245 = ~1'b0 ;
  assign y8246 = ~n19475 ;
  assign y8247 = ~n19476 ;
  assign y8248 = ~n19477 ;
  assign y8249 = n8029 ;
  assign y8250 = ~n19478 ;
  assign y8251 = ~n14619 ;
  assign y8252 = ~1'b0 ;
  assign y8253 = ~n19481 ;
  assign y8254 = ~n19482 ;
  assign y8255 = ~1'b0 ;
  assign y8256 = ~n19483 ;
  assign y8257 = ~n19486 ;
  assign y8258 = ~1'b0 ;
  assign y8259 = ~n19489 ;
  assign y8260 = ~n19492 ;
  assign y8261 = ~n19495 ;
  assign y8262 = ~n19508 ;
  assign y8263 = n19512 ;
  assign y8264 = n19513 ;
  assign y8265 = ~1'b0 ;
  assign y8266 = n19516 ;
  assign y8267 = n13925 ;
  assign y8268 = ~1'b0 ;
  assign y8269 = ~n19517 ;
  assign y8270 = n19521 ;
  assign y8271 = ~1'b0 ;
  assign y8272 = ~n19522 ;
  assign y8273 = ~1'b0 ;
  assign y8274 = n19528 ;
  assign y8275 = ~n19532 ;
  assign y8276 = ~n1255 ;
  assign y8277 = ~n19540 ;
  assign y8278 = ~n19542 ;
  assign y8279 = ~1'b0 ;
  assign y8280 = ~n19545 ;
  assign y8281 = ~1'b0 ;
  assign y8282 = ~1'b0 ;
  assign y8283 = ~n19553 ;
  assign y8284 = ~n19556 ;
  assign y8285 = n19561 ;
  assign y8286 = n19562 ;
  assign y8287 = n19563 ;
  assign y8288 = n19564 ;
  assign y8289 = ~n19568 ;
  assign y8290 = ~n19569 ;
  assign y8291 = n19570 ;
  assign y8292 = n19574 ;
  assign y8293 = ~n16126 ;
  assign y8294 = n19575 ;
  assign y8295 = ~n19582 ;
  assign y8296 = ~n19591 ;
  assign y8297 = ~n19593 ;
  assign y8298 = ~1'b0 ;
  assign y8299 = ~n19596 ;
  assign y8300 = n19599 ;
  assign y8301 = n19600 ;
  assign y8302 = ~n19606 ;
  assign y8303 = ~1'b0 ;
  assign y8304 = ~1'b0 ;
  assign y8305 = ~1'b0 ;
  assign y8306 = ~1'b0 ;
  assign y8307 = n19607 ;
  assign y8308 = ~n19608 ;
  assign y8309 = ~1'b0 ;
  assign y8310 = ~1'b0 ;
  assign y8311 = 1'b0 ;
  assign y8312 = ~n19609 ;
  assign y8313 = ~1'b0 ;
  assign y8314 = ~1'b0 ;
  assign y8315 = ~n19613 ;
  assign y8316 = ~1'b0 ;
  assign y8317 = ~n19614 ;
  assign y8318 = ~n19619 ;
  assign y8319 = n19620 ;
  assign y8320 = n19622 ;
  assign y8321 = ~1'b0 ;
  assign y8322 = ~1'b0 ;
  assign y8323 = ~n19626 ;
  assign y8324 = ~n3343 ;
  assign y8325 = n19627 ;
  assign y8326 = ~1'b0 ;
  assign y8327 = ~n19634 ;
  assign y8328 = ~n19643 ;
  assign y8329 = n19647 ;
  assign y8330 = n19648 ;
  assign y8331 = ~n19650 ;
  assign y8332 = ~n19651 ;
  assign y8333 = ~1'b0 ;
  assign y8334 = ~n19654 ;
  assign y8335 = n19657 ;
  assign y8336 = ~n19661 ;
  assign y8337 = ~n19662 ;
  assign y8338 = n19666 ;
  assign y8339 = n19667 ;
  assign y8340 = ~1'b0 ;
  assign y8341 = ~1'b0 ;
  assign y8342 = ~1'b0 ;
  assign y8343 = ~n19668 ;
  assign y8344 = ~n19669 ;
  assign y8345 = ~n19672 ;
  assign y8346 = ~n19675 ;
  assign y8347 = n19678 ;
  assign y8348 = n19683 ;
  assign y8349 = ~n19687 ;
  assign y8350 = ~1'b0 ;
  assign y8351 = n19690 ;
  assign y8352 = n19692 ;
  assign y8353 = ~n10364 ;
  assign y8354 = n19697 ;
  assign y8355 = ~1'b0 ;
  assign y8356 = ~n19699 ;
  assign y8357 = ~n19701 ;
  assign y8358 = ~n11587 ;
  assign y8359 = n19703 ;
  assign y8360 = ~n19706 ;
  assign y8361 = ~1'b0 ;
  assign y8362 = ~1'b0 ;
  assign y8363 = n19710 ;
  assign y8364 = n19712 ;
  assign y8365 = n19718 ;
  assign y8366 = n19719 ;
  assign y8367 = n19720 ;
  assign y8368 = ~n19725 ;
  assign y8369 = n19727 ;
  assign y8370 = n19728 ;
  assign y8371 = ~n19729 ;
  assign y8372 = ~n19734 ;
  assign y8373 = n19737 ;
  assign y8374 = n19738 ;
  assign y8375 = n19739 ;
  assign y8376 = ~1'b0 ;
  assign y8377 = ~n19741 ;
  assign y8378 = ~n19744 ;
  assign y8379 = ~n19746 ;
  assign y8380 = ~n19747 ;
  assign y8381 = ~n19750 ;
  assign y8382 = ~n19751 ;
  assign y8383 = n19760 ;
  assign y8384 = ~n19761 ;
  assign y8385 = n19762 ;
  assign y8386 = ~1'b0 ;
  assign y8387 = n19767 ;
  assign y8388 = n19768 ;
  assign y8389 = n19781 ;
  assign y8390 = ~1'b0 ;
  assign y8391 = n19787 ;
  assign y8392 = ~1'b0 ;
  assign y8393 = n19788 ;
  assign y8394 = ~n19791 ;
  assign y8395 = ~n19794 ;
  assign y8396 = n19796 ;
  assign y8397 = ~n19803 ;
  assign y8398 = n19806 ;
  assign y8399 = ~n19811 ;
  assign y8400 = ~1'b0 ;
  assign y8401 = n19813 ;
  assign y8402 = n19816 ;
  assign y8403 = n16891 ;
  assign y8404 = n19818 ;
  assign y8405 = ~1'b0 ;
  assign y8406 = n19823 ;
  assign y8407 = ~1'b0 ;
  assign y8408 = ~1'b0 ;
  assign y8409 = n19831 ;
  assign y8410 = ~n19839 ;
  assign y8411 = ~n19842 ;
  assign y8412 = ~n19844 ;
  assign y8413 = n19852 ;
  assign y8414 = ~n19854 ;
  assign y8415 = ~n19857 ;
  assign y8416 = n19859 ;
  assign y8417 = ~1'b0 ;
  assign y8418 = ~1'b0 ;
  assign y8419 = ~n19864 ;
  assign y8420 = n19869 ;
  assign y8421 = ~n19870 ;
  assign y8422 = n19871 ;
  assign y8423 = ~1'b0 ;
  assign y8424 = ~n19876 ;
  assign y8425 = ~n19878 ;
  assign y8426 = n19881 ;
  assign y8427 = n19895 ;
  assign y8428 = ~1'b0 ;
  assign y8429 = ~1'b0 ;
  assign y8430 = ~n19896 ;
  assign y8431 = ~1'b0 ;
  assign y8432 = ~1'b0 ;
  assign y8433 = ~1'b0 ;
  assign y8434 = ~n456 ;
  assign y8435 = n19900 ;
  assign y8436 = n19901 ;
  assign y8437 = ~n19903 ;
  assign y8438 = n19904 ;
  assign y8439 = ~n19906 ;
  assign y8440 = ~1'b0 ;
  assign y8441 = ~n15070 ;
  assign y8442 = ~1'b0 ;
  assign y8443 = n19911 ;
  assign y8444 = ~1'b0 ;
  assign y8445 = ~1'b0 ;
  assign y8446 = ~n19915 ;
  assign y8447 = ~n11380 ;
  assign y8448 = n19916 ;
  assign y8449 = ~1'b0 ;
  assign y8450 = ~n19920 ;
  assign y8451 = ~1'b0 ;
  assign y8452 = ~1'b0 ;
  assign y8453 = ~1'b0 ;
  assign y8454 = ~n19923 ;
  assign y8455 = ~n19925 ;
  assign y8456 = ~n19929 ;
  assign y8457 = ~1'b0 ;
  assign y8458 = n19931 ;
  assign y8459 = ~1'b0 ;
  assign y8460 = ~n19934 ;
  assign y8461 = ~n19935 ;
  assign y8462 = n19939 ;
  assign y8463 = n19950 ;
  assign y8464 = ~n19957 ;
  assign y8465 = ~n19958 ;
  assign y8466 = ~n19960 ;
  assign y8467 = ~1'b0 ;
  assign y8468 = ~n19966 ;
  assign y8469 = ~n19970 ;
  assign y8470 = n19976 ;
  assign y8471 = ~n18323 ;
  assign y8472 = ~n19978 ;
  assign y8473 = ~n19980 ;
  assign y8474 = n19985 ;
  assign y8475 = ~n19986 ;
  assign y8476 = ~n19988 ;
  assign y8477 = ~n19991 ;
  assign y8478 = ~n19994 ;
  assign y8479 = ~n19995 ;
  assign y8480 = n19996 ;
  assign y8481 = n20001 ;
  assign y8482 = n20006 ;
  assign y8483 = ~n20012 ;
  assign y8484 = n20013 ;
  assign y8485 = n20015 ;
  assign y8486 = n20021 ;
  assign y8487 = ~n20023 ;
  assign y8488 = n20024 ;
  assign y8489 = n20028 ;
  assign y8490 = ~n20029 ;
  assign y8491 = ~n20033 ;
  assign y8492 = ~n20035 ;
  assign y8493 = ~1'b0 ;
  assign y8494 = n20037 ;
  assign y8495 = n20040 ;
  assign y8496 = n20042 ;
  assign y8497 = n20049 ;
  assign y8498 = ~n20053 ;
  assign y8499 = ~n20058 ;
  assign y8500 = ~1'b0 ;
  assign y8501 = ~1'b0 ;
  assign y8502 = n18953 ;
  assign y8503 = n18850 ;
  assign y8504 = n20059 ;
  assign y8505 = ~n20061 ;
  assign y8506 = n17532 ;
  assign y8507 = ~n20062 ;
  assign y8508 = ~n20064 ;
  assign y8509 = n20065 ;
  assign y8510 = ~n20066 ;
  assign y8511 = n20068 ;
  assign y8512 = ~1'b0 ;
  assign y8513 = ~1'b0 ;
  assign y8514 = n20070 ;
  assign y8515 = ~1'b0 ;
  assign y8516 = n20071 ;
  assign y8517 = ~n3965 ;
  assign y8518 = ~n20074 ;
  assign y8519 = ~n20077 ;
  assign y8520 = ~n20078 ;
  assign y8521 = n20079 ;
  assign y8522 = n2488 ;
  assign y8523 = ~1'b0 ;
  assign y8524 = ~n20087 ;
  assign y8525 = ~1'b0 ;
  assign y8526 = ~n20091 ;
  assign y8527 = ~n20093 ;
  assign y8528 = n20099 ;
  assign y8529 = n20109 ;
  assign y8530 = ~1'b0 ;
  assign y8531 = ~1'b0 ;
  assign y8532 = ~n20114 ;
  assign y8533 = ~n20119 ;
  assign y8534 = ~1'b0 ;
  assign y8535 = ~n20120 ;
  assign y8536 = ~1'b0 ;
  assign y8537 = n20121 ;
  assign y8538 = n20122 ;
  assign y8539 = ~n20123 ;
  assign y8540 = ~n20133 ;
  assign y8541 = ~1'b0 ;
  assign y8542 = n20134 ;
  assign y8543 = n20135 ;
  assign y8544 = n5378 ;
  assign y8545 = ~n20138 ;
  assign y8546 = n20140 ;
  assign y8547 = 1'b0 ;
  assign y8548 = ~n20144 ;
  assign y8549 = ~1'b0 ;
  assign y8550 = ~1'b0 ;
  assign y8551 = n20148 ;
  assign y8552 = ~n20150 ;
  assign y8553 = ~n20151 ;
  assign y8554 = ~n20152 ;
  assign y8555 = n20153 ;
  assign y8556 = ~n20155 ;
  assign y8557 = n20157 ;
  assign y8558 = n20160 ;
  assign y8559 = ~1'b0 ;
  assign y8560 = ~1'b0 ;
  assign y8561 = ~n20162 ;
  assign y8562 = n20168 ;
  assign y8563 = ~n20169 ;
  assign y8564 = n20173 ;
  assign y8565 = ~n20175 ;
  assign y8566 = ~n20177 ;
  assign y8567 = ~n20179 ;
  assign y8568 = ~n20181 ;
  assign y8569 = ~n20183 ;
  assign y8570 = ~1'b0 ;
  assign y8571 = ~n20187 ;
  assign y8572 = ~1'b0 ;
  assign y8573 = ~n20195 ;
  assign y8574 = n20196 ;
  assign y8575 = ~n20197 ;
  assign y8576 = n20202 ;
  assign y8577 = n20208 ;
  assign y8578 = n20221 ;
  assign y8579 = ~n20224 ;
  assign y8580 = n20226 ;
  assign y8581 = ~n20234 ;
  assign y8582 = ~1'b0 ;
  assign y8583 = ~n20235 ;
  assign y8584 = n20237 ;
  assign y8585 = n13926 ;
  assign y8586 = ~n20240 ;
  assign y8587 = ~1'b0 ;
  assign y8588 = ~n20254 ;
  assign y8589 = ~1'b0 ;
  assign y8590 = n20255 ;
  assign y8591 = ~n20261 ;
  assign y8592 = n20262 ;
  assign y8593 = ~n20267 ;
  assign y8594 = ~n20268 ;
  assign y8595 = ~n20270 ;
  assign y8596 = ~n20275 ;
  assign y8597 = ~1'b0 ;
  assign y8598 = n20277 ;
  assign y8599 = n20283 ;
  assign y8600 = ~n20288 ;
  assign y8601 = ~1'b0 ;
  assign y8602 = ~1'b0 ;
  assign y8603 = n20291 ;
  assign y8604 = ~n20292 ;
  assign y8605 = n20295 ;
  assign y8606 = n10203 ;
  assign y8607 = ~n8690 ;
  assign y8608 = ~n20298 ;
  assign y8609 = ~n20299 ;
  assign y8610 = ~n20301 ;
  assign y8611 = n20302 ;
  assign y8612 = ~n20308 ;
  assign y8613 = ~1'b0 ;
  assign y8614 = ~1'b0 ;
  assign y8615 = ~n20317 ;
  assign y8616 = n20320 ;
  assign y8617 = ~n20322 ;
  assign y8618 = ~1'b0 ;
  assign y8619 = ~1'b0 ;
  assign y8620 = n20326 ;
  assign y8621 = ~1'b0 ;
  assign y8622 = ~n20331 ;
  assign y8623 = n20337 ;
  assign y8624 = ~n8927 ;
  assign y8625 = ~n20340 ;
  assign y8626 = ~1'b0 ;
  assign y8627 = ~1'b0 ;
  assign y8628 = n20341 ;
  assign y8629 = ~n20349 ;
  assign y8630 = ~n20350 ;
  assign y8631 = n20355 ;
  assign y8632 = ~1'b0 ;
  assign y8633 = ~1'b0 ;
  assign y8634 = n20357 ;
  assign y8635 = ~n20361 ;
  assign y8636 = n20367 ;
  assign y8637 = ~1'b0 ;
  assign y8638 = n20370 ;
  assign y8639 = n20371 ;
  assign y8640 = n20380 ;
  assign y8641 = n20385 ;
  assign y8642 = n20388 ;
  assign y8643 = n20389 ;
  assign y8644 = n20390 ;
  assign y8645 = ~n20393 ;
  assign y8646 = ~n20394 ;
  assign y8647 = ~1'b0 ;
  assign y8648 = n20398 ;
  assign y8649 = ~n20401 ;
  assign y8650 = ~1'b0 ;
  assign y8651 = n20405 ;
  assign y8652 = n6711 ;
  assign y8653 = ~n6647 ;
  assign y8654 = n20413 ;
  assign y8655 = ~n13161 ;
  assign y8656 = n20414 ;
  assign y8657 = ~1'b0 ;
  assign y8658 = n20415 ;
  assign y8659 = ~1'b0 ;
  assign y8660 = ~n20416 ;
  assign y8661 = n20424 ;
  assign y8662 = ~n4144 ;
  assign y8663 = n2118 ;
  assign y8664 = ~n20429 ;
  assign y8665 = ~1'b0 ;
  assign y8666 = ~n20435 ;
  assign y8667 = ~n20436 ;
  assign y8668 = n20437 ;
  assign y8669 = n20442 ;
  assign y8670 = ~1'b0 ;
  assign y8671 = ~n20445 ;
  assign y8672 = ~n20448 ;
  assign y8673 = n12131 ;
  assign y8674 = ~n20453 ;
  assign y8675 = n20458 ;
  assign y8676 = 1'b0 ;
  assign y8677 = ~n20459 ;
  assign y8678 = ~n20460 ;
  assign y8679 = ~n20461 ;
  assign y8680 = n19583 ;
  assign y8681 = n20462 ;
  assign y8682 = ~n20463 ;
  assign y8683 = ~n20469 ;
  assign y8684 = ~1'b0 ;
  assign y8685 = ~n20471 ;
  assign y8686 = n20478 ;
  assign y8687 = n20484 ;
  assign y8688 = ~1'b0 ;
  assign y8689 = ~1'b0 ;
  assign y8690 = ~1'b0 ;
  assign y8691 = n20486 ;
  assign y8692 = n20494 ;
  assign y8693 = ~n20501 ;
  assign y8694 = ~1'b0 ;
  assign y8695 = n20502 ;
  assign y8696 = n20504 ;
  assign y8697 = ~1'b0 ;
  assign y8698 = ~1'b0 ;
  assign y8699 = ~n20505 ;
  assign y8700 = ~n20506 ;
  assign y8701 = n20507 ;
  assign y8702 = n20512 ;
  assign y8703 = n20519 ;
  assign y8704 = ~1'b0 ;
  assign y8705 = ~1'b0 ;
  assign y8706 = n20521 ;
  assign y8707 = ~n20523 ;
  assign y8708 = ~1'b0 ;
  assign y8709 = ~n20525 ;
  assign y8710 = ~1'b0 ;
  assign y8711 = ~n20528 ;
  assign y8712 = ~n20529 ;
  assign y8713 = ~1'b0 ;
  assign y8714 = n5348 ;
  assign y8715 = ~1'b0 ;
  assign y8716 = n20537 ;
  assign y8717 = ~1'b0 ;
  assign y8718 = ~n20539 ;
  assign y8719 = ~n20551 ;
  assign y8720 = n20552 ;
  assign y8721 = n20556 ;
  assign y8722 = n7306 ;
  assign y8723 = ~1'b0 ;
  assign y8724 = n20557 ;
  assign y8725 = ~n20565 ;
  assign y8726 = ~1'b0 ;
  assign y8727 = n20567 ;
  assign y8728 = ~1'b0 ;
  assign y8729 = ~n20569 ;
  assign y8730 = ~n14483 ;
  assign y8731 = n20572 ;
  assign y8732 = n11844 ;
  assign y8733 = n20575 ;
  assign y8734 = ~n20577 ;
  assign y8735 = n20578 ;
  assign y8736 = n20580 ;
  assign y8737 = ~n20589 ;
  assign y8738 = n20590 ;
  assign y8739 = ~n20593 ;
  assign y8740 = n20596 ;
  assign y8741 = ~n20597 ;
  assign y8742 = ~n20598 ;
  assign y8743 = n20600 ;
  assign y8744 = n20602 ;
  assign y8745 = n20607 ;
  assign y8746 = n20608 ;
  assign y8747 = ~n20610 ;
  assign y8748 = n20613 ;
  assign y8749 = ~n20621 ;
  assign y8750 = ~1'b0 ;
  assign y8751 = n20622 ;
  assign y8752 = ~n20623 ;
  assign y8753 = n20629 ;
  assign y8754 = ~1'b0 ;
  assign y8755 = ~n20633 ;
  assign y8756 = n20638 ;
  assign y8757 = ~1'b0 ;
  assign y8758 = ~1'b0 ;
  assign y8759 = n20640 ;
  assign y8760 = ~n20642 ;
  assign y8761 = ~1'b0 ;
  assign y8762 = n20647 ;
  assign y8763 = n20652 ;
  assign y8764 = ~n20654 ;
  assign y8765 = n20656 ;
  assign y8766 = ~n20660 ;
  assign y8767 = ~n20663 ;
  assign y8768 = n20668 ;
  assign y8769 = ~n20669 ;
  assign y8770 = ~n20673 ;
  assign y8771 = ~n20677 ;
  assign y8772 = ~n20680 ;
  assign y8773 = ~n20681 ;
  assign y8774 = ~1'b0 ;
  assign y8775 = 1'b0 ;
  assign y8776 = n20690 ;
  assign y8777 = n20691 ;
  assign y8778 = x7 ;
  assign y8779 = ~1'b0 ;
  assign y8780 = ~1'b0 ;
  assign y8781 = ~1'b0 ;
  assign y8782 = ~1'b0 ;
  assign y8783 = ~n20692 ;
  assign y8784 = n14171 ;
  assign y8785 = n20694 ;
  assign y8786 = ~n20697 ;
  assign y8787 = ~1'b0 ;
  assign y8788 = ~1'b0 ;
  assign y8789 = ~1'b0 ;
  assign y8790 = n20699 ;
  assign y8791 = ~n20701 ;
  assign y8792 = n20702 ;
  assign y8793 = ~n20704 ;
  assign y8794 = ~1'b0 ;
  assign y8795 = ~1'b0 ;
  assign y8796 = n20709 ;
  assign y8797 = n20710 ;
  assign y8798 = ~1'b0 ;
  assign y8799 = ~n20713 ;
  assign y8800 = ~n20715 ;
  assign y8801 = ~n20716 ;
  assign y8802 = n20717 ;
  assign y8803 = ~1'b0 ;
  assign y8804 = ~n20722 ;
  assign y8805 = n20725 ;
  assign y8806 = ~n20728 ;
  assign y8807 = ~n20734 ;
  assign y8808 = ~1'b0 ;
  assign y8809 = n20736 ;
  assign y8810 = ~n7552 ;
  assign y8811 = ~n20740 ;
  assign y8812 = ~n20745 ;
  assign y8813 = ~n20746 ;
  assign y8814 = n20747 ;
  assign y8815 = n9752 ;
  assign y8816 = n20750 ;
  assign y8817 = n20757 ;
  assign y8818 = 1'b0 ;
  assign y8819 = ~n20760 ;
  assign y8820 = ~1'b0 ;
  assign y8821 = n20764 ;
  assign y8822 = n20766 ;
  assign y8823 = ~n20773 ;
  assign y8824 = ~n20776 ;
  assign y8825 = n20785 ;
  assign y8826 = ~n20786 ;
  assign y8827 = ~1'b0 ;
  assign y8828 = ~n20787 ;
  assign y8829 = ~1'b0 ;
  assign y8830 = ~1'b0 ;
  assign y8831 = n20788 ;
  assign y8832 = ~1'b0 ;
  assign y8833 = ~1'b0 ;
  assign y8834 = n20792 ;
  assign y8835 = n20798 ;
  assign y8836 = ~n20799 ;
  assign y8837 = ~n20803 ;
  assign y8838 = ~n20807 ;
  assign y8839 = ~n20810 ;
  assign y8840 = ~n20811 ;
  assign y8841 = ~n20813 ;
  assign y8842 = n20815 ;
  assign y8843 = ~n20817 ;
  assign y8844 = ~n20819 ;
  assign y8845 = ~1'b0 ;
  assign y8846 = ~n20820 ;
  assign y8847 = n20826 ;
  assign y8848 = n15985 ;
  assign y8849 = n20827 ;
  assign y8850 = ~n20828 ;
  assign y8851 = n20829 ;
  assign y8852 = n20831 ;
  assign y8853 = ~n20834 ;
  assign y8854 = ~n20836 ;
  assign y8855 = ~1'b0 ;
  assign y8856 = ~1'b0 ;
  assign y8857 = ~n20840 ;
  assign y8858 = ~1'b0 ;
  assign y8859 = ~1'b0 ;
  assign y8860 = n8058 ;
  assign y8861 = n20841 ;
  assign y8862 = ~n20844 ;
  assign y8863 = ~n20848 ;
  assign y8864 = ~n20857 ;
  assign y8865 = n20858 ;
  assign y8866 = n20859 ;
  assign y8867 = n20861 ;
  assign y8868 = ~n9133 ;
  assign y8869 = ~n20862 ;
  assign y8870 = ~n20867 ;
  assign y8871 = ~n20871 ;
  assign y8872 = ~1'b0 ;
  assign y8873 = ~n20873 ;
  assign y8874 = ~1'b0 ;
  assign y8875 = ~1'b0 ;
  assign y8876 = ~n20878 ;
  assign y8877 = ~1'b0 ;
  assign y8878 = n20879 ;
  assign y8879 = n20881 ;
  assign y8880 = ~n20884 ;
  assign y8881 = ~1'b0 ;
  assign y8882 = n20891 ;
  assign y8883 = n20897 ;
  assign y8884 = ~1'b0 ;
  assign y8885 = n20898 ;
  assign y8886 = n20900 ;
  assign y8887 = ~n20901 ;
  assign y8888 = n20906 ;
  assign y8889 = ~1'b0 ;
  assign y8890 = n20913 ;
  assign y8891 = n20916 ;
  assign y8892 = ~n20920 ;
  assign y8893 = ~1'b0 ;
  assign y8894 = ~n20924 ;
  assign y8895 = n20928 ;
  assign y8896 = ~n20929 ;
  assign y8897 = n20930 ;
  assign y8898 = ~n20936 ;
  assign y8899 = n20940 ;
  assign y8900 = n20942 ;
  assign y8901 = ~n20948 ;
  assign y8902 = ~n20949 ;
  assign y8903 = ~1'b0 ;
  assign y8904 = 1'b0 ;
  assign y8905 = n20951 ;
  assign y8906 = ~n20954 ;
  assign y8907 = ~n20962 ;
  assign y8908 = n20963 ;
  assign y8909 = ~1'b0 ;
  assign y8910 = n20967 ;
  assign y8911 = ~n20971 ;
  assign y8912 = ~1'b0 ;
  assign y8913 = ~1'b0 ;
  assign y8914 = ~1'b0 ;
  assign y8915 = n20975 ;
  assign y8916 = n20977 ;
  assign y8917 = n20978 ;
  assign y8918 = ~1'b0 ;
  assign y8919 = ~n20982 ;
  assign y8920 = ~n20986 ;
  assign y8921 = ~1'b0 ;
  assign y8922 = n20989 ;
  assign y8923 = ~n20992 ;
  assign y8924 = ~n20997 ;
  assign y8925 = ~n20998 ;
  assign y8926 = n21002 ;
  assign y8927 = n21003 ;
  assign y8928 = n21004 ;
  assign y8929 = n21006 ;
  assign y8930 = n21007 ;
  assign y8931 = ~1'b0 ;
  assign y8932 = ~1'b0 ;
  assign y8933 = n21009 ;
  assign y8934 = n21011 ;
  assign y8935 = ~1'b0 ;
  assign y8936 = ~1'b0 ;
  assign y8937 = ~1'b0 ;
  assign y8938 = ~1'b0 ;
  assign y8939 = ~n8993 ;
  assign y8940 = ~n21013 ;
  assign y8941 = n21019 ;
  assign y8942 = ~n21027 ;
  assign y8943 = n21031 ;
  assign y8944 = n21038 ;
  assign y8945 = ~1'b0 ;
  assign y8946 = ~1'b0 ;
  assign y8947 = ~n21042 ;
  assign y8948 = n21043 ;
  assign y8949 = ~n21044 ;
  assign y8950 = ~n21046 ;
  assign y8951 = ~n21059 ;
  assign y8952 = n21065 ;
  assign y8953 = ~n21070 ;
  assign y8954 = ~n21073 ;
  assign y8955 = n21074 ;
  assign y8956 = ~1'b0 ;
  assign y8957 = ~1'b0 ;
  assign y8958 = n21078 ;
  assign y8959 = n21081 ;
  assign y8960 = ~n21086 ;
  assign y8961 = ~n21087 ;
  assign y8962 = n21090 ;
  assign y8963 = ~1'b0 ;
  assign y8964 = n21095 ;
  assign y8965 = n2201 ;
  assign y8966 = ~1'b0 ;
  assign y8967 = n1158 ;
  assign y8968 = n21098 ;
  assign y8969 = ~n21110 ;
  assign y8970 = ~n21114 ;
  assign y8971 = ~n21116 ;
  assign y8972 = n21118 ;
  assign y8973 = n21125 ;
  assign y8974 = ~1'b0 ;
  assign y8975 = n21127 ;
  assign y8976 = ~n21129 ;
  assign y8977 = ~n21132 ;
  assign y8978 = ~1'b0 ;
  assign y8979 = n21137 ;
  assign y8980 = ~1'b0 ;
  assign y8981 = n21140 ;
  assign y8982 = ~1'b0 ;
  assign y8983 = ~n21141 ;
  assign y8984 = ~n21143 ;
  assign y8985 = ~n21144 ;
  assign y8986 = ~n21145 ;
  assign y8987 = ~n21147 ;
  assign y8988 = ~1'b0 ;
  assign y8989 = n21150 ;
  assign y8990 = n12408 ;
  assign y8991 = n21152 ;
  assign y8992 = n21153 ;
  assign y8993 = n21154 ;
  assign y8994 = ~1'b0 ;
  assign y8995 = n21156 ;
  assign y8996 = n21158 ;
  assign y8997 = n21162 ;
  assign y8998 = n21163 ;
  assign y8999 = ~1'b0 ;
  assign y9000 = n21167 ;
  assign y9001 = ~n21169 ;
  assign y9002 = ~n21172 ;
  assign y9003 = ~1'b0 ;
  assign y9004 = ~n21174 ;
  assign y9005 = n8459 ;
  assign y9006 = ~n21176 ;
  assign y9007 = ~1'b0 ;
  assign y9008 = ~1'b0 ;
  assign y9009 = n21179 ;
  assign y9010 = n21180 ;
  assign y9011 = ~n21185 ;
  assign y9012 = ~1'b0 ;
  assign y9013 = ~n21186 ;
  assign y9014 = ~n21187 ;
  assign y9015 = ~1'b0 ;
  assign y9016 = ~1'b0 ;
  assign y9017 = ~1'b0 ;
  assign y9018 = ~n21189 ;
  assign y9019 = ~1'b0 ;
  assign y9020 = n21191 ;
  assign y9021 = ~n21194 ;
  assign y9022 = n21199 ;
  assign y9023 = n21204 ;
  assign y9024 = ~n21207 ;
  assign y9025 = n21208 ;
  assign y9026 = ~n21212 ;
  assign y9027 = n21214 ;
  assign y9028 = n21218 ;
  assign y9029 = n21219 ;
  assign y9030 = n21223 ;
  assign y9031 = ~1'b0 ;
  assign y9032 = ~1'b0 ;
  assign y9033 = ~n21225 ;
  assign y9034 = n21232 ;
  assign y9035 = ~1'b0 ;
  assign y9036 = ~1'b0 ;
  assign y9037 = ~n21236 ;
  assign y9038 = ~1'b0 ;
  assign y9039 = ~n21237 ;
  assign y9040 = n21238 ;
  assign y9041 = ~n21240 ;
  assign y9042 = n21243 ;
  assign y9043 = ~1'b0 ;
  assign y9044 = n21244 ;
  assign y9045 = ~1'b0 ;
  assign y9046 = ~n21247 ;
  assign y9047 = n21249 ;
  assign y9048 = n21250 ;
  assign y9049 = n21251 ;
  assign y9050 = ~n21260 ;
  assign y9051 = ~1'b0 ;
  assign y9052 = ~1'b0 ;
  assign y9053 = n21261 ;
  assign y9054 = ~1'b0 ;
  assign y9055 = n21262 ;
  assign y9056 = ~1'b0 ;
  assign y9057 = ~n21266 ;
  assign y9058 = n21275 ;
  assign y9059 = ~1'b0 ;
  assign y9060 = ~1'b0 ;
  assign y9061 = n21276 ;
  assign y9062 = ~n21279 ;
  assign y9063 = ~n21280 ;
  assign y9064 = n21281 ;
  assign y9065 = ~n21285 ;
  assign y9066 = n2561 ;
  assign y9067 = ~1'b0 ;
  assign y9068 = ~n21288 ;
  assign y9069 = n21289 ;
  assign y9070 = n21290 ;
  assign y9071 = 1'b0 ;
  assign y9072 = n21291 ;
  assign y9073 = ~1'b0 ;
  assign y9074 = ~n21292 ;
  assign y9075 = n21294 ;
  assign y9076 = n21295 ;
  assign y9077 = ~n21298 ;
  assign y9078 = n21300 ;
  assign y9079 = ~n21302 ;
  assign y9080 = n21303 ;
  assign y9081 = n21304 ;
  assign y9082 = ~n21305 ;
  assign y9083 = ~n21306 ;
  assign y9084 = ~n21311 ;
  assign y9085 = ~1'b0 ;
  assign y9086 = ~1'b0 ;
  assign y9087 = ~n3199 ;
  assign y9088 = n21312 ;
  assign y9089 = n21313 ;
  assign y9090 = ~1'b0 ;
  assign y9091 = ~n21317 ;
  assign y9092 = ~1'b0 ;
  assign y9093 = n21318 ;
  assign y9094 = n21321 ;
  assign y9095 = n21323 ;
  assign y9096 = ~n21326 ;
  assign y9097 = ~n21328 ;
  assign y9098 = ~n21331 ;
  assign y9099 = n21332 ;
  assign y9100 = ~n21340 ;
  assign y9101 = ~n21352 ;
  assign y9102 = 1'b0 ;
  assign y9103 = ~n21353 ;
  assign y9104 = ~1'b0 ;
  assign y9105 = n21355 ;
  assign y9106 = ~n21356 ;
  assign y9107 = ~n21357 ;
  assign y9108 = n21359 ;
  assign y9109 = ~1'b0 ;
  assign y9110 = ~1'b0 ;
  assign y9111 = n21369 ;
  assign y9112 = 1'b0 ;
  assign y9113 = n21372 ;
  assign y9114 = ~n21375 ;
  assign y9115 = ~1'b0 ;
  assign y9116 = n21379 ;
  assign y9117 = ~n21383 ;
  assign y9118 = n21384 ;
  assign y9119 = n21386 ;
  assign y9120 = ~n21394 ;
  assign y9121 = n12834 ;
  assign y9122 = ~n21395 ;
  assign y9123 = n21398 ;
  assign y9124 = n21400 ;
  assign y9125 = n21402 ;
  assign y9126 = ~1'b0 ;
  assign y9127 = ~n21404 ;
  assign y9128 = ~n21406 ;
  assign y9129 = n5542 ;
  assign y9130 = ~1'b0 ;
  assign y9131 = n21407 ;
  assign y9132 = ~n21409 ;
  assign y9133 = ~1'b0 ;
  assign y9134 = ~n1239 ;
  assign y9135 = ~n21410 ;
  assign y9136 = n21415 ;
  assign y9137 = ~n21418 ;
  assign y9138 = ~n21420 ;
  assign y9139 = n21421 ;
  assign y9140 = n21426 ;
  assign y9141 = n21432 ;
  assign y9142 = ~n21437 ;
  assign y9143 = ~n21439 ;
  assign y9144 = ~n21441 ;
  assign y9145 = n21442 ;
  assign y9146 = n21443 ;
  assign y9147 = n21445 ;
  assign y9148 = ~n21448 ;
  assign y9149 = ~1'b0 ;
  assign y9150 = n21451 ;
  assign y9151 = ~n21454 ;
  assign y9152 = ~1'b0 ;
  assign y9153 = n21455 ;
  assign y9154 = ~n21459 ;
  assign y9155 = n305 ;
  assign y9156 = ~1'b0 ;
  assign y9157 = ~n21465 ;
  assign y9158 = ~1'b0 ;
  assign y9159 = ~n21469 ;
  assign y9160 = ~n21471 ;
  assign y9161 = ~1'b0 ;
  assign y9162 = ~n21472 ;
  assign y9163 = ~n21473 ;
  assign y9164 = n21476 ;
  assign y9165 = ~1'b0 ;
  assign y9166 = ~n21478 ;
  assign y9167 = ~n21479 ;
  assign y9168 = n21480 ;
  assign y9169 = ~1'b0 ;
  assign y9170 = n21483 ;
  assign y9171 = n21486 ;
  assign y9172 = ~1'b0 ;
  assign y9173 = n21489 ;
  assign y9174 = n14587 ;
  assign y9175 = ~1'b0 ;
  assign y9176 = n21496 ;
  assign y9177 = n21499 ;
  assign y9178 = ~n21500 ;
  assign y9179 = n21501 ;
  assign y9180 = ~1'b0 ;
  assign y9181 = ~n21502 ;
  assign y9182 = ~n21503 ;
  assign y9183 = ~n13982 ;
  assign y9184 = n21512 ;
  assign y9185 = ~1'b0 ;
  assign y9186 = ~1'b0 ;
  assign y9187 = n21513 ;
  assign y9188 = n21517 ;
  assign y9189 = ~n21519 ;
  assign y9190 = n21522 ;
  assign y9191 = n21529 ;
  assign y9192 = ~n21530 ;
  assign y9193 = ~1'b0 ;
  assign y9194 = ~1'b0 ;
  assign y9195 = ~1'b0 ;
  assign y9196 = n21534 ;
  assign y9197 = ~n21538 ;
  assign y9198 = ~1'b0 ;
  assign y9199 = n18327 ;
  assign y9200 = ~x61 ;
  assign y9201 = ~1'b0 ;
  assign y9202 = ~n21547 ;
  assign y9203 = ~1'b0 ;
  assign y9204 = n21553 ;
  assign y9205 = n21558 ;
  assign y9206 = n21559 ;
  assign y9207 = ~n21563 ;
  assign y9208 = ~n21567 ;
  assign y9209 = ~1'b0 ;
  assign y9210 = ~n15649 ;
  assign y9211 = n21569 ;
  assign y9212 = n21571 ;
  assign y9213 = ~n21577 ;
  assign y9214 = ~n21578 ;
  assign y9215 = n21586 ;
  assign y9216 = ~n21587 ;
  assign y9217 = ~n21593 ;
  assign y9218 = n21595 ;
  assign y9219 = n21597 ;
  assign y9220 = ~n21598 ;
  assign y9221 = ~n21599 ;
  assign y9222 = ~1'b0 ;
  assign y9223 = ~1'b0 ;
  assign y9224 = n21601 ;
  assign y9225 = ~1'b0 ;
  assign y9226 = n21605 ;
  assign y9227 = ~n21607 ;
  assign y9228 = ~n21610 ;
  assign y9229 = ~1'b0 ;
  assign y9230 = ~n21612 ;
  assign y9231 = ~n21614 ;
  assign y9232 = n21618 ;
  assign y9233 = ~n21621 ;
  assign y9234 = n21623 ;
  assign y9235 = ~n21624 ;
  assign y9236 = n21625 ;
  assign y9237 = ~1'b0 ;
  assign y9238 = ~1'b0 ;
  assign y9239 = ~n21632 ;
  assign y9240 = n21635 ;
  assign y9241 = ~n17994 ;
  assign y9242 = ~n21639 ;
  assign y9243 = ~n21641 ;
  assign y9244 = n21644 ;
  assign y9245 = ~n21647 ;
  assign y9246 = ~n21651 ;
  assign y9247 = ~n21658 ;
  assign y9248 = ~n21660 ;
  assign y9249 = ~1'b0 ;
  assign y9250 = n7777 ;
  assign y9251 = n21661 ;
  assign y9252 = ~1'b0 ;
  assign y9253 = ~n21662 ;
  assign y9254 = ~n21664 ;
  assign y9255 = ~n21666 ;
  assign y9256 = n21667 ;
  assign y9257 = ~n21669 ;
  assign y9258 = ~1'b0 ;
  assign y9259 = ~1'b0 ;
  assign y9260 = ~n21673 ;
  assign y9261 = n21678 ;
  assign y9262 = ~n21683 ;
  assign y9263 = ~n21690 ;
  assign y9264 = ~n21692 ;
  assign y9265 = ~n21694 ;
  assign y9266 = n21699 ;
  assign y9267 = n21700 ;
  assign y9268 = ~1'b0 ;
  assign y9269 = ~n21703 ;
  assign y9270 = n21706 ;
  assign y9271 = ~n8122 ;
  assign y9272 = ~1'b0 ;
  assign y9273 = ~n21730 ;
  assign y9274 = ~1'b0 ;
  assign y9275 = n21736 ;
  assign y9276 = ~1'b0 ;
  assign y9277 = ~x132 ;
  assign y9278 = ~n21742 ;
  assign y9279 = ~n7607 ;
  assign y9280 = ~n21745 ;
  assign y9281 = ~n21748 ;
  assign y9282 = ~n21752 ;
  assign y9283 = ~n21759 ;
  assign y9284 = ~n21762 ;
  assign y9285 = n21766 ;
  assign y9286 = n21776 ;
  assign y9287 = ~1'b0 ;
  assign y9288 = ~n21779 ;
  assign y9289 = n21786 ;
  assign y9290 = ~1'b0 ;
  assign y9291 = n21789 ;
  assign y9292 = ~n21791 ;
  assign y9293 = ~1'b0 ;
  assign y9294 = ~1'b0 ;
  assign y9295 = n21792 ;
  assign y9296 = n12080 ;
  assign y9297 = ~n21794 ;
  assign y9298 = n21795 ;
  assign y9299 = n21797 ;
  assign y9300 = ~n21800 ;
  assign y9301 = ~1'b0 ;
  assign y9302 = ~n21803 ;
  assign y9303 = ~1'b0 ;
  assign y9304 = n21805 ;
  assign y9305 = n21806 ;
  assign y9306 = n21807 ;
  assign y9307 = n21809 ;
  assign y9308 = ~1'b0 ;
  assign y9309 = ~n21812 ;
  assign y9310 = ~1'b0 ;
  assign y9311 = 1'b0 ;
  assign y9312 = n21813 ;
  assign y9313 = n21818 ;
  assign y9314 = ~n21820 ;
  assign y9315 = ~1'b0 ;
  assign y9316 = ~1'b0 ;
  assign y9317 = x30 ;
  assign y9318 = ~n21824 ;
  assign y9319 = 1'b0 ;
  assign y9320 = n21826 ;
  assign y9321 = n21827 ;
  assign y9322 = n21828 ;
  assign y9323 = n21829 ;
  assign y9324 = n21835 ;
  assign y9325 = ~n21837 ;
  assign y9326 = n21841 ;
  assign y9327 = ~n21842 ;
  assign y9328 = n21844 ;
  assign y9329 = ~1'b0 ;
  assign y9330 = n21847 ;
  assign y9331 = ~1'b0 ;
  assign y9332 = ~n21848 ;
  assign y9333 = ~1'b0 ;
  assign y9334 = n21855 ;
  assign y9335 = ~n5584 ;
  assign y9336 = ~n21856 ;
  assign y9337 = ~1'b0 ;
  assign y9338 = n21858 ;
  assign y9339 = n21860 ;
  assign y9340 = ~n21863 ;
  assign y9341 = ~n21867 ;
  assign y9342 = n21870 ;
  assign y9343 = ~1'b0 ;
  assign y9344 = n21872 ;
  assign y9345 = ~n21882 ;
  assign y9346 = ~1'b0 ;
  assign y9347 = ~n21884 ;
  assign y9348 = ~n21886 ;
  assign y9349 = ~n21888 ;
  assign y9350 = ~1'b0 ;
  assign y9351 = ~n21890 ;
  assign y9352 = ~1'b0 ;
  assign y9353 = ~n21892 ;
  assign y9354 = n21893 ;
  assign y9355 = ~1'b0 ;
  assign y9356 = n21896 ;
  assign y9357 = ~1'b0 ;
  assign y9358 = n21897 ;
  assign y9359 = ~1'b0 ;
  assign y9360 = ~n21900 ;
  assign y9361 = 1'b0 ;
  assign y9362 = ~n21903 ;
  assign y9363 = ~n2437 ;
  assign y9364 = ~n21908 ;
  assign y9365 = n21913 ;
  assign y9366 = ~1'b0 ;
  assign y9367 = n21914 ;
  assign y9368 = ~n21917 ;
  assign y9369 = n21919 ;
  assign y9370 = n21920 ;
  assign y9371 = n21923 ;
  assign y9372 = ~n21924 ;
  assign y9373 = n21925 ;
  assign y9374 = ~1'b0 ;
  assign y9375 = n21929 ;
  assign y9376 = ~1'b0 ;
  assign y9377 = ~n21935 ;
  assign y9378 = ~n21937 ;
  assign y9379 = n21938 ;
  assign y9380 = ~1'b0 ;
  assign y9381 = n21939 ;
  assign y9382 = ~1'b0 ;
  assign y9383 = ~n21941 ;
  assign y9384 = ~n21943 ;
  assign y9385 = ~1'b0 ;
  assign y9386 = ~1'b0 ;
  assign y9387 = ~n21946 ;
  assign y9388 = n21948 ;
  assign y9389 = ~1'b0 ;
  assign y9390 = ~n21955 ;
  assign y9391 = n21957 ;
  assign y9392 = ~n21972 ;
  assign y9393 = n21974 ;
  assign y9394 = ~n21975 ;
  assign y9395 = ~n21980 ;
  assign y9396 = n21983 ;
  assign y9397 = ~n21984 ;
  assign y9398 = ~n21985 ;
  assign y9399 = n21986 ;
  assign y9400 = n21992 ;
  assign y9401 = ~n21997 ;
  assign y9402 = ~n22001 ;
  assign y9403 = ~n22004 ;
  assign y9404 = n22006 ;
  assign y9405 = ~n22010 ;
  assign y9406 = n22011 ;
  assign y9407 = n22012 ;
  assign y9408 = ~1'b0 ;
  assign y9409 = ~1'b0 ;
  assign y9410 = ~1'b0 ;
  assign y9411 = n22014 ;
  assign y9412 = n22015 ;
  assign y9413 = n4977 ;
  assign y9414 = ~n22019 ;
  assign y9415 = ~n13020 ;
  assign y9416 = ~1'b0 ;
  assign y9417 = ~1'b0 ;
  assign y9418 = ~n22021 ;
  assign y9419 = ~n22023 ;
  assign y9420 = ~1'b0 ;
  assign y9421 = ~1'b0 ;
  assign y9422 = ~n20845 ;
  assign y9423 = ~n22028 ;
  assign y9424 = ~1'b0 ;
  assign y9425 = n22030 ;
  assign y9426 = ~1'b0 ;
  assign y9427 = n22039 ;
  assign y9428 = ~n22041 ;
  assign y9429 = ~n22043 ;
  assign y9430 = n22044 ;
  assign y9431 = ~n22046 ;
  assign y9432 = ~n22050 ;
  assign y9433 = n21822 ;
  assign y9434 = n22053 ;
  assign y9435 = ~n22057 ;
  assign y9436 = ~n22065 ;
  assign y9437 = n22075 ;
  assign y9438 = ~n22076 ;
  assign y9439 = ~n22083 ;
  assign y9440 = ~n22086 ;
  assign y9441 = n22089 ;
  assign y9442 = ~n22101 ;
  assign y9443 = n22104 ;
  assign y9444 = ~n22105 ;
  assign y9445 = n22107 ;
  assign y9446 = n22111 ;
  assign y9447 = ~n22113 ;
  assign y9448 = ~1'b0 ;
  assign y9449 = ~n22116 ;
  assign y9450 = ~n22117 ;
  assign y9451 = ~n22119 ;
  assign y9452 = n4489 ;
  assign y9453 = ~n22120 ;
  assign y9454 = ~n22125 ;
  assign y9455 = ~1'b0 ;
  assign y9456 = n22129 ;
  assign y9457 = ~n22130 ;
  assign y9458 = n22131 ;
  assign y9459 = ~n22136 ;
  assign y9460 = ~n22137 ;
  assign y9461 = ~1'b0 ;
  assign y9462 = n22141 ;
  assign y9463 = ~1'b0 ;
  assign y9464 = n22144 ;
  assign y9465 = ~n22145 ;
  assign y9466 = ~n22146 ;
  assign y9467 = ~n22148 ;
  assign y9468 = ~n22154 ;
  assign y9469 = n5302 ;
  assign y9470 = n22155 ;
  assign y9471 = ~1'b0 ;
  assign y9472 = n22156 ;
  assign y9473 = ~n22158 ;
  assign y9474 = ~n22161 ;
  assign y9475 = ~1'b0 ;
  assign y9476 = ~n22162 ;
  assign y9477 = n22165 ;
  assign y9478 = n22166 ;
  assign y9479 = n22174 ;
  assign y9480 = ~n22179 ;
  assign y9481 = n22180 ;
  assign y9482 = ~n22182 ;
  assign y9483 = ~1'b0 ;
  assign y9484 = 1'b0 ;
  assign y9485 = ~n22193 ;
  assign y9486 = n22197 ;
  assign y9487 = n17219 ;
  assign y9488 = ~n22199 ;
  assign y9489 = ~1'b0 ;
  assign y9490 = n22202 ;
  assign y9491 = n22207 ;
  assign y9492 = n22208 ;
  assign y9493 = ~1'b0 ;
  assign y9494 = ~n22212 ;
  assign y9495 = n22213 ;
  assign y9496 = ~n22217 ;
  assign y9497 = ~n22218 ;
  assign y9498 = ~n22221 ;
  assign y9499 = n22223 ;
  assign y9500 = ~1'b0 ;
  assign y9501 = n22225 ;
  assign y9502 = n22226 ;
  assign y9503 = 1'b0 ;
  assign y9504 = n22228 ;
  assign y9505 = ~n22229 ;
  assign y9506 = n22231 ;
  assign y9507 = n22232 ;
  assign y9508 = n22235 ;
  assign y9509 = ~1'b0 ;
  assign y9510 = ~n22237 ;
  assign y9511 = ~n22240 ;
  assign y9512 = ~1'b0 ;
  assign y9513 = ~1'b0 ;
  assign y9514 = n22243 ;
  assign y9515 = ~1'b0 ;
  assign y9516 = n22255 ;
  assign y9517 = ~n22258 ;
  assign y9518 = n22259 ;
  assign y9519 = n22262 ;
  assign y9520 = n22263 ;
  assign y9521 = ~1'b0 ;
  assign y9522 = ~n22265 ;
  assign y9523 = ~n22266 ;
  assign y9524 = ~1'b0 ;
  assign y9525 = n22270 ;
  assign y9526 = ~n22271 ;
  assign y9527 = ~n22272 ;
  assign y9528 = ~n22275 ;
  assign y9529 = ~n22278 ;
  assign y9530 = ~1'b0 ;
  assign y9531 = n22283 ;
  assign y9532 = n22288 ;
  assign y9533 = ~n22292 ;
  assign y9534 = ~n22293 ;
  assign y9535 = n10092 ;
  assign y9536 = 1'b0 ;
  assign y9537 = n22297 ;
  assign y9538 = n22299 ;
  assign y9539 = n22300 ;
  assign y9540 = n22301 ;
  assign y9541 = ~n12002 ;
  assign y9542 = ~n21251 ;
  assign y9543 = n22303 ;
  assign y9544 = ~1'b0 ;
  assign y9545 = ~1'b0 ;
  assign y9546 = ~n5468 ;
  assign y9547 = ~n22304 ;
  assign y9548 = n22310 ;
  assign y9549 = ~n22311 ;
  assign y9550 = n22315 ;
  assign y9551 = n22319 ;
  assign y9552 = ~n22320 ;
  assign y9553 = ~n22322 ;
  assign y9554 = n22324 ;
  assign y9555 = ~n22331 ;
  assign y9556 = n22334 ;
  assign y9557 = n22336 ;
  assign y9558 = ~n22338 ;
  assign y9559 = n22344 ;
  assign y9560 = ~n22346 ;
  assign y9561 = ~n22349 ;
  assign y9562 = ~n22350 ;
  assign y9563 = ~1'b0 ;
  assign y9564 = ~1'b0 ;
  assign y9565 = ~1'b0 ;
  assign y9566 = ~1'b0 ;
  assign y9567 = ~1'b0 ;
  assign y9568 = ~n22355 ;
  assign y9569 = ~n22356 ;
  assign y9570 = ~1'b0 ;
  assign y9571 = ~1'b0 ;
  assign y9572 = ~n22358 ;
  assign y9573 = ~1'b0 ;
  assign y9574 = n22363 ;
  assign y9575 = ~1'b0 ;
  assign y9576 = ~1'b0 ;
  assign y9577 = ~n22364 ;
  assign y9578 = ~1'b0 ;
  assign y9579 = n22372 ;
  assign y9580 = n22376 ;
  assign y9581 = n22381 ;
  assign y9582 = n22383 ;
  assign y9583 = ~n22385 ;
  assign y9584 = ~n22386 ;
  assign y9585 = n22387 ;
  assign y9586 = n22388 ;
  assign y9587 = 1'b0 ;
  assign y9588 = n22393 ;
  assign y9589 = n22399 ;
  assign y9590 = ~1'b0 ;
  assign y9591 = n22402 ;
  assign y9592 = ~n22404 ;
  assign y9593 = n22406 ;
  assign y9594 = ~1'b0 ;
  assign y9595 = n22413 ;
  assign y9596 = n22418 ;
  assign y9597 = ~1'b0 ;
  assign y9598 = ~1'b0 ;
  assign y9599 = n22421 ;
  assign y9600 = ~n22422 ;
  assign y9601 = 1'b0 ;
  assign y9602 = ~n22425 ;
  assign y9603 = n22426 ;
  assign y9604 = ~1'b0 ;
  assign y9605 = ~n22428 ;
  assign y9606 = ~1'b0 ;
  assign y9607 = ~1'b0 ;
  assign y9608 = n22431 ;
  assign y9609 = ~n842 ;
  assign y9610 = ~n22436 ;
  assign y9611 = ~n22441 ;
  assign y9612 = ~1'b0 ;
  assign y9613 = ~1'b0 ;
  assign y9614 = ~n22444 ;
  assign y9615 = n22446 ;
  assign y9616 = ~n22449 ;
  assign y9617 = ~1'b0 ;
  assign y9618 = ~1'b0 ;
  assign y9619 = ~n22450 ;
  assign y9620 = ~n22454 ;
  assign y9621 = ~1'b0 ;
  assign y9622 = ~n22457 ;
  assign y9623 = n22459 ;
  assign y9624 = 1'b0 ;
  assign y9625 = n22463 ;
  assign y9626 = n22465 ;
  assign y9627 = ~1'b0 ;
  assign y9628 = ~n22467 ;
  assign y9629 = n22470 ;
  assign y9630 = n22471 ;
  assign y9631 = ~1'b0 ;
  assign y9632 = ~n16810 ;
  assign y9633 = ~n22476 ;
  assign y9634 = n22479 ;
  assign y9635 = ~1'b0 ;
  assign y9636 = n22481 ;
  assign y9637 = n22482 ;
  assign y9638 = n22483 ;
  assign y9639 = ~1'b0 ;
  assign y9640 = ~n22484 ;
  assign y9641 = ~n22489 ;
  assign y9642 = n22493 ;
  assign y9643 = ~n22494 ;
  assign y9644 = ~n22496 ;
  assign y9645 = n22499 ;
  assign y9646 = ~1'b0 ;
  assign y9647 = 1'b0 ;
  assign y9648 = n22509 ;
  assign y9649 = n22511 ;
  assign y9650 = ~1'b0 ;
  assign y9651 = ~1'b0 ;
  assign y9652 = ~n22512 ;
  assign y9653 = n22515 ;
  assign y9654 = n22518 ;
  assign y9655 = n22519 ;
  assign y9656 = ~1'b0 ;
  assign y9657 = ~n22521 ;
  assign y9658 = n22522 ;
  assign y9659 = ~n22524 ;
  assign y9660 = n22527 ;
  assign y9661 = n22528 ;
  assign y9662 = ~n22531 ;
  assign y9663 = ~1'b0 ;
  assign y9664 = ~n22534 ;
  assign y9665 = ~n8665 ;
  assign y9666 = ~1'b0 ;
  assign y9667 = ~n1401 ;
  assign y9668 = n22536 ;
  assign y9669 = ~n22539 ;
  assign y9670 = ~1'b0 ;
  assign y9671 = ~n22540 ;
  assign y9672 = ~n22541 ;
  assign y9673 = ~n22542 ;
  assign y9674 = ~n22544 ;
  assign y9675 = ~n15462 ;
  assign y9676 = ~n22547 ;
  assign y9677 = n22548 ;
  assign y9678 = ~n22550 ;
  assign y9679 = ~n22552 ;
  assign y9680 = n22554 ;
  assign y9681 = ~n22556 ;
  assign y9682 = ~1'b0 ;
  assign y9683 = n22557 ;
  assign y9684 = ~1'b0 ;
  assign y9685 = ~n22558 ;
  assign y9686 = ~n22560 ;
  assign y9687 = ~n22562 ;
  assign y9688 = ~1'b0 ;
  assign y9689 = 1'b0 ;
  assign y9690 = ~1'b0 ;
  assign y9691 = ~n22576 ;
  assign y9692 = 1'b0 ;
  assign y9693 = ~n22577 ;
  assign y9694 = n22578 ;
  assign y9695 = n22579 ;
  assign y9696 = ~n22580 ;
  assign y9697 = ~1'b0 ;
  assign y9698 = ~n22581 ;
  assign y9699 = n4630 ;
  assign y9700 = ~1'b0 ;
  assign y9701 = n22584 ;
  assign y9702 = ~n22588 ;
  assign y9703 = ~1'b0 ;
  assign y9704 = n22590 ;
  assign y9705 = ~1'b0 ;
  assign y9706 = ~1'b0 ;
  assign y9707 = n22591 ;
  assign y9708 = ~n22596 ;
  assign y9709 = n22601 ;
  assign y9710 = n22602 ;
  assign y9711 = n22608 ;
  assign y9712 = ~n22612 ;
  assign y9713 = n22613 ;
  assign y9714 = n22614 ;
  assign y9715 = n22615 ;
  assign y9716 = n22618 ;
  assign y9717 = ~n22622 ;
  assign y9718 = ~n22624 ;
  assign y9719 = ~1'b0 ;
  assign y9720 = n22627 ;
  assign y9721 = ~n22631 ;
  assign y9722 = ~n22633 ;
  assign y9723 = n22634 ;
  assign y9724 = n22636 ;
  assign y9725 = n22638 ;
  assign y9726 = ~n22641 ;
  assign y9727 = n22650 ;
  assign y9728 = ~n22652 ;
  assign y9729 = n22656 ;
  assign y9730 = ~n22662 ;
  assign y9731 = ~1'b0 ;
  assign y9732 = n22672 ;
  assign y9733 = n22676 ;
  assign y9734 = ~1'b0 ;
  assign y9735 = n22679 ;
  assign y9736 = ~1'b0 ;
  assign y9737 = ~n22680 ;
  assign y9738 = ~1'b0 ;
  assign y9739 = ~n22683 ;
  assign y9740 = n22684 ;
  assign y9741 = ~1'b0 ;
  assign y9742 = ~n22686 ;
  assign y9743 = ~1'b0 ;
  assign y9744 = ~1'b0 ;
  assign y9745 = n22690 ;
  assign y9746 = ~1'b0 ;
  assign y9747 = n22695 ;
  assign y9748 = ~n22698 ;
  assign y9749 = ~n22700 ;
  assign y9750 = ~1'b0 ;
  assign y9751 = ~n22701 ;
  assign y9752 = n22702 ;
  assign y9753 = ~n22703 ;
  assign y9754 = n22707 ;
  assign y9755 = ~n22711 ;
  assign y9756 = ~n22714 ;
  assign y9757 = ~1'b0 ;
  assign y9758 = ~n22718 ;
  assign y9759 = ~n22721 ;
  assign y9760 = n22723 ;
  assign y9761 = ~1'b0 ;
  assign y9762 = ~n22726 ;
  assign y9763 = n22728 ;
  assign y9764 = n11053 ;
  assign y9765 = ~n22730 ;
  assign y9766 = ~1'b0 ;
  assign y9767 = ~n22732 ;
  assign y9768 = n22736 ;
  assign y9769 = ~1'b0 ;
  assign y9770 = n22737 ;
  assign y9771 = ~n7401 ;
  assign y9772 = n22739 ;
  assign y9773 = ~1'b0 ;
  assign y9774 = ~1'b0 ;
  assign y9775 = ~1'b0 ;
  assign y9776 = n22748 ;
  assign y9777 = ~n22752 ;
  assign y9778 = ~n22755 ;
  assign y9779 = n4264 ;
  assign y9780 = n22756 ;
  assign y9781 = n17708 ;
  assign y9782 = ~n22757 ;
  assign y9783 = ~1'b0 ;
  assign y9784 = n22761 ;
  assign y9785 = n22762 ;
  assign y9786 = ~1'b0 ;
  assign y9787 = ~n22769 ;
  assign y9788 = ~1'b0 ;
  assign y9789 = ~1'b0 ;
  assign y9790 = ~n22770 ;
  assign y9791 = ~1'b0 ;
  assign y9792 = ~n22774 ;
  assign y9793 = ~1'b0 ;
  assign y9794 = ~1'b0 ;
  assign y9795 = ~n22776 ;
  assign y9796 = ~1'b0 ;
  assign y9797 = ~n22777 ;
  assign y9798 = n22783 ;
  assign y9799 = ~1'b0 ;
  assign y9800 = ~n22793 ;
  assign y9801 = 1'b0 ;
  assign y9802 = ~n22797 ;
  assign y9803 = ~n22799 ;
  assign y9804 = ~n22802 ;
  assign y9805 = ~1'b0 ;
  assign y9806 = ~n22804 ;
  assign y9807 = n22807 ;
  assign y9808 = ~1'b0 ;
  assign y9809 = ~1'b0 ;
  assign y9810 = ~1'b0 ;
  assign y9811 = ~n2460 ;
  assign y9812 = ~n22808 ;
  assign y9813 = n22810 ;
  assign y9814 = n22812 ;
  assign y9815 = ~1'b0 ;
  assign y9816 = ~1'b0 ;
  assign y9817 = n22819 ;
  assign y9818 = ~1'b0 ;
  assign y9819 = ~1'b0 ;
  assign y9820 = ~n22820 ;
  assign y9821 = n22821 ;
  assign y9822 = ~n22823 ;
  assign y9823 = ~1'b0 ;
  assign y9824 = ~n22826 ;
  assign y9825 = ~1'b0 ;
  assign y9826 = ~n22830 ;
  assign y9827 = n22834 ;
  assign y9828 = n22837 ;
  assign y9829 = ~n22842 ;
  assign y9830 = n22843 ;
  assign y9831 = 1'b0 ;
  assign y9832 = n22845 ;
  assign y9833 = ~n22847 ;
  assign y9834 = ~1'b0 ;
  assign y9835 = ~n22849 ;
  assign y9836 = n22854 ;
  assign y9837 = n22857 ;
  assign y9838 = ~1'b0 ;
  assign y9839 = n22861 ;
  assign y9840 = ~n22863 ;
  assign y9841 = ~1'b0 ;
  assign y9842 = n22866 ;
  assign y9843 = n22871 ;
  assign y9844 = ~1'b0 ;
  assign y9845 = ~n22875 ;
  assign y9846 = n22877 ;
  assign y9847 = n22882 ;
  assign y9848 = n22887 ;
  assign y9849 = n17258 ;
  assign y9850 = ~n22891 ;
  assign y9851 = n22896 ;
  assign y9852 = n22900 ;
  assign y9853 = ~n22904 ;
  assign y9854 = ~1'b0 ;
  assign y9855 = ~1'b0 ;
  assign y9856 = n22905 ;
  assign y9857 = n22912 ;
  assign y9858 = ~1'b0 ;
  assign y9859 = n22915 ;
  assign y9860 = ~n22917 ;
  assign y9861 = ~n22919 ;
  assign y9862 = ~n22921 ;
  assign y9863 = ~n22922 ;
  assign y9864 = n22928 ;
  assign y9865 = ~n22934 ;
  assign y9866 = ~1'b0 ;
  assign y9867 = n22937 ;
  assign y9868 = n22939 ;
  assign y9869 = ~n22941 ;
  assign y9870 = ~n22943 ;
  assign y9871 = ~1'b0 ;
  assign y9872 = ~1'b0 ;
  assign y9873 = ~1'b0 ;
  assign y9874 = ~n22948 ;
  assign y9875 = n22950 ;
  assign y9876 = n22953 ;
  assign y9877 = ~n22955 ;
  assign y9878 = ~n22964 ;
  assign y9879 = ~n22968 ;
  assign y9880 = n3310 ;
  assign y9881 = n22974 ;
  assign y9882 = ~n22977 ;
  assign y9883 = n22981 ;
  assign y9884 = ~n11131 ;
  assign y9885 = ~1'b0 ;
  assign y9886 = ~1'b0 ;
  assign y9887 = ~1'b0 ;
  assign y9888 = n22982 ;
  assign y9889 = ~n22983 ;
  assign y9890 = ~n22984 ;
  assign y9891 = ~1'b0 ;
  assign y9892 = ~n22990 ;
  assign y9893 = ~1'b0 ;
  assign y9894 = ~n22993 ;
  assign y9895 = ~n22995 ;
  assign y9896 = ~1'b0 ;
  assign y9897 = n22997 ;
  assign y9898 = n22998 ;
  assign y9899 = n23006 ;
  assign y9900 = ~n7696 ;
  assign y9901 = ~1'b0 ;
  assign y9902 = n23009 ;
  assign y9903 = ~1'b0 ;
  assign y9904 = n23012 ;
  assign y9905 = ~n23015 ;
  assign y9906 = n23017 ;
  assign y9907 = n23020 ;
  assign y9908 = ~1'b0 ;
  assign y9909 = ~1'b0 ;
  assign y9910 = ~1'b0 ;
  assign y9911 = n23022 ;
  assign y9912 = n23025 ;
  assign y9913 = ~n23028 ;
  assign y9914 = ~1'b0 ;
  assign y9915 = n5425 ;
  assign y9916 = n23033 ;
  assign y9917 = ~n23044 ;
  assign y9918 = ~n23047 ;
  assign y9919 = ~1'b0 ;
  assign y9920 = n23049 ;
  assign y9921 = ~n23053 ;
  assign y9922 = ~n23058 ;
  assign y9923 = ~n23061 ;
  assign y9924 = ~1'b0 ;
  assign y9925 = n1619 ;
  assign y9926 = ~1'b0 ;
  assign y9927 = ~n23063 ;
  assign y9928 = ~n23069 ;
  assign y9929 = ~1'b0 ;
  assign y9930 = n23078 ;
  assign y9931 = ~1'b0 ;
  assign y9932 = ~1'b0 ;
  assign y9933 = ~n23079 ;
  assign y9934 = ~n23082 ;
  assign y9935 = ~n23084 ;
  assign y9936 = ~1'b0 ;
  assign y9937 = ~1'b0 ;
  assign y9938 = ~n23085 ;
  assign y9939 = ~1'b0 ;
  assign y9940 = ~1'b0 ;
  assign y9941 = n1991 ;
  assign y9942 = ~n23090 ;
  assign y9943 = ~n15803 ;
  assign y9944 = n23091 ;
  assign y9945 = ~1'b0 ;
  assign y9946 = ~n23097 ;
  assign y9947 = n23099 ;
  assign y9948 = ~1'b0 ;
  assign y9949 = n23104 ;
  assign y9950 = ~n23105 ;
  assign y9951 = ~1'b0 ;
  assign y9952 = ~n23108 ;
  assign y9953 = n23112 ;
  assign y9954 = n23114 ;
  assign y9955 = ~1'b0 ;
  assign y9956 = ~n23117 ;
  assign y9957 = ~1'b0 ;
  assign y9958 = ~n23118 ;
  assign y9959 = ~n23119 ;
  assign y9960 = n23121 ;
  assign y9961 = 1'b0 ;
  assign y9962 = n23122 ;
  assign y9963 = ~1'b0 ;
  assign y9964 = ~n21559 ;
  assign y9965 = n23139 ;
  assign y9966 = ~n23141 ;
  assign y9967 = n23149 ;
  assign y9968 = n23150 ;
  assign y9969 = ~1'b0 ;
  assign y9970 = n23151 ;
  assign y9971 = n23157 ;
  assign y9972 = ~n23159 ;
  assign y9973 = ~n8834 ;
  assign y9974 = ~1'b0 ;
  assign y9975 = n23163 ;
  assign y9976 = ~n23165 ;
  assign y9977 = ~1'b0 ;
  assign y9978 = ~n23169 ;
  assign y9979 = ~n23170 ;
  assign y9980 = ~1'b0 ;
  assign y9981 = ~n23175 ;
  assign y9982 = n23179 ;
  assign y9983 = ~1'b0 ;
  assign y9984 = ~1'b0 ;
  assign y9985 = ~1'b0 ;
  assign y9986 = ~n23180 ;
  assign y9987 = ~n23183 ;
  assign y9988 = ~n23185 ;
  assign y9989 = n23190 ;
  assign y9990 = n23193 ;
  assign y9991 = n23196 ;
  assign y9992 = ~n23201 ;
  assign y9993 = n23205 ;
  assign y9994 = n23212 ;
  assign y9995 = ~n23217 ;
  assign y9996 = ~1'b0 ;
  assign y9997 = n23218 ;
  assign y9998 = ~1'b0 ;
  assign y9999 = ~1'b0 ;
  assign y10000 = n23219 ;
  assign y10001 = n23220 ;
  assign y10002 = n23223 ;
  assign y10003 = n23225 ;
  assign y10004 = ~n23228 ;
  assign y10005 = ~n23236 ;
  assign y10006 = n23238 ;
  assign y10007 = ~1'b0 ;
  assign y10008 = ~n23246 ;
  assign y10009 = ~n23247 ;
  assign y10010 = ~1'b0 ;
  assign y10011 = n23249 ;
  assign y10012 = ~n23250 ;
  assign y10013 = ~1'b0 ;
  assign y10014 = ~1'b0 ;
  assign y10015 = ~1'b0 ;
  assign y10016 = ~1'b0 ;
  assign y10017 = n23251 ;
  assign y10018 = n23257 ;
  assign y10019 = ~1'b0 ;
  assign y10020 = ~1'b0 ;
  assign y10021 = n23258 ;
  assign y10022 = ~n23262 ;
  assign y10023 = ~n23266 ;
  assign y10024 = ~n23267 ;
  assign y10025 = n23268 ;
  assign y10026 = n23269 ;
  assign y10027 = ~1'b0 ;
  assign y10028 = n23271 ;
  assign y10029 = ~n23275 ;
  assign y10030 = ~1'b0 ;
  assign y10031 = ~1'b0 ;
  assign y10032 = ~n23283 ;
  assign y10033 = ~n23284 ;
  assign y10034 = n23287 ;
  assign y10035 = n23295 ;
  assign y10036 = ~1'b0 ;
  assign y10037 = ~n23299 ;
  assign y10038 = ~n23301 ;
  assign y10039 = n23302 ;
  assign y10040 = ~n23303 ;
  assign y10041 = ~n23304 ;
  assign y10042 = ~n23309 ;
  assign y10043 = ~n23313 ;
  assign y10044 = n23314 ;
  assign y10045 = ~n23319 ;
  assign y10046 = 1'b0 ;
  assign y10047 = ~n23320 ;
  assign y10048 = ~1'b0 ;
  assign y10049 = ~n23323 ;
  assign y10050 = ~n23327 ;
  assign y10051 = 1'b0 ;
  assign y10052 = ~1'b0 ;
  assign y10053 = n23329 ;
  assign y10054 = ~1'b0 ;
  assign y10055 = ~1'b0 ;
  assign y10056 = ~1'b0 ;
  assign y10057 = n23331 ;
  assign y10058 = ~n12869 ;
  assign y10059 = ~n23340 ;
  assign y10060 = n23344 ;
  assign y10061 = n23345 ;
  assign y10062 = ~1'b0 ;
  assign y10063 = ~n23346 ;
  assign y10064 = n23347 ;
  assign y10065 = n23348 ;
  assign y10066 = ~n23350 ;
  assign y10067 = n23357 ;
  assign y10068 = ~1'b0 ;
  assign y10069 = ~1'b0 ;
  assign y10070 = ~n23359 ;
  assign y10071 = ~1'b0 ;
  assign y10072 = ~n23369 ;
  assign y10073 = ~n23371 ;
  assign y10074 = n23374 ;
  assign y10075 = n23376 ;
  assign y10076 = n23378 ;
  assign y10077 = ~n23379 ;
  assign y10078 = ~n23382 ;
  assign y10079 = ~1'b0 ;
  assign y10080 = ~1'b0 ;
  assign y10081 = n23385 ;
  assign y10082 = ~n23386 ;
  assign y10083 = ~n23387 ;
  assign y10084 = n23393 ;
  assign y10085 = ~n23395 ;
  assign y10086 = ~n23398 ;
  assign y10087 = ~n23410 ;
  assign y10088 = ~n23411 ;
  assign y10089 = n5678 ;
  assign y10090 = ~n23416 ;
  assign y10091 = n23417 ;
  assign y10092 = ~1'b0 ;
  assign y10093 = n23419 ;
  assign y10094 = ~n23420 ;
  assign y10095 = ~n23424 ;
  assign y10096 = ~1'b0 ;
  assign y10097 = n23427 ;
  assign y10098 = n23430 ;
  assign y10099 = ~n23434 ;
  assign y10100 = ~1'b0 ;
  assign y10101 = ~1'b0 ;
  assign y10102 = 1'b0 ;
  assign y10103 = ~n23439 ;
  assign y10104 = ~n23441 ;
  assign y10105 = x55 ;
  assign y10106 = ~n23444 ;
  assign y10107 = ~1'b0 ;
  assign y10108 = n23446 ;
  assign y10109 = n23447 ;
  assign y10110 = ~n23448 ;
  assign y10111 = ~n23450 ;
  assign y10112 = n23451 ;
  assign y10113 = ~1'b0 ;
  assign y10114 = ~n23454 ;
  assign y10115 = 1'b0 ;
  assign y10116 = ~n23455 ;
  assign y10117 = ~n23456 ;
  assign y10118 = ~n23458 ;
  assign y10119 = n12635 ;
  assign y10120 = n23469 ;
  assign y10121 = ~1'b0 ;
  assign y10122 = n23471 ;
  assign y10123 = ~1'b0 ;
  assign y10124 = ~1'b0 ;
  assign y10125 = ~n23472 ;
  assign y10126 = ~1'b0 ;
  assign y10127 = n23475 ;
  assign y10128 = ~n23477 ;
  assign y10129 = n23482 ;
  assign y10130 = ~1'b0 ;
  assign y10131 = n23483 ;
  assign y10132 = ~1'b0 ;
  assign y10133 = ~n23487 ;
  assign y10134 = ~1'b0 ;
  assign y10135 = ~1'b0 ;
  assign y10136 = ~1'b0 ;
  assign y10137 = ~n23497 ;
  assign y10138 = ~n23503 ;
  assign y10139 = n23504 ;
  assign y10140 = ~n23508 ;
  assign y10141 = ~n23509 ;
  assign y10142 = ~1'b0 ;
  assign y10143 = n23513 ;
  assign y10144 = ~n23515 ;
  assign y10145 = n23517 ;
  assign y10146 = ~1'b0 ;
  assign y10147 = ~n23524 ;
  assign y10148 = n23526 ;
  assign y10149 = ~n23530 ;
  assign y10150 = n20706 ;
  assign y10151 = ~1'b0 ;
  assign y10152 = ~n4775 ;
  assign y10153 = ~1'b0 ;
  assign y10154 = ~n23531 ;
  assign y10155 = n23533 ;
  assign y10156 = ~n21713 ;
  assign y10157 = ~n23534 ;
  assign y10158 = ~1'b0 ;
  assign y10159 = n23536 ;
  assign y10160 = n23537 ;
  assign y10161 = ~n22816 ;
  assign y10162 = n23539 ;
  assign y10163 = ~n23543 ;
  assign y10164 = n23545 ;
  assign y10165 = ~n23550 ;
  assign y10166 = ~1'b0 ;
  assign y10167 = ~n23555 ;
  assign y10168 = n23556 ;
  assign y10169 = ~n23558 ;
  assign y10170 = n23561 ;
  assign y10171 = n23563 ;
  assign y10172 = ~n23567 ;
  assign y10173 = ~n23570 ;
  assign y10174 = ~1'b0 ;
  assign y10175 = ~n23571 ;
  assign y10176 = n23572 ;
  assign y10177 = n23574 ;
  assign y10178 = ~n23575 ;
  assign y10179 = n23576 ;
  assign y10180 = n23577 ;
  assign y10181 = n23581 ;
  assign y10182 = ~n704 ;
  assign y10183 = ~n23584 ;
  assign y10184 = ~n23590 ;
  assign y10185 = n23591 ;
  assign y10186 = ~1'b0 ;
  assign y10187 = ~n10940 ;
  assign y10188 = n23596 ;
  assign y10189 = ~n23598 ;
  assign y10190 = ~n23599 ;
  assign y10191 = ~n23601 ;
  assign y10192 = ~n23603 ;
  assign y10193 = ~n23604 ;
  assign y10194 = ~n23608 ;
  assign y10195 = ~1'b0 ;
  assign y10196 = ~1'b0 ;
  assign y10197 = ~1'b0 ;
  assign y10198 = n23609 ;
  assign y10199 = n23610 ;
  assign y10200 = n23620 ;
  assign y10201 = n23621 ;
  assign y10202 = ~n23623 ;
  assign y10203 = n23625 ;
  assign y10204 = ~1'b0 ;
  assign y10205 = n23628 ;
  assign y10206 = n23630 ;
  assign y10207 = ~n23635 ;
  assign y10208 = ~1'b0 ;
  assign y10209 = ~1'b0 ;
  assign y10210 = ~1'b0 ;
  assign y10211 = n23636 ;
  assign y10212 = ~n23641 ;
  assign y10213 = ~n23646 ;
  assign y10214 = ~1'b0 ;
  assign y10215 = ~n23649 ;
  assign y10216 = n23650 ;
  assign y10217 = n23652 ;
  assign y10218 = ~n23655 ;
  assign y10219 = ~n23656 ;
  assign y10220 = n11718 ;
  assign y10221 = n23659 ;
  assign y10222 = n23660 ;
  assign y10223 = ~1'b0 ;
  assign y10224 = ~1'b0 ;
  assign y10225 = n23663 ;
  assign y10226 = ~n23668 ;
  assign y10227 = ~1'b0 ;
  assign y10228 = ~n23672 ;
  assign y10229 = ~n23674 ;
  assign y10230 = ~n23676 ;
  assign y10231 = ~n5304 ;
  assign y10232 = ~1'b0 ;
  assign y10233 = ~1'b0 ;
  assign y10234 = ~1'b0 ;
  assign y10235 = ~n23679 ;
  assign y10236 = ~1'b0 ;
  assign y10237 = n23683 ;
  assign y10238 = n23684 ;
  assign y10239 = ~1'b0 ;
  assign y10240 = ~1'b0 ;
  assign y10241 = ~n23687 ;
  assign y10242 = n23689 ;
  assign y10243 = ~n23693 ;
  assign y10244 = n6613 ;
  assign y10245 = n23694 ;
  assign y10246 = n23696 ;
  assign y10247 = n23697 ;
  assign y10248 = ~n23708 ;
  assign y10249 = ~1'b0 ;
  assign y10250 = n23712 ;
  assign y10251 = ~n21626 ;
  assign y10252 = ~1'b0 ;
  assign y10253 = n6885 ;
  assign y10254 = ~1'b0 ;
  assign y10255 = n23713 ;
  assign y10256 = n23717 ;
  assign y10257 = n23730 ;
  assign y10258 = n23733 ;
  assign y10259 = n23737 ;
  assign y10260 = ~n23738 ;
  assign y10261 = ~n23743 ;
  assign y10262 = n23749 ;
  assign y10263 = n23752 ;
  assign y10264 = ~1'b0 ;
  assign y10265 = ~n23754 ;
  assign y10266 = ~n23758 ;
  assign y10267 = ~n23759 ;
  assign y10268 = n23761 ;
  assign y10269 = n17557 ;
  assign y10270 = ~1'b0 ;
  assign y10271 = n23763 ;
  assign y10272 = ~1'b0 ;
  assign y10273 = ~1'b0 ;
  assign y10274 = ~1'b0 ;
  assign y10275 = ~1'b0 ;
  assign y10276 = ~n23768 ;
  assign y10277 = n23771 ;
  assign y10278 = n23774 ;
  assign y10279 = 1'b0 ;
  assign y10280 = n23777 ;
  assign y10281 = ~1'b0 ;
  assign y10282 = n23783 ;
  assign y10283 = ~n23787 ;
  assign y10284 = ~n23790 ;
  assign y10285 = ~n23792 ;
  assign y10286 = n23794 ;
  assign y10287 = ~1'b0 ;
  assign y10288 = n23796 ;
  assign y10289 = 1'b0 ;
  assign y10290 = n23797 ;
  assign y10291 = n23800 ;
  assign y10292 = ~n23803 ;
  assign y10293 = ~n23807 ;
  assign y10294 = n8949 ;
  assign y10295 = n23809 ;
  assign y10296 = n23810 ;
  assign y10297 = ~1'b0 ;
  assign y10298 = ~n23815 ;
  assign y10299 = ~1'b0 ;
  assign y10300 = n23817 ;
  assign y10301 = n23818 ;
  assign y10302 = ~1'b0 ;
  assign y10303 = 1'b0 ;
  assign y10304 = ~n23819 ;
  assign y10305 = ~n23820 ;
  assign y10306 = ~1'b0 ;
  assign y10307 = n23823 ;
  assign y10308 = ~1'b0 ;
  assign y10309 = n23827 ;
  assign y10310 = ~1'b0 ;
  assign y10311 = ~n23830 ;
  assign y10312 = ~n7360 ;
  assign y10313 = ~n23832 ;
  assign y10314 = ~n23836 ;
  assign y10315 = ~n23838 ;
  assign y10316 = ~1'b0 ;
  assign y10317 = n23839 ;
  assign y10318 = ~n23840 ;
  assign y10319 = n23841 ;
  assign y10320 = ~1'b0 ;
  assign y10321 = ~1'b0 ;
  assign y10322 = n21034 ;
  assign y10323 = ~n23843 ;
  assign y10324 = ~n23844 ;
  assign y10325 = ~1'b0 ;
  assign y10326 = ~n23846 ;
  assign y10327 = n5387 ;
  assign y10328 = n23847 ;
  assign y10329 = ~n13634 ;
  assign y10330 = n23849 ;
  assign y10331 = n23850 ;
  assign y10332 = n4770 ;
  assign y10333 = n23853 ;
  assign y10334 = n23854 ;
  assign y10335 = ~n15197 ;
  assign y10336 = n23858 ;
  assign y10337 = ~n23862 ;
  assign y10338 = ~n23864 ;
  assign y10339 = ~n23868 ;
  assign y10340 = n23871 ;
  assign y10341 = n23873 ;
  assign y10342 = ~n23874 ;
  assign y10343 = n23879 ;
  assign y10344 = ~n23882 ;
  assign y10345 = ~n23884 ;
  assign y10346 = ~n23887 ;
  assign y10347 = n23889 ;
  assign y10348 = ~n23895 ;
  assign y10349 = ~1'b0 ;
  assign y10350 = n23899 ;
  assign y10351 = ~1'b0 ;
  assign y10352 = n23900 ;
  assign y10353 = n23904 ;
  assign y10354 = ~1'b0 ;
  assign y10355 = ~1'b0 ;
  assign y10356 = ~n23905 ;
  assign y10357 = ~1'b0 ;
  assign y10358 = n23906 ;
  assign y10359 = ~1'b0 ;
  assign y10360 = n1872 ;
  assign y10361 = ~1'b0 ;
  assign y10362 = ~n23907 ;
  assign y10363 = ~1'b0 ;
  assign y10364 = ~1'b0 ;
  assign y10365 = n23909 ;
  assign y10366 = ~1'b0 ;
  assign y10367 = ~n23911 ;
  assign y10368 = n23914 ;
  assign y10369 = n23916 ;
  assign y10370 = n23918 ;
  assign y10371 = ~1'b0 ;
  assign y10372 = ~n23921 ;
  assign y10373 = ~1'b0 ;
  assign y10374 = n23923 ;
  assign y10375 = ~n23924 ;
  assign y10376 = ~n23930 ;
  assign y10377 = ~1'b0 ;
  assign y10378 = ~n23934 ;
  assign y10379 = n744 ;
  assign y10380 = ~n23935 ;
  assign y10381 = ~1'b0 ;
  assign y10382 = ~n23938 ;
  assign y10383 = ~n23941 ;
  assign y10384 = ~1'b0 ;
  assign y10385 = ~1'b0 ;
  assign y10386 = ~1'b0 ;
  assign y10387 = ~1'b0 ;
  assign y10388 = ~1'b0 ;
  assign y10389 = ~n23943 ;
  assign y10390 = ~1'b0 ;
  assign y10391 = ~n23945 ;
  assign y10392 = ~n23951 ;
  assign y10393 = ~1'b0 ;
  assign y10394 = ~n23953 ;
  assign y10395 = ~n23956 ;
  assign y10396 = ~1'b0 ;
  assign y10397 = ~1'b0 ;
  assign y10398 = ~n23957 ;
  assign y10399 = ~1'b0 ;
  assign y10400 = ~1'b0 ;
  assign y10401 = ~n6274 ;
  assign y10402 = ~1'b0 ;
  assign y10403 = ~1'b0 ;
  assign y10404 = ~n23964 ;
  assign y10405 = ~n23965 ;
  assign y10406 = n23975 ;
  assign y10407 = ~n23977 ;
  assign y10408 = ~1'b0 ;
  assign y10409 = ~1'b0 ;
  assign y10410 = n23979 ;
  assign y10411 = ~n23980 ;
  assign y10412 = n23985 ;
  assign y10413 = ~1'b0 ;
  assign y10414 = ~n23986 ;
  assign y10415 = n23989 ;
  assign y10416 = ~n20188 ;
  assign y10417 = n23992 ;
  assign y10418 = n23995 ;
  assign y10419 = n23997 ;
  assign y10420 = ~n24000 ;
  assign y10421 = ~n24002 ;
  assign y10422 = n24003 ;
  assign y10423 = n24004 ;
  assign y10424 = ~n24005 ;
  assign y10425 = ~n24010 ;
  assign y10426 = ~n24011 ;
  assign y10427 = n5939 ;
  assign y10428 = ~n24013 ;
  assign y10429 = ~n24015 ;
  assign y10430 = ~n10886 ;
  assign y10431 = ~n24016 ;
  assign y10432 = ~1'b0 ;
  assign y10433 = n24020 ;
  assign y10434 = n24023 ;
  assign y10435 = ~n24026 ;
  assign y10436 = n24027 ;
  assign y10437 = ~1'b0 ;
  assign y10438 = ~n24029 ;
  assign y10439 = ~n24033 ;
  assign y10440 = ~1'b0 ;
  assign y10441 = n24034 ;
  assign y10442 = ~n21681 ;
  assign y10443 = n24036 ;
  assign y10444 = ~1'b0 ;
  assign y10445 = ~n21317 ;
  assign y10446 = ~n24044 ;
  assign y10447 = n24047 ;
  assign y10448 = ~1'b0 ;
  assign y10449 = n24050 ;
  assign y10450 = n24057 ;
  assign y10451 = n24059 ;
  assign y10452 = ~1'b0 ;
  assign y10453 = ~n24061 ;
  assign y10454 = n24065 ;
  assign y10455 = ~1'b0 ;
  assign y10456 = ~n24069 ;
  assign y10457 = n24070 ;
  assign y10458 = ~n24073 ;
  assign y10459 = n24077 ;
  assign y10460 = n24090 ;
  assign y10461 = n24093 ;
  assign y10462 = ~n24099 ;
  assign y10463 = n24104 ;
  assign y10464 = ~1'b0 ;
  assign y10465 = ~n24105 ;
  assign y10466 = n19157 ;
  assign y10467 = n24107 ;
  assign y10468 = ~n24108 ;
  assign y10469 = n24109 ;
  assign y10470 = n24112 ;
  assign y10471 = ~1'b0 ;
  assign y10472 = ~1'b0 ;
  assign y10473 = n24115 ;
  assign y10474 = n24117 ;
  assign y10475 = n24122 ;
  assign y10476 = ~1'b0 ;
  assign y10477 = n24123 ;
  assign y10478 = n24125 ;
  assign y10479 = ~n24127 ;
  assign y10480 = ~1'b0 ;
  assign y10481 = n3052 ;
  assign y10482 = ~1'b0 ;
  assign y10483 = n24132 ;
  assign y10484 = ~n24133 ;
  assign y10485 = ~n24138 ;
  assign y10486 = n24139 ;
  assign y10487 = n24141 ;
  assign y10488 = ~n24142 ;
  assign y10489 = n24144 ;
  assign y10490 = ~n24146 ;
  assign y10491 = n24149 ;
  assign y10492 = n24159 ;
  assign y10493 = ~1'b0 ;
  assign y10494 = 1'b0 ;
  assign y10495 = ~1'b0 ;
  assign y10496 = ~1'b0 ;
  assign y10497 = ~n24160 ;
  assign y10498 = n24161 ;
  assign y10499 = 1'b0 ;
  assign y10500 = n21836 ;
  assign y10501 = n24163 ;
  assign y10502 = ~1'b0 ;
  assign y10503 = ~1'b0 ;
  assign y10504 = n24164 ;
  assign y10505 = n24167 ;
  assign y10506 = ~n24168 ;
  assign y10507 = n19773 ;
  assign y10508 = ~n24171 ;
  assign y10509 = n24173 ;
  assign y10510 = n24175 ;
  assign y10511 = n24179 ;
  assign y10512 = n24182 ;
  assign y10513 = ~n24187 ;
  assign y10514 = n24188 ;
  assign y10515 = ~n24190 ;
  assign y10516 = n24195 ;
  assign y10517 = ~n24201 ;
  assign y10518 = ~n24202 ;
  assign y10519 = n24206 ;
  assign y10520 = ~n24207 ;
  assign y10521 = ~n24208 ;
  assign y10522 = ~n24216 ;
  assign y10523 = ~n24225 ;
  assign y10524 = ~n24230 ;
  assign y10525 = ~n24231 ;
  assign y10526 = ~n24232 ;
  assign y10527 = ~n24235 ;
  assign y10528 = ~n24236 ;
  assign y10529 = ~n24238 ;
  assign y10530 = ~1'b0 ;
  assign y10531 = ~1'b0 ;
  assign y10532 = ~n24239 ;
  assign y10533 = n24240 ;
  assign y10534 = n24249 ;
  assign y10535 = ~n24251 ;
  assign y10536 = ~1'b0 ;
  assign y10537 = n24253 ;
  assign y10538 = ~1'b0 ;
  assign y10539 = ~1'b0 ;
  assign y10540 = ~1'b0 ;
  assign y10541 = n24257 ;
  assign y10542 = n24260 ;
  assign y10543 = n24266 ;
  assign y10544 = ~1'b0 ;
  assign y10545 = ~n24268 ;
  assign y10546 = ~n24274 ;
  assign y10547 = ~n24280 ;
  assign y10548 = n24283 ;
  assign y10549 = ~n24284 ;
  assign y10550 = ~1'b0 ;
  assign y10551 = ~n24293 ;
  assign y10552 = ~1'b0 ;
  assign y10553 = ~n24297 ;
  assign y10554 = n24299 ;
  assign y10555 = ~1'b0 ;
  assign y10556 = ~n24300 ;
  assign y10557 = n2774 ;
  assign y10558 = ~n24303 ;
  assign y10559 = ~n24305 ;
  assign y10560 = n24306 ;
  assign y10561 = n24308 ;
  assign y10562 = ~1'b0 ;
  assign y10563 = 1'b0 ;
  assign y10564 = n24313 ;
  assign y10565 = ~1'b0 ;
  assign y10566 = ~1'b0 ;
  assign y10567 = ~n24316 ;
  assign y10568 = ~n24317 ;
  assign y10569 = ~n24319 ;
  assign y10570 = ~1'b0 ;
  assign y10571 = n24320 ;
  assign y10572 = ~1'b0 ;
  assign y10573 = ~n24322 ;
  assign y10574 = ~n24325 ;
  assign y10575 = ~1'b0 ;
  assign y10576 = n24326 ;
  assign y10577 = ~n24329 ;
  assign y10578 = n24330 ;
  assign y10579 = ~n24333 ;
  assign y10580 = ~n24335 ;
  assign y10581 = ~1'b0 ;
  assign y10582 = ~n24336 ;
  assign y10583 = n24338 ;
  assign y10584 = n24345 ;
  assign y10585 = ~1'b0 ;
  assign y10586 = ~1'b0 ;
  assign y10587 = n24346 ;
  assign y10588 = ~1'b0 ;
  assign y10589 = ~n24351 ;
  assign y10590 = ~n24352 ;
  assign y10591 = n24356 ;
  assign y10592 = n24359 ;
  assign y10593 = ~n24361 ;
  assign y10594 = n24363 ;
  assign y10595 = ~1'b0 ;
  assign y10596 = n24365 ;
  assign y10597 = n24367 ;
  assign y10598 = ~n8432 ;
  assign y10599 = n24371 ;
  assign y10600 = ~n24377 ;
  assign y10601 = ~1'b0 ;
  assign y10602 = ~1'b0 ;
  assign y10603 = n24378 ;
  assign y10604 = ~1'b0 ;
  assign y10605 = ~1'b0 ;
  assign y10606 = n24380 ;
  assign y10607 = n24381 ;
  assign y10608 = ~n24385 ;
  assign y10609 = ~n24386 ;
  assign y10610 = ~n24388 ;
  assign y10611 = 1'b0 ;
  assign y10612 = ~1'b0 ;
  assign y10613 = ~n24390 ;
  assign y10614 = ~n24395 ;
  assign y10615 = n24396 ;
  assign y10616 = ~n4058 ;
  assign y10617 = ~n24397 ;
  assign y10618 = n24400 ;
  assign y10619 = ~n24401 ;
  assign y10620 = ~1'b0 ;
  assign y10621 = n24402 ;
  assign y10622 = ~n24404 ;
  assign y10623 = n24405 ;
  assign y10624 = ~1'b0 ;
  assign y10625 = ~n24406 ;
  assign y10626 = ~n24407 ;
  assign y10627 = ~n24409 ;
  assign y10628 = ~1'b0 ;
  assign y10629 = n24410 ;
  assign y10630 = ~n24411 ;
  assign y10631 = ~n24412 ;
  assign y10632 = ~1'b0 ;
  assign y10633 = ~n24413 ;
  assign y10634 = ~n24417 ;
  assign y10635 = n24423 ;
  assign y10636 = n24427 ;
  assign y10637 = ~n24428 ;
  assign y10638 = ~1'b0 ;
  assign y10639 = ~1'b0 ;
  assign y10640 = n24430 ;
  assign y10641 = n24431 ;
  assign y10642 = ~n24434 ;
  assign y10643 = 1'b0 ;
  assign y10644 = ~1'b0 ;
  assign y10645 = ~1'b0 ;
  assign y10646 = n24447 ;
  assign y10647 = ~1'b0 ;
  assign y10648 = n17007 ;
  assign y10649 = n24448 ;
  assign y10650 = ~n24449 ;
  assign y10651 = n24452 ;
  assign y10652 = ~1'b0 ;
  assign y10653 = ~1'b0 ;
  assign y10654 = n24460 ;
  assign y10655 = n24461 ;
  assign y10656 = n24463 ;
  assign y10657 = ~1'b0 ;
  assign y10658 = n24466 ;
  assign y10659 = ~n24470 ;
  assign y10660 = ~1'b0 ;
  assign y10661 = n24473 ;
  assign y10662 = ~1'b0 ;
  assign y10663 = ~n24477 ;
  assign y10664 = ~1'b0 ;
  assign y10665 = ~1'b0 ;
  assign y10666 = n24487 ;
  assign y10667 = ~n24490 ;
  assign y10668 = ~1'b0 ;
  assign y10669 = n24492 ;
  assign y10670 = ~n24494 ;
  assign y10671 = ~n24495 ;
  assign y10672 = n24497 ;
  assign y10673 = ~1'b0 ;
  assign y10674 = ~n24500 ;
  assign y10675 = 1'b0 ;
  assign y10676 = ~n24507 ;
  assign y10677 = n24509 ;
  assign y10678 = n24514 ;
  assign y10679 = n24516 ;
  assign y10680 = n24518 ;
  assign y10681 = ~n24521 ;
  assign y10682 = ~n24522 ;
  assign y10683 = n24528 ;
  assign y10684 = n24530 ;
  assign y10685 = ~n24533 ;
  assign y10686 = n24535 ;
  assign y10687 = n24541 ;
  assign y10688 = n24545 ;
  assign y10689 = ~1'b0 ;
  assign y10690 = n24550 ;
  assign y10691 = n24554 ;
  assign y10692 = n14550 ;
  assign y10693 = ~1'b0 ;
  assign y10694 = ~1'b0 ;
  assign y10695 = n24557 ;
  assign y10696 = ~n24567 ;
  assign y10697 = ~n24568 ;
  assign y10698 = ~n23511 ;
  assign y10699 = ~n24569 ;
  assign y10700 = ~n10582 ;
  assign y10701 = ~n24572 ;
  assign y10702 = ~n24573 ;
  assign y10703 = n24577 ;
  assign y10704 = ~1'b0 ;
  assign y10705 = n24578 ;
  assign y10706 = ~n24579 ;
  assign y10707 = n24581 ;
  assign y10708 = ~1'b0 ;
  assign y10709 = ~1'b0 ;
  assign y10710 = ~n24583 ;
  assign y10711 = ~n24585 ;
  assign y10712 = ~1'b0 ;
  assign y10713 = n24586 ;
  assign y10714 = ~n24589 ;
  assign y10715 = ~n24591 ;
  assign y10716 = n24592 ;
  assign y10717 = n24594 ;
  assign y10718 = ~1'b0 ;
  assign y10719 = ~n24595 ;
  assign y10720 = ~1'b0 ;
  assign y10721 = ~1'b0 ;
  assign y10722 = n24597 ;
  assign y10723 = ~1'b0 ;
  assign y10724 = n24601 ;
  assign y10725 = ~n24604 ;
  assign y10726 = ~n24608 ;
  assign y10727 = n24615 ;
  assign y10728 = ~1'b0 ;
  assign y10729 = ~n24621 ;
  assign y10730 = ~n24622 ;
  assign y10731 = n24626 ;
  assign y10732 = n24632 ;
  assign y10733 = ~1'b0 ;
  assign y10734 = ~n24638 ;
  assign y10735 = ~n24640 ;
  assign y10736 = ~1'b0 ;
  assign y10737 = ~1'b0 ;
  assign y10738 = ~1'b0 ;
  assign y10739 = n24641 ;
  assign y10740 = n24642 ;
  assign y10741 = n24643 ;
  assign y10742 = n24645 ;
  assign y10743 = n24648 ;
  assign y10744 = ~n24651 ;
  assign y10745 = ~n24653 ;
  assign y10746 = ~n24655 ;
  assign y10747 = ~1'b0 ;
  assign y10748 = ~n24660 ;
  assign y10749 = ~1'b0 ;
  assign y10750 = ~n24663 ;
  assign y10751 = n24664 ;
  assign y10752 = ~n24671 ;
  assign y10753 = ~n24676 ;
  assign y10754 = n24175 ;
  assign y10755 = 1'b0 ;
  assign y10756 = 1'b0 ;
  assign y10757 = n24680 ;
  assign y10758 = ~n24681 ;
  assign y10759 = ~n24682 ;
  assign y10760 = n24683 ;
  assign y10761 = n24684 ;
  assign y10762 = ~1'b0 ;
  assign y10763 = n24687 ;
  assign y10764 = ~n24311 ;
  assign y10765 = n24691 ;
  assign y10766 = n24693 ;
  assign y10767 = ~1'b0 ;
  assign y10768 = n24694 ;
  assign y10769 = n24696 ;
  assign y10770 = ~n24697 ;
  assign y10771 = n24700 ;
  assign y10772 = ~n24701 ;
  assign y10773 = ~1'b0 ;
  assign y10774 = n24702 ;
  assign y10775 = ~n24704 ;
  assign y10776 = ~1'b0 ;
  assign y10777 = ~1'b0 ;
  assign y10778 = ~1'b0 ;
  assign y10779 = ~n24706 ;
  assign y10780 = n24710 ;
  assign y10781 = ~n24713 ;
  assign y10782 = ~n24715 ;
  assign y10783 = n24717 ;
  assign y10784 = n24719 ;
  assign y10785 = ~n24722 ;
  assign y10786 = 1'b0 ;
  assign y10787 = ~n24723 ;
  assign y10788 = n9482 ;
  assign y10789 = ~n24724 ;
  assign y10790 = ~n24728 ;
  assign y10791 = n24730 ;
  assign y10792 = n24732 ;
  assign y10793 = n24735 ;
  assign y10794 = n24738 ;
  assign y10795 = n24745 ;
  assign y10796 = ~n24749 ;
  assign y10797 = n24750 ;
  assign y10798 = n24751 ;
  assign y10799 = ~1'b0 ;
  assign y10800 = n24752 ;
  assign y10801 = ~n24755 ;
  assign y10802 = ~n24758 ;
  assign y10803 = ~n24759 ;
  assign y10804 = ~n24760 ;
  assign y10805 = n24761 ;
  assign y10806 = ~1'b0 ;
  assign y10807 = ~n24763 ;
  assign y10808 = n24767 ;
  assign y10809 = ~1'b0 ;
  assign y10810 = n24768 ;
  assign y10811 = ~n24769 ;
  assign y10812 = ~n24770 ;
  assign y10813 = ~1'b0 ;
  assign y10814 = n24776 ;
  assign y10815 = ~n22006 ;
  assign y10816 = n4509 ;
  assign y10817 = ~1'b0 ;
  assign y10818 = ~1'b0 ;
  assign y10819 = n14046 ;
  assign y10820 = n11426 ;
  assign y10821 = 1'b0 ;
  assign y10822 = ~1'b0 ;
  assign y10823 = ~1'b0 ;
  assign y10824 = n24781 ;
  assign y10825 = ~n24782 ;
  assign y10826 = n1506 ;
  assign y10827 = n24785 ;
  assign y10828 = ~1'b0 ;
  assign y10829 = n24787 ;
  assign y10830 = n24788 ;
  assign y10831 = ~n24792 ;
  assign y10832 = n24795 ;
  assign y10833 = ~1'b0 ;
  assign y10834 = ~1'b0 ;
  assign y10835 = n24796 ;
  assign y10836 = n9836 ;
  assign y10837 = ~x156 ;
  assign y10838 = ~n24801 ;
  assign y10839 = ~1'b0 ;
  assign y10840 = ~1'b0 ;
  assign y10841 = n24804 ;
  assign y10842 = ~1'b0 ;
  assign y10843 = ~n24805 ;
  assign y10844 = ~n24810 ;
  assign y10845 = ~n24811 ;
  assign y10846 = ~1'b0 ;
  assign y10847 = n24813 ;
  assign y10848 = ~n12221 ;
  assign y10849 = ~n18508 ;
  assign y10850 = ~n24815 ;
  assign y10851 = ~n24816 ;
  assign y10852 = n24819 ;
  assign y10853 = ~n24822 ;
  assign y10854 = n24825 ;
  assign y10855 = ~1'b0 ;
  assign y10856 = ~n24826 ;
  assign y10857 = ~n24830 ;
  assign y10858 = ~1'b0 ;
  assign y10859 = n24831 ;
  assign y10860 = ~1'b0 ;
  assign y10861 = ~n24834 ;
  assign y10862 = ~n24838 ;
  assign y10863 = ~1'b0 ;
  assign y10864 = n24839 ;
  assign y10865 = n24841 ;
  assign y10866 = n24842 ;
  assign y10867 = ~n24845 ;
  assign y10868 = n24846 ;
  assign y10869 = ~n24850 ;
  assign y10870 = n24851 ;
  assign y10871 = n24853 ;
  assign y10872 = ~n24856 ;
  assign y10873 = ~1'b0 ;
  assign y10874 = ~n24863 ;
  assign y10875 = ~n24867 ;
  assign y10876 = ~n24869 ;
  assign y10877 = ~x157 ;
  assign y10878 = n24871 ;
  assign y10879 = n24874 ;
  assign y10880 = ~n24876 ;
  assign y10881 = ~n24877 ;
  assign y10882 = n24878 ;
  assign y10883 = ~n24885 ;
  assign y10884 = n24886 ;
  assign y10885 = ~n24894 ;
  assign y10886 = ~1'b0 ;
  assign y10887 = ~n24896 ;
  assign y10888 = ~n24898 ;
  assign y10889 = n24899 ;
  assign y10890 = n24903 ;
  assign y10891 = ~1'b0 ;
  assign y10892 = ~1'b0 ;
  assign y10893 = n24908 ;
  assign y10894 = n24912 ;
  assign y10895 = n24917 ;
  assign y10896 = n24920 ;
  assign y10897 = ~1'b0 ;
  assign y10898 = ~n24924 ;
  assign y10899 = ~1'b0 ;
  assign y10900 = ~n24934 ;
  assign y10901 = ~n24935 ;
  assign y10902 = ~1'b0 ;
  assign y10903 = ~1'b0 ;
  assign y10904 = ~1'b0 ;
  assign y10905 = ~1'b0 ;
  assign y10906 = ~n24943 ;
  assign y10907 = ~1'b0 ;
  assign y10908 = n24948 ;
  assign y10909 = n24950 ;
  assign y10910 = n24951 ;
  assign y10911 = ~n24955 ;
  assign y10912 = ~1'b0 ;
  assign y10913 = n24956 ;
  assign y10914 = n24959 ;
  assign y10915 = n24961 ;
  assign y10916 = n24965 ;
  assign y10917 = ~n24969 ;
  assign y10918 = ~1'b0 ;
  assign y10919 = ~n24980 ;
  assign y10920 = n24982 ;
  assign y10921 = n24983 ;
  assign y10922 = ~n24988 ;
  assign y10923 = n24991 ;
  assign y10924 = n24993 ;
  assign y10925 = ~n24996 ;
  assign y10926 = ~1'b0 ;
  assign y10927 = n24999 ;
  assign y10928 = ~1'b0 ;
  assign y10929 = n25001 ;
  assign y10930 = ~1'b0 ;
  assign y10931 = ~n25004 ;
  assign y10932 = n25011 ;
  assign y10933 = ~1'b0 ;
  assign y10934 = x57 ;
  assign y10935 = n25013 ;
  assign y10936 = ~n25016 ;
  assign y10937 = n25017 ;
  assign y10938 = ~n25021 ;
  assign y10939 = n25024 ;
  assign y10940 = ~1'b0 ;
  assign y10941 = n25027 ;
  assign y10942 = ~1'b0 ;
  assign y10943 = n25030 ;
  assign y10944 = ~n25031 ;
  assign y10945 = ~n25033 ;
  assign y10946 = ~1'b0 ;
  assign y10947 = 1'b0 ;
  assign y10948 = n25036 ;
  assign y10949 = ~n25041 ;
  assign y10950 = n25042 ;
  assign y10951 = ~n5059 ;
  assign y10952 = n25043 ;
  assign y10953 = ~1'b0 ;
  assign y10954 = ~n21701 ;
  assign y10955 = n12546 ;
  assign y10956 = ~n25050 ;
  assign y10957 = ~n25054 ;
  assign y10958 = ~n6665 ;
  assign y10959 = n25057 ;
  assign y10960 = ~n25063 ;
  assign y10961 = ~1'b0 ;
  assign y10962 = ~n25064 ;
  assign y10963 = ~n25072 ;
  assign y10964 = ~n25073 ;
  assign y10965 = n25076 ;
  assign y10966 = ~1'b0 ;
  assign y10967 = n25077 ;
  assign y10968 = ~1'b0 ;
  assign y10969 = n25081 ;
  assign y10970 = ~n25084 ;
  assign y10971 = n25086 ;
  assign y10972 = n25087 ;
  assign y10973 = ~n25100 ;
  assign y10974 = n25102 ;
  assign y10975 = ~1'b0 ;
  assign y10976 = n25113 ;
  assign y10977 = ~1'b0 ;
  assign y10978 = ~1'b0 ;
  assign y10979 = ~1'b0 ;
  assign y10980 = ~n25114 ;
  assign y10981 = ~n25116 ;
  assign y10982 = ~1'b0 ;
  assign y10983 = n25118 ;
  assign y10984 = ~1'b0 ;
  assign y10985 = n25119 ;
  assign y10986 = ~n25122 ;
  assign y10987 = n10621 ;
  assign y10988 = ~n25125 ;
  assign y10989 = ~n25127 ;
  assign y10990 = ~n25128 ;
  assign y10991 = ~n25130 ;
  assign y10992 = ~n25132 ;
  assign y10993 = ~n25139 ;
  assign y10994 = ~1'b0 ;
  assign y10995 = ~n25140 ;
  assign y10996 = n25145 ;
  assign y10997 = n25147 ;
  assign y10998 = n25149 ;
  assign y10999 = n25152 ;
  assign y11000 = ~n25153 ;
  assign y11001 = n25154 ;
  assign y11002 = ~n25158 ;
  assign y11003 = n25163 ;
  assign y11004 = n25169 ;
  assign y11005 = ~n25179 ;
  assign y11006 = n25182 ;
  assign y11007 = ~n21777 ;
  assign y11008 = n25185 ;
  assign y11009 = ~n25191 ;
  assign y11010 = n25195 ;
  assign y11011 = n5689 ;
  assign y11012 = ~1'b0 ;
  assign y11013 = n6249 ;
  assign y11014 = ~n25198 ;
  assign y11015 = n25201 ;
  assign y11016 = n25207 ;
  assign y11017 = n25208 ;
  assign y11018 = ~n25209 ;
  assign y11019 = ~1'b0 ;
  assign y11020 = ~1'b0 ;
  assign y11021 = ~1'b0 ;
  assign y11022 = ~1'b0 ;
  assign y11023 = 1'b0 ;
  assign y11024 = n19532 ;
  assign y11025 = n25216 ;
  assign y11026 = ~1'b0 ;
  assign y11027 = ~n25226 ;
  assign y11028 = ~n25229 ;
  assign y11029 = n25231 ;
  assign y11030 = n25233 ;
  assign y11031 = n25234 ;
  assign y11032 = ~n25236 ;
  assign y11033 = n25240 ;
  assign y11034 = n25242 ;
  assign y11035 = ~1'b0 ;
  assign y11036 = ~1'b0 ;
  assign y11037 = ~n22400 ;
  assign y11038 = n25245 ;
  assign y11039 = ~n25246 ;
  assign y11040 = ~n25247 ;
  assign y11041 = ~1'b0 ;
  assign y11042 = ~1'b0 ;
  assign y11043 = n25248 ;
  assign y11044 = ~1'b0 ;
  assign y11045 = ~n25254 ;
  assign y11046 = n25255 ;
  assign y11047 = n23005 ;
  assign y11048 = n25256 ;
  assign y11049 = n25257 ;
  assign y11050 = ~n25258 ;
  assign y11051 = ~n25262 ;
  assign y11052 = n25264 ;
  assign y11053 = n25266 ;
  assign y11054 = ~1'b0 ;
  assign y11055 = n25268 ;
  assign y11056 = n25270 ;
  assign y11057 = ~n25273 ;
  assign y11058 = ~1'b0 ;
  assign y11059 = ~n25280 ;
  assign y11060 = n25282 ;
  assign y11061 = n25285 ;
  assign y11062 = ~n25287 ;
  assign y11063 = n25293 ;
  assign y11064 = ~1'b0 ;
  assign y11065 = ~n25301 ;
  assign y11066 = ~n25308 ;
  assign y11067 = n25312 ;
  assign y11068 = n25319 ;
  assign y11069 = n25320 ;
  assign y11070 = ~n25321 ;
  assign y11071 = n25322 ;
  assign y11072 = ~n25324 ;
  assign y11073 = ~n25325 ;
  assign y11074 = n25328 ;
  assign y11075 = ~n25333 ;
  assign y11076 = n565 ;
  assign y11077 = ~1'b0 ;
  assign y11078 = n25334 ;
  assign y11079 = n25339 ;
  assign y11080 = ~n25341 ;
  assign y11081 = ~n25342 ;
  assign y11082 = ~1'b0 ;
  assign y11083 = ~n25345 ;
  assign y11084 = ~n11123 ;
  assign y11085 = ~1'b0 ;
  assign y11086 = ~1'b0 ;
  assign y11087 = ~n25347 ;
  assign y11088 = n25348 ;
  assign y11089 = n25354 ;
  assign y11090 = ~n25359 ;
  assign y11091 = ~1'b0 ;
  assign y11092 = n25362 ;
  assign y11093 = n25365 ;
  assign y11094 = 1'b0 ;
  assign y11095 = ~n25372 ;
  assign y11096 = n25373 ;
  assign y11097 = n25376 ;
  assign y11098 = n25378 ;
  assign y11099 = n25382 ;
  assign y11100 = ~n25388 ;
  assign y11101 = n25392 ;
  assign y11102 = ~n25394 ;
  assign y11103 = ~1'b0 ;
  assign y11104 = ~1'b0 ;
  assign y11105 = ~1'b0 ;
  assign y11106 = n25395 ;
  assign y11107 = n25397 ;
  assign y11108 = n1651 ;
  assign y11109 = ~1'b0 ;
  assign y11110 = n25402 ;
  assign y11111 = ~n25405 ;
  assign y11112 = n25408 ;
  assign y11113 = n25411 ;
  assign y11114 = n25414 ;
  assign y11115 = ~1'b0 ;
  assign y11116 = n25416 ;
  assign y11117 = ~n25418 ;
  assign y11118 = ~n25419 ;
  assign y11119 = ~n25423 ;
  assign y11120 = n25424 ;
  assign y11121 = n25429 ;
  assign y11122 = ~1'b0 ;
  assign y11123 = n25430 ;
  assign y11124 = ~1'b0 ;
  assign y11125 = n25433 ;
  assign y11126 = n23205 ;
  assign y11127 = ~n25437 ;
  assign y11128 = 1'b0 ;
  assign y11129 = n18307 ;
  assign y11130 = ~1'b0 ;
  assign y11131 = n25444 ;
  assign y11132 = n25447 ;
  assign y11133 = n25453 ;
  assign y11134 = n25457 ;
  assign y11135 = n25459 ;
  assign y11136 = n25462 ;
  assign y11137 = ~n25464 ;
  assign y11138 = ~n25474 ;
  assign y11139 = n25477 ;
  assign y11140 = ~1'b0 ;
  assign y11141 = ~n21930 ;
  assign y11142 = ~n25481 ;
  assign y11143 = ~1'b0 ;
  assign y11144 = ~n5816 ;
  assign y11145 = n25482 ;
  assign y11146 = n25487 ;
  assign y11147 = n25499 ;
  assign y11148 = ~n25501 ;
  assign y11149 = ~n25503 ;
  assign y11150 = ~n25514 ;
  assign y11151 = ~1'b0 ;
  assign y11152 = ~n25521 ;
  assign y11153 = ~1'b0 ;
  assign y11154 = n25525 ;
  assign y11155 = ~n9556 ;
  assign y11156 = ~n25529 ;
  assign y11157 = ~n25532 ;
  assign y11158 = n25533 ;
  assign y11159 = ~n25535 ;
  assign y11160 = ~1'b0 ;
  assign y11161 = ~n25539 ;
  assign y11162 = ~1'b0 ;
  assign y11163 = ~1'b0 ;
  assign y11164 = ~n25543 ;
  assign y11165 = ~n25544 ;
  assign y11166 = ~n25547 ;
  assign y11167 = ~n25553 ;
  assign y11168 = ~n25554 ;
  assign y11169 = ~1'b0 ;
  assign y11170 = n25556 ;
  assign y11171 = n25557 ;
  assign y11172 = n25559 ;
  assign y11173 = ~1'b0 ;
  assign y11174 = ~1'b0 ;
  assign y11175 = ~1'b0 ;
  assign y11176 = ~n25566 ;
  assign y11177 = ~1'b0 ;
  assign y11178 = n25568 ;
  assign y11179 = ~n25573 ;
  assign y11180 = ~1'b0 ;
  assign y11181 = n25574 ;
  assign y11182 = ~n25575 ;
  assign y11183 = ~1'b0 ;
  assign y11184 = 1'b0 ;
  assign y11185 = ~1'b0 ;
  assign y11186 = ~n25579 ;
  assign y11187 = n25585 ;
  assign y11188 = ~1'b0 ;
  assign y11189 = ~1'b0 ;
  assign y11190 = n25586 ;
  assign y11191 = n25587 ;
  assign y11192 = ~n25592 ;
  assign y11193 = ~n25594 ;
  assign y11194 = n25597 ;
  assign y11195 = ~1'b0 ;
  assign y11196 = ~1'b0 ;
  assign y11197 = ~n25599 ;
  assign y11198 = ~1'b0 ;
  assign y11199 = ~1'b0 ;
  assign y11200 = n25600 ;
  assign y11201 = ~n25602 ;
  assign y11202 = n25606 ;
  assign y11203 = ~1'b0 ;
  assign y11204 = n25608 ;
  assign y11205 = ~n25610 ;
  assign y11206 = ~1'b0 ;
  assign y11207 = n25613 ;
  assign y11208 = ~1'b0 ;
  assign y11209 = 1'b0 ;
  assign y11210 = ~n25629 ;
  assign y11211 = n25634 ;
  assign y11212 = ~1'b0 ;
  assign y11213 = ~1'b0 ;
  assign y11214 = n25639 ;
  assign y11215 = ~n25643 ;
  assign y11216 = ~n25645 ;
  assign y11217 = n25647 ;
  assign y11218 = n25648 ;
  assign y11219 = ~n25652 ;
  assign y11220 = ~n25653 ;
  assign y11221 = ~1'b0 ;
  assign y11222 = ~1'b0 ;
  assign y11223 = n25657 ;
  assign y11224 = n25665 ;
  assign y11225 = 1'b0 ;
  assign y11226 = ~1'b0 ;
  assign y11227 = ~n25667 ;
  assign y11228 = ~n25672 ;
  assign y11229 = ~1'b0 ;
  assign y11230 = ~1'b0 ;
  assign y11231 = ~n25675 ;
  assign y11232 = ~n25677 ;
  assign y11233 = n25680 ;
  assign y11234 = ~n25681 ;
  assign y11235 = n25683 ;
  assign y11236 = n25689 ;
  assign y11237 = ~1'b0 ;
  assign y11238 = n25691 ;
  assign y11239 = ~n25698 ;
  assign y11240 = n25700 ;
  assign y11241 = ~1'b0 ;
  assign y11242 = n25702 ;
  assign y11243 = n16577 ;
  assign y11244 = ~n25703 ;
  assign y11245 = n25705 ;
  assign y11246 = n25706 ;
  assign y11247 = n25711 ;
  assign y11248 = ~n25716 ;
  assign y11249 = ~n25719 ;
  assign y11250 = ~1'b0 ;
  assign y11251 = n25721 ;
  assign y11252 = ~1'b0 ;
  assign y11253 = n25723 ;
  assign y11254 = ~n25724 ;
  assign y11255 = ~1'b0 ;
  assign y11256 = n25725 ;
  assign y11257 = ~n25727 ;
  assign y11258 = ~n25728 ;
  assign y11259 = n25731 ;
  assign y11260 = ~n25735 ;
  assign y11261 = n25736 ;
  assign y11262 = ~n25741 ;
  assign y11263 = n25742 ;
  assign y11264 = n25745 ;
  assign y11265 = n25752 ;
  assign y11266 = n25753 ;
  assign y11267 = n25757 ;
  assign y11268 = ~n25759 ;
  assign y11269 = n25762 ;
  assign y11270 = ~n25768 ;
  assign y11271 = ~n25769 ;
  assign y11272 = ~1'b0 ;
  assign y11273 = n906 ;
  assign y11274 = ~1'b0 ;
  assign y11275 = ~n25777 ;
  assign y11276 = ~n25779 ;
  assign y11277 = n25785 ;
  assign y11278 = ~n25786 ;
  assign y11279 = ~n25787 ;
  assign y11280 = ~n25789 ;
  assign y11281 = ~n24706 ;
  assign y11282 = n25794 ;
  assign y11283 = ~n25795 ;
  assign y11284 = ~n25796 ;
  assign y11285 = ~n25804 ;
  assign y11286 = ~1'b0 ;
  assign y11287 = ~n25805 ;
  assign y11288 = n25809 ;
  assign y11289 = n25810 ;
  assign y11290 = ~n25815 ;
  assign y11291 = ~n25816 ;
  assign y11292 = ~n25818 ;
  assign y11293 = ~1'b0 ;
  assign y11294 = n538 ;
  assign y11295 = n25819 ;
  assign y11296 = ~1'b0 ;
  assign y11297 = ~n25821 ;
  assign y11298 = n25822 ;
  assign y11299 = ~n25824 ;
  assign y11300 = ~1'b0 ;
  assign y11301 = n25826 ;
  assign y11302 = ~1'b0 ;
  assign y11303 = ~1'b0 ;
  assign y11304 = ~n25830 ;
  assign y11305 = ~n25831 ;
  assign y11306 = n4582 ;
  assign y11307 = 1'b0 ;
  assign y11308 = ~n25834 ;
  assign y11309 = n25320 ;
  assign y11310 = n25838 ;
  assign y11311 = ~1'b0 ;
  assign y11312 = ~n7756 ;
  assign y11313 = n25841 ;
  assign y11314 = ~n25845 ;
  assign y11315 = ~1'b0 ;
  assign y11316 = ~1'b0 ;
  assign y11317 = ~n25854 ;
  assign y11318 = n25855 ;
  assign y11319 = ~n18464 ;
  assign y11320 = n25856 ;
  assign y11321 = ~n25857 ;
  assign y11322 = n25860 ;
  assign y11323 = ~n25861 ;
  assign y11324 = ~n25862 ;
  assign y11325 = ~1'b0 ;
  assign y11326 = ~1'b0 ;
  assign y11327 = 1'b0 ;
  assign y11328 = ~n25863 ;
  assign y11329 = n25864 ;
  assign y11330 = ~n15124 ;
  assign y11331 = ~n25868 ;
  assign y11332 = ~n25869 ;
  assign y11333 = ~1'b0 ;
  assign y11334 = n25870 ;
  assign y11335 = ~n25872 ;
  assign y11336 = n25875 ;
  assign y11337 = n25878 ;
  assign y11338 = n6648 ;
  assign y11339 = n25882 ;
  assign y11340 = 1'b0 ;
  assign y11341 = ~n25884 ;
  assign y11342 = ~1'b0 ;
  assign y11343 = ~n25885 ;
  assign y11344 = n23588 ;
  assign y11345 = ~n25886 ;
  assign y11346 = n25888 ;
  assign y11347 = n25892 ;
  assign y11348 = ~n25893 ;
  assign y11349 = ~1'b0 ;
  assign y11350 = ~1'b0 ;
  assign y11351 = n25898 ;
  assign y11352 = n25900 ;
  assign y11353 = ~n25901 ;
  assign y11354 = ~1'b0 ;
  assign y11355 = ~n25903 ;
  assign y11356 = n25904 ;
  assign y11357 = ~1'b0 ;
  assign y11358 = ~1'b0 ;
  assign y11359 = n25908 ;
  assign y11360 = n25911 ;
  assign y11361 = ~n25912 ;
  assign y11362 = ~1'b0 ;
  assign y11363 = n25917 ;
  assign y11364 = ~n25921 ;
  assign y11365 = n25923 ;
  assign y11366 = ~n25924 ;
  assign y11367 = n25926 ;
  assign y11368 = n25934 ;
  assign y11369 = n25937 ;
  assign y11370 = n25938 ;
  assign y11371 = n25940 ;
  assign y11372 = n25955 ;
  assign y11373 = ~n25957 ;
  assign y11374 = n25958 ;
  assign y11375 = n25962 ;
  assign y11376 = n25966 ;
  assign y11377 = n25972 ;
  assign y11378 = ~n25976 ;
  assign y11379 = ~n25977 ;
  assign y11380 = ~1'b0 ;
  assign y11381 = ~1'b0 ;
  assign y11382 = n25978 ;
  assign y11383 = ~n25980 ;
  assign y11384 = ~n25981 ;
  assign y11385 = ~n25984 ;
  assign y11386 = ~1'b0 ;
  assign y11387 = n25985 ;
  assign y11388 = n25987 ;
  assign y11389 = ~n25991 ;
  assign y11390 = ~n25992 ;
  assign y11391 = ~n25998 ;
  assign y11392 = n26002 ;
  assign y11393 = n26012 ;
  assign y11394 = ~n26013 ;
  assign y11395 = ~1'b0 ;
  assign y11396 = ~n26015 ;
  assign y11397 = n26016 ;
  assign y11398 = ~n26017 ;
  assign y11399 = n26018 ;
  assign y11400 = n26020 ;
  assign y11401 = ~n26022 ;
  assign y11402 = ~n26023 ;
  assign y11403 = ~n26025 ;
  assign y11404 = 1'b0 ;
  assign y11405 = n26027 ;
  assign y11406 = n26028 ;
  assign y11407 = ~1'b0 ;
  assign y11408 = n26033 ;
  assign y11409 = n26034 ;
  assign y11410 = ~n26036 ;
  assign y11411 = ~n26041 ;
  assign y11412 = ~n26043 ;
  assign y11413 = n26049 ;
  assign y11414 = n26050 ;
  assign y11415 = ~1'b0 ;
  assign y11416 = n26051 ;
  assign y11417 = ~n26053 ;
  assign y11418 = ~1'b0 ;
  assign y11419 = n26056 ;
  assign y11420 = ~n26061 ;
  assign y11421 = n26063 ;
  assign y11422 = n26064 ;
  assign y11423 = ~1'b0 ;
  assign y11424 = ~n26065 ;
  assign y11425 = ~n26066 ;
  assign y11426 = n26067 ;
  assign y11427 = n26070 ;
  assign y11428 = n26072 ;
  assign y11429 = ~1'b0 ;
  assign y11430 = n26073 ;
  assign y11431 = n26076 ;
  assign y11432 = ~1'b0 ;
  assign y11433 = n26078 ;
  assign y11434 = n26086 ;
  assign y11435 = ~n26091 ;
  assign y11436 = n26093 ;
  assign y11437 = n26098 ;
  assign y11438 = 1'b0 ;
  assign y11439 = ~1'b0 ;
  assign y11440 = n26101 ;
  assign y11441 = ~1'b0 ;
  assign y11442 = ~n26102 ;
  assign y11443 = ~n26105 ;
  assign y11444 = ~n26106 ;
  assign y11445 = n26108 ;
  assign y11446 = n26109 ;
  assign y11447 = n26114 ;
  assign y11448 = ~n12393 ;
  assign y11449 = ~n26116 ;
  assign y11450 = ~n26117 ;
  assign y11451 = ~1'b0 ;
  assign y11452 = ~1'b0 ;
  assign y11453 = n26121 ;
  assign y11454 = ~1'b0 ;
  assign y11455 = ~1'b0 ;
  assign y11456 = n24175 ;
  assign y11457 = n26123 ;
  assign y11458 = ~n26127 ;
  assign y11459 = n26130 ;
  assign y11460 = ~n26134 ;
  assign y11461 = ~n26136 ;
  assign y11462 = ~n26140 ;
  assign y11463 = ~1'b0 ;
  assign y11464 = ~n26142 ;
  assign y11465 = ~1'b0 ;
  assign y11466 = ~n26147 ;
  assign y11467 = ~1'b0 ;
  assign y11468 = ~n26149 ;
  assign y11469 = n26151 ;
  assign y11470 = ~n26153 ;
  assign y11471 = n26159 ;
  assign y11472 = n26165 ;
  assign y11473 = n26166 ;
  assign y11474 = ~n26173 ;
  assign y11475 = ~n26176 ;
  assign y11476 = ~n26182 ;
  assign y11477 = ~1'b0 ;
  assign y11478 = n26188 ;
  assign y11479 = ~n26189 ;
  assign y11480 = ~n26206 ;
  assign y11481 = ~n26208 ;
  assign y11482 = ~1'b0 ;
  assign y11483 = n26211 ;
  assign y11484 = ~n26212 ;
  assign y11485 = ~1'b0 ;
  assign y11486 = 1'b0 ;
  assign y11487 = ~1'b0 ;
  assign y11488 = n26215 ;
  assign y11489 = n26216 ;
  assign y11490 = ~1'b0 ;
  assign y11491 = n22854 ;
  assign y11492 = n26221 ;
  assign y11493 = n26222 ;
  assign y11494 = ~n26225 ;
  assign y11495 = n26228 ;
  assign y11496 = n14599 ;
  assign y11497 = ~1'b0 ;
  assign y11498 = n26230 ;
  assign y11499 = n26231 ;
  assign y11500 = ~n26233 ;
  assign y11501 = n26237 ;
  assign y11502 = ~n26239 ;
  assign y11503 = ~1'b0 ;
  assign y11504 = ~n26241 ;
  assign y11505 = n26242 ;
  assign y11506 = ~1'b0 ;
  assign y11507 = ~1'b0 ;
  assign y11508 = ~n26244 ;
  assign y11509 = n26246 ;
  assign y11510 = ~1'b0 ;
  assign y11511 = ~1'b0 ;
  assign y11512 = n26250 ;
  assign y11513 = n26252 ;
  assign y11514 = n26253 ;
  assign y11515 = ~n26256 ;
  assign y11516 = n26257 ;
  assign y11517 = ~1'b0 ;
  assign y11518 = ~n26261 ;
  assign y11519 = ~n26263 ;
  assign y11520 = ~n26267 ;
  assign y11521 = ~1'b0 ;
  assign y11522 = n26269 ;
  assign y11523 = n26270 ;
  assign y11524 = ~n26271 ;
  assign y11525 = ~1'b0 ;
  assign y11526 = ~1'b0 ;
  assign y11527 = n26277 ;
  assign y11528 = n26280 ;
  assign y11529 = ~n26284 ;
  assign y11530 = ~n26286 ;
  assign y11531 = n26288 ;
  assign y11532 = n26292 ;
  assign y11533 = ~1'b0 ;
  assign y11534 = n26293 ;
  assign y11535 = ~1'b0 ;
  assign y11536 = ~1'b0 ;
  assign y11537 = n26295 ;
  assign y11538 = n26303 ;
  assign y11539 = 1'b0 ;
  assign y11540 = n24532 ;
  assign y11541 = ~n26307 ;
  assign y11542 = n26310 ;
  assign y11543 = ~1'b0 ;
  assign y11544 = ~1'b0 ;
  assign y11545 = ~n26311 ;
  assign y11546 = ~n26313 ;
  assign y11547 = n26315 ;
  assign y11548 = ~1'b0 ;
  assign y11549 = ~1'b0 ;
  assign y11550 = n26319 ;
  assign y11551 = ~n26322 ;
  assign y11552 = n9224 ;
  assign y11553 = ~n26323 ;
  assign y11554 = ~n14703 ;
  assign y11555 = n26325 ;
  assign y11556 = ~1'b0 ;
  assign y11557 = 1'b0 ;
  assign y11558 = n26327 ;
  assign y11559 = n26329 ;
  assign y11560 = ~n26331 ;
  assign y11561 = ~1'b0 ;
  assign y11562 = n26332 ;
  assign y11563 = ~1'b0 ;
  assign y11564 = ~n26337 ;
  assign y11565 = ~n26338 ;
  assign y11566 = ~n26342 ;
  assign y11567 = ~1'b0 ;
  assign y11568 = n26343 ;
  assign y11569 = ~n26344 ;
  assign y11570 = 1'b0 ;
  assign y11571 = n26346 ;
  assign y11572 = ~1'b0 ;
  assign y11573 = ~n26349 ;
  assign y11574 = ~n26355 ;
  assign y11575 = n26357 ;
  assign y11576 = n26364 ;
  assign y11577 = ~n5300 ;
  assign y11578 = ~n26365 ;
  assign y11579 = n26369 ;
  assign y11580 = ~n26370 ;
  assign y11581 = ~1'b0 ;
  assign y11582 = ~n26378 ;
  assign y11583 = ~n26380 ;
  assign y11584 = n26382 ;
  assign y11585 = ~n26384 ;
  assign y11586 = ~n26389 ;
  assign y11587 = ~1'b0 ;
  assign y11588 = ~1'b0 ;
  assign y11589 = ~1'b0 ;
  assign y11590 = ~n26390 ;
  assign y11591 = n6361 ;
  assign y11592 = ~n26393 ;
  assign y11593 = ~1'b0 ;
  assign y11594 = ~1'b0 ;
  assign y11595 = n26397 ;
  assign y11596 = ~n26399 ;
  assign y11597 = 1'b0 ;
  assign y11598 = ~n26401 ;
  assign y11599 = n1164 ;
  assign y11600 = ~1'b0 ;
  assign y11601 = ~1'b0 ;
  assign y11602 = ~n26408 ;
  assign y11603 = n26411 ;
  assign y11604 = n26412 ;
  assign y11605 = n26414 ;
  assign y11606 = ~n26418 ;
  assign y11607 = n26419 ;
  assign y11608 = n26421 ;
  assign y11609 = n16006 ;
  assign y11610 = n26423 ;
  assign y11611 = ~1'b0 ;
  assign y11612 = ~n26428 ;
  assign y11613 = n26429 ;
  assign y11614 = ~1'b0 ;
  assign y11615 = n26431 ;
  assign y11616 = n26432 ;
  assign y11617 = ~1'b0 ;
  assign y11618 = ~n26434 ;
  assign y11619 = n26436 ;
  assign y11620 = ~n26437 ;
  assign y11621 = ~n26438 ;
  assign y11622 = ~1'b0 ;
  assign y11623 = n26439 ;
  assign y11624 = n26444 ;
  assign y11625 = n9974 ;
  assign y11626 = ~1'b0 ;
  assign y11627 = n26452 ;
  assign y11628 = ~n26454 ;
  assign y11629 = ~1'b0 ;
  assign y11630 = ~n26459 ;
  assign y11631 = n26464 ;
  assign y11632 = n26472 ;
  assign y11633 = ~n26474 ;
  assign y11634 = ~1'b0 ;
  assign y11635 = ~1'b0 ;
  assign y11636 = n26475 ;
  assign y11637 = n25729 ;
  assign y11638 = n26476 ;
  assign y11639 = n26479 ;
  assign y11640 = ~n26481 ;
  assign y11641 = n26486 ;
  assign y11642 = ~n26497 ;
  assign y11643 = ~n26498 ;
  assign y11644 = n26499 ;
  assign y11645 = ~1'b0 ;
  assign y11646 = ~1'b0 ;
  assign y11647 = ~n26500 ;
  assign y11648 = ~n26502 ;
  assign y11649 = ~n26506 ;
  assign y11650 = n26511 ;
  assign y11651 = ~1'b0 ;
  assign y11652 = n26512 ;
  assign y11653 = ~n26513 ;
  assign y11654 = n26514 ;
  assign y11655 = n26516 ;
  assign y11656 = ~1'b0 ;
  assign y11657 = ~1'b0 ;
  assign y11658 = n26517 ;
  assign y11659 = n26521 ;
  assign y11660 = n26528 ;
  assign y11661 = n26530 ;
  assign y11662 = ~n26537 ;
  assign y11663 = ~n26543 ;
  assign y11664 = n26551 ;
  assign y11665 = n26552 ;
  assign y11666 = n26553 ;
  assign y11667 = ~n26555 ;
  assign y11668 = n26569 ;
  assign y11669 = ~1'b0 ;
  assign y11670 = ~n26572 ;
  assign y11671 = ~n26582 ;
  assign y11672 = n26583 ;
  assign y11673 = ~n26585 ;
  assign y11674 = ~n26587 ;
  assign y11675 = n26589 ;
  assign y11676 = n26597 ;
  assign y11677 = ~n26599 ;
  assign y11678 = ~n26608 ;
  assign y11679 = 1'b0 ;
  assign y11680 = n26611 ;
  assign y11681 = ~n26624 ;
  assign y11682 = n26625 ;
  assign y11683 = ~n12474 ;
  assign y11684 = ~1'b0 ;
  assign y11685 = ~1'b0 ;
  assign y11686 = n26627 ;
  assign y11687 = n26630 ;
  assign y11688 = ~1'b0 ;
  assign y11689 = ~n26631 ;
  assign y11690 = ~n26633 ;
  assign y11691 = ~1'b0 ;
  assign y11692 = 1'b0 ;
  assign y11693 = n26634 ;
  assign y11694 = n26638 ;
  assign y11695 = ~n1707 ;
  assign y11696 = ~1'b0 ;
  assign y11697 = ~1'b0 ;
  assign y11698 = ~1'b0 ;
  assign y11699 = 1'b0 ;
  assign y11700 = n26639 ;
  assign y11701 = ~n26644 ;
  assign y11702 = n26648 ;
  assign y11703 = n26651 ;
  assign y11704 = ~n26654 ;
  assign y11705 = n26655 ;
  assign y11706 = n7846 ;
  assign y11707 = ~1'b0 ;
  assign y11708 = ~n26662 ;
  assign y11709 = ~n26670 ;
  assign y11710 = ~1'b0 ;
  assign y11711 = ~n26672 ;
  assign y11712 = n26673 ;
  assign y11713 = ~n26675 ;
  assign y11714 = ~n26677 ;
  assign y11715 = ~n26679 ;
  assign y11716 = n26682 ;
  assign y11717 = ~n26686 ;
  assign y11718 = ~n15657 ;
  assign y11719 = ~1'b0 ;
  assign y11720 = n26687 ;
  assign y11721 = ~1'b0 ;
  assign y11722 = ~n26695 ;
  assign y11723 = ~n26697 ;
  assign y11724 = ~1'b0 ;
  assign y11725 = ~n26699 ;
  assign y11726 = ~n26708 ;
  assign y11727 = n26710 ;
  assign y11728 = n26712 ;
  assign y11729 = ~n26714 ;
  assign y11730 = ~1'b0 ;
  assign y11731 = ~n26715 ;
  assign y11732 = ~1'b0 ;
  assign y11733 = 1'b0 ;
  assign y11734 = ~n26717 ;
  assign y11735 = n26719 ;
  assign y11736 = n26721 ;
  assign y11737 = n26734 ;
  assign y11738 = n26735 ;
  assign y11739 = n26736 ;
  assign y11740 = n19151 ;
  assign y11741 = ~n26738 ;
  assign y11742 = n26742 ;
  assign y11743 = ~n26745 ;
  assign y11744 = ~n26747 ;
  assign y11745 = ~n26748 ;
  assign y11746 = ~1'b0 ;
  assign y11747 = ~1'b0 ;
  assign y11748 = ~n26753 ;
  assign y11749 = ~1'b0 ;
  assign y11750 = n26755 ;
  assign y11751 = ~n26756 ;
  assign y11752 = n26759 ;
  assign y11753 = ~n19486 ;
  assign y11754 = ~n26761 ;
  assign y11755 = n7937 ;
  assign y11756 = ~n26763 ;
  assign y11757 = ~n26766 ;
  assign y11758 = n26770 ;
  assign y11759 = ~1'b0 ;
  assign y11760 = ~n26772 ;
  assign y11761 = ~1'b0 ;
  assign y11762 = n26775 ;
  assign y11763 = ~n26776 ;
  assign y11764 = n26785 ;
  assign y11765 = ~1'b0 ;
  assign y11766 = n26786 ;
  assign y11767 = n26795 ;
  assign y11768 = ~n26796 ;
  assign y11769 = n26797 ;
  assign y11770 = n26802 ;
  assign y11771 = ~n26807 ;
  assign y11772 = ~n26808 ;
  assign y11773 = ~n26812 ;
  assign y11774 = ~n26819 ;
  assign y11775 = n26820 ;
  assign y11776 = ~n26824 ;
  assign y11777 = ~1'b0 ;
  assign y11778 = ~1'b0 ;
  assign y11779 = ~1'b0 ;
  assign y11780 = ~1'b0 ;
  assign y11781 = ~1'b0 ;
  assign y11782 = ~n26826 ;
  assign y11783 = n26828 ;
  assign y11784 = ~1'b0 ;
  assign y11785 = ~n26831 ;
  assign y11786 = ~n26832 ;
  assign y11787 = ~1'b0 ;
  assign y11788 = n14629 ;
  assign y11789 = ~1'b0 ;
  assign y11790 = ~n26833 ;
  assign y11791 = ~n26835 ;
  assign y11792 = ~n26840 ;
  assign y11793 = n26841 ;
  assign y11794 = ~n26845 ;
  assign y11795 = n26847 ;
  assign y11796 = n26849 ;
  assign y11797 = n26856 ;
  assign y11798 = n26857 ;
  assign y11799 = n26858 ;
  assign y11800 = ~1'b0 ;
  assign y11801 = n26860 ;
  assign y11802 = n26861 ;
  assign y11803 = n5509 ;
  assign y11804 = n26862 ;
  assign y11805 = ~n26864 ;
  assign y11806 = ~n26865 ;
  assign y11807 = ~1'b0 ;
  assign y11808 = ~1'b0 ;
  assign y11809 = ~n26869 ;
  assign y11810 = ~1'b0 ;
  assign y11811 = ~n26881 ;
  assign y11812 = n26886 ;
  assign y11813 = ~n26891 ;
  assign y11814 = ~n26901 ;
  assign y11815 = ~n26902 ;
  assign y11816 = ~n26904 ;
  assign y11817 = 1'b0 ;
  assign y11818 = ~n26914 ;
  assign y11819 = ~n26915 ;
  assign y11820 = ~1'b0 ;
  assign y11821 = ~n26919 ;
  assign y11822 = ~n26920 ;
  assign y11823 = ~n2142 ;
  assign y11824 = n26923 ;
  assign y11825 = ~1'b0 ;
  assign y11826 = ~n26925 ;
  assign y11827 = ~n26927 ;
  assign y11828 = n26929 ;
  assign y11829 = n26931 ;
  assign y11830 = n26936 ;
  assign y11831 = n26938 ;
  assign y11832 = n26941 ;
  assign y11833 = n26942 ;
  assign y11834 = n26943 ;
  assign y11835 = ~n26947 ;
  assign y11836 = n26949 ;
  assign y11837 = ~n26954 ;
  assign y11838 = ~1'b0 ;
  assign y11839 = ~1'b0 ;
  assign y11840 = ~n26957 ;
  assign y11841 = ~n26960 ;
  assign y11842 = n26965 ;
  assign y11843 = ~n26967 ;
  assign y11844 = ~n26971 ;
  assign y11845 = n26973 ;
  assign y11846 = n26974 ;
  assign y11847 = n26978 ;
  assign y11848 = ~1'b0 ;
  assign y11849 = ~n26979 ;
  assign y11850 = ~1'b0 ;
  assign y11851 = n26981 ;
  assign y11852 = n14424 ;
  assign y11853 = ~n26983 ;
  assign y11854 = ~n26984 ;
  assign y11855 = ~n26985 ;
  assign y11856 = ~n26986 ;
  assign y11857 = ~n26989 ;
  assign y11858 = ~n26993 ;
  assign y11859 = ~n13903 ;
  assign y11860 = ~n26994 ;
  assign y11861 = ~n26995 ;
  assign y11862 = ~1'b0 ;
  assign y11863 = ~n26996 ;
  assign y11864 = ~1'b0 ;
  assign y11865 = ~n27004 ;
  assign y11866 = ~n27005 ;
  assign y11867 = ~n27006 ;
  assign y11868 = ~1'b0 ;
  assign y11869 = ~1'b0 ;
  assign y11870 = ~1'b0 ;
  assign y11871 = ~n27009 ;
  assign y11872 = n19934 ;
  assign y11873 = ~n27017 ;
  assign y11874 = n27018 ;
  assign y11875 = ~n27022 ;
  assign y11876 = n9810 ;
  assign y11877 = n27023 ;
  assign y11878 = n27026 ;
  assign y11879 = ~1'b0 ;
  assign y11880 = ~n27027 ;
  assign y11881 = ~1'b0 ;
  assign y11882 = ~1'b0 ;
  assign y11883 = 1'b0 ;
  assign y11884 = ~n10543 ;
  assign y11885 = ~n27028 ;
  assign y11886 = ~n27032 ;
  assign y11887 = n27035 ;
  assign y11888 = n25193 ;
  assign y11889 = n27037 ;
  assign y11890 = n27039 ;
  assign y11891 = ~n27047 ;
  assign y11892 = n27050 ;
  assign y11893 = ~n27054 ;
  assign y11894 = ~1'b0 ;
  assign y11895 = ~n27059 ;
  assign y11896 = ~1'b0 ;
  assign y11897 = ~n27060 ;
  assign y11898 = ~n27063 ;
  assign y11899 = n27064 ;
  assign y11900 = ~n27066 ;
  assign y11901 = ~1'b0 ;
  assign y11902 = ~n27069 ;
  assign y11903 = ~n27073 ;
  assign y11904 = ~n27077 ;
  assign y11905 = ~1'b0 ;
  assign y11906 = n27079 ;
  assign y11907 = ~1'b0 ;
  assign y11908 = ~1'b0 ;
  assign y11909 = ~1'b0 ;
  assign y11910 = ~1'b0 ;
  assign y11911 = ~n5229 ;
  assign y11912 = ~n27080 ;
  assign y11913 = ~1'b0 ;
  assign y11914 = n27082 ;
  assign y11915 = ~1'b0 ;
  assign y11916 = ~1'b0 ;
  assign y11917 = n27088 ;
  assign y11918 = n27091 ;
  assign y11919 = ~n27093 ;
  assign y11920 = ~n27102 ;
  assign y11921 = n27103 ;
  assign y11922 = ~n27105 ;
  assign y11923 = ~n27107 ;
  assign y11924 = n27109 ;
  assign y11925 = n27115 ;
  assign y11926 = n27118 ;
  assign y11927 = n27122 ;
  assign y11928 = n27128 ;
  assign y11929 = ~n27129 ;
  assign y11930 = ~n27132 ;
  assign y11931 = n27138 ;
  assign y11932 = ~1'b0 ;
  assign y11933 = ~1'b0 ;
  assign y11934 = ~n27139 ;
  assign y11935 = ~1'b0 ;
  assign y11936 = ~1'b0 ;
  assign y11937 = ~n27146 ;
  assign y11938 = ~1'b0 ;
  assign y11939 = ~1'b0 ;
  assign y11940 = ~n27149 ;
  assign y11941 = ~1'b0 ;
  assign y11942 = n27150 ;
  assign y11943 = ~1'b0 ;
  assign y11944 = n27152 ;
  assign y11945 = ~1'b0 ;
  assign y11946 = ~n27157 ;
  assign y11947 = 1'b0 ;
  assign y11948 = n27162 ;
  assign y11949 = n27164 ;
  assign y11950 = n27168 ;
  assign y11951 = ~1'b0 ;
  assign y11952 = n27172 ;
  assign y11953 = n27174 ;
  assign y11954 = ~n27176 ;
  assign y11955 = n27178 ;
  assign y11956 = ~n27179 ;
  assign y11957 = ~1'b0 ;
  assign y11958 = n27180 ;
  assign y11959 = n27186 ;
  assign y11960 = ~n27188 ;
  assign y11961 = n14777 ;
  assign y11962 = ~n11926 ;
  assign y11963 = ~n27189 ;
  assign y11964 = n27192 ;
  assign y11965 = n27200 ;
  assign y11966 = n27201 ;
  assign y11967 = ~1'b0 ;
  assign y11968 = ~1'b0 ;
  assign y11969 = ~1'b0 ;
  assign y11970 = ~1'b0 ;
  assign y11971 = ~1'b0 ;
  assign y11972 = ~n27209 ;
  assign y11973 = n27211 ;
  assign y11974 = n27212 ;
  assign y11975 = ~n27217 ;
  assign y11976 = ~1'b0 ;
  assign y11977 = ~1'b0 ;
  assign y11978 = ~n27218 ;
  assign y11979 = n17954 ;
  assign y11980 = n27221 ;
  assign y11981 = ~1'b0 ;
  assign y11982 = n27225 ;
  assign y11983 = ~n27227 ;
  assign y11984 = ~1'b0 ;
  assign y11985 = ~n27228 ;
  assign y11986 = ~n27229 ;
  assign y11987 = n27232 ;
  assign y11988 = ~n27237 ;
  assign y11989 = ~1'b0 ;
  assign y11990 = n27240 ;
  assign y11991 = ~n2067 ;
  assign y11992 = n27242 ;
  assign y11993 = n27247 ;
  assign y11994 = ~1'b0 ;
  assign y11995 = ~n27250 ;
  assign y11996 = ~n27251 ;
  assign y11997 = ~1'b0 ;
  assign y11998 = n27255 ;
  assign y11999 = ~n27256 ;
  assign y12000 = n27257 ;
  assign y12001 = n27259 ;
  assign y12002 = ~n27262 ;
  assign y12003 = ~1'b0 ;
  assign y12004 = n27263 ;
  assign y12005 = n27269 ;
  assign y12006 = n27273 ;
  assign y12007 = n27280 ;
  assign y12008 = ~1'b0 ;
  assign y12009 = n22756 ;
  assign y12010 = n27281 ;
  assign y12011 = n27285 ;
  assign y12012 = ~1'b0 ;
  assign y12013 = ~n27293 ;
  assign y12014 = ~n27296 ;
  assign y12015 = ~n27297 ;
  assign y12016 = ~n27301 ;
  assign y12017 = ~1'b0 ;
  assign y12018 = n24862 ;
  assign y12019 = ~1'b0 ;
  assign y12020 = ~1'b0 ;
  assign y12021 = ~1'b0 ;
  assign y12022 = ~n27302 ;
  assign y12023 = ~1'b0 ;
  assign y12024 = ~n27303 ;
  assign y12025 = n27304 ;
  assign y12026 = n27305 ;
  assign y12027 = n27316 ;
  assign y12028 = n27320 ;
  assign y12029 = n27323 ;
  assign y12030 = n27324 ;
  assign y12031 = ~n27326 ;
  assign y12032 = ~n27327 ;
  assign y12033 = n27336 ;
  assign y12034 = ~1'b0 ;
  assign y12035 = ~n27337 ;
  assign y12036 = ~1'b0 ;
  assign y12037 = ~n27339 ;
  assign y12038 = ~n27341 ;
  assign y12039 = n27344 ;
  assign y12040 = ~n27348 ;
  assign y12041 = n27349 ;
  assign y12042 = ~1'b0 ;
  assign y12043 = ~n27351 ;
  assign y12044 = ~1'b0 ;
  assign y12045 = ~1'b0 ;
  assign y12046 = ~n27355 ;
  assign y12047 = ~n27357 ;
  assign y12048 = n11531 ;
  assign y12049 = n27360 ;
  assign y12050 = ~n27362 ;
  assign y12051 = ~1'b0 ;
  assign y12052 = ~n27363 ;
  assign y12053 = ~n27366 ;
  assign y12054 = ~n27368 ;
  assign y12055 = ~1'b0 ;
  assign y12056 = n27369 ;
  assign y12057 = ~n27370 ;
  assign y12058 = ~n27372 ;
  assign y12059 = ~1'b0 ;
  assign y12060 = n27373 ;
  assign y12061 = n27377 ;
  assign y12062 = n27379 ;
  assign y12063 = ~n27382 ;
  assign y12064 = ~n27387 ;
  assign y12065 = n27388 ;
  assign y12066 = n27391 ;
  assign y12067 = ~1'b0 ;
  assign y12068 = ~1'b0 ;
  assign y12069 = ~n27397 ;
  assign y12070 = n27399 ;
  assign y12071 = n27403 ;
  assign y12072 = ~1'b0 ;
  assign y12073 = n27404 ;
  assign y12074 = n27407 ;
  assign y12075 = n27410 ;
  assign y12076 = n27416 ;
  assign y12077 = ~n27419 ;
  assign y12078 = ~n27420 ;
  assign y12079 = ~n27427 ;
  assign y12080 = n27429 ;
  assign y12081 = n27430 ;
  assign y12082 = n27431 ;
  assign y12083 = ~n27434 ;
  assign y12084 = ~1'b0 ;
  assign y12085 = ~n27436 ;
  assign y12086 = n27440 ;
  assign y12087 = n27442 ;
  assign y12088 = ~n27448 ;
  assign y12089 = ~n27449 ;
  assign y12090 = ~1'b0 ;
  assign y12091 = ~n5620 ;
  assign y12092 = ~1'b0 ;
  assign y12093 = n27450 ;
  assign y12094 = ~1'b0 ;
  assign y12095 = ~1'b0 ;
  assign y12096 = ~n27451 ;
  assign y12097 = ~1'b0 ;
  assign y12098 = ~n27452 ;
  assign y12099 = ~n27454 ;
  assign y12100 = ~1'b0 ;
  assign y12101 = ~1'b0 ;
  assign y12102 = n27463 ;
  assign y12103 = n27467 ;
  assign y12104 = n27470 ;
  assign y12105 = 1'b0 ;
  assign y12106 = ~1'b0 ;
  assign y12107 = n27472 ;
  assign y12108 = ~n27473 ;
  assign y12109 = ~n27475 ;
  assign y12110 = n27476 ;
  assign y12111 = ~1'b0 ;
  assign y12112 = ~1'b0 ;
  assign y12113 = ~n27479 ;
  assign y12114 = ~n27483 ;
  assign y12115 = ~1'b0 ;
  assign y12116 = n27489 ;
  assign y12117 = ~1'b0 ;
  assign y12118 = n27490 ;
  assign y12119 = n27492 ;
  assign y12120 = ~1'b0 ;
  assign y12121 = n27494 ;
  assign y12122 = n27495 ;
  assign y12123 = ~n27498 ;
  assign y12124 = ~n27501 ;
  assign y12125 = n27502 ;
  assign y12126 = n27504 ;
  assign y12127 = 1'b0 ;
  assign y12128 = ~n27506 ;
  assign y12129 = ~n27509 ;
  assign y12130 = ~1'b0 ;
  assign y12131 = n27511 ;
  assign y12132 = n27512 ;
  assign y12133 = ~n27515 ;
  assign y12134 = ~n27516 ;
  assign y12135 = ~n27521 ;
  assign y12136 = ~1'b0 ;
  assign y12137 = 1'b0 ;
  assign y12138 = n27522 ;
  assign y12139 = ~1'b0 ;
  assign y12140 = ~n6690 ;
  assign y12141 = n27528 ;
  assign y12142 = n27530 ;
  assign y12143 = n27534 ;
  assign y12144 = ~n27535 ;
  assign y12145 = ~n27538 ;
  assign y12146 = ~1'b0 ;
  assign y12147 = ~1'b0 ;
  assign y12148 = ~n27539 ;
  assign y12149 = ~n27544 ;
  assign y12150 = n27550 ;
  assign y12151 = n27551 ;
  assign y12152 = n27552 ;
  assign y12153 = ~1'b0 ;
  assign y12154 = ~n27554 ;
  assign y12155 = n9442 ;
  assign y12156 = ~n27557 ;
  assign y12157 = ~1'b0 ;
  assign y12158 = ~1'b0 ;
  assign y12159 = n27559 ;
  assign y12160 = n27565 ;
  assign y12161 = ~n27566 ;
  assign y12162 = ~1'b0 ;
  assign y12163 = ~1'b0 ;
  assign y12164 = ~n27568 ;
  assign y12165 = ~n27573 ;
  assign y12166 = n27576 ;
  assign y12167 = ~n27580 ;
  assign y12168 = n27583 ;
  assign y12169 = ~1'b0 ;
  assign y12170 = ~n27584 ;
  assign y12171 = ~n23978 ;
  assign y12172 = ~1'b0 ;
  assign y12173 = ~n8945 ;
  assign y12174 = n25102 ;
  assign y12175 = ~n27585 ;
  assign y12176 = n27586 ;
  assign y12177 = ~1'b0 ;
  assign y12178 = ~n27587 ;
  assign y12179 = ~1'b0 ;
  assign y12180 = n27597 ;
  assign y12181 = n27599 ;
  assign y12182 = ~n27602 ;
  assign y12183 = n27607 ;
  assign y12184 = ~n27609 ;
  assign y12185 = n27610 ;
  assign y12186 = n27615 ;
  assign y12187 = ~1'b0 ;
  assign y12188 = ~n27616 ;
  assign y12189 = n27617 ;
  assign y12190 = ~1'b0 ;
  assign y12191 = n27618 ;
  assign y12192 = ~n27619 ;
  assign y12193 = n1805 ;
  assign y12194 = n27621 ;
  assign y12195 = ~n27624 ;
  assign y12196 = ~n9173 ;
  assign y12197 = ~n27631 ;
  assign y12198 = ~1'b0 ;
  assign y12199 = ~1'b0 ;
  assign y12200 = ~n27632 ;
  assign y12201 = n9055 ;
  assign y12202 = n24476 ;
  assign y12203 = ~1'b0 ;
  assign y12204 = ~n27635 ;
  assign y12205 = n27637 ;
  assign y12206 = ~1'b0 ;
  assign y12207 = n27644 ;
  assign y12208 = n27645 ;
  assign y12209 = ~n27648 ;
  assign y12210 = n27649 ;
  assign y12211 = ~1'b0 ;
  assign y12212 = ~n27655 ;
  assign y12213 = ~n27656 ;
  assign y12214 = n27664 ;
  assign y12215 = ~1'b0 ;
  assign y12216 = n27667 ;
  assign y12217 = ~n27668 ;
  assign y12218 = ~n27672 ;
  assign y12219 = ~1'b0 ;
  assign y12220 = n27673 ;
  assign y12221 = ~n27674 ;
  assign y12222 = ~n27676 ;
  assign y12223 = n23461 ;
  assign y12224 = 1'b0 ;
  assign y12225 = n27681 ;
  assign y12226 = ~n27683 ;
  assign y12227 = n27688 ;
  assign y12228 = ~n27690 ;
  assign y12229 = ~n27693 ;
  assign y12230 = ~1'b0 ;
  assign y12231 = ~1'b0 ;
  assign y12232 = ~1'b0 ;
  assign y12233 = ~n27694 ;
  assign y12234 = 1'b0 ;
  assign y12235 = ~n27701 ;
  assign y12236 = ~1'b0 ;
  assign y12237 = ~n27705 ;
  assign y12238 = ~1'b0 ;
  assign y12239 = ~n27708 ;
  assign y12240 = n27709 ;
  assign y12241 = ~1'b0 ;
  assign y12242 = ~n27710 ;
  assign y12243 = ~n27717 ;
  assign y12244 = ~n27719 ;
  assign y12245 = ~1'b0 ;
  assign y12246 = ~1'b0 ;
  assign y12247 = n27723 ;
  assign y12248 = ~1'b0 ;
  assign y12249 = 1'b0 ;
  assign y12250 = n27724 ;
  assign y12251 = ~n27725 ;
  assign y12252 = n27726 ;
  assign y12253 = ~n27727 ;
  assign y12254 = n27730 ;
  assign y12255 = ~n5822 ;
  assign y12256 = n27731 ;
  assign y12257 = ~1'b0 ;
  assign y12258 = n27734 ;
  assign y12259 = ~n27736 ;
  assign y12260 = n27737 ;
  assign y12261 = n27738 ;
  assign y12262 = ~n27742 ;
  assign y12263 = n27743 ;
  assign y12264 = ~n27745 ;
  assign y12265 = ~n27751 ;
  assign y12266 = ~n27755 ;
  assign y12267 = n27761 ;
  assign y12268 = n5102 ;
  assign y12269 = n26199 ;
  assign y12270 = ~n18868 ;
  assign y12271 = ~1'b0 ;
  assign y12272 = ~1'b0 ;
  assign y12273 = ~1'b0 ;
  assign y12274 = ~n27763 ;
  assign y12275 = ~1'b0 ;
  assign y12276 = n27764 ;
  assign y12277 = ~n27765 ;
  assign y12278 = ~n27767 ;
  assign y12279 = ~n27771 ;
  assign y12280 = n27773 ;
  assign y12281 = ~n27774 ;
  assign y12282 = n27775 ;
  assign y12283 = ~n27781 ;
  assign y12284 = ~n27786 ;
  assign y12285 = n27787 ;
  assign y12286 = n27790 ;
  assign y12287 = n27792 ;
  assign y12288 = ~n27796 ;
  assign y12289 = ~1'b0 ;
  assign y12290 = ~1'b0 ;
  assign y12291 = ~1'b0 ;
  assign y12292 = ~n27798 ;
  assign y12293 = ~n27800 ;
  assign y12294 = n27802 ;
  assign y12295 = ~n27804 ;
  assign y12296 = ~n27806 ;
  assign y12297 = ~1'b0 ;
  assign y12298 = ~1'b0 ;
  assign y12299 = ~n27809 ;
  assign y12300 = ~n27811 ;
  assign y12301 = n27815 ;
  assign y12302 = ~n27816 ;
  assign y12303 = ~n27820 ;
  assign y12304 = ~1'b0 ;
  assign y12305 = ~n27824 ;
  assign y12306 = ~n27825 ;
  assign y12307 = n27826 ;
  assign y12308 = n27827 ;
  assign y12309 = ~n27828 ;
  assign y12310 = ~n27830 ;
  assign y12311 = ~n27835 ;
  assign y12312 = ~n12850 ;
  assign y12313 = ~1'b0 ;
  assign y12314 = ~1'b0 ;
  assign y12315 = ~n27836 ;
  assign y12316 = ~1'b0 ;
  assign y12317 = n27838 ;
  assign y12318 = ~n27841 ;
  assign y12319 = ~1'b0 ;
  assign y12320 = n27843 ;
  assign y12321 = n27845 ;
  assign y12322 = n27846 ;
  assign y12323 = ~n27847 ;
  assign y12324 = n27848 ;
  assign y12325 = n27853 ;
  assign y12326 = ~1'b0 ;
  assign y12327 = ~n27855 ;
  assign y12328 = ~n27856 ;
  assign y12329 = n27858 ;
  assign y12330 = n27859 ;
  assign y12331 = n27862 ;
  assign y12332 = n27863 ;
  assign y12333 = ~n27867 ;
  assign y12334 = ~1'b0 ;
  assign y12335 = ~1'b0 ;
  assign y12336 = n27868 ;
  assign y12337 = n27870 ;
  assign y12338 = n27874 ;
  assign y12339 = n27875 ;
  assign y12340 = ~n27883 ;
  assign y12341 = ~n27884 ;
  assign y12342 = n27887 ;
  assign y12343 = n27891 ;
  assign y12344 = ~1'b0 ;
  assign y12345 = n27892 ;
  assign y12346 = ~n27899 ;
  assign y12347 = ~n27900 ;
  assign y12348 = ~n27912 ;
  assign y12349 = ~1'b0 ;
  assign y12350 = ~1'b0 ;
  assign y12351 = ~1'b0 ;
  assign y12352 = n27913 ;
  assign y12353 = ~n27919 ;
  assign y12354 = ~n27922 ;
  assign y12355 = ~1'b0 ;
  assign y12356 = n27924 ;
  assign y12357 = n27926 ;
  assign y12358 = ~1'b0 ;
  assign y12359 = ~1'b0 ;
  assign y12360 = n27927 ;
  assign y12361 = n27934 ;
  assign y12362 = ~1'b0 ;
  assign y12363 = ~1'b0 ;
  assign y12364 = n27935 ;
  assign y12365 = ~n27936 ;
  assign y12366 = n27938 ;
  assign y12367 = n27941 ;
  assign y12368 = n27948 ;
  assign y12369 = ~n27949 ;
  assign y12370 = n27954 ;
  assign y12371 = 1'b0 ;
  assign y12372 = n27958 ;
  assign y12373 = ~1'b0 ;
  assign y12374 = ~1'b0 ;
  assign y12375 = n21671 ;
  assign y12376 = n27959 ;
  assign y12377 = n27960 ;
  assign y12378 = n27961 ;
  assign y12379 = ~n27962 ;
  assign y12380 = ~1'b0 ;
  assign y12381 = ~1'b0 ;
  assign y12382 = ~n27965 ;
  assign y12383 = ~n27968 ;
  assign y12384 = n27971 ;
  assign y12385 = n2890 ;
  assign y12386 = ~1'b0 ;
  assign y12387 = ~n27975 ;
  assign y12388 = n27980 ;
  assign y12389 = ~1'b0 ;
  assign y12390 = n27983 ;
  assign y12391 = ~1'b0 ;
  assign y12392 = n27985 ;
  assign y12393 = n27986 ;
  assign y12394 = n27989 ;
  assign y12395 = ~n27990 ;
  assign y12396 = ~n27994 ;
  assign y12397 = n27995 ;
  assign y12398 = 1'b0 ;
  assign y12399 = ~n27997 ;
  assign y12400 = ~n27998 ;
  assign y12401 = ~n27999 ;
  assign y12402 = ~1'b0 ;
  assign y12403 = ~n28001 ;
  assign y12404 = n28002 ;
  assign y12405 = n28007 ;
  assign y12406 = ~n28010 ;
  assign y12407 = ~n28011 ;
  assign y12408 = ~1'b0 ;
  assign y12409 = n28012 ;
  assign y12410 = n28013 ;
  assign y12411 = ~n28014 ;
  assign y12412 = ~n28015 ;
  assign y12413 = ~n28018 ;
  assign y12414 = 1'b0 ;
  assign y12415 = ~1'b0 ;
  assign y12416 = ~n28021 ;
  assign y12417 = n28023 ;
  assign y12418 = ~n28026 ;
  assign y12419 = ~n28028 ;
  assign y12420 = n28029 ;
  assign y12421 = 1'b0 ;
  assign y12422 = n21377 ;
  assign y12423 = ~n28035 ;
  assign y12424 = ~n7374 ;
  assign y12425 = n28037 ;
  assign y12426 = ~1'b0 ;
  assign y12427 = n28038 ;
  assign y12428 = ~1'b0 ;
  assign y12429 = n3073 ;
  assign y12430 = n28048 ;
  assign y12431 = ~n28049 ;
  assign y12432 = ~n28050 ;
  assign y12433 = ~1'b0 ;
  assign y12434 = ~1'b0 ;
  assign y12435 = ~1'b0 ;
  assign y12436 = ~n28054 ;
  assign y12437 = n3626 ;
  assign y12438 = ~1'b0 ;
  assign y12439 = n28057 ;
  assign y12440 = ~n28060 ;
  assign y12441 = ~n28062 ;
  assign y12442 = ~n28064 ;
  assign y12443 = n28068 ;
  assign y12444 = ~n28074 ;
  assign y12445 = ~n23035 ;
  assign y12446 = ~1'b0 ;
  assign y12447 = n28078 ;
  assign y12448 = ~1'b0 ;
  assign y12449 = ~n28082 ;
  assign y12450 = n28093 ;
  assign y12451 = n28105 ;
  assign y12452 = ~n28111 ;
  assign y12453 = n28112 ;
  assign y12454 = ~1'b0 ;
  assign y12455 = ~1'b0 ;
  assign y12456 = n28115 ;
  assign y12457 = ~1'b0 ;
  assign y12458 = n28116 ;
  assign y12459 = ~n28119 ;
  assign y12460 = ~n28121 ;
  assign y12461 = n28122 ;
  assign y12462 = ~n28126 ;
  assign y12463 = ~n28128 ;
  assign y12464 = n28136 ;
  assign y12465 = n28139 ;
  assign y12466 = n28141 ;
  assign y12467 = ~1'b0 ;
  assign y12468 = ~n28144 ;
  assign y12469 = ~1'b0 ;
  assign y12470 = ~1'b0 ;
  assign y12471 = ~n28149 ;
  assign y12472 = ~n28152 ;
  assign y12473 = n28154 ;
  assign y12474 = ~n28161 ;
  assign y12475 = n28164 ;
  assign y12476 = ~n28166 ;
  assign y12477 = n28167 ;
  assign y12478 = n28171 ;
  assign y12479 = n28172 ;
  assign y12480 = n28173 ;
  assign y12481 = n28175 ;
  assign y12482 = ~n28176 ;
  assign y12483 = n28179 ;
  assign y12484 = ~n28182 ;
  assign y12485 = n28184 ;
  assign y12486 = ~1'b0 ;
  assign y12487 = ~n28187 ;
  assign y12488 = n28189 ;
  assign y12489 = n28191 ;
  assign y12490 = n28192 ;
  assign y12491 = n28193 ;
  assign y12492 = ~n28194 ;
  assign y12493 = ~1'b0 ;
  assign y12494 = ~1'b0 ;
  assign y12495 = ~1'b0 ;
  assign y12496 = n28196 ;
  assign y12497 = n28203 ;
  assign y12498 = n28204 ;
  assign y12499 = n28205 ;
  assign y12500 = ~1'b0 ;
  assign y12501 = ~1'b0 ;
  assign y12502 = ~n28206 ;
  assign y12503 = ~1'b0 ;
  assign y12504 = ~n28210 ;
  assign y12505 = ~n28213 ;
  assign y12506 = n28214 ;
  assign y12507 = ~1'b0 ;
  assign y12508 = ~n28215 ;
  assign y12509 = ~n6613 ;
  assign y12510 = ~n28219 ;
  assign y12511 = ~n28220 ;
  assign y12512 = n28221 ;
  assign y12513 = ~n28223 ;
  assign y12514 = ~n28224 ;
  assign y12515 = n28226 ;
  assign y12516 = ~n28228 ;
  assign y12517 = n28229 ;
  assign y12518 = ~n28230 ;
  assign y12519 = ~n28234 ;
  assign y12520 = ~n28236 ;
  assign y12521 = 1'b0 ;
  assign y12522 = n28240 ;
  assign y12523 = ~n28242 ;
  assign y12524 = ~1'b0 ;
  assign y12525 = n28244 ;
  assign y12526 = ~n28247 ;
  assign y12527 = ~n7460 ;
  assign y12528 = ~1'b0 ;
  assign y12529 = ~n28254 ;
  assign y12530 = n28256 ;
  assign y12531 = n28262 ;
  assign y12532 = ~1'b0 ;
  assign y12533 = n28264 ;
  assign y12534 = ~n28266 ;
  assign y12535 = ~n28267 ;
  assign y12536 = ~n28269 ;
  assign y12537 = ~n27951 ;
  assign y12538 = ~1'b0 ;
  assign y12539 = ~n28279 ;
  assign y12540 = n28280 ;
  assign y12541 = n28288 ;
  assign y12542 = n28293 ;
  assign y12543 = n28305 ;
  assign y12544 = n28308 ;
  assign y12545 = n28311 ;
  assign y12546 = n28313 ;
  assign y12547 = ~n28317 ;
  assign y12548 = n28318 ;
  assign y12549 = n7781 ;
  assign y12550 = n28322 ;
  assign y12551 = ~n28326 ;
  assign y12552 = n28332 ;
  assign y12553 = ~n28333 ;
  assign y12554 = ~1'b0 ;
  assign y12555 = ~n12157 ;
  assign y12556 = ~n28335 ;
  assign y12557 = ~n28336 ;
  assign y12558 = ~n28337 ;
  assign y12559 = ~1'b0 ;
  assign y12560 = ~n28343 ;
  assign y12561 = ~1'b0 ;
  assign y12562 = ~1'b0 ;
  assign y12563 = n28348 ;
  assign y12564 = ~n28351 ;
  assign y12565 = ~n28352 ;
  assign y12566 = n271 ;
  assign y12567 = 1'b0 ;
  assign y12568 = ~n28353 ;
  assign y12569 = ~1'b0 ;
  assign y12570 = ~n28354 ;
  assign y12571 = n28355 ;
  assign y12572 = n28356 ;
  assign y12573 = ~n28357 ;
  assign y12574 = ~n28359 ;
  assign y12575 = ~1'b0 ;
  assign y12576 = ~n28360 ;
  assign y12577 = n28362 ;
  assign y12578 = ~n28363 ;
  assign y12579 = n28366 ;
  assign y12580 = ~n28369 ;
  assign y12581 = n28371 ;
  assign y12582 = n28373 ;
  assign y12583 = n28374 ;
  assign y12584 = n26043 ;
  assign y12585 = n28378 ;
  assign y12586 = ~n28379 ;
  assign y12587 = ~n28381 ;
  assign y12588 = n5327 ;
  assign y12589 = ~n28382 ;
  assign y12590 = ~n28387 ;
  assign y12591 = ~n28388 ;
  assign y12592 = 1'b0 ;
  assign y12593 = ~1'b0 ;
  assign y12594 = ~n28390 ;
  assign y12595 = ~n28392 ;
  assign y12596 = ~n28393 ;
  assign y12597 = n28398 ;
  assign y12598 = ~n28401 ;
  assign y12599 = n28403 ;
  assign y12600 = ~n28405 ;
  assign y12601 = ~1'b0 ;
  assign y12602 = ~n806 ;
  assign y12603 = n28406 ;
  assign y12604 = n28412 ;
  assign y12605 = ~n28414 ;
  assign y12606 = ~n6683 ;
  assign y12607 = n28415 ;
  assign y12608 = ~n28416 ;
  assign y12609 = ~1'b0 ;
  assign y12610 = n28423 ;
  assign y12611 = ~n28424 ;
  assign y12612 = 1'b0 ;
  assign y12613 = ~n28428 ;
  assign y12614 = ~n28430 ;
  assign y12615 = ~1'b0 ;
  assign y12616 = ~1'b0 ;
  assign y12617 = n28431 ;
  assign y12618 = n28434 ;
  assign y12619 = n28439 ;
  assign y12620 = ~n28441 ;
  assign y12621 = n28444 ;
  assign y12622 = ~n28445 ;
  assign y12623 = ~1'b0 ;
  assign y12624 = ~n28446 ;
  assign y12625 = ~n28448 ;
  assign y12626 = ~1'b0 ;
  assign y12627 = ~n28450 ;
  assign y12628 = ~n28451 ;
  assign y12629 = ~n28454 ;
  assign y12630 = ~n28459 ;
  assign y12631 = ~1'b0 ;
  assign y12632 = ~n28465 ;
  assign y12633 = n28467 ;
  assign y12634 = ~1'b0 ;
  assign y12635 = ~1'b0 ;
  assign y12636 = n28468 ;
  assign y12637 = n28469 ;
  assign y12638 = n28472 ;
  assign y12639 = ~1'b0 ;
  assign y12640 = ~n28475 ;
  assign y12641 = ~1'b0 ;
  assign y12642 = ~n28477 ;
  assign y12643 = n28483 ;
  assign y12644 = n28484 ;
  assign y12645 = n28487 ;
  assign y12646 = n28491 ;
  assign y12647 = 1'b0 ;
  assign y12648 = n28492 ;
  assign y12649 = ~n28493 ;
  assign y12650 = n28497 ;
  assign y12651 = ~1'b0 ;
  assign y12652 = n5304 ;
  assign y12653 = n28498 ;
  assign y12654 = ~n28499 ;
  assign y12655 = n28502 ;
  assign y12656 = ~n28504 ;
  assign y12657 = n28513 ;
  assign y12658 = n28514 ;
  assign y12659 = ~n28515 ;
  assign y12660 = n28518 ;
  assign y12661 = ~n28522 ;
  assign y12662 = ~n28523 ;
  assign y12663 = ~1'b0 ;
  assign y12664 = ~1'b0 ;
  assign y12665 = ~n28524 ;
  assign y12666 = n28527 ;
  assign y12667 = ~1'b0 ;
  assign y12668 = ~n28533 ;
  assign y12669 = n28537 ;
  assign y12670 = n28539 ;
  assign y12671 = ~1'b0 ;
  assign y12672 = ~n28543 ;
  assign y12673 = ~1'b0 ;
  assign y12674 = n28546 ;
  assign y12675 = n28547 ;
  assign y12676 = ~n28551 ;
  assign y12677 = ~n28556 ;
  assign y12678 = ~1'b0 ;
  assign y12679 = ~1'b0 ;
  assign y12680 = n28559 ;
  assign y12681 = ~n28563 ;
  assign y12682 = ~n28565 ;
  assign y12683 = ~1'b0 ;
  assign y12684 = ~n28567 ;
  assign y12685 = ~n28569 ;
  assign y12686 = ~n28571 ;
  assign y12687 = ~n28573 ;
  assign y12688 = ~1'b0 ;
  assign y12689 = n28574 ;
  assign y12690 = n28578 ;
  assign y12691 = ~1'b0 ;
  assign y12692 = n28580 ;
  assign y12693 = ~1'b0 ;
  assign y12694 = ~n28582 ;
  assign y12695 = ~n1455 ;
  assign y12696 = ~n28583 ;
  assign y12697 = ~n28586 ;
  assign y12698 = n28590 ;
  assign y12699 = ~1'b0 ;
  assign y12700 = 1'b0 ;
  assign y12701 = ~n17891 ;
  assign y12702 = n28593 ;
  assign y12703 = ~n9482 ;
  assign y12704 = n28595 ;
  assign y12705 = ~n28597 ;
  assign y12706 = ~n28599 ;
  assign y12707 = ~n28600 ;
  assign y12708 = ~n28602 ;
  assign y12709 = 1'b0 ;
  assign y12710 = ~1'b0 ;
  assign y12711 = ~n28609 ;
  assign y12712 = ~n28610 ;
  assign y12713 = n28614 ;
  assign y12714 = ~1'b0 ;
  assign y12715 = ~n28615 ;
  assign y12716 = ~n28622 ;
  assign y12717 = n28623 ;
  assign y12718 = ~n28624 ;
  assign y12719 = ~n28625 ;
  assign y12720 = ~1'b0 ;
  assign y12721 = n28628 ;
  assign y12722 = n28629 ;
  assign y12723 = ~1'b0 ;
  assign y12724 = ~1'b0 ;
  assign y12725 = ~n28630 ;
  assign y12726 = n28634 ;
  assign y12727 = ~n28635 ;
  assign y12728 = n28639 ;
  assign y12729 = n28645 ;
  assign y12730 = ~1'b0 ;
  assign y12731 = ~1'b0 ;
  assign y12732 = 1'b0 ;
  assign y12733 = ~n28651 ;
  assign y12734 = n28652 ;
  assign y12735 = ~n28655 ;
  assign y12736 = ~1'b0 ;
  assign y12737 = n28658 ;
  assign y12738 = ~1'b0 ;
  assign y12739 = ~n28662 ;
  assign y12740 = ~n28665 ;
  assign y12741 = n28667 ;
  assign y12742 = n28668 ;
  assign y12743 = n28679 ;
  assign y12744 = ~n28686 ;
  assign y12745 = 1'b0 ;
  assign y12746 = ~n28691 ;
  assign y12747 = ~n28693 ;
  assign y12748 = ~n28699 ;
  assign y12749 = ~n28701 ;
  assign y12750 = ~n20257 ;
  assign y12751 = n28707 ;
  assign y12752 = n28709 ;
  assign y12753 = ~n28715 ;
  assign y12754 = n28717 ;
  assign y12755 = ~n28718 ;
  assign y12756 = n28721 ;
  assign y12757 = n28723 ;
  assign y12758 = ~n28724 ;
  assign y12759 = ~n28726 ;
  assign y12760 = n28728 ;
  assign y12761 = ~n28733 ;
  assign y12762 = ~n28736 ;
  assign y12763 = ~n28738 ;
  assign y12764 = ~n28741 ;
  assign y12765 = n28742 ;
  assign y12766 = ~n28743 ;
  assign y12767 = ~n28749 ;
  assign y12768 = ~n28750 ;
  assign y12769 = ~1'b0 ;
  assign y12770 = ~n18948 ;
  assign y12771 = ~1'b0 ;
  assign y12772 = n7464 ;
  assign y12773 = ~n12462 ;
  assign y12774 = ~n28752 ;
  assign y12775 = n28753 ;
  assign y12776 = ~n28759 ;
  assign y12777 = ~1'b0 ;
  assign y12778 = ~n28761 ;
  assign y12779 = ~1'b0 ;
  assign y12780 = ~n28762 ;
  assign y12781 = n28763 ;
  assign y12782 = ~n28765 ;
  assign y12783 = ~1'b0 ;
  assign y12784 = ~1'b0 ;
  assign y12785 = n28766 ;
  assign y12786 = ~n28768 ;
  assign y12787 = ~1'b0 ;
  assign y12788 = n28769 ;
  assign y12789 = n28770 ;
  assign y12790 = ~n28771 ;
  assign y12791 = ~n28772 ;
  assign y12792 = n28774 ;
  assign y12793 = n28776 ;
  assign y12794 = n28778 ;
  assign y12795 = ~n28782 ;
  assign y12796 = n28787 ;
  assign y12797 = ~n28790 ;
  assign y12798 = n28792 ;
  assign y12799 = n28795 ;
  assign y12800 = n28797 ;
  assign y12801 = ~1'b0 ;
  assign y12802 = n28802 ;
  assign y12803 = ~1'b0 ;
  assign y12804 = ~1'b0 ;
  assign y12805 = ~n28807 ;
  assign y12806 = ~n28809 ;
  assign y12807 = n28811 ;
  assign y12808 = ~n3773 ;
  assign y12809 = ~1'b0 ;
  assign y12810 = ~n28815 ;
  assign y12811 = n28816 ;
  assign y12812 = n28817 ;
  assign y12813 = ~n28818 ;
  assign y12814 = n28821 ;
  assign y12815 = ~n28825 ;
  assign y12816 = ~n28830 ;
  assign y12817 = ~n28836 ;
  assign y12818 = n28839 ;
  assign y12819 = ~1'b0 ;
  assign y12820 = ~n28840 ;
  assign y12821 = ~1'b0 ;
  assign y12822 = ~n28842 ;
  assign y12823 = ~n12778 ;
  assign y12824 = ~n28844 ;
  assign y12825 = n28849 ;
  assign y12826 = ~1'b0 ;
  assign y12827 = ~n28851 ;
  assign y12828 = ~n28852 ;
  assign y12829 = ~n28853 ;
  assign y12830 = ~n28855 ;
  assign y12831 = n28860 ;
  assign y12832 = n28868 ;
  assign y12833 = ~1'b0 ;
  assign y12834 = ~1'b0 ;
  assign y12835 = ~1'b0 ;
  assign y12836 = n27496 ;
  assign y12837 = n28871 ;
  assign y12838 = ~n28879 ;
  assign y12839 = ~n28882 ;
  assign y12840 = ~1'b0 ;
  assign y12841 = ~n28883 ;
  assign y12842 = 1'b0 ;
  assign y12843 = n28887 ;
  assign y12844 = ~n28895 ;
  assign y12845 = n28897 ;
  assign y12846 = ~n28900 ;
  assign y12847 = n28902 ;
  assign y12848 = n28905 ;
  assign y12849 = ~n28908 ;
  assign y12850 = n28913 ;
  assign y12851 = ~1'b0 ;
  assign y12852 = ~1'b0 ;
  assign y12853 = ~n28916 ;
  assign y12854 = n28920 ;
  assign y12855 = n28921 ;
  assign y12856 = n28923 ;
  assign y12857 = n8914 ;
  assign y12858 = ~1'b0 ;
  assign y12859 = ~n28926 ;
  assign y12860 = n28929 ;
  assign y12861 = n28930 ;
  assign y12862 = ~n28931 ;
  assign y12863 = ~n28938 ;
  assign y12864 = ~1'b0 ;
  assign y12865 = ~n28940 ;
  assign y12866 = ~1'b0 ;
  assign y12867 = n28947 ;
  assign y12868 = ~n28950 ;
  assign y12869 = ~1'b0 ;
  assign y12870 = ~n9331 ;
  assign y12871 = ~1'b0 ;
  assign y12872 = ~1'b0 ;
  assign y12873 = ~n28953 ;
  assign y12874 = ~n28955 ;
  assign y12875 = n28956 ;
  assign y12876 = ~1'b0 ;
  assign y12877 = ~1'b0 ;
  assign y12878 = ~n28958 ;
  assign y12879 = ~n28960 ;
  assign y12880 = n28967 ;
  assign y12881 = ~n22394 ;
  assign y12882 = ~n28970 ;
  assign y12883 = n12661 ;
  assign y12884 = ~1'b0 ;
  assign y12885 = ~n28978 ;
  assign y12886 = ~1'b0 ;
  assign y12887 = n28980 ;
  assign y12888 = ~n28983 ;
  assign y12889 = n28984 ;
  assign y12890 = ~n28986 ;
  assign y12891 = ~n28988 ;
  assign y12892 = n28993 ;
  assign y12893 = ~n28994 ;
  assign y12894 = n28999 ;
  assign y12895 = ~1'b0 ;
  assign y12896 = n12882 ;
  assign y12897 = ~1'b0 ;
  assign y12898 = ~n29000 ;
  assign y12899 = n29001 ;
  assign y12900 = n29003 ;
  assign y12901 = ~n29005 ;
  assign y12902 = ~1'b0 ;
  assign y12903 = ~n27449 ;
  assign y12904 = ~1'b0 ;
  assign y12905 = n29015 ;
  assign y12906 = ~n29016 ;
  assign y12907 = n29021 ;
  assign y12908 = ~1'b0 ;
  assign y12909 = ~n29023 ;
  assign y12910 = n28445 ;
  assign y12911 = n29024 ;
  assign y12912 = ~n29029 ;
  assign y12913 = ~n29032 ;
  assign y12914 = ~1'b0 ;
  assign y12915 = ~n29035 ;
  assign y12916 = ~1'b0 ;
  assign y12917 = n29037 ;
  assign y12918 = ~n29039 ;
  assign y12919 = ~n29044 ;
  assign y12920 = 1'b0 ;
  assign y12921 = ~n29047 ;
  assign y12922 = ~1'b0 ;
  assign y12923 = n29049 ;
  assign y12924 = ~n29051 ;
  assign y12925 = ~n29053 ;
  assign y12926 = ~n29057 ;
  assign y12927 = n29058 ;
  assign y12928 = ~n29059 ;
  assign y12929 = ~1'b0 ;
  assign y12930 = ~n29061 ;
  assign y12931 = n29063 ;
  assign y12932 = ~n29064 ;
  assign y12933 = ~1'b0 ;
  assign y12934 = ~1'b0 ;
  assign y12935 = n29068 ;
  assign y12936 = n29069 ;
  assign y12937 = n29072 ;
  assign y12938 = n4260 ;
  assign y12939 = ~n29078 ;
  assign y12940 = ~1'b0 ;
  assign y12941 = ~1'b0 ;
  assign y12942 = ~n3775 ;
  assign y12943 = n29083 ;
  assign y12944 = ~n29085 ;
  assign y12945 = n29087 ;
  assign y12946 = n29089 ;
  assign y12947 = n29102 ;
  assign y12948 = ~1'b0 ;
  assign y12949 = ~n29105 ;
  assign y12950 = ~1'b0 ;
  assign y12951 = n29110 ;
  assign y12952 = n29111 ;
  assign y12953 = n29114 ;
  assign y12954 = n29117 ;
  assign y12955 = ~n29118 ;
  assign y12956 = 1'b0 ;
  assign y12957 = n29124 ;
  assign y12958 = n29127 ;
  assign y12959 = ~1'b0 ;
  assign y12960 = n29129 ;
  assign y12961 = ~1'b0 ;
  assign y12962 = ~n29131 ;
  assign y12963 = n29133 ;
  assign y12964 = ~n29135 ;
  assign y12965 = n29139 ;
  assign y12966 = n29144 ;
  assign y12967 = n29149 ;
  assign y12968 = ~n29152 ;
  assign y12969 = n29153 ;
  assign y12970 = n29159 ;
  assign y12971 = n29164 ;
  assign y12972 = ~n29167 ;
  assign y12973 = n4865 ;
  assign y12974 = ~1'b0 ;
  assign y12975 = 1'b0 ;
  assign y12976 = ~1'b0 ;
  assign y12977 = ~1'b0 ;
  assign y12978 = ~1'b0 ;
  assign y12979 = 1'b0 ;
  assign y12980 = ~1'b0 ;
  assign y12981 = n21787 ;
  assign y12982 = n15542 ;
  assign y12983 = ~n29172 ;
  assign y12984 = ~n29176 ;
  assign y12985 = n29178 ;
  assign y12986 = ~1'b0 ;
  assign y12987 = ~n29180 ;
  assign y12988 = ~n29182 ;
  assign y12989 = n29185 ;
  assign y12990 = ~n29189 ;
  assign y12991 = ~n29190 ;
  assign y12992 = ~1'b0 ;
  assign y12993 = ~1'b0 ;
  assign y12994 = n29192 ;
  assign y12995 = ~1'b0 ;
  assign y12996 = ~1'b0 ;
  assign y12997 = ~n29193 ;
  assign y12998 = n29194 ;
  assign y12999 = n29196 ;
  assign y13000 = n29201 ;
  assign y13001 = ~n27518 ;
  assign y13002 = ~n29203 ;
  assign y13003 = ~1'b0 ;
  assign y13004 = n29205 ;
  assign y13005 = ~n29214 ;
  assign y13006 = ~n29216 ;
  assign y13007 = ~n29218 ;
  assign y13008 = n29224 ;
  assign y13009 = n29226 ;
  assign y13010 = ~1'b0 ;
  assign y13011 = ~n29228 ;
  assign y13012 = ~1'b0 ;
  assign y13013 = ~n29230 ;
  assign y13014 = ~n29232 ;
  assign y13015 = ~n5598 ;
  assign y13016 = ~1'b0 ;
  assign y13017 = ~1'b0 ;
  assign y13018 = ~n29234 ;
  assign y13019 = n29235 ;
  assign y13020 = ~n29236 ;
  assign y13021 = ~1'b0 ;
  assign y13022 = n29239 ;
  assign y13023 = n29243 ;
  assign y13024 = ~n29245 ;
  assign y13025 = ~n29254 ;
  assign y13026 = ~1'b0 ;
  assign y13027 = ~1'b0 ;
  assign y13028 = ~1'b0 ;
  assign y13029 = ~1'b0 ;
  assign y13030 = ~n29258 ;
  assign y13031 = n29259 ;
  assign y13032 = ~n29260 ;
  assign y13033 = n29262 ;
  assign y13034 = ~n29264 ;
  assign y13035 = ~n29266 ;
  assign y13036 = ~n29268 ;
  assign y13037 = 1'b0 ;
  assign y13038 = ~1'b0 ;
  assign y13039 = ~1'b0 ;
  assign y13040 = ~n29270 ;
  assign y13041 = n29272 ;
  assign y13042 = n29274 ;
  assign y13043 = ~1'b0 ;
  assign y13044 = n16735 ;
  assign y13045 = ~n29278 ;
  assign y13046 = n29281 ;
  assign y13047 = n1086 ;
  assign y13048 = ~n4686 ;
  assign y13049 = n29284 ;
  assign y13050 = ~n29292 ;
  assign y13051 = n29293 ;
  assign y13052 = ~1'b0 ;
  assign y13053 = n29295 ;
  assign y13054 = ~1'b0 ;
  assign y13055 = ~1'b0 ;
  assign y13056 = n29296 ;
  assign y13057 = n2309 ;
  assign y13058 = ~1'b0 ;
  assign y13059 = ~n1760 ;
  assign y13060 = ~n29314 ;
  assign y13061 = ~n29315 ;
  assign y13062 = ~n29316 ;
  assign y13063 = n5229 ;
  assign y13064 = ~1'b0 ;
  assign y13065 = ~n29317 ;
  assign y13066 = n29319 ;
  assign y13067 = ~1'b0 ;
  assign y13068 = ~n29320 ;
  assign y13069 = ~1'b0 ;
  assign y13070 = ~n29321 ;
  assign y13071 = ~1'b0 ;
  assign y13072 = ~1'b0 ;
  assign y13073 = ~n29323 ;
  assign y13074 = n29328 ;
  assign y13075 = n29329 ;
  assign y13076 = n29330 ;
  assign y13077 = n29333 ;
  assign y13078 = n29337 ;
  assign y13079 = ~n29339 ;
  assign y13080 = ~n29341 ;
  assign y13081 = ~n29342 ;
  assign y13082 = ~n29349 ;
  assign y13083 = n29353 ;
  assign y13084 = ~n29355 ;
  assign y13085 = n29357 ;
  assign y13086 = 1'b0 ;
  assign y13087 = n29358 ;
  assign y13088 = ~n29359 ;
  assign y13089 = ~1'b0 ;
  assign y13090 = ~1'b0 ;
  assign y13091 = ~n29360 ;
  assign y13092 = ~1'b0 ;
  assign y13093 = n29363 ;
  assign y13094 = n29364 ;
  assign y13095 = ~n29366 ;
  assign y13096 = ~n29367 ;
  assign y13097 = ~1'b0 ;
  assign y13098 = ~1'b0 ;
  assign y13099 = n29372 ;
  assign y13100 = n29377 ;
  assign y13101 = ~1'b0 ;
  assign y13102 = n29379 ;
  assign y13103 = n29380 ;
  assign y13104 = n29389 ;
  assign y13105 = ~n29393 ;
  assign y13106 = n29396 ;
  assign y13107 = ~n29400 ;
  assign y13108 = ~1'b0 ;
  assign y13109 = ~1'b0 ;
  assign y13110 = ~1'b0 ;
  assign y13111 = ~n29404 ;
  assign y13112 = ~1'b0 ;
  assign y13113 = ~1'b0 ;
  assign y13114 = ~n29406 ;
  assign y13115 = ~n28382 ;
  assign y13116 = n29409 ;
  assign y13117 = n29411 ;
  assign y13118 = ~1'b0 ;
  assign y13119 = n29412 ;
  assign y13120 = n29414 ;
  assign y13121 = n29416 ;
  assign y13122 = ~n29417 ;
  assign y13123 = n29418 ;
  assign y13124 = ~1'b0 ;
  assign y13125 = ~1'b0 ;
  assign y13126 = n29421 ;
  assign y13127 = ~n29426 ;
  assign y13128 = n29429 ;
  assign y13129 = ~n29430 ;
  assign y13130 = ~n29433 ;
  assign y13131 = ~n29435 ;
  assign y13132 = ~n29437 ;
  assign y13133 = ~1'b0 ;
  assign y13134 = ~1'b0 ;
  assign y13135 = ~n7337 ;
  assign y13136 = n29443 ;
  assign y13137 = ~1'b0 ;
  assign y13138 = n29020 ;
  assign y13139 = ~n29449 ;
  assign y13140 = n29452 ;
  assign y13141 = ~1'b0 ;
  assign y13142 = n29453 ;
  assign y13143 = n29456 ;
  assign y13144 = ~n29460 ;
  assign y13145 = 1'b0 ;
  assign y13146 = n29462 ;
  assign y13147 = ~1'b0 ;
  assign y13148 = ~n29468 ;
  assign y13149 = n29472 ;
  assign y13150 = ~n13614 ;
  assign y13151 = ~n29474 ;
  assign y13152 = n29475 ;
  assign y13153 = n29478 ;
  assign y13154 = n25748 ;
  assign y13155 = n7916 ;
  assign y13156 = n29484 ;
  assign y13157 = ~n29487 ;
  assign y13158 = ~1'b0 ;
  assign y13159 = ~n29488 ;
  assign y13160 = ~n29496 ;
  assign y13161 = ~1'b0 ;
  assign y13162 = ~1'b0 ;
  assign y13163 = ~1'b0 ;
  assign y13164 = ~1'b0 ;
  assign y13165 = n29500 ;
  assign y13166 = ~n29502 ;
  assign y13167 = n29504 ;
  assign y13168 = ~n29511 ;
  assign y13169 = n29514 ;
  assign y13170 = ~1'b0 ;
  assign y13171 = n29517 ;
  assign y13172 = ~n29518 ;
  assign y13173 = ~n29520 ;
  assign y13174 = ~n29522 ;
  assign y13175 = ~1'b0 ;
  assign y13176 = ~n29524 ;
  assign y13177 = ~n29526 ;
  assign y13178 = n29527 ;
  assign y13179 = n29528 ;
  assign y13180 = n29529 ;
  assign y13181 = ~n29532 ;
  assign y13182 = ~n29536 ;
  assign y13183 = n29539 ;
  assign y13184 = n29545 ;
  assign y13185 = ~n29547 ;
  assign y13186 = ~1'b0 ;
  assign y13187 = n29549 ;
  assign y13188 = ~1'b0 ;
  assign y13189 = ~n29550 ;
  assign y13190 = n29554 ;
  assign y13191 = ~1'b0 ;
  assign y13192 = ~1'b0 ;
  assign y13193 = n29560 ;
  assign y13194 = n29563 ;
  assign y13195 = n29565 ;
  assign y13196 = ~n29568 ;
  assign y13197 = ~1'b0 ;
  assign y13198 = ~1'b0 ;
  assign y13199 = ~n29571 ;
  assign y13200 = n29578 ;
  assign y13201 = n29580 ;
  assign y13202 = ~n29581 ;
  assign y13203 = ~1'b0 ;
  assign y13204 = n29584 ;
  assign y13205 = ~1'b0 ;
  assign y13206 = ~1'b0 ;
  assign y13207 = n29585 ;
  assign y13208 = n29589 ;
  assign y13209 = n29595 ;
  assign y13210 = ~n29600 ;
  assign y13211 = ~1'b0 ;
  assign y13212 = ~n29603 ;
  assign y13213 = ~n29605 ;
  assign y13214 = ~n29609 ;
  assign y13215 = ~n29614 ;
  assign y13216 = ~1'b0 ;
  assign y13217 = ~1'b0 ;
  assign y13218 = ~n29619 ;
  assign y13219 = ~n29621 ;
  assign y13220 = ~n29623 ;
  assign y13221 = ~1'b0 ;
  assign y13222 = ~n29624 ;
  assign y13223 = ~n29625 ;
  assign y13224 = ~n6363 ;
  assign y13225 = ~n29629 ;
  assign y13226 = ~1'b0 ;
  assign y13227 = n29632 ;
  assign y13228 = n29635 ;
  assign y13229 = n29636 ;
  assign y13230 = n7024 ;
  assign y13231 = n29643 ;
  assign y13232 = ~n29647 ;
  assign y13233 = ~n29649 ;
  assign y13234 = n7485 ;
  assign y13235 = n29650 ;
  assign y13236 = n29653 ;
  assign y13237 = ~n29657 ;
  assign y13238 = ~n29659 ;
  assign y13239 = n29661 ;
  assign y13240 = n29662 ;
  assign y13241 = ~n29663 ;
  assign y13242 = ~n29666 ;
  assign y13243 = ~1'b0 ;
  assign y13244 = n29670 ;
  assign y13245 = n29673 ;
  assign y13246 = n29675 ;
  assign y13247 = n20899 ;
  assign y13248 = n29676 ;
  assign y13249 = ~1'b0 ;
  assign y13250 = ~n29680 ;
  assign y13251 = ~1'b0 ;
  assign y13252 = ~1'b0 ;
  assign y13253 = ~n29682 ;
  assign y13254 = ~1'b0 ;
  assign y13255 = n14715 ;
  assign y13256 = ~n29685 ;
  assign y13257 = ~n29690 ;
  assign y13258 = ~n29695 ;
  assign y13259 = ~n29696 ;
  assign y13260 = ~1'b0 ;
  assign y13261 = ~n29697 ;
  assign y13262 = ~1'b0 ;
  assign y13263 = n29699 ;
  assign y13264 = ~n7281 ;
  assign y13265 = n29702 ;
  assign y13266 = ~n29704 ;
  assign y13267 = ~n29706 ;
  assign y13268 = n13687 ;
  assign y13269 = ~n29708 ;
  assign y13270 = n29710 ;
  assign y13271 = ~1'b0 ;
  assign y13272 = ~n29713 ;
  assign y13273 = n29715 ;
  assign y13274 = n29716 ;
  assign y13275 = n14262 ;
  assign y13276 = n29718 ;
  assign y13277 = ~1'b0 ;
  assign y13278 = n29719 ;
  assign y13279 = ~n29722 ;
  assign y13280 = ~1'b0 ;
  assign y13281 = 1'b0 ;
  assign y13282 = ~n29729 ;
  assign y13283 = n29732 ;
  assign y13284 = ~1'b0 ;
  assign y13285 = n9783 ;
  assign y13286 = n29734 ;
  assign y13287 = n29736 ;
  assign y13288 = n29738 ;
  assign y13289 = n29739 ;
  assign y13290 = ~n29743 ;
  assign y13291 = n29745 ;
  assign y13292 = ~1'b0 ;
  assign y13293 = ~1'b0 ;
  assign y13294 = ~1'b0 ;
  assign y13295 = ~n29746 ;
  assign y13296 = n10019 ;
  assign y13297 = n29748 ;
  assign y13298 = ~1'b0 ;
  assign y13299 = ~1'b0 ;
  assign y13300 = ~1'b0 ;
  assign y13301 = ~1'b0 ;
  assign y13302 = ~n26321 ;
  assign y13303 = ~1'b0 ;
  assign y13304 = ~n29750 ;
  assign y13305 = ~1'b0 ;
  assign y13306 = ~n29753 ;
  assign y13307 = n29756 ;
  assign y13308 = n29758 ;
  assign y13309 = n29759 ;
  assign y13310 = ~n29760 ;
  assign y13311 = n29761 ;
  assign y13312 = n29763 ;
  assign y13313 = ~n29765 ;
  assign y13314 = ~n29767 ;
  assign y13315 = ~n6253 ;
  assign y13316 = n29769 ;
  assign y13317 = n29770 ;
  assign y13318 = ~1'b0 ;
  assign y13319 = n29772 ;
  assign y13320 = ~n29773 ;
  assign y13321 = n29775 ;
  assign y13322 = ~n29783 ;
  assign y13323 = n29784 ;
  assign y13324 = ~n29786 ;
  assign y13325 = ~1'b0 ;
  assign y13326 = n29787 ;
  assign y13327 = n29790 ;
  assign y13328 = ~1'b0 ;
  assign y13329 = n29799 ;
  assign y13330 = n29800 ;
  assign y13331 = ~1'b0 ;
  assign y13332 = n29802 ;
  assign y13333 = ~1'b0 ;
  assign y13334 = ~n29805 ;
  assign y13335 = ~n26130 ;
  assign y13336 = ~1'b0 ;
  assign y13337 = ~n29807 ;
  assign y13338 = 1'b0 ;
  assign y13339 = n29810 ;
  assign y13340 = n29814 ;
  assign y13341 = ~n29816 ;
  assign y13342 = ~n29817 ;
  assign y13343 = n29820 ;
  assign y13344 = ~1'b0 ;
  assign y13345 = n29822 ;
  assign y13346 = n29824 ;
  assign y13347 = n29825 ;
  assign y13348 = n29826 ;
  assign y13349 = n29827 ;
  assign y13350 = ~1'b0 ;
  assign y13351 = ~n29832 ;
  assign y13352 = n29835 ;
  assign y13353 = n29836 ;
  assign y13354 = n29843 ;
  assign y13355 = n29845 ;
  assign y13356 = ~n29846 ;
  assign y13357 = n29856 ;
  assign y13358 = ~1'b0 ;
  assign y13359 = n29859 ;
  assign y13360 = n29860 ;
  assign y13361 = ~n29864 ;
  assign y13362 = n29865 ;
  assign y13363 = ~n29868 ;
  assign y13364 = n29870 ;
  assign y13365 = n29874 ;
  assign y13366 = n29878 ;
  assign y13367 = ~1'b0 ;
  assign y13368 = ~n29880 ;
  assign y13369 = ~1'b0 ;
  assign y13370 = ~n29882 ;
  assign y13371 = n29884 ;
  assign y13372 = ~n29889 ;
  assign y13373 = n7027 ;
  assign y13374 = n29890 ;
  assign y13375 = ~1'b0 ;
  assign y13376 = ~n29891 ;
  assign y13377 = ~n29893 ;
  assign y13378 = n29894 ;
  assign y13379 = ~1'b0 ;
  assign y13380 = ~n29897 ;
  assign y13381 = ~n29898 ;
  assign y13382 = n29905 ;
  assign y13383 = ~1'b0 ;
  assign y13384 = ~1'b0 ;
  assign y13385 = n29906 ;
  assign y13386 = ~n29912 ;
  assign y13387 = ~n29913 ;
  assign y13388 = n29916 ;
  assign y13389 = n29920 ;
  assign y13390 = ~n22716 ;
  assign y13391 = n29921 ;
  assign y13392 = ~n3183 ;
  assign y13393 = ~n29923 ;
  assign y13394 = ~n29924 ;
  assign y13395 = n29930 ;
  assign y13396 = n15227 ;
  assign y13397 = n29933 ;
  assign y13398 = n29934 ;
  assign y13399 = ~n29939 ;
  assign y13400 = ~1'b0 ;
  assign y13401 = n29940 ;
  assign y13402 = n29941 ;
  assign y13403 = n29942 ;
  assign y13404 = n29943 ;
  assign y13405 = ~1'b0 ;
  assign y13406 = ~n29944 ;
  assign y13407 = ~1'b0 ;
  assign y13408 = ~n29949 ;
  assign y13409 = ~n29950 ;
  assign y13410 = n29952 ;
  assign y13411 = n29953 ;
  assign y13412 = n29956 ;
  assign y13413 = ~n29957 ;
  assign y13414 = ~n29961 ;
  assign y13415 = ~n29963 ;
  assign y13416 = n29966 ;
  assign y13417 = ~n29967 ;
  assign y13418 = n29973 ;
  assign y13419 = n29974 ;
  assign y13420 = ~1'b0 ;
  assign y13421 = n29975 ;
  assign y13422 = n29977 ;
  assign y13423 = ~n29980 ;
  assign y13424 = ~n29984 ;
  assign y13425 = n29985 ;
  assign y13426 = ~n29987 ;
  assign y13427 = ~n29990 ;
  assign y13428 = n29992 ;
  assign y13429 = n21785 ;
  assign y13430 = ~n29994 ;
  assign y13431 = n29996 ;
  assign y13432 = 1'b0 ;
  assign y13433 = ~n29998 ;
  assign y13434 = n4286 ;
  assign y13435 = n30003 ;
  assign y13436 = ~n30004 ;
  assign y13437 = ~n30005 ;
  assign y13438 = ~n30008 ;
  assign y13439 = ~1'b0 ;
  assign y13440 = ~n30011 ;
  assign y13441 = ~n30013 ;
  assign y13442 = n30014 ;
  assign y13443 = ~1'b0 ;
  assign y13444 = n30017 ;
  assign y13445 = ~1'b0 ;
  assign y13446 = ~1'b0 ;
  assign y13447 = ~n30021 ;
  assign y13448 = n30022 ;
  assign y13449 = ~n30023 ;
  assign y13450 = n30029 ;
  assign y13451 = n30030 ;
  assign y13452 = ~1'b0 ;
  assign y13453 = ~1'b0 ;
  assign y13454 = n30033 ;
  assign y13455 = ~n30040 ;
  assign y13456 = ~1'b0 ;
  assign y13457 = ~1'b0 ;
  assign y13458 = ~n30042 ;
  assign y13459 = n30045 ;
  assign y13460 = ~n30050 ;
  assign y13461 = ~n30052 ;
  assign y13462 = ~n4378 ;
  assign y13463 = ~n30062 ;
  assign y13464 = ~n30065 ;
  assign y13465 = ~n30068 ;
  assign y13466 = ~1'b0 ;
  assign y13467 = ~1'b0 ;
  assign y13468 = n30069 ;
  assign y13469 = n30070 ;
  assign y13470 = n30071 ;
  assign y13471 = n30076 ;
  assign y13472 = n30077 ;
  assign y13473 = ~n30080 ;
  assign y13474 = n30082 ;
  assign y13475 = n30084 ;
  assign y13476 = ~n30086 ;
  assign y13477 = ~n30090 ;
  assign y13478 = n30091 ;
  assign y13479 = ~1'b0 ;
  assign y13480 = n30092 ;
  assign y13481 = ~n30096 ;
  assign y13482 = ~n30098 ;
  assign y13483 = ~n30102 ;
  assign y13484 = ~n30104 ;
  assign y13485 = n11267 ;
  assign y13486 = ~1'b0 ;
  assign y13487 = ~n30106 ;
  assign y13488 = ~n30108 ;
  assign y13489 = n5474 ;
  assign y13490 = n30111 ;
  assign y13491 = ~n30114 ;
  assign y13492 = n30115 ;
  assign y13493 = ~1'b0 ;
  assign y13494 = ~n30117 ;
  assign y13495 = ~n30118 ;
  assign y13496 = ~1'b0 ;
  assign y13497 = ~1'b0 ;
  assign y13498 = n30120 ;
  assign y13499 = n30121 ;
  assign y13500 = ~n30123 ;
  assign y13501 = ~n30125 ;
  assign y13502 = ~1'b0 ;
  assign y13503 = ~1'b0 ;
  assign y13504 = ~n30129 ;
  assign y13505 = ~n30132 ;
  assign y13506 = ~1'b0 ;
  assign y13507 = ~n30134 ;
  assign y13508 = ~n30136 ;
  assign y13509 = ~1'b0 ;
  assign y13510 = ~1'b0 ;
  assign y13511 = n30138 ;
  assign y13512 = n30139 ;
  assign y13513 = n30140 ;
  assign y13514 = ~n30142 ;
  assign y13515 = ~1'b0 ;
  assign y13516 = ~n30143 ;
  assign y13517 = n30145 ;
  assign y13518 = ~n30149 ;
  assign y13519 = ~n30151 ;
  assign y13520 = n30153 ;
  assign y13521 = n30155 ;
  assign y13522 = ~1'b0 ;
  assign y13523 = ~n30156 ;
  assign y13524 = n30157 ;
  assign y13525 = n11055 ;
  assign y13526 = ~n30162 ;
  assign y13527 = ~1'b0 ;
  assign y13528 = ~1'b0 ;
  assign y13529 = n30165 ;
  assign y13530 = ~n30167 ;
  assign y13531 = ~n30173 ;
  assign y13532 = n30177 ;
  assign y13533 = 1'b0 ;
  assign y13534 = n30181 ;
  assign y13535 = n26705 ;
  assign y13536 = ~n30183 ;
  assign y13537 = n30187 ;
  assign y13538 = n30191 ;
  assign y13539 = n30193 ;
  assign y13540 = ~n30200 ;
  assign y13541 = ~n30203 ;
  assign y13542 = n30206 ;
  assign y13543 = ~1'b0 ;
  assign y13544 = ~1'b0 ;
  assign y13545 = n30210 ;
  assign y13546 = n30212 ;
  assign y13547 = ~n30218 ;
  assign y13548 = n30220 ;
  assign y13549 = n30222 ;
  assign y13550 = n30223 ;
  assign y13551 = n30230 ;
  assign y13552 = n30231 ;
  assign y13553 = ~n30235 ;
  assign y13554 = n30237 ;
  assign y13555 = ~1'b0 ;
  assign y13556 = ~n30239 ;
  assign y13557 = n30240 ;
  assign y13558 = ~n30242 ;
  assign y13559 = ~1'b0 ;
  assign y13560 = ~n30247 ;
  assign y13561 = n30248 ;
  assign y13562 = ~n11129 ;
  assign y13563 = ~1'b0 ;
  assign y13564 = n30252 ;
  assign y13565 = ~1'b0 ;
  assign y13566 = ~1'b0 ;
  assign y13567 = ~n30254 ;
  assign y13568 = ~n3376 ;
  assign y13569 = n30256 ;
  assign y13570 = ~n30259 ;
  assign y13571 = n30262 ;
  assign y13572 = ~n16999 ;
  assign y13573 = n30264 ;
  assign y13574 = ~n30267 ;
  assign y13575 = ~n30269 ;
  assign y13576 = n30271 ;
  assign y13577 = n30272 ;
  assign y13578 = ~n30275 ;
  assign y13579 = ~n30276 ;
  assign y13580 = ~n30277 ;
  assign y13581 = ~1'b0 ;
  assign y13582 = ~1'b0 ;
  assign y13583 = n30279 ;
  assign y13584 = ~n1712 ;
  assign y13585 = n17009 ;
  assign y13586 = ~n30281 ;
  assign y13587 = ~1'b0 ;
  assign y13588 = ~n30283 ;
  assign y13589 = ~n30285 ;
  assign y13590 = ~n30286 ;
  assign y13591 = ~1'b0 ;
  assign y13592 = ~n30287 ;
  assign y13593 = n30288 ;
  assign y13594 = n30289 ;
  assign y13595 = ~n30291 ;
  assign y13596 = n30293 ;
  assign y13597 = n30294 ;
  assign y13598 = n30297 ;
  assign y13599 = ~1'b0 ;
  assign y13600 = n30298 ;
  assign y13601 = ~n30299 ;
  assign y13602 = n30300 ;
  assign y13603 = n30302 ;
  assign y13604 = n30304 ;
  assign y13605 = ~1'b0 ;
  assign y13606 = 1'b0 ;
  assign y13607 = n30305 ;
  assign y13608 = n30306 ;
  assign y13609 = n30307 ;
  assign y13610 = ~n30312 ;
  assign y13611 = n30316 ;
  assign y13612 = ~1'b0 ;
  assign y13613 = 1'b0 ;
  assign y13614 = ~n4658 ;
  assign y13615 = ~n30318 ;
  assign y13616 = n30319 ;
  assign y13617 = ~n30322 ;
  assign y13618 = ~n30323 ;
  assign y13619 = n30324 ;
  assign y13620 = ~1'b0 ;
  assign y13621 = ~n30325 ;
  assign y13622 = ~1'b0 ;
  assign y13623 = ~n30326 ;
  assign y13624 = n30327 ;
  assign y13625 = ~1'b0 ;
  assign y13626 = n30328 ;
  assign y13627 = ~n30329 ;
  assign y13628 = ~n30330 ;
  assign y13629 = ~n7518 ;
  assign y13630 = ~n30331 ;
  assign y13631 = n13830 ;
  assign y13632 = ~n30333 ;
  assign y13633 = n30334 ;
  assign y13634 = n6885 ;
  assign y13635 = n30336 ;
  assign y13636 = n30340 ;
  assign y13637 = n30341 ;
  assign y13638 = ~n30342 ;
  assign y13639 = ~1'b0 ;
  assign y13640 = ~n30345 ;
  assign y13641 = ~n30346 ;
  assign y13642 = n30347 ;
  assign y13643 = n30352 ;
  assign y13644 = ~1'b0 ;
  assign y13645 = n30353 ;
  assign y13646 = n30358 ;
  assign y13647 = ~n30360 ;
  assign y13648 = ~n30362 ;
  assign y13649 = ~n30364 ;
  assign y13650 = n30368 ;
  assign y13651 = ~n30369 ;
  assign y13652 = ~n30371 ;
  assign y13653 = n30372 ;
  assign y13654 = ~n30378 ;
  assign y13655 = ~n30379 ;
  assign y13656 = n30380 ;
  assign y13657 = ~n30382 ;
  assign y13658 = ~n19393 ;
  assign y13659 = ~1'b0 ;
  assign y13660 = ~n30392 ;
  assign y13661 = ~1'b0 ;
  assign y13662 = n30395 ;
  assign y13663 = ~n15390 ;
  assign y13664 = n30403 ;
  assign y13665 = n30405 ;
  assign y13666 = ~1'b0 ;
  assign y13667 = n30408 ;
  assign y13668 = n20392 ;
  assign y13669 = ~1'b0 ;
  assign y13670 = ~1'b0 ;
  assign y13671 = n30411 ;
  assign y13672 = ~n30412 ;
  assign y13673 = ~n30413 ;
  assign y13674 = n30414 ;
  assign y13675 = ~n30415 ;
  assign y13676 = ~n11004 ;
  assign y13677 = ~n30416 ;
  assign y13678 = n30418 ;
  assign y13679 = n30421 ;
  assign y13680 = ~1'b0 ;
  assign y13681 = n30425 ;
  assign y13682 = ~1'b0 ;
  assign y13683 = ~n30426 ;
  assign y13684 = ~n30429 ;
  assign y13685 = ~1'b0 ;
  assign y13686 = ~n30433 ;
  assign y13687 = ~1'b0 ;
  assign y13688 = ~n30436 ;
  assign y13689 = ~1'b0 ;
  assign y13690 = n30437 ;
  assign y13691 = n30439 ;
  assign y13692 = ~1'b0 ;
  assign y13693 = ~1'b0 ;
  assign y13694 = n30440 ;
  assign y13695 = ~1'b0 ;
  assign y13696 = ~1'b0 ;
  assign y13697 = n30444 ;
  assign y13698 = ~n30446 ;
  assign y13699 = ~1'b0 ;
  assign y13700 = ~n30448 ;
  assign y13701 = ~1'b0 ;
  assign y13702 = n30450 ;
  assign y13703 = ~1'b0 ;
  assign y13704 = n28588 ;
  assign y13705 = ~n30452 ;
  assign y13706 = ~n30453 ;
  assign y13707 = ~1'b0 ;
  assign y13708 = ~n30454 ;
  assign y13709 = ~n30458 ;
  assign y13710 = ~1'b0 ;
  assign y13711 = ~1'b0 ;
  assign y13712 = ~n30460 ;
  assign y13713 = ~1'b0 ;
  assign y13714 = ~n30467 ;
  assign y13715 = n9513 ;
  assign y13716 = ~n30470 ;
  assign y13717 = ~1'b0 ;
  assign y13718 = ~1'b0 ;
  assign y13719 = ~n30471 ;
  assign y13720 = n5491 ;
  assign y13721 = n30472 ;
  assign y13722 = n30475 ;
  assign y13723 = ~n30476 ;
  assign y13724 = ~1'b0 ;
  assign y13725 = ~n30477 ;
  assign y13726 = ~1'b0 ;
  assign y13727 = n30478 ;
  assign y13728 = ~n30484 ;
  assign y13729 = n30487 ;
  assign y13730 = ~n30489 ;
  assign y13731 = ~n16902 ;
  assign y13732 = n30492 ;
  assign y13733 = ~n25318 ;
  assign y13734 = ~n30493 ;
  assign y13735 = ~n30494 ;
  assign y13736 = ~n30495 ;
  assign y13737 = ~1'b0 ;
  assign y13738 = n30496 ;
  assign y13739 = n30498 ;
  assign y13740 = n30502 ;
  assign y13741 = n30503 ;
  assign y13742 = ~1'b0 ;
  assign y13743 = n30507 ;
  assign y13744 = ~n30509 ;
  assign y13745 = n30511 ;
  assign y13746 = ~n30514 ;
  assign y13747 = ~n30521 ;
  assign y13748 = n30523 ;
  assign y13749 = n30526 ;
  assign y13750 = ~1'b0 ;
  assign y13751 = ~1'b0 ;
  assign y13752 = ~n30527 ;
  assign y13753 = ~1'b0 ;
  assign y13754 = ~n30528 ;
  assign y13755 = ~n30534 ;
  assign y13756 = ~1'b0 ;
  assign y13757 = ~1'b0 ;
  assign y13758 = ~1'b0 ;
  assign y13759 = ~n30537 ;
  assign y13760 = ~1'b0 ;
  assign y13761 = n30542 ;
  assign y13762 = ~n30546 ;
  assign y13763 = ~n30550 ;
  assign y13764 = ~1'b0 ;
  assign y13765 = n30551 ;
  assign y13766 = ~1'b0 ;
  assign y13767 = n30552 ;
  assign y13768 = n30553 ;
  assign y13769 = ~n22283 ;
  assign y13770 = ~1'b0 ;
  assign y13771 = ~1'b0 ;
  assign y13772 = n30569 ;
  assign y13773 = ~1'b0 ;
  assign y13774 = n30571 ;
  assign y13775 = n13628 ;
  assign y13776 = ~n30575 ;
  assign y13777 = n30579 ;
  assign y13778 = n30580 ;
  assign y13779 = n20723 ;
  assign y13780 = ~1'b0 ;
  assign y13781 = ~1'b0 ;
  assign y13782 = ~n30581 ;
  assign y13783 = n30582 ;
  assign y13784 = n30584 ;
  assign y13785 = ~n30585 ;
  assign y13786 = ~n30588 ;
  assign y13787 = ~n30589 ;
  assign y13788 = n30591 ;
  assign y13789 = n30593 ;
  assign y13790 = ~1'b0 ;
  assign y13791 = ~n30596 ;
  assign y13792 = ~1'b0 ;
  assign y13793 = ~n30603 ;
  assign y13794 = ~1'b0 ;
  assign y13795 = ~1'b0 ;
  assign y13796 = ~n30604 ;
  assign y13797 = n30609 ;
  assign y13798 = ~n30610 ;
  assign y13799 = ~n30611 ;
  assign y13800 = ~1'b0 ;
  assign y13801 = ~n30614 ;
  assign y13802 = n30616 ;
  assign y13803 = n30618 ;
  assign y13804 = ~n30620 ;
  assign y13805 = ~1'b0 ;
  assign y13806 = ~1'b0 ;
  assign y13807 = ~1'b0 ;
  assign y13808 = ~n30622 ;
  assign y13809 = ~1'b0 ;
  assign y13810 = ~1'b0 ;
  assign y13811 = n30624 ;
  assign y13812 = ~1'b0 ;
  assign y13813 = ~1'b0 ;
  assign y13814 = n30626 ;
  assign y13815 = ~1'b0 ;
  assign y13816 = n9086 ;
  assign y13817 = n30629 ;
  assign y13818 = ~n30630 ;
  assign y13819 = n30631 ;
  assign y13820 = ~1'b0 ;
  assign y13821 = ~n30633 ;
  assign y13822 = ~1'b0 ;
  assign y13823 = ~n30635 ;
  assign y13824 = ~1'b0 ;
  assign y13825 = n30636 ;
  assign y13826 = ~n30638 ;
  assign y13827 = n30639 ;
  assign y13828 = n30640 ;
  assign y13829 = ~n30641 ;
  assign y13830 = n30643 ;
  assign y13831 = ~n30645 ;
  assign y13832 = n30646 ;
  assign y13833 = ~n30654 ;
  assign y13834 = ~1'b0 ;
  assign y13835 = n30659 ;
  assign y13836 = ~n30660 ;
  assign y13837 = ~1'b0 ;
  assign y13838 = ~1'b0 ;
  assign y13839 = n30661 ;
  assign y13840 = ~1'b0 ;
  assign y13841 = n30665 ;
  assign y13842 = ~n30668 ;
  assign y13843 = ~n30670 ;
  assign y13844 = ~n30672 ;
  assign y13845 = n30674 ;
  assign y13846 = n30676 ;
  assign y13847 = ~1'b0 ;
  assign y13848 = n30683 ;
  assign y13849 = ~n30684 ;
  assign y13850 = n4538 ;
  assign y13851 = ~n30686 ;
  assign y13852 = n30687 ;
  assign y13853 = ~1'b0 ;
  assign y13854 = ~1'b0 ;
  assign y13855 = ~n30691 ;
  assign y13856 = ~n30693 ;
  assign y13857 = ~1'b0 ;
  assign y13858 = n30694 ;
  assign y13859 = n30698 ;
  assign y13860 = ~1'b0 ;
  assign y13861 = ~n30701 ;
  assign y13862 = ~n30702 ;
  assign y13863 = n30703 ;
  assign y13864 = n30708 ;
  assign y13865 = n30709 ;
  assign y13866 = ~1'b0 ;
  assign y13867 = ~n30710 ;
  assign y13868 = ~n30712 ;
  assign y13869 = ~n30714 ;
  assign y13870 = n30716 ;
  assign y13871 = ~n30719 ;
  assign y13872 = n30720 ;
  assign y13873 = ~1'b0 ;
  assign y13874 = ~n11449 ;
  assign y13875 = n30721 ;
  assign y13876 = ~n30723 ;
  assign y13877 = ~n30729 ;
  assign y13878 = ~n30732 ;
  assign y13879 = n30733 ;
  assign y13880 = ~1'b0 ;
  assign y13881 = ~n30735 ;
  assign y13882 = ~n30736 ;
  assign y13883 = ~n30741 ;
  assign y13884 = n30745 ;
  assign y13885 = ~n30746 ;
  assign y13886 = ~n30747 ;
  assign y13887 = ~n30750 ;
  assign y13888 = ~n30756 ;
  assign y13889 = n30762 ;
  assign y13890 = n30765 ;
  assign y13891 = n30769 ;
  assign y13892 = n30771 ;
  assign y13893 = ~1'b0 ;
  assign y13894 = n30776 ;
  assign y13895 = ~n30778 ;
  assign y13896 = n10863 ;
  assign y13897 = ~n30779 ;
  assign y13898 = ~n19721 ;
  assign y13899 = ~n30782 ;
  assign y13900 = ~n30786 ;
  assign y13901 = ~1'b0 ;
  assign y13902 = n30787 ;
  assign y13903 = ~n30790 ;
  assign y13904 = n30791 ;
  assign y13905 = ~n30795 ;
  assign y13906 = ~n17168 ;
  assign y13907 = ~1'b0 ;
  assign y13908 = n30798 ;
  assign y13909 = n30799 ;
  assign y13910 = ~n30804 ;
  assign y13911 = ~1'b0 ;
  assign y13912 = ~n30805 ;
  assign y13913 = ~1'b0 ;
  assign y13914 = n30812 ;
  assign y13915 = ~1'b0 ;
  assign y13916 = n3308 ;
  assign y13917 = n30815 ;
  assign y13918 = n30816 ;
  assign y13919 = n30818 ;
  assign y13920 = n30819 ;
  assign y13921 = n30820 ;
  assign y13922 = n30822 ;
  assign y13923 = ~n30823 ;
  assign y13924 = n20956 ;
  assign y13925 = ~n30826 ;
  assign y13926 = n30829 ;
  assign y13927 = n30830 ;
  assign y13928 = n30832 ;
  assign y13929 = ~n30834 ;
  assign y13930 = n30840 ;
  assign y13931 = ~n30847 ;
  assign y13932 = n30850 ;
  assign y13933 = n30852 ;
  assign y13934 = n30854 ;
  assign y13935 = n30856 ;
  assign y13936 = ~n30868 ;
  assign y13937 = ~n30874 ;
  assign y13938 = n30878 ;
  assign y13939 = ~1'b0 ;
  assign y13940 = ~n30880 ;
  assign y13941 = n30886 ;
  assign y13942 = n30888 ;
  assign y13943 = ~n30889 ;
  assign y13944 = ~1'b0 ;
  assign y13945 = n30890 ;
  assign y13946 = ~n30892 ;
  assign y13947 = ~n30894 ;
  assign y13948 = ~n30897 ;
  assign y13949 = n30900 ;
  assign y13950 = ~n20300 ;
  assign y13951 = ~n30903 ;
  assign y13952 = ~1'b0 ;
  assign y13953 = ~1'b0 ;
  assign y13954 = ~n30905 ;
  assign y13955 = 1'b0 ;
  assign y13956 = n30907 ;
  assign y13957 = ~n30908 ;
  assign y13958 = n30909 ;
  assign y13959 = ~n30910 ;
  assign y13960 = n30913 ;
  assign y13961 = ~n30914 ;
  assign y13962 = ~1'b0 ;
  assign y13963 = ~1'b0 ;
  assign y13964 = ~1'b0 ;
  assign y13965 = ~n2955 ;
  assign y13966 = n30915 ;
  assign y13967 = ~n30920 ;
  assign y13968 = n30921 ;
  assign y13969 = n30923 ;
  assign y13970 = ~1'b0 ;
  assign y13971 = n30931 ;
  assign y13972 = n30932 ;
  assign y13973 = ~1'b0 ;
  assign y13974 = ~1'b0 ;
  assign y13975 = n14251 ;
  assign y13976 = ~n30934 ;
  assign y13977 = ~n30939 ;
  assign y13978 = ~1'b0 ;
  assign y13979 = n30941 ;
  assign y13980 = ~n30943 ;
  assign y13981 = ~n30947 ;
  assign y13982 = n30949 ;
  assign y13983 = ~1'b0 ;
  assign y13984 = ~1'b0 ;
  assign y13985 = n30951 ;
  assign y13986 = ~1'b0 ;
  assign y13987 = n30985 ;
  assign y13988 = ~n30986 ;
  assign y13989 = ~1'b0 ;
  assign y13990 = ~n30987 ;
  assign y13991 = ~n30989 ;
  assign y13992 = ~1'b0 ;
  assign y13993 = n30990 ;
  assign y13994 = ~n30994 ;
  assign y13995 = ~n30997 ;
  assign y13996 = ~n30999 ;
  assign y13997 = ~1'b0 ;
  assign y13998 = n31001 ;
  assign y13999 = ~n31002 ;
  assign y14000 = n31005 ;
  assign y14001 = n31010 ;
  assign y14002 = ~n31014 ;
  assign y14003 = ~1'b0 ;
  assign y14004 = ~1'b0 ;
  assign y14005 = n31015 ;
  assign y14006 = n31018 ;
  assign y14007 = ~1'b0 ;
  assign y14008 = n31022 ;
  assign y14009 = 1'b0 ;
  assign y14010 = ~1'b0 ;
  assign y14011 = ~n31025 ;
  assign y14012 = n17118 ;
  assign y14013 = ~n31026 ;
  assign y14014 = n31030 ;
  assign y14015 = ~n31031 ;
  assign y14016 = ~n31033 ;
  assign y14017 = ~1'b0 ;
  assign y14018 = n31034 ;
  assign y14019 = ~n6481 ;
  assign y14020 = n27085 ;
  assign y14021 = n31035 ;
  assign y14022 = n31037 ;
  assign y14023 = ~n31039 ;
  assign y14024 = ~n31041 ;
  assign y14025 = n31043 ;
  assign y14026 = n31057 ;
  assign y14027 = ~n31060 ;
  assign y14028 = n31066 ;
  assign y14029 = ~1'b0 ;
  assign y14030 = ~1'b0 ;
  assign y14031 = n31068 ;
  assign y14032 = ~n31074 ;
  assign y14033 = ~n31075 ;
  assign y14034 = ~n31076 ;
  assign y14035 = ~n31077 ;
  assign y14036 = ~n31079 ;
  assign y14037 = n31080 ;
  assign y14038 = ~1'b0 ;
  assign y14039 = ~n31086 ;
  assign y14040 = n31088 ;
  assign y14041 = ~1'b0 ;
  assign y14042 = ~n31089 ;
  assign y14043 = ~n31091 ;
  assign y14044 = n31093 ;
  assign y14045 = n31094 ;
  assign y14046 = n31098 ;
  assign y14047 = ~1'b0 ;
  assign y14048 = n31100 ;
  assign y14049 = n31102 ;
  assign y14050 = ~n31103 ;
  assign y14051 = n31104 ;
  assign y14052 = n31106 ;
  assign y14053 = ~1'b0 ;
  assign y14054 = ~1'b0 ;
  assign y14055 = ~1'b0 ;
  assign y14056 = ~1'b0 ;
  assign y14057 = ~n31109 ;
  assign y14058 = ~n26838 ;
  assign y14059 = n31111 ;
  assign y14060 = ~1'b0 ;
  assign y14061 = ~n31113 ;
  assign y14062 = n31116 ;
  assign y14063 = n31118 ;
  assign y14064 = n31119 ;
  assign y14065 = n31120 ;
  assign y14066 = ~n31121 ;
  assign y14067 = ~n31122 ;
  assign y14068 = ~n31127 ;
  assign y14069 = n31130 ;
  assign y14070 = ~1'b0 ;
  assign y14071 = n31131 ;
  assign y14072 = ~n31148 ;
  assign y14073 = ~n31151 ;
  assign y14074 = ~1'b0 ;
  assign y14075 = ~n31152 ;
  assign y14076 = ~1'b0 ;
  assign y14077 = ~1'b0 ;
  assign y14078 = n31157 ;
  assign y14079 = ~1'b0 ;
  assign y14080 = n31158 ;
  assign y14081 = ~n31160 ;
  assign y14082 = ~n31161 ;
  assign y14083 = n31163 ;
  assign y14084 = n31166 ;
  assign y14085 = ~n31169 ;
  assign y14086 = ~n31170 ;
  assign y14087 = ~n31173 ;
  assign y14088 = ~n17001 ;
  assign y14089 = ~n31177 ;
  assign y14090 = n31179 ;
  assign y14091 = ~n31182 ;
  assign y14092 = ~n31184 ;
  assign y14093 = ~n31186 ;
  assign y14094 = ~n31190 ;
  assign y14095 = n31191 ;
  assign y14096 = n31192 ;
  assign y14097 = ~n31195 ;
  assign y14098 = ~n31197 ;
  assign y14099 = ~n31199 ;
  assign y14100 = n26410 ;
  assign y14101 = ~n31206 ;
  assign y14102 = ~1'b0 ;
  assign y14103 = ~1'b0 ;
  assign y14104 = n31208 ;
  assign y14105 = ~1'b0 ;
  assign y14106 = ~1'b0 ;
  assign y14107 = ~n31210 ;
  assign y14108 = ~n22803 ;
  assign y14109 = ~1'b0 ;
  assign y14110 = n31211 ;
  assign y14111 = ~n31213 ;
  assign y14112 = n31214 ;
  assign y14113 = n2024 ;
  assign y14114 = ~n31218 ;
  assign y14115 = n31223 ;
  assign y14116 = ~1'b0 ;
  assign y14117 = ~1'b0 ;
  assign y14118 = n31224 ;
  assign y14119 = ~n6244 ;
  assign y14120 = ~n31227 ;
  assign y14121 = n31229 ;
  assign y14122 = ~n31232 ;
  assign y14123 = ~1'b0 ;
  assign y14124 = ~1'b0 ;
  assign y14125 = n31233 ;
  assign y14126 = ~n31235 ;
  assign y14127 = n31237 ;
  assign y14128 = ~n31239 ;
  assign y14129 = ~1'b0 ;
  assign y14130 = ~1'b0 ;
  assign y14131 = ~1'b0 ;
  assign y14132 = n31241 ;
  assign y14133 = ~n686 ;
  assign y14134 = ~n31245 ;
  assign y14135 = n31247 ;
  assign y14136 = ~1'b0 ;
  assign y14137 = ~1'b0 ;
  assign y14138 = ~n31253 ;
  assign y14139 = n31254 ;
  assign y14140 = n31260 ;
  assign y14141 = n31264 ;
  assign y14142 = ~1'b0 ;
  assign y14143 = n14165 ;
  assign y14144 = ~n22475 ;
  assign y14145 = ~1'b0 ;
  assign y14146 = n31265 ;
  assign y14147 = n31266 ;
  assign y14148 = ~n31270 ;
  assign y14149 = ~n31272 ;
  assign y14150 = ~1'b0 ;
  assign y14151 = ~1'b0 ;
  assign y14152 = ~1'b0 ;
  assign y14153 = n31273 ;
  assign y14154 = ~n31277 ;
  assign y14155 = n31280 ;
  assign y14156 = n31284 ;
  assign y14157 = 1'b0 ;
  assign y14158 = ~1'b0 ;
  assign y14159 = n31286 ;
  assign y14160 = n31287 ;
  assign y14161 = ~1'b0 ;
  assign y14162 = n31291 ;
  assign y14163 = n31292 ;
  assign y14164 = ~n31300 ;
  assign y14165 = ~1'b0 ;
  assign y14166 = n31303 ;
  assign y14167 = 1'b0 ;
  assign y14168 = n31306 ;
  assign y14169 = ~n397 ;
  assign y14170 = ~1'b0 ;
  assign y14171 = ~1'b0 ;
  assign y14172 = ~n31308 ;
  assign y14173 = ~1'b0 ;
  assign y14174 = n31313 ;
  assign y14175 = n31316 ;
  assign y14176 = n31318 ;
  assign y14177 = n31320 ;
  assign y14178 = ~1'b0 ;
  assign y14179 = n23471 ;
  assign y14180 = ~n31321 ;
  assign y14181 = n31327 ;
  assign y14182 = n31330 ;
  assign y14183 = ~1'b0 ;
  assign y14184 = n31331 ;
  assign y14185 = n31336 ;
  assign y14186 = ~1'b0 ;
  assign y14187 = ~1'b0 ;
  assign y14188 = ~1'b0 ;
  assign y14189 = ~n31340 ;
  assign y14190 = ~n31344 ;
  assign y14191 = ~n31345 ;
  assign y14192 = ~1'b0 ;
  assign y14193 = ~1'b0 ;
  assign y14194 = ~n31348 ;
  assign y14195 = ~n31355 ;
  assign y14196 = n31357 ;
  assign y14197 = ~n31359 ;
  assign y14198 = ~1'b0 ;
  assign y14199 = ~n31362 ;
  assign y14200 = ~1'b0 ;
  assign y14201 = n31367 ;
  assign y14202 = n31368 ;
  assign y14203 = ~n31369 ;
  assign y14204 = ~n31371 ;
  assign y14205 = n31372 ;
  assign y14206 = ~1'b0 ;
  assign y14207 = ~n31373 ;
  assign y14208 = ~1'b0 ;
  assign y14209 = n31375 ;
  assign y14210 = ~n31377 ;
  assign y14211 = n31378 ;
  assign y14212 = ~n31379 ;
  assign y14213 = ~1'b0 ;
  assign y14214 = ~n31385 ;
  assign y14215 = n31386 ;
  assign y14216 = n31390 ;
  assign y14217 = ~n31392 ;
  assign y14218 = ~n31394 ;
  assign y14219 = n31395 ;
  assign y14220 = n31399 ;
  assign y14221 = ~n31401 ;
  assign y14222 = ~n31402 ;
  assign y14223 = ~n31406 ;
  assign y14224 = ~n31409 ;
  assign y14225 = ~1'b0 ;
  assign y14226 = n31410 ;
  assign y14227 = n31413 ;
  assign y14228 = ~n31423 ;
  assign y14229 = n31424 ;
  assign y14230 = n31426 ;
  assign y14231 = ~1'b0 ;
  assign y14232 = ~n31428 ;
  assign y14233 = ~1'b0 ;
  assign y14234 = ~1'b0 ;
  assign y14235 = ~n31430 ;
  assign y14236 = ~n31434 ;
  assign y14237 = ~n31435 ;
  assign y14238 = ~1'b0 ;
  assign y14239 = ~1'b0 ;
  assign y14240 = ~1'b0 ;
  assign y14241 = n31436 ;
  assign y14242 = ~n31437 ;
  assign y14243 = n31438 ;
  assign y14244 = ~n31441 ;
  assign y14245 = ~n31445 ;
  assign y14246 = n31446 ;
  assign y14247 = ~n31449 ;
  assign y14248 = n31450 ;
  assign y14249 = n31452 ;
  assign y14250 = ~n12411 ;
  assign y14251 = n31455 ;
  assign y14252 = n31457 ;
  assign y14253 = ~n31459 ;
  assign y14254 = ~1'b0 ;
  assign y14255 = ~n29720 ;
  assign y14256 = n31460 ;
  assign y14257 = ~n31462 ;
  assign y14258 = n31465 ;
  assign y14259 = ~n31470 ;
  assign y14260 = ~n31473 ;
  assign y14261 = ~n31477 ;
  assign y14262 = 1'b0 ;
  assign y14263 = ~n31482 ;
  assign y14264 = n31484 ;
  assign y14265 = ~1'b0 ;
  assign y14266 = n31489 ;
  assign y14267 = ~1'b0 ;
  assign y14268 = ~n17296 ;
  assign y14269 = ~1'b0 ;
  assign y14270 = ~1'b0 ;
  assign y14271 = ~n31491 ;
  assign y14272 = ~n31494 ;
  assign y14273 = ~n31495 ;
  assign y14274 = n31498 ;
  assign y14275 = n31499 ;
  assign y14276 = ~1'b0 ;
  assign y14277 = ~n21790 ;
  assign y14278 = n31500 ;
  assign y14279 = ~1'b0 ;
  assign y14280 = ~n31511 ;
  assign y14281 = ~n31513 ;
  assign y14282 = n31515 ;
  assign y14283 = ~1'b0 ;
  assign y14284 = ~1'b0 ;
  assign y14285 = ~n31516 ;
  assign y14286 = ~1'b0 ;
  assign y14287 = n28982 ;
  assign y14288 = n5822 ;
  assign y14289 = n31520 ;
  assign y14290 = ~n31521 ;
  assign y14291 = n31523 ;
  assign y14292 = ~1'b0 ;
  assign y14293 = n31527 ;
  assign y14294 = ~n31529 ;
  assign y14295 = n31531 ;
  assign y14296 = ~n31536 ;
  assign y14297 = ~n31541 ;
  assign y14298 = ~n31543 ;
  assign y14299 = ~1'b0 ;
  assign y14300 = ~n31546 ;
  assign y14301 = n31547 ;
  assign y14302 = n31550 ;
  assign y14303 = ~n31552 ;
  assign y14304 = ~n9074 ;
  assign y14305 = ~n31554 ;
  assign y14306 = ~1'b0 ;
  assign y14307 = n31555 ;
  assign y14308 = ~1'b0 ;
  assign y14309 = ~1'b0 ;
  assign y14310 = ~n31561 ;
  assign y14311 = n31562 ;
  assign y14312 = ~n31563 ;
  assign y14313 = ~1'b0 ;
  assign y14314 = ~n31564 ;
  assign y14315 = ~1'b0 ;
  assign y14316 = ~n31566 ;
  assign y14317 = ~1'b0 ;
  assign y14318 = ~1'b0 ;
  assign y14319 = ~n31567 ;
  assign y14320 = ~n31568 ;
  assign y14321 = ~n16054 ;
  assign y14322 = ~n31569 ;
  assign y14323 = ~n31571 ;
  assign y14324 = ~1'b0 ;
  assign y14325 = ~1'b0 ;
  assign y14326 = n31572 ;
  assign y14327 = n31575 ;
  assign y14328 = ~n31578 ;
  assign y14329 = n31580 ;
  assign y14330 = ~n31583 ;
  assign y14331 = ~1'b0 ;
  assign y14332 = n31584 ;
  assign y14333 = n31586 ;
  assign y14334 = n31587 ;
  assign y14335 = n31589 ;
  assign y14336 = ~1'b0 ;
  assign y14337 = ~n31590 ;
  assign y14338 = n26986 ;
  assign y14339 = ~n31592 ;
  assign y14340 = ~n31594 ;
  assign y14341 = 1'b0 ;
  assign y14342 = ~1'b0 ;
  assign y14343 = ~1'b0 ;
  assign y14344 = ~n31596 ;
  assign y14345 = n31597 ;
  assign y14346 = ~n31598 ;
  assign y14347 = ~n31601 ;
  assign y14348 = ~n31602 ;
  assign y14349 = ~n31606 ;
  assign y14350 = n31609 ;
  assign y14351 = ~n31614 ;
  assign y14352 = ~1'b0 ;
  assign y14353 = ~1'b0 ;
  assign y14354 = ~n31615 ;
  assign y14355 = n31616 ;
  assign y14356 = ~1'b0 ;
  assign y14357 = ~n31618 ;
  assign y14358 = n31620 ;
  assign y14359 = ~n31621 ;
  assign y14360 = ~n31631 ;
  assign y14361 = ~1'b0 ;
  assign y14362 = n31632 ;
  assign y14363 = ~n31637 ;
  assign y14364 = ~n31642 ;
  assign y14365 = ~1'b0 ;
  assign y14366 = n31644 ;
  assign y14367 = ~1'b0 ;
  assign y14368 = ~1'b0 ;
  assign y14369 = n31647 ;
  assign y14370 = n31651 ;
  assign y14371 = ~1'b0 ;
  assign y14372 = n31652 ;
  assign y14373 = ~n31658 ;
  assign y14374 = n31659 ;
  assign y14375 = ~n31661 ;
  assign y14376 = n31663 ;
  assign y14377 = ~n31664 ;
  assign y14378 = ~n31665 ;
  assign y14379 = ~n31666 ;
  assign y14380 = ~1'b0 ;
  assign y14381 = ~1'b0 ;
  assign y14382 = ~1'b0 ;
  assign y14383 = n31670 ;
  assign y14384 = n31672 ;
  assign y14385 = ~n31673 ;
  assign y14386 = ~n31674 ;
  assign y14387 = ~1'b0 ;
  assign y14388 = ~n31677 ;
  assign y14389 = ~n31678 ;
  assign y14390 = ~n1976 ;
  assign y14391 = ~n31680 ;
  assign y14392 = n5375 ;
  assign y14393 = ~n23960 ;
  assign y14394 = ~n31684 ;
  assign y14395 = n31685 ;
  assign y14396 = n31690 ;
  assign y14397 = ~n31691 ;
  assign y14398 = n31695 ;
  assign y14399 = n18289 ;
  assign y14400 = n31697 ;
  assign y14401 = ~n31701 ;
  assign y14402 = ~1'b0 ;
  assign y14403 = ~1'b0 ;
  assign y14404 = ~1'b0 ;
  assign y14405 = n31703 ;
  assign y14406 = ~n31704 ;
  assign y14407 = n31706 ;
  assign y14408 = ~n31707 ;
  assign y14409 = ~1'b0 ;
  assign y14410 = n31708 ;
  assign y14411 = ~1'b0 ;
  assign y14412 = n31712 ;
  assign y14413 = ~1'b0 ;
  assign y14414 = ~1'b0 ;
  assign y14415 = n31714 ;
  assign y14416 = ~n31715 ;
  assign y14417 = n31717 ;
  assign y14418 = n31719 ;
  assign y14419 = ~n31723 ;
  assign y14420 = ~1'b0 ;
  assign y14421 = ~1'b0 ;
  assign y14422 = n31725 ;
  assign y14423 = ~n31727 ;
  assign y14424 = ~1'b0 ;
  assign y14425 = ~n31730 ;
  assign y14426 = ~n31731 ;
  assign y14427 = ~n31732 ;
  assign y14428 = ~1'b0 ;
  assign y14429 = ~1'b0 ;
  assign y14430 = 1'b0 ;
  assign y14431 = n31733 ;
  assign y14432 = ~1'b0 ;
  assign y14433 = n31734 ;
  assign y14434 = ~n31735 ;
  assign y14435 = n31736 ;
  assign y14436 = n31743 ;
  assign y14437 = ~1'b0 ;
  assign y14438 = n31744 ;
  assign y14439 = ~n31745 ;
  assign y14440 = n31746 ;
  assign y14441 = n31748 ;
  assign y14442 = ~n31749 ;
  assign y14443 = ~n31755 ;
  assign y14444 = 1'b0 ;
  assign y14445 = ~n31758 ;
  assign y14446 = n31760 ;
  assign y14447 = ~n31761 ;
  assign y14448 = ~1'b0 ;
  assign y14449 = ~n31762 ;
  assign y14450 = ~n31763 ;
  assign y14451 = ~n31765 ;
  assign y14452 = ~1'b0 ;
  assign y14453 = ~n31772 ;
  assign y14454 = n31776 ;
  assign y14455 = n31777 ;
  assign y14456 = ~n31779 ;
  assign y14457 = n31780 ;
  assign y14458 = ~n17486 ;
  assign y14459 = n31781 ;
  assign y14460 = ~1'b0 ;
  assign y14461 = ~1'b0 ;
  assign y14462 = n31785 ;
  assign y14463 = ~n22674 ;
  assign y14464 = ~n31786 ;
  assign y14465 = n31787 ;
  assign y14466 = ~n31788 ;
  assign y14467 = ~1'b0 ;
  assign y14468 = ~n31790 ;
  assign y14469 = n31793 ;
  assign y14470 = ~n31795 ;
  assign y14471 = n31797 ;
  assign y14472 = ~n31799 ;
  assign y14473 = n31801 ;
  assign y14474 = n27270 ;
  assign y14475 = n31803 ;
  assign y14476 = ~1'b0 ;
  assign y14477 = ~1'b0 ;
  assign y14478 = ~n31804 ;
  assign y14479 = n31805 ;
  assign y14480 = ~1'b0 ;
  assign y14481 = ~n31807 ;
  assign y14482 = ~n31811 ;
  assign y14483 = n31814 ;
  assign y14484 = n31826 ;
  assign y14485 = n31827 ;
  assign y14486 = ~n31828 ;
  assign y14487 = n31829 ;
  assign y14488 = n31830 ;
  assign y14489 = ~1'b0 ;
  assign y14490 = ~n31835 ;
  assign y14491 = n31841 ;
  assign y14492 = n31843 ;
  assign y14493 = ~n11446 ;
  assign y14494 = 1'b0 ;
  assign y14495 = ~n31844 ;
  assign y14496 = ~n10360 ;
  assign y14497 = n31848 ;
  assign y14498 = ~1'b0 ;
  assign y14499 = n31849 ;
  assign y14500 = ~n3711 ;
  assign y14501 = n31852 ;
  assign y14502 = ~n31856 ;
  assign y14503 = ~n31859 ;
  assign y14504 = ~1'b0 ;
  assign y14505 = ~1'b0 ;
  assign y14506 = ~n31863 ;
  assign y14507 = ~n31867 ;
  assign y14508 = ~n31868 ;
  assign y14509 = ~1'b0 ;
  assign y14510 = ~n31873 ;
  assign y14511 = 1'b0 ;
  assign y14512 = n31875 ;
  assign y14513 = ~1'b0 ;
  assign y14514 = ~1'b0 ;
  assign y14515 = n31878 ;
  assign y14516 = n31879 ;
  assign y14517 = ~n31883 ;
  assign y14518 = ~1'b0 ;
  assign y14519 = n31884 ;
  assign y14520 = n31886 ;
  assign y14521 = ~1'b0 ;
  assign y14522 = ~n31888 ;
  assign y14523 = n31889 ;
  assign y14524 = n31891 ;
  assign y14525 = n31893 ;
  assign y14526 = ~n31894 ;
  assign y14527 = n31896 ;
  assign y14528 = ~n31897 ;
  assign y14529 = ~1'b0 ;
  assign y14530 = 1'b0 ;
  assign y14531 = ~n31900 ;
  assign y14532 = ~n31901 ;
  assign y14533 = n31902 ;
  assign y14534 = n31905 ;
  assign y14535 = ~n31907 ;
  assign y14536 = n31909 ;
  assign y14537 = n31917 ;
  assign y14538 = ~n31920 ;
  assign y14539 = ~1'b0 ;
  assign y14540 = ~n4679 ;
  assign y14541 = n31922 ;
  assign y14542 = ~n31924 ;
  assign y14543 = n31929 ;
  assign y14544 = ~1'b0 ;
  assign y14545 = ~n31932 ;
  assign y14546 = ~n31941 ;
  assign y14547 = n31945 ;
  assign y14548 = ~n31947 ;
  assign y14549 = ~n31951 ;
  assign y14550 = ~1'b0 ;
  assign y14551 = n31954 ;
  assign y14552 = n31960 ;
  assign y14553 = n31961 ;
  assign y14554 = ~n1595 ;
  assign y14555 = ~n19966 ;
  assign y14556 = ~1'b0 ;
  assign y14557 = ~1'b0 ;
  assign y14558 = n31970 ;
  assign y14559 = n31973 ;
  assign y14560 = n31974 ;
  assign y14561 = n31978 ;
  assign y14562 = ~n31980 ;
  assign y14563 = n31985 ;
  assign y14564 = n31989 ;
  assign y14565 = ~n31990 ;
  assign y14566 = n31991 ;
  assign y14567 = ~n31996 ;
  assign y14568 = ~n32000 ;
  assign y14569 = ~n32003 ;
  assign y14570 = ~n32004 ;
  assign y14571 = ~n32014 ;
  assign y14572 = ~n32016 ;
  assign y14573 = n32021 ;
  assign y14574 = ~n32024 ;
  assign y14575 = ~n32028 ;
  assign y14576 = n14980 ;
  assign y14577 = ~1'b0 ;
  assign y14578 = 1'b0 ;
  assign y14579 = ~n32029 ;
  assign y14580 = n32030 ;
  assign y14581 = ~n32033 ;
  assign y14582 = ~1'b0 ;
  assign y14583 = n32037 ;
  assign y14584 = ~n32041 ;
  assign y14585 = n32042 ;
  assign y14586 = ~n32055 ;
  assign y14587 = ~n32056 ;
  assign y14588 = ~n32061 ;
  assign y14589 = n32064 ;
  assign y14590 = n32068 ;
  assign y14591 = n32071 ;
  assign y14592 = ~n32075 ;
  assign y14593 = ~1'b0 ;
  assign y14594 = ~n32077 ;
  assign y14595 = ~n32078 ;
  assign y14596 = ~n32082 ;
  assign y14597 = n32083 ;
  assign y14598 = ~1'b0 ;
  assign y14599 = ~n32086 ;
  assign y14600 = ~n32089 ;
  assign y14601 = ~1'b0 ;
  assign y14602 = ~1'b0 ;
  assign y14603 = n32090 ;
  assign y14604 = ~1'b0 ;
  assign y14605 = ~1'b0 ;
  assign y14606 = ~1'b0 ;
  assign y14607 = n32091 ;
  assign y14608 = n32093 ;
  assign y14609 = ~n32094 ;
  assign y14610 = n32097 ;
  assign y14611 = n32101 ;
  assign y14612 = ~1'b0 ;
  assign y14613 = n32106 ;
  assign y14614 = n32112 ;
  assign y14615 = n32115 ;
  assign y14616 = n32119 ;
  assign y14617 = n32120 ;
  assign y14618 = 1'b0 ;
  assign y14619 = n32121 ;
  assign y14620 = n32122 ;
  assign y14621 = ~n32127 ;
  assign y14622 = ~1'b0 ;
  assign y14623 = ~1'b0 ;
  assign y14624 = ~1'b0 ;
  assign y14625 = n32129 ;
  assign y14626 = ~1'b0 ;
  assign y14627 = n32134 ;
  assign y14628 = ~n32137 ;
  assign y14629 = ~1'b0 ;
  assign y14630 = n32139 ;
  assign y14631 = n32143 ;
  assign y14632 = ~n32144 ;
  assign y14633 = n32145 ;
  assign y14634 = ~n32148 ;
  assign y14635 = ~n32151 ;
  assign y14636 = ~n32152 ;
  assign y14637 = ~1'b0 ;
  assign y14638 = ~n32155 ;
  assign y14639 = n32158 ;
  assign y14640 = n32162 ;
  assign y14641 = ~n32166 ;
  assign y14642 = ~n32167 ;
  assign y14643 = n32168 ;
  assign y14644 = ~n32174 ;
  assign y14645 = ~n32178 ;
  assign y14646 = n32180 ;
  assign y14647 = n32181 ;
  assign y14648 = n32182 ;
  assign y14649 = n32184 ;
  assign y14650 = n32194 ;
  assign y14651 = ~1'b0 ;
  assign y14652 = n32195 ;
  assign y14653 = n32199 ;
  assign y14654 = n32200 ;
  assign y14655 = ~n32203 ;
  assign y14656 = ~n32204 ;
  assign y14657 = n32214 ;
  assign y14658 = ~n32223 ;
  assign y14659 = 1'b0 ;
  assign y14660 = n32227 ;
  assign y14661 = n32231 ;
  assign y14662 = ~1'b0 ;
  assign y14663 = n32233 ;
  assign y14664 = n32238 ;
  assign y14665 = ~n32242 ;
  assign y14666 = ~n32243 ;
  assign y14667 = ~1'b0 ;
  assign y14668 = ~1'b0 ;
  assign y14669 = n14468 ;
  assign y14670 = ~1'b0 ;
  assign y14671 = n32245 ;
  assign y14672 = n32246 ;
  assign y14673 = ~n32248 ;
  assign y14674 = ~1'b0 ;
  assign y14675 = n32254 ;
  assign y14676 = n32255 ;
  assign y14677 = ~1'b0 ;
  assign y14678 = n32258 ;
  assign y14679 = ~n32261 ;
  assign y14680 = ~1'b0 ;
  assign y14681 = ~n32265 ;
  assign y14682 = n32267 ;
  assign y14683 = n32271 ;
  assign y14684 = ~1'b0 ;
  assign y14685 = ~1'b0 ;
  assign y14686 = n32272 ;
  assign y14687 = n32273 ;
  assign y14688 = ~n32276 ;
  assign y14689 = n32278 ;
  assign y14690 = ~n32283 ;
  assign y14691 = ~1'b0 ;
  assign y14692 = ~n32285 ;
  assign y14693 = ~1'b0 ;
  assign y14694 = n32286 ;
  assign y14695 = ~n32287 ;
  assign y14696 = ~n32289 ;
  assign y14697 = n32291 ;
  assign y14698 = ~n32295 ;
  assign y14699 = ~n32297 ;
  assign y14700 = n32299 ;
  assign y14701 = n32300 ;
  assign y14702 = ~n32302 ;
  assign y14703 = ~1'b0 ;
  assign y14704 = ~n32307 ;
  assign y14705 = ~n32315 ;
  assign y14706 = n32319 ;
  assign y14707 = ~n32321 ;
  assign y14708 = n32324 ;
  assign y14709 = ~1'b0 ;
  assign y14710 = 1'b0 ;
  assign y14711 = ~n32326 ;
  assign y14712 = ~1'b0 ;
  assign y14713 = n1952 ;
  assign y14714 = ~n32330 ;
  assign y14715 = ~1'b0 ;
  assign y14716 = n32333 ;
  assign y14717 = n32334 ;
  assign y14718 = n32335 ;
  assign y14719 = n32336 ;
  assign y14720 = ~n32337 ;
  assign y14721 = n32340 ;
  assign y14722 = n32344 ;
  assign y14723 = n32346 ;
  assign y14724 = ~1'b0 ;
  assign y14725 = ~n32353 ;
  assign y14726 = ~1'b0 ;
  assign y14727 = ~n32355 ;
  assign y14728 = ~n32356 ;
  assign y14729 = ~n32357 ;
  assign y14730 = ~n32360 ;
  assign y14731 = ~n32361 ;
  assign y14732 = ~1'b0 ;
  assign y14733 = n6833 ;
  assign y14734 = ~n32364 ;
  assign y14735 = n32366 ;
  assign y14736 = ~n32368 ;
  assign y14737 = n32370 ;
  assign y14738 = n32374 ;
  assign y14739 = n32376 ;
  assign y14740 = ~n32377 ;
  assign y14741 = ~n32379 ;
  assign y14742 = n32380 ;
  assign y14743 = n32381 ;
  assign y14744 = ~n32383 ;
  assign y14745 = ~1'b0 ;
  assign y14746 = ~1'b0 ;
  assign y14747 = ~1'b0 ;
  assign y14748 = n32386 ;
  assign y14749 = ~n32396 ;
  assign y14750 = ~1'b0 ;
  assign y14751 = n32400 ;
  assign y14752 = n32402 ;
  assign y14753 = n32404 ;
  assign y14754 = ~n32408 ;
  assign y14755 = ~n32410 ;
  assign y14756 = ~n32411 ;
  assign y14757 = ~1'b0 ;
  assign y14758 = ~n32415 ;
  assign y14759 = n32416 ;
  assign y14760 = ~1'b0 ;
  assign y14761 = ~n32419 ;
  assign y14762 = n32423 ;
  assign y14763 = ~1'b0 ;
  assign y14764 = ~n32425 ;
  assign y14765 = n32427 ;
  assign y14766 = n32428 ;
  assign y14767 = n32429 ;
  assign y14768 = n32437 ;
  assign y14769 = ~n32439 ;
  assign y14770 = n32442 ;
  assign y14771 = ~1'b0 ;
  assign y14772 = ~n32444 ;
  assign y14773 = ~1'b0 ;
  assign y14774 = ~n32447 ;
  assign y14775 = n32448 ;
  assign y14776 = ~n32450 ;
  assign y14777 = ~n32452 ;
  assign y14778 = n32453 ;
  assign y14779 = ~n32456 ;
  assign y14780 = ~1'b0 ;
  assign y14781 = ~n32460 ;
  assign y14782 = ~n32464 ;
  assign y14783 = n32466 ;
  assign y14784 = ~n32469 ;
  assign y14785 = ~n32470 ;
  assign y14786 = n32472 ;
  assign y14787 = ~n32475 ;
  assign y14788 = n32479 ;
  assign y14789 = n32481 ;
  assign y14790 = n32485 ;
  assign y14791 = n2447 ;
  assign y14792 = ~1'b0 ;
  assign y14793 = n18694 ;
  assign y14794 = ~1'b0 ;
  assign y14795 = ~n32489 ;
  assign y14796 = ~n26834 ;
  assign y14797 = n32493 ;
  assign y14798 = ~n7617 ;
  assign y14799 = n32503 ;
  assign y14800 = ~n32505 ;
  assign y14801 = ~n32509 ;
  assign y14802 = n32511 ;
  assign y14803 = ~n32513 ;
  assign y14804 = ~n32515 ;
  assign y14805 = ~n32516 ;
  assign y14806 = ~n32520 ;
  assign y14807 = ~1'b0 ;
  assign y14808 = ~1'b0 ;
  assign y14809 = ~1'b0 ;
  assign y14810 = n32528 ;
  assign y14811 = ~n32529 ;
  assign y14812 = ~1'b0 ;
  assign y14813 = ~1'b0 ;
  assign y14814 = n32531 ;
  assign y14815 = n32532 ;
  assign y14816 = ~n32535 ;
  assign y14817 = ~n32537 ;
  assign y14818 = n32539 ;
  assign y14819 = n32540 ;
  assign y14820 = ~1'b0 ;
  assign y14821 = ~1'b0 ;
  assign y14822 = ~n32542 ;
  assign y14823 = n32551 ;
  assign y14824 = ~n32552 ;
  assign y14825 = ~n32553 ;
  assign y14826 = ~n32556 ;
  assign y14827 = ~n32557 ;
  assign y14828 = ~1'b0 ;
  assign y14829 = ~1'b0 ;
  assign y14830 = ~n32559 ;
  assign y14831 = n32560 ;
  assign y14832 = n32561 ;
  assign y14833 = n32565 ;
  assign y14834 = ~n32566 ;
  assign y14835 = ~n32572 ;
  assign y14836 = ~1'b0 ;
  assign y14837 = n32573 ;
  assign y14838 = ~1'b0 ;
  assign y14839 = ~n32574 ;
  assign y14840 = ~n32579 ;
  assign y14841 = n32581 ;
  assign y14842 = ~1'b0 ;
  assign y14843 = ~1'b0 ;
  assign y14844 = n32582 ;
  assign y14845 = n32584 ;
  assign y14846 = n32590 ;
  assign y14847 = n32591 ;
  assign y14848 = n32593 ;
  assign y14849 = n32597 ;
  assign y14850 = n32598 ;
  assign y14851 = ~1'b0 ;
  assign y14852 = ~1'b0 ;
  assign y14853 = ~n32600 ;
  assign y14854 = n32601 ;
  assign y14855 = ~n32603 ;
  assign y14856 = ~n32605 ;
  assign y14857 = ~n32606 ;
  assign y14858 = n29129 ;
  assign y14859 = ~1'b0 ;
  assign y14860 = ~n32608 ;
  assign y14861 = n32612 ;
  assign y14862 = ~1'b0 ;
  assign y14863 = n32613 ;
  assign y14864 = ~n32614 ;
  assign y14865 = ~n32617 ;
  assign y14866 = ~n32623 ;
  assign y14867 = n32624 ;
  assign y14868 = n32629 ;
  assign y14869 = n32630 ;
  assign y14870 = ~1'b0 ;
  assign y14871 = ~n32633 ;
  assign y14872 = ~1'b0 ;
  assign y14873 = n12718 ;
  assign y14874 = ~n32635 ;
  assign y14875 = n32636 ;
  assign y14876 = ~x123 ;
  assign y14877 = n32638 ;
  assign y14878 = ~1'b0 ;
  assign y14879 = n32640 ;
  assign y14880 = n32641 ;
  assign y14881 = n32643 ;
  assign y14882 = ~n32644 ;
  assign y14883 = ~n20339 ;
  assign y14884 = ~1'b0 ;
  assign y14885 = n32649 ;
  assign y14886 = n32650 ;
  assign y14887 = ~1'b0 ;
  assign y14888 = n32651 ;
  assign y14889 = n32654 ;
  assign y14890 = n32655 ;
  assign y14891 = ~n20359 ;
  assign y14892 = n32662 ;
  assign y14893 = ~1'b0 ;
  assign y14894 = ~n32667 ;
  assign y14895 = ~n32670 ;
  assign y14896 = n32676 ;
  assign y14897 = ~n32677 ;
  assign y14898 = ~n16964 ;
  assign y14899 = ~1'b0 ;
  assign y14900 = n32680 ;
  assign y14901 = n32683 ;
  assign y14902 = n32685 ;
  assign y14903 = ~n32688 ;
  assign y14904 = n32689 ;
  assign y14905 = ~n32693 ;
  assign y14906 = ~1'b0 ;
  assign y14907 = n32694 ;
  assign y14908 = n32701 ;
  assign y14909 = n32703 ;
  assign y14910 = 1'b0 ;
  assign y14911 = n32710 ;
  assign y14912 = n32711 ;
  assign y14913 = ~n32716 ;
  assign y14914 = ~1'b0 ;
  assign y14915 = ~n28222 ;
  assign y14916 = ~1'b0 ;
  assign y14917 = ~n32719 ;
  assign y14918 = ~1'b0 ;
  assign y14919 = ~n32720 ;
  assign y14920 = n32722 ;
  assign y14921 = ~n32723 ;
  assign y14922 = n32724 ;
  assign y14923 = ~n32725 ;
  assign y14924 = ~n32726 ;
  assign y14925 = ~1'b0 ;
  assign y14926 = ~n32727 ;
  assign y14927 = n32728 ;
  assign y14928 = n32730 ;
  assign y14929 = ~n5365 ;
  assign y14930 = n32733 ;
  assign y14931 = ~1'b0 ;
  assign y14932 = ~n32740 ;
  assign y14933 = ~1'b0 ;
  assign y14934 = n32742 ;
  assign y14935 = 1'b0 ;
  assign y14936 = ~n32743 ;
  assign y14937 = n32746 ;
  assign y14938 = n32747 ;
  assign y14939 = n28038 ;
  assign y14940 = ~1'b0 ;
  assign y14941 = ~1'b0 ;
  assign y14942 = n32750 ;
  assign y14943 = ~1'b0 ;
  assign y14944 = n32751 ;
  assign y14945 = ~1'b0 ;
  assign y14946 = ~n32754 ;
  assign y14947 = n32757 ;
  assign y14948 = n32760 ;
  assign y14949 = ~n32763 ;
  assign y14950 = ~n1922 ;
  assign y14951 = ~n32764 ;
  assign y14952 = ~n32765 ;
  assign y14953 = n9639 ;
  assign y14954 = ~1'b0 ;
  assign y14955 = ~n32767 ;
  assign y14956 = ~n32769 ;
  assign y14957 = n32771 ;
  assign y14958 = ~n32773 ;
  assign y14959 = ~1'b0 ;
  assign y14960 = ~1'b0 ;
  assign y14961 = ~1'b0 ;
  assign y14962 = n32774 ;
  assign y14963 = ~n32775 ;
  assign y14964 = ~n32776 ;
  assign y14965 = n32778 ;
  assign y14966 = n32780 ;
  assign y14967 = ~1'b0 ;
  assign y14968 = ~n32782 ;
  assign y14969 = ~n32784 ;
  assign y14970 = ~1'b0 ;
  assign y14971 = ~n32785 ;
  assign y14972 = n32787 ;
  assign y14973 = ~n32789 ;
  assign y14974 = ~n32793 ;
  assign y14975 = ~1'b0 ;
  assign y14976 = ~n32796 ;
  assign y14977 = ~n32797 ;
  assign y14978 = ~n32800 ;
  assign y14979 = ~n32802 ;
  assign y14980 = n32803 ;
  assign y14981 = n32806 ;
  assign y14982 = n32810 ;
  assign y14983 = n19631 ;
  assign y14984 = n32812 ;
  assign y14985 = ~1'b0 ;
  assign y14986 = n32815 ;
  assign y14987 = ~1'b0 ;
  assign y14988 = ~n32820 ;
  assign y14989 = ~n32822 ;
  assign y14990 = n32823 ;
  assign y14991 = ~n32827 ;
  assign y14992 = ~n32829 ;
  assign y14993 = ~1'b0 ;
  assign y14994 = ~n20397 ;
  assign y14995 = ~1'b0 ;
  assign y14996 = n32830 ;
  assign y14997 = ~1'b0 ;
  assign y14998 = ~n32834 ;
  assign y14999 = ~n32839 ;
  assign y15000 = ~n1681 ;
  assign y15001 = ~n32841 ;
  assign y15002 = n32843 ;
  assign y15003 = ~1'b0 ;
  assign y15004 = n32844 ;
  assign y15005 = n32846 ;
  assign y15006 = n32848 ;
  assign y15007 = n32850 ;
  assign y15008 = ~1'b0 ;
  assign y15009 = n32852 ;
  assign y15010 = n32854 ;
  assign y15011 = n32856 ;
  assign y15012 = ~n32863 ;
  assign y15013 = ~n32864 ;
  assign y15014 = ~n32867 ;
  assign y15015 = n32869 ;
  assign y15016 = ~n32880 ;
  assign y15017 = ~1'b0 ;
  assign y15018 = 1'b0 ;
  assign y15019 = ~n32882 ;
  assign y15020 = ~1'b0 ;
  assign y15021 = n32885 ;
  assign y15022 = n32886 ;
  assign y15023 = n32890 ;
  assign y15024 = ~n32892 ;
  assign y15025 = ~1'b0 ;
  assign y15026 = n32894 ;
  assign y15027 = n32896 ;
  assign y15028 = n32897 ;
  assign y15029 = n32900 ;
  assign y15030 = n32901 ;
  assign y15031 = n32742 ;
  assign y15032 = ~n32907 ;
  assign y15033 = n32909 ;
  assign y15034 = n11275 ;
  assign y15035 = n32911 ;
  assign y15036 = ~1'b0 ;
  assign y15037 = ~1'b0 ;
  assign y15038 = ~n32913 ;
  assign y15039 = ~1'b0 ;
  assign y15040 = ~n32915 ;
  assign y15041 = n32916 ;
  assign y15042 = n32918 ;
  assign y15043 = ~1'b0 ;
  assign y15044 = ~n32920 ;
  assign y15045 = ~1'b0 ;
  assign y15046 = ~n11593 ;
  assign y15047 = ~1'b0 ;
  assign y15048 = ~n32928 ;
  assign y15049 = ~n32930 ;
  assign y15050 = ~n32931 ;
  assign y15051 = ~n32934 ;
  assign y15052 = n32935 ;
  assign y15053 = n32938 ;
  assign y15054 = ~1'b0 ;
  assign y15055 = n32940 ;
  assign y15056 = n32942 ;
  assign y15057 = n32944 ;
  assign y15058 = ~1'b0 ;
  assign y15059 = n2441 ;
  assign y15060 = ~n32947 ;
  assign y15061 = ~1'b0 ;
  assign y15062 = n32948 ;
  assign y15063 = ~1'b0 ;
  assign y15064 = ~n32950 ;
  assign y15065 = n32952 ;
  assign y15066 = ~1'b0 ;
  assign y15067 = ~n32954 ;
  assign y15068 = n32955 ;
  assign y15069 = ~1'b0 ;
  assign y15070 = ~1'b0 ;
  assign y15071 = ~n32963 ;
  assign y15072 = n32964 ;
  assign y15073 = ~n32965 ;
  assign y15074 = ~1'b0 ;
  assign y15075 = n32970 ;
  assign y15076 = ~n32972 ;
  assign y15077 = ~1'b0 ;
  assign y15078 = ~1'b0 ;
  assign y15079 = n32976 ;
  assign y15080 = n32982 ;
  assign y15081 = ~n32983 ;
  assign y15082 = ~n32986 ;
  assign y15083 = n32987 ;
  assign y15084 = n32989 ;
  assign y15085 = ~n32991 ;
  assign y15086 = n32992 ;
  assign y15087 = n32993 ;
  assign y15088 = n32994 ;
  assign y15089 = ~1'b0 ;
  assign y15090 = n32997 ;
  assign y15091 = n32998 ;
  assign y15092 = n32999 ;
  assign y15093 = ~n33002 ;
  assign y15094 = ~1'b0 ;
  assign y15095 = ~1'b0 ;
  assign y15096 = ~1'b0 ;
  assign y15097 = ~n33004 ;
  assign y15098 = ~n12986 ;
  assign y15099 = ~1'b0 ;
  assign y15100 = n33005 ;
  assign y15101 = ~n33010 ;
  assign y15102 = n33014 ;
  assign y15103 = n33017 ;
  assign y15104 = 1'b0 ;
  assign y15105 = ~1'b0 ;
  assign y15106 = n33019 ;
  assign y15107 = ~1'b0 ;
  assign y15108 = ~1'b0 ;
  assign y15109 = ~n33020 ;
  assign y15110 = ~n33021 ;
  assign y15111 = ~n33022 ;
  assign y15112 = ~1'b0 ;
  assign y15113 = n33024 ;
  assign y15114 = ~1'b0 ;
  assign y15115 = ~n33027 ;
  assign y15116 = ~n33031 ;
  assign y15117 = ~n33036 ;
  assign y15118 = ~1'b0 ;
  assign y15119 = ~1'b0 ;
  assign y15120 = n33037 ;
  assign y15121 = n17657 ;
  assign y15122 = n33042 ;
  assign y15123 = ~1'b0 ;
  assign y15124 = ~1'b0 ;
  assign y15125 = ~n33046 ;
  assign y15126 = n33047 ;
  assign y15127 = ~1'b0 ;
  assign y15128 = n33050 ;
  assign y15129 = n33052 ;
  assign y15130 = ~n33053 ;
  assign y15131 = n33060 ;
  assign y15132 = n33064 ;
  assign y15133 = ~1'b0 ;
  assign y15134 = n19224 ;
  assign y15135 = n33068 ;
  assign y15136 = n33069 ;
  assign y15137 = ~n33070 ;
  assign y15138 = ~1'b0 ;
  assign y15139 = ~n7785 ;
  assign y15140 = ~n33075 ;
  assign y15141 = n33077 ;
  assign y15142 = ~n33086 ;
  assign y15143 = n33088 ;
  assign y15144 = n16163 ;
  assign y15145 = n33089 ;
  assign y15146 = n33092 ;
  assign y15147 = ~n33094 ;
  assign y15148 = n33096 ;
  assign y15149 = 1'b0 ;
  assign y15150 = ~1'b0 ;
  assign y15151 = ~n9330 ;
  assign y15152 = ~n33098 ;
  assign y15153 = ~1'b0 ;
  assign y15154 = n33101 ;
  assign y15155 = ~1'b0 ;
  assign y15156 = ~1'b0 ;
  assign y15157 = n33102 ;
  assign y15158 = n33103 ;
  assign y15159 = n33104 ;
  assign y15160 = 1'b0 ;
  assign y15161 = n33112 ;
  assign y15162 = n33114 ;
  assign y15163 = ~n33118 ;
  assign y15164 = ~1'b0 ;
  assign y15165 = ~n33121 ;
  assign y15166 = ~1'b0 ;
  assign y15167 = 1'b0 ;
  assign y15168 = ~1'b0 ;
  assign y15169 = ~n33124 ;
  assign y15170 = ~n33125 ;
  assign y15171 = ~1'b0 ;
  assign y15172 = ~n33126 ;
  assign y15173 = n33128 ;
  assign y15174 = ~n33129 ;
  assign y15175 = n33130 ;
  assign y15176 = ~1'b0 ;
  assign y15177 = ~n10445 ;
  assign y15178 = n33135 ;
  assign y15179 = n33137 ;
  assign y15180 = n33139 ;
  assign y15181 = ~1'b0 ;
  assign y15182 = n33140 ;
  assign y15183 = ~n33146 ;
  assign y15184 = 1'b0 ;
  assign y15185 = n33150 ;
  assign y15186 = ~n33151 ;
  assign y15187 = ~1'b0 ;
  assign y15188 = ~1'b0 ;
  assign y15189 = ~n33152 ;
  assign y15190 = ~n33153 ;
  assign y15191 = n33154 ;
  assign y15192 = ~1'b0 ;
  assign y15193 = ~n33155 ;
  assign y15194 = ~n13048 ;
  assign y15195 = n33157 ;
  assign y15196 = ~1'b0 ;
  assign y15197 = ~1'b0 ;
  assign y15198 = ~n33160 ;
  assign y15199 = ~1'b0 ;
  assign y15200 = ~n9595 ;
  assign y15201 = n33166 ;
  assign y15202 = ~n33167 ;
  assign y15203 = n33171 ;
  assign y15204 = n33172 ;
  assign y15205 = n33174 ;
  assign y15206 = ~n1129 ;
  assign y15207 = ~1'b0 ;
  assign y15208 = ~n8623 ;
  assign y15209 = ~1'b0 ;
  assign y15210 = ~1'b0 ;
  assign y15211 = n33180 ;
  assign y15212 = ~n33185 ;
  assign y15213 = n33189 ;
  assign y15214 = ~1'b0 ;
  assign y15215 = ~n33191 ;
  assign y15216 = ~1'b0 ;
  assign y15217 = n33193 ;
  assign y15218 = ~n33195 ;
  assign y15219 = ~n33199 ;
  assign y15220 = ~n33204 ;
  assign y15221 = n33210 ;
  assign y15222 = n33211 ;
  assign y15223 = n33212 ;
  assign y15224 = n33216 ;
  assign y15225 = n33218 ;
  assign y15226 = ~n33219 ;
  assign y15227 = ~n33221 ;
  assign y15228 = ~1'b0 ;
  assign y15229 = ~n33225 ;
  assign y15230 = ~1'b0 ;
  assign y15231 = n33228 ;
  assign y15232 = ~n18711 ;
  assign y15233 = n33230 ;
  assign y15234 = ~1'b0 ;
  assign y15235 = ~n33232 ;
  assign y15236 = n33233 ;
  assign y15237 = ~n33237 ;
  assign y15238 = ~1'b0 ;
  assign y15239 = n33238 ;
  assign y15240 = n33241 ;
  assign y15241 = ~1'b0 ;
  assign y15242 = ~n33244 ;
  assign y15243 = ~1'b0 ;
  assign y15244 = ~n33261 ;
  assign y15245 = ~1'b0 ;
  assign y15246 = ~n33262 ;
  assign y15247 = ~n33265 ;
  assign y15248 = ~n33267 ;
  assign y15249 = n33271 ;
  assign y15250 = ~1'b0 ;
  assign y15251 = ~n33273 ;
  assign y15252 = n33275 ;
  assign y15253 = ~n33276 ;
  assign y15254 = n33277 ;
  assign y15255 = ~1'b0 ;
  assign y15256 = ~n33280 ;
  assign y15257 = ~n33284 ;
  assign y15258 = n33287 ;
  assign y15259 = ~1'b0 ;
  assign y15260 = ~1'b0 ;
  assign y15261 = n33293 ;
  assign y15262 = 1'b0 ;
  assign y15263 = n33294 ;
  assign y15264 = n33297 ;
  assign y15265 = ~n33298 ;
  assign y15266 = n33299 ;
  assign y15267 = ~1'b0 ;
  assign y15268 = n6232 ;
  assign y15269 = ~1'b0 ;
  assign y15270 = ~n33302 ;
  assign y15271 = n33303 ;
  assign y15272 = n33308 ;
  assign y15273 = n33309 ;
  assign y15274 = ~n33312 ;
  assign y15275 = n33314 ;
  assign y15276 = ~n33317 ;
  assign y15277 = ~1'b0 ;
  assign y15278 = n33320 ;
  assign y15279 = 1'b0 ;
  assign y15280 = n33324 ;
  assign y15281 = n33325 ;
  assign y15282 = ~n33327 ;
  assign y15283 = n33330 ;
  assign y15284 = n33333 ;
  assign y15285 = ~n5164 ;
  assign y15286 = ~1'b0 ;
  assign y15287 = ~n33338 ;
  assign y15288 = n33343 ;
  assign y15289 = ~1'b0 ;
  assign y15290 = ~1'b0 ;
  assign y15291 = ~1'b0 ;
  assign y15292 = ~n33352 ;
  assign y15293 = ~n33355 ;
  assign y15294 = ~n33363 ;
  assign y15295 = ~n33365 ;
  assign y15296 = ~1'b0 ;
  assign y15297 = ~1'b0 ;
  assign y15298 = ~n33369 ;
  assign y15299 = n33371 ;
  assign y15300 = ~1'b0 ;
  assign y15301 = ~1'b0 ;
  assign y15302 = ~1'b0 ;
  assign y15303 = ~1'b0 ;
  assign y15304 = ~n33378 ;
  assign y15305 = ~n33386 ;
  assign y15306 = ~n33388 ;
  assign y15307 = n33389 ;
  assign y15308 = n33394 ;
  assign y15309 = ~n33399 ;
  assign y15310 = ~n9338 ;
  assign y15311 = ~1'b0 ;
  assign y15312 = ~n33401 ;
  assign y15313 = n33402 ;
  assign y15314 = ~1'b0 ;
  assign y15315 = ~n33408 ;
  assign y15316 = n33411 ;
  assign y15317 = ~n33415 ;
  assign y15318 = ~1'b0 ;
  assign y15319 = ~n33419 ;
  assign y15320 = ~n33420 ;
  assign y15321 = n33421 ;
  assign y15322 = ~n15618 ;
  assign y15323 = n33433 ;
  assign y15324 = ~1'b0 ;
  assign y15325 = ~1'b0 ;
  assign y15326 = n33441 ;
  assign y15327 = n33445 ;
  assign y15328 = ~1'b0 ;
  assign y15329 = ~1'b0 ;
  assign y15330 = n33448 ;
  assign y15331 = n33450 ;
  assign y15332 = n33451 ;
  assign y15333 = ~n33453 ;
  assign y15334 = n33457 ;
  assign y15335 = n33459 ;
  assign y15336 = ~n23968 ;
  assign y15337 = ~n33461 ;
  assign y15338 = ~1'b0 ;
  assign y15339 = ~n33464 ;
  assign y15340 = ~n33466 ;
  assign y15341 = n33473 ;
  assign y15342 = ~n33475 ;
  assign y15343 = ~1'b0 ;
  assign y15344 = ~1'b0 ;
  assign y15345 = ~1'b0 ;
  assign y15346 = n33478 ;
  assign y15347 = ~1'b0 ;
  assign y15348 = ~n33482 ;
  assign y15349 = n33483 ;
  assign y15350 = ~n33486 ;
  assign y15351 = ~n33489 ;
  assign y15352 = ~1'b0 ;
  assign y15353 = ~1'b0 ;
  assign y15354 = ~n31742 ;
  assign y15355 = n33490 ;
  assign y15356 = n3253 ;
  assign y15357 = ~n33493 ;
  assign y15358 = n33494 ;
  assign y15359 = ~1'b0 ;
  assign y15360 = n33496 ;
  assign y15361 = ~1'b0 ;
  assign y15362 = ~1'b0 ;
  assign y15363 = n33497 ;
  assign y15364 = n33502 ;
  assign y15365 = ~n33504 ;
  assign y15366 = n33505 ;
  assign y15367 = ~1'b0 ;
  assign y15368 = ~n33508 ;
  assign y15369 = ~n33509 ;
  assign y15370 = n742 ;
  assign y15371 = ~n33510 ;
  assign y15372 = ~1'b0 ;
  assign y15373 = n33514 ;
  assign y15374 = ~n33516 ;
  assign y15375 = n33521 ;
  assign y15376 = ~1'b0 ;
  assign y15377 = ~1'b0 ;
  assign y15378 = ~1'b0 ;
  assign y15379 = ~n33525 ;
  assign y15380 = n33526 ;
  assign y15381 = n33528 ;
  assign y15382 = ~n33533 ;
  assign y15383 = ~n33537 ;
  assign y15384 = ~n33542 ;
  assign y15385 = ~n33547 ;
  assign y15386 = n33548 ;
  assign y15387 = ~n33550 ;
  assign y15388 = n33551 ;
  assign y15389 = ~1'b0 ;
  assign y15390 = ~1'b0 ;
  assign y15391 = ~n33552 ;
  assign y15392 = n23625 ;
  assign y15393 = n14949 ;
  assign y15394 = ~1'b0 ;
  assign y15395 = ~1'b0 ;
  assign y15396 = ~1'b0 ;
  assign y15397 = ~n33554 ;
  assign y15398 = ~n33555 ;
  assign y15399 = ~1'b0 ;
  assign y15400 = ~n33558 ;
  assign y15401 = n33562 ;
  assign y15402 = ~n33563 ;
  assign y15403 = ~n33569 ;
  assign y15404 = ~n10243 ;
  assign y15405 = n33573 ;
  assign y15406 = n33577 ;
  assign y15407 = ~1'b0 ;
  assign y15408 = ~n33582 ;
  assign y15409 = ~n33584 ;
  assign y15410 = ~n33585 ;
  assign y15411 = ~n33587 ;
  assign y15412 = ~1'b0 ;
  assign y15413 = n33589 ;
  assign y15414 = ~1'b0 ;
  assign y15415 = n33590 ;
  assign y15416 = ~n33592 ;
  assign y15417 = ~n33595 ;
  assign y15418 = ~1'b0 ;
  assign y15419 = n33599 ;
  assign y15420 = ~1'b0 ;
  assign y15421 = ~n33601 ;
  assign y15422 = ~n33603 ;
  assign y15423 = n33605 ;
  assign y15424 = ~n33606 ;
  assign y15425 = ~n33608 ;
  assign y15426 = ~n33611 ;
  assign y15427 = ~n33613 ;
  assign y15428 = ~n31983 ;
  assign y15429 = n33614 ;
  assign y15430 = ~n21491 ;
  assign y15431 = ~n14662 ;
  assign y15432 = ~n33615 ;
  assign y15433 = ~1'b0 ;
  assign y15434 = ~n33616 ;
  assign y15435 = n33617 ;
  assign y15436 = n33620 ;
  assign y15437 = ~n33625 ;
  assign y15438 = ~1'b0 ;
  assign y15439 = ~n33629 ;
  assign y15440 = ~1'b0 ;
  assign y15441 = ~1'b0 ;
  assign y15442 = ~1'b0 ;
  assign y15443 = ~1'b0 ;
  assign y15444 = n33631 ;
  assign y15445 = n33632 ;
  assign y15446 = ~n33634 ;
  assign y15447 = n33635 ;
  assign y15448 = n33640 ;
  assign y15449 = ~n33644 ;
  assign y15450 = n33647 ;
  assign y15451 = ~1'b0 ;
  assign y15452 = n33655 ;
  assign y15453 = ~1'b0 ;
  assign y15454 = ~1'b0 ;
  assign y15455 = n33658 ;
  assign y15456 = ~n33662 ;
  assign y15457 = n33664 ;
  assign y15458 = ~1'b0 ;
  assign y15459 = ~1'b0 ;
  assign y15460 = n33665 ;
  assign y15461 = ~n33673 ;
  assign y15462 = ~n33674 ;
  assign y15463 = 1'b0 ;
  assign y15464 = ~n33676 ;
  assign y15465 = ~n33682 ;
  assign y15466 = n33684 ;
  assign y15467 = ~1'b0 ;
  assign y15468 = ~n33687 ;
  assign y15469 = n33691 ;
  assign y15470 = n12169 ;
  assign y15471 = ~1'b0 ;
  assign y15472 = ~n33693 ;
  assign y15473 = n33702 ;
  assign y15474 = ~1'b0 ;
  assign y15475 = ~n33707 ;
  assign y15476 = ~n33713 ;
  assign y15477 = ~n33714 ;
  assign y15478 = ~1'b0 ;
  assign y15479 = ~1'b0 ;
  assign y15480 = ~1'b0 ;
  assign y15481 = ~n17571 ;
  assign y15482 = n33717 ;
  assign y15483 = n33718 ;
  assign y15484 = ~n33725 ;
  assign y15485 = ~n33726 ;
  assign y15486 = ~n33729 ;
  assign y15487 = ~n33730 ;
  assign y15488 = ~n33734 ;
  assign y15489 = n33742 ;
  assign y15490 = n33745 ;
  assign y15491 = n33749 ;
  assign y15492 = n33753 ;
  assign y15493 = ~n33755 ;
  assign y15494 = n33758 ;
  assign y15495 = n33759 ;
  assign y15496 = n33760 ;
  assign y15497 = ~n33763 ;
  assign y15498 = ~n33764 ;
  assign y15499 = ~1'b0 ;
  assign y15500 = ~n33766 ;
  assign y15501 = ~n33767 ;
  assign y15502 = ~1'b0 ;
  assign y15503 = n33770 ;
  assign y15504 = n33774 ;
  assign y15505 = n33779 ;
  assign y15506 = ~n33781 ;
  assign y15507 = n33783 ;
  assign y15508 = n33784 ;
  assign y15509 = ~n33787 ;
  assign y15510 = ~n33790 ;
  assign y15511 = n33791 ;
  assign y15512 = ~n33792 ;
  assign y15513 = ~1'b0 ;
  assign y15514 = ~n33793 ;
  assign y15515 = ~n33795 ;
  assign y15516 = ~1'b0 ;
  assign y15517 = ~1'b0 ;
  assign y15518 = ~1'b0 ;
  assign y15519 = ~n33800 ;
  assign y15520 = n33810 ;
  assign y15521 = ~1'b0 ;
  assign y15522 = ~n33812 ;
  assign y15523 = ~n33813 ;
  assign y15524 = ~n33814 ;
  assign y15525 = ~n33815 ;
  assign y15526 = n33818 ;
  assign y15527 = ~n33819 ;
  assign y15528 = ~1'b0 ;
  assign y15529 = ~n33822 ;
  assign y15530 = ~1'b0 ;
  assign y15531 = ~n33824 ;
  assign y15532 = n33825 ;
  assign y15533 = ~n33829 ;
  assign y15534 = n33831 ;
  assign y15535 = n33834 ;
  assign y15536 = n3554 ;
  assign y15537 = ~n33836 ;
  assign y15538 = n33838 ;
  assign y15539 = ~n33842 ;
  assign y15540 = ~1'b0 ;
  assign y15541 = 1'b0 ;
  assign y15542 = n33843 ;
  assign y15543 = n33844 ;
  assign y15544 = n33847 ;
  assign y15545 = n33852 ;
  assign y15546 = ~n33857 ;
  assign y15547 = ~n33859 ;
  assign y15548 = n33860 ;
  assign y15549 = 1'b0 ;
  assign y15550 = ~n18367 ;
  assign y15551 = ~n33862 ;
  assign y15552 = n33864 ;
  assign y15553 = 1'b0 ;
  assign y15554 = ~n33872 ;
  assign y15555 = ~n33873 ;
  assign y15556 = ~n33876 ;
  assign y15557 = n33877 ;
  assign y15558 = ~n33880 ;
  assign y15559 = ~n33884 ;
  assign y15560 = ~n33885 ;
  assign y15561 = ~1'b0 ;
  assign y15562 = ~1'b0 ;
  assign y15563 = ~n33892 ;
  assign y15564 = ~n33896 ;
  assign y15565 = ~1'b0 ;
  assign y15566 = ~n33897 ;
  assign y15567 = n33901 ;
  assign y15568 = ~n33905 ;
  assign y15569 = ~1'b0 ;
  assign y15570 = ~n31817 ;
  assign y15571 = n9267 ;
  assign y15572 = ~n33906 ;
  assign y15573 = ~n33908 ;
  assign y15574 = ~n33909 ;
  assign y15575 = ~n33910 ;
  assign y15576 = ~1'b0 ;
  assign y15577 = ~1'b0 ;
  assign y15578 = ~1'b0 ;
  assign y15579 = ~n33928 ;
  assign y15580 = ~n33931 ;
  assign y15581 = ~1'b0 ;
  assign y15582 = ~1'b0 ;
  assign y15583 = n33935 ;
  assign y15584 = ~n33941 ;
  assign y15585 = n33944 ;
  assign y15586 = n33946 ;
  assign y15587 = ~1'b0 ;
  assign y15588 = n33950 ;
  assign y15589 = ~1'b0 ;
  assign y15590 = n33955 ;
  assign y15591 = ~n33956 ;
  assign y15592 = ~n2757 ;
  assign y15593 = n33960 ;
  assign y15594 = ~n33961 ;
  assign y15595 = ~n33962 ;
  assign y15596 = n33967 ;
  assign y15597 = n33969 ;
  assign y15598 = n33973 ;
  assign y15599 = ~1'b0 ;
  assign y15600 = n33976 ;
  assign y15601 = ~n33982 ;
  assign y15602 = ~n33985 ;
  assign y15603 = ~1'b0 ;
  assign y15604 = n33987 ;
  assign y15605 = n33990 ;
  assign y15606 = n33993 ;
  assign y15607 = n33994 ;
  assign y15608 = n33996 ;
  assign y15609 = n33998 ;
  assign y15610 = n33999 ;
  assign y15611 = n34003 ;
  assign y15612 = ~n34004 ;
  assign y15613 = ~1'b0 ;
  assign y15614 = n34005 ;
  assign y15615 = n34006 ;
  assign y15616 = ~n34008 ;
  assign y15617 = ~n34010 ;
  assign y15618 = n34012 ;
  assign y15619 = n34013 ;
  assign y15620 = ~n34021 ;
  assign y15621 = ~n15734 ;
  assign y15622 = n34025 ;
  assign y15623 = ~n9331 ;
  assign y15624 = ~1'b0 ;
  assign y15625 = ~n34027 ;
  assign y15626 = n34029 ;
  assign y15627 = ~n34043 ;
  assign y15628 = ~1'b0 ;
  assign y15629 = n34048 ;
  assign y15630 = ~n34049 ;
  assign y15631 = n34053 ;
  assign y15632 = n34057 ;
  assign y15633 = ~n6196 ;
  assign y15634 = n34058 ;
  assign y15635 = n34060 ;
  assign y15636 = ~1'b0 ;
  assign y15637 = ~n32782 ;
  assign y15638 = ~n34064 ;
  assign y15639 = ~n34065 ;
  assign y15640 = n34067 ;
  assign y15641 = ~n34070 ;
  assign y15642 = ~n34071 ;
  assign y15643 = n34074 ;
  assign y15644 = ~1'b0 ;
  assign y15645 = ~n34076 ;
  assign y15646 = n34078 ;
  assign y15647 = ~n34082 ;
  assign y15648 = 1'b0 ;
  assign y15649 = n34086 ;
  assign y15650 = n34091 ;
  assign y15651 = ~n6390 ;
  assign y15652 = n34094 ;
  assign y15653 = ~1'b0 ;
  assign y15654 = ~n34096 ;
  assign y15655 = ~n34105 ;
  assign y15656 = ~n34108 ;
  assign y15657 = ~n34112 ;
  assign y15658 = n34115 ;
  assign y15659 = ~n19957 ;
  assign y15660 = ~1'b0 ;
  assign y15661 = ~1'b0 ;
  assign y15662 = n34116 ;
  assign y15663 = ~1'b0 ;
  assign y15664 = ~1'b0 ;
  assign y15665 = ~1'b0 ;
  assign y15666 = n34118 ;
  assign y15667 = n34120 ;
  assign y15668 = n34122 ;
  assign y15669 = ~1'b0 ;
  assign y15670 = ~1'b0 ;
  assign y15671 = n34123 ;
  assign y15672 = n34124 ;
  assign y15673 = ~1'b0 ;
  assign y15674 = n34125 ;
  assign y15675 = ~x206 ;
  assign y15676 = ~1'b0 ;
  assign y15677 = ~1'b0 ;
  assign y15678 = ~n34126 ;
  assign y15679 = n34134 ;
  assign y15680 = ~n34139 ;
  assign y15681 = ~n34140 ;
  assign y15682 = n34144 ;
  assign y15683 = ~n34146 ;
  assign y15684 = ~1'b0 ;
  assign y15685 = n34148 ;
  assign y15686 = ~1'b0 ;
  assign y15687 = n34153 ;
  assign y15688 = n34155 ;
  assign y15689 = ~n34158 ;
  assign y15690 = n34160 ;
  assign y15691 = ~n34194 ;
  assign y15692 = ~n34199 ;
  assign y15693 = n34203 ;
  assign y15694 = 1'b0 ;
  assign y15695 = n34205 ;
  assign y15696 = n34208 ;
  assign y15697 = ~1'b0 ;
  assign y15698 = n824 ;
  assign y15699 = ~n34209 ;
  assign y15700 = n34210 ;
  assign y15701 = n34216 ;
  assign y15702 = n3316 ;
  assign y15703 = n34219 ;
  assign y15704 = ~n34221 ;
  assign y15705 = n34222 ;
  assign y15706 = 1'b0 ;
  assign y15707 = ~n12172 ;
  assign y15708 = n34224 ;
  assign y15709 = ~n34226 ;
  assign y15710 = n34229 ;
  assign y15711 = ~1'b0 ;
  assign y15712 = ~1'b0 ;
  assign y15713 = n34230 ;
  assign y15714 = ~n34233 ;
  assign y15715 = n34234 ;
  assign y15716 = ~n34235 ;
  assign y15717 = n34237 ;
  assign y15718 = ~n34239 ;
  assign y15719 = n34246 ;
  assign y15720 = ~n34254 ;
  assign y15721 = n34256 ;
  assign y15722 = ~n34259 ;
  assign y15723 = n34265 ;
  assign y15724 = n34267 ;
  assign y15725 = ~n34268 ;
  assign y15726 = ~n34271 ;
  assign y15727 = ~n34274 ;
  assign y15728 = ~n34275 ;
  assign y15729 = ~1'b0 ;
  assign y15730 = n34277 ;
  assign y15731 = ~n34278 ;
  assign y15732 = ~n34281 ;
  assign y15733 = n34282 ;
  assign y15734 = 1'b0 ;
  assign y15735 = ~n34285 ;
  assign y15736 = ~n34288 ;
  assign y15737 = ~n34293 ;
  assign y15738 = n34297 ;
  assign y15739 = n34298 ;
  assign y15740 = n34299 ;
  assign y15741 = ~1'b0 ;
  assign y15742 = n34304 ;
  assign y15743 = n34305 ;
  assign y15744 = ~n34307 ;
  assign y15745 = ~1'b0 ;
  assign y15746 = ~n1239 ;
  assign y15747 = n34308 ;
  assign y15748 = ~n34309 ;
  assign y15749 = ~1'b0 ;
  assign y15750 = ~n34315 ;
  assign y15751 = ~n34317 ;
  assign y15752 = ~n34318 ;
  assign y15753 = ~1'b0 ;
  assign y15754 = n34321 ;
  assign y15755 = n34323 ;
  assign y15756 = ~n34324 ;
  assign y15757 = ~n34326 ;
  assign y15758 = ~1'b0 ;
  assign y15759 = n34327 ;
  assign y15760 = n34332 ;
  assign y15761 = ~n34334 ;
  assign y15762 = ~1'b0 ;
  assign y15763 = n34336 ;
  assign y15764 = n25464 ;
  assign y15765 = ~1'b0 ;
  assign y15766 = n34339 ;
  assign y15767 = ~n34341 ;
  assign y15768 = ~1'b0 ;
  assign y15769 = n34344 ;
  assign y15770 = n34346 ;
  assign y15771 = ~n34351 ;
  assign y15772 = ~n34360 ;
  assign y15773 = n34368 ;
  assign y15774 = ~1'b0 ;
  assign y15775 = ~1'b0 ;
  assign y15776 = ~n34372 ;
  assign y15777 = ~1'b0 ;
  assign y15778 = n34374 ;
  assign y15779 = ~n34376 ;
  assign y15780 = n28231 ;
  assign y15781 = n34378 ;
  assign y15782 = n34380 ;
  assign y15783 = ~n34382 ;
  assign y15784 = ~1'b0 ;
  assign y15785 = ~n34386 ;
  assign y15786 = ~n34388 ;
  assign y15787 = ~n34390 ;
  assign y15788 = ~1'b0 ;
  assign y15789 = ~n34392 ;
  assign y15790 = ~1'b0 ;
  assign y15791 = ~n34396 ;
  assign y15792 = ~1'b0 ;
  assign y15793 = n34399 ;
  assign y15794 = ~n34401 ;
  assign y15795 = n34402 ;
  assign y15796 = ~n34405 ;
  assign y15797 = ~1'b0 ;
  assign y15798 = ~n34407 ;
  assign y15799 = ~1'b0 ;
  assign y15800 = n34409 ;
  assign y15801 = ~1'b0 ;
  assign y15802 = ~n34412 ;
  assign y15803 = ~n34413 ;
  assign y15804 = n20010 ;
  assign y15805 = ~n34415 ;
  assign y15806 = n34416 ;
  assign y15807 = n34417 ;
  assign y15808 = n34418 ;
  assign y15809 = ~1'b0 ;
  assign y15810 = ~1'b0 ;
  assign y15811 = ~1'b0 ;
  assign y15812 = ~n34423 ;
  assign y15813 = ~n34424 ;
  assign y15814 = ~n34425 ;
  assign y15815 = n34427 ;
  assign y15816 = n34430 ;
  assign y15817 = ~n34432 ;
  assign y15818 = n34433 ;
  assign y15819 = n34434 ;
  assign y15820 = ~1'b0 ;
  assign y15821 = n34436 ;
  assign y15822 = n34442 ;
  assign y15823 = ~1'b0 ;
  assign y15824 = ~n34446 ;
  assign y15825 = n34448 ;
  assign y15826 = ~1'b0 ;
  assign y15827 = ~n34450 ;
  assign y15828 = n34455 ;
  assign y15829 = ~n34458 ;
  assign y15830 = ~n34460 ;
  assign y15831 = ~n6408 ;
  assign y15832 = ~n34461 ;
  assign y15833 = ~n34462 ;
  assign y15834 = ~n34464 ;
  assign y15835 = ~1'b0 ;
  assign y15836 = ~n34465 ;
  assign y15837 = ~n34468 ;
  assign y15838 = ~n34470 ;
  assign y15839 = n34475 ;
  assign y15840 = n17861 ;
  assign y15841 = n34477 ;
  assign y15842 = ~n34479 ;
  assign y15843 = ~1'b0 ;
  assign y15844 = ~n34480 ;
  assign y15845 = ~1'b0 ;
  assign y15846 = ~n34484 ;
  assign y15847 = ~n34486 ;
  assign y15848 = n14262 ;
  assign y15849 = n34488 ;
  assign y15850 = ~1'b0 ;
  assign y15851 = n34489 ;
  assign y15852 = n34490 ;
  assign y15853 = n34493 ;
  assign y15854 = ~1'b0 ;
  assign y15855 = ~n34496 ;
  assign y15856 = n34499 ;
  assign y15857 = n34501 ;
  assign y15858 = ~n34507 ;
  assign y15859 = n34508 ;
  assign y15860 = n3308 ;
  assign y15861 = ~n34510 ;
  assign y15862 = ~n34513 ;
  assign y15863 = ~n34516 ;
  assign y15864 = ~n34518 ;
  assign y15865 = n29188 ;
  assign y15866 = ~1'b0 ;
  assign y15867 = ~1'b0 ;
  assign y15868 = ~1'b0 ;
  assign y15869 = n34523 ;
  assign y15870 = ~n34528 ;
  assign y15871 = n34530 ;
  assign y15872 = ~1'b0 ;
  assign y15873 = ~1'b0 ;
  assign y15874 = ~1'b0 ;
  assign y15875 = ~1'b0 ;
  assign y15876 = ~n34532 ;
  assign y15877 = n34533 ;
  assign y15878 = n34534 ;
  assign y15879 = ~1'b0 ;
  assign y15880 = ~n34535 ;
  assign y15881 = ~n34537 ;
  assign y15882 = ~n34543 ;
  assign y15883 = ~1'b0 ;
  assign y15884 = n34547 ;
  assign y15885 = n34548 ;
  assign y15886 = n34555 ;
  assign y15887 = ~1'b0 ;
  assign y15888 = n34558 ;
  assign y15889 = n34559 ;
  assign y15890 = ~1'b0 ;
  assign y15891 = n34565 ;
  assign y15892 = ~1'b0 ;
  assign y15893 = n34567 ;
  assign y15894 = ~n34568 ;
  assign y15895 = n34569 ;
  assign y15896 = ~1'b0 ;
  assign y15897 = ~n34570 ;
  assign y15898 = ~n34573 ;
  assign y15899 = ~1'b0 ;
  assign y15900 = ~n34576 ;
  assign y15901 = n34581 ;
  assign y15902 = n34583 ;
  assign y15903 = ~n34587 ;
  assign y15904 = ~n34590 ;
  assign y15905 = ~1'b0 ;
  assign y15906 = ~1'b0 ;
  assign y15907 = ~n34593 ;
  assign y15908 = ~n34595 ;
  assign y15909 = n34597 ;
  assign y15910 = n34599 ;
  assign y15911 = n18070 ;
  assign y15912 = ~1'b0 ;
  assign y15913 = ~n34602 ;
  assign y15914 = n34604 ;
  assign y15915 = ~n34606 ;
  assign y15916 = ~n34611 ;
  assign y15917 = n34612 ;
  assign y15918 = ~1'b0 ;
  assign y15919 = ~n34616 ;
  assign y15920 = ~n4294 ;
  assign y15921 = ~n34618 ;
  assign y15922 = n34620 ;
  assign y15923 = n34622 ;
  assign y15924 = ~1'b0 ;
  assign y15925 = n34624 ;
  assign y15926 = n34625 ;
  assign y15927 = n34626 ;
  assign y15928 = n34627 ;
  assign y15929 = ~n34629 ;
  assign y15930 = ~1'b0 ;
  assign y15931 = n34633 ;
  assign y15932 = n34636 ;
  assign y15933 = n34637 ;
  assign y15934 = n34638 ;
  assign y15935 = ~n34641 ;
  assign y15936 = ~1'b0 ;
  assign y15937 = ~n30229 ;
  assign y15938 = ~1'b0 ;
  assign y15939 = ~1'b0 ;
  assign y15940 = ~n34643 ;
  assign y15941 = ~1'b0 ;
  assign y15942 = n34647 ;
  assign y15943 = ~1'b0 ;
  assign y15944 = ~1'b0 ;
  assign y15945 = n34652 ;
  assign y15946 = ~1'b0 ;
  assign y15947 = ~n34658 ;
  assign y15948 = ~n34661 ;
  assign y15949 = n34662 ;
  assign y15950 = ~1'b0 ;
  assign y15951 = n34666 ;
  assign y15952 = 1'b0 ;
  assign y15953 = n34669 ;
  assign y15954 = ~1'b0 ;
  assign y15955 = ~1'b0 ;
  assign y15956 = n34671 ;
  assign y15957 = n34672 ;
  assign y15958 = n34676 ;
  assign y15959 = ~1'b0 ;
  assign y15960 = ~1'b0 ;
  assign y15961 = ~1'b0 ;
  assign y15962 = ~1'b0 ;
  assign y15963 = ~1'b0 ;
  assign y15964 = ~1'b0 ;
  assign y15965 = n34685 ;
  assign y15966 = ~n34687 ;
  assign y15967 = ~n34689 ;
  assign y15968 = ~n34690 ;
  assign y15969 = n34699 ;
  assign y15970 = ~1'b0 ;
  assign y15971 = ~1'b0 ;
  assign y15972 = n34700 ;
  assign y15973 = ~n34705 ;
  assign y15974 = ~n34708 ;
  assign y15975 = n34710 ;
  assign y15976 = ~n34714 ;
  assign y15977 = ~1'b0 ;
  assign y15978 = n34715 ;
  assign y15979 = ~n34716 ;
  assign y15980 = ~n34722 ;
  assign y15981 = ~1'b0 ;
  assign y15982 = ~1'b0 ;
  assign y15983 = ~n34724 ;
  assign y15984 = n34729 ;
  assign y15985 = ~n6611 ;
  assign y15986 = ~n34730 ;
  assign y15987 = ~1'b0 ;
  assign y15988 = ~n34732 ;
  assign y15989 = n34739 ;
  assign y15990 = n34740 ;
  assign y15991 = n34743 ;
  assign y15992 = ~n34744 ;
  assign y15993 = ~n34748 ;
  assign y15994 = ~n34755 ;
  assign y15995 = n34759 ;
  assign y15996 = ~1'b0 ;
  assign y15997 = ~n34768 ;
  assign y15998 = ~1'b0 ;
  assign y15999 = ~1'b0 ;
  assign y16000 = ~n34769 ;
  assign y16001 = n34771 ;
  assign y16002 = ~n34772 ;
  assign y16003 = n34775 ;
  assign y16004 = ~1'b0 ;
  assign y16005 = n34776 ;
  assign y16006 = n34777 ;
  assign y16007 = n34778 ;
  assign y16008 = ~n34780 ;
  assign y16009 = n34781 ;
  assign y16010 = n34782 ;
  assign y16011 = n16825 ;
  assign y16012 = n34783 ;
  assign y16013 = n34785 ;
  assign y16014 = ~n34787 ;
  assign y16015 = ~n34791 ;
  assign y16016 = ~1'b0 ;
  assign y16017 = n8750 ;
  assign y16018 = ~1'b0 ;
  assign y16019 = n34795 ;
  assign y16020 = ~n34800 ;
  assign y16021 = n34804 ;
  assign y16022 = n34808 ;
  assign y16023 = n34810 ;
  assign y16024 = ~n34813 ;
  assign y16025 = ~n34814 ;
  assign y16026 = ~n34816 ;
  assign y16027 = ~n34821 ;
  assign y16028 = n34823 ;
  assign y16029 = ~n21526 ;
  assign y16030 = ~1'b0 ;
  assign y16031 = n34828 ;
  assign y16032 = n34829 ;
  assign y16033 = n34832 ;
  assign y16034 = n34835 ;
  assign y16035 = ~1'b0 ;
  assign y16036 = ~1'b0 ;
  assign y16037 = ~n34837 ;
  assign y16038 = n34839 ;
  assign y16039 = n34840 ;
  assign y16040 = ~1'b0 ;
  assign y16041 = n34842 ;
  assign y16042 = ~1'b0 ;
  assign y16043 = n34846 ;
  assign y16044 = ~n34853 ;
  assign y16045 = 1'b0 ;
  assign y16046 = ~1'b0 ;
  assign y16047 = n34855 ;
  assign y16048 = ~n34858 ;
  assign y16049 = n34859 ;
  assign y16050 = ~n34861 ;
  assign y16051 = ~1'b0 ;
  assign y16052 = ~1'b0 ;
  assign y16053 = ~n8634 ;
  assign y16054 = ~n34862 ;
  assign y16055 = ~1'b0 ;
  assign y16056 = ~1'b0 ;
  assign y16057 = ~n34864 ;
  assign y16058 = n34865 ;
  assign y16059 = ~n34868 ;
  assign y16060 = ~1'b0 ;
  assign y16061 = ~n34875 ;
  assign y16062 = ~1'b0 ;
  assign y16063 = ~1'b0 ;
  assign y16064 = ~n34879 ;
  assign y16065 = ~n34883 ;
  assign y16066 = n34884 ;
  assign y16067 = ~n30931 ;
  assign y16068 = n34888 ;
  assign y16069 = ~1'b0 ;
  assign y16070 = ~n34890 ;
  assign y16071 = n34896 ;
  assign y16072 = ~1'b0 ;
  assign y16073 = ~1'b0 ;
  assign y16074 = ~1'b0 ;
  assign y16075 = n34900 ;
  assign y16076 = ~n34902 ;
  assign y16077 = n34905 ;
  assign y16078 = n34906 ;
  assign y16079 = ~n34909 ;
  assign y16080 = ~1'b0 ;
  assign y16081 = n34910 ;
  assign y16082 = ~n34912 ;
  assign y16083 = ~n34914 ;
  assign y16084 = n34915 ;
  assign y16085 = n34916 ;
  assign y16086 = ~n34919 ;
  assign y16087 = 1'b0 ;
  assign y16088 = n34920 ;
  assign y16089 = ~1'b0 ;
  assign y16090 = 1'b0 ;
  assign y16091 = ~n34921 ;
  assign y16092 = ~n34922 ;
  assign y16093 = ~1'b0 ;
  assign y16094 = ~1'b0 ;
  assign y16095 = n34924 ;
  assign y16096 = n34925 ;
  assign y16097 = ~1'b0 ;
  assign y16098 = n34931 ;
  assign y16099 = ~n34932 ;
  assign y16100 = n34942 ;
  assign y16101 = 1'b0 ;
  assign y16102 = ~n34943 ;
  assign y16103 = ~1'b0 ;
  assign y16104 = ~1'b0 ;
  assign y16105 = n34946 ;
  assign y16106 = ~n34947 ;
  assign y16107 = ~1'b0 ;
  assign y16108 = ~1'b0 ;
  assign y16109 = ~1'b0 ;
  assign y16110 = n34948 ;
  assign y16111 = ~n34949 ;
  assign y16112 = ~1'b0 ;
  assign y16113 = n34953 ;
  assign y16114 = ~1'b0 ;
  assign y16115 = n34958 ;
  assign y16116 = ~n34959 ;
  assign y16117 = ~n34960 ;
  assign y16118 = ~n34961 ;
  assign y16119 = n12665 ;
  assign y16120 = ~n34963 ;
  assign y16121 = ~n22999 ;
  assign y16122 = ~1'b0 ;
  assign y16123 = n34966 ;
  assign y16124 = n34968 ;
  assign y16125 = n34969 ;
  assign y16126 = ~n34974 ;
  assign y16127 = n34975 ;
  assign y16128 = n34978 ;
  assign y16129 = ~n34985 ;
  assign y16130 = ~1'b0 ;
  assign y16131 = n12687 ;
  assign y16132 = ~x210 ;
  assign y16133 = ~1'b0 ;
  assign y16134 = ~n34987 ;
  assign y16135 = n34989 ;
  assign y16136 = ~n34991 ;
  assign y16137 = ~1'b0 ;
  assign y16138 = ~n34993 ;
  assign y16139 = n34998 ;
  assign y16140 = ~1'b0 ;
  assign y16141 = n34999 ;
  assign y16142 = n35001 ;
  assign y16143 = ~n35008 ;
  assign y16144 = ~n35011 ;
  assign y16145 = ~n35012 ;
  assign y16146 = ~n35014 ;
  assign y16147 = ~1'b0 ;
  assign y16148 = ~1'b0 ;
  assign y16149 = ~n35015 ;
  assign y16150 = n35018 ;
  assign y16151 = n35023 ;
  assign y16152 = n35027 ;
  assign y16153 = n35029 ;
  assign y16154 = n35031 ;
  assign y16155 = 1'b0 ;
  assign y16156 = ~n35035 ;
  assign y16157 = ~n35036 ;
  assign y16158 = ~1'b0 ;
  assign y16159 = n35037 ;
  assign y16160 = n35039 ;
  assign y16161 = n35040 ;
  assign y16162 = n35041 ;
  assign y16163 = ~1'b0 ;
  assign y16164 = ~1'b0 ;
  assign y16165 = ~n35044 ;
  assign y16166 = n35045 ;
  assign y16167 = ~n35047 ;
  assign y16168 = ~1'b0 ;
  assign y16169 = n35049 ;
  assign y16170 = n35052 ;
  assign y16171 = ~n35054 ;
  assign y16172 = n35056 ;
  assign y16173 = ~n35065 ;
  assign y16174 = n35067 ;
  assign y16175 = ~n35070 ;
  assign y16176 = n35073 ;
  assign y16177 = n35074 ;
  assign y16178 = ~1'b0 ;
  assign y16179 = n35075 ;
  assign y16180 = n35078 ;
  assign y16181 = n35079 ;
  assign y16182 = ~n35082 ;
  assign y16183 = ~1'b0 ;
  assign y16184 = n35088 ;
  assign y16185 = ~n35093 ;
  assign y16186 = n35095 ;
  assign y16187 = ~n35098 ;
  assign y16188 = n35100 ;
  assign y16189 = n35101 ;
  assign y16190 = ~n35107 ;
  assign y16191 = n35109 ;
  assign y16192 = ~n35115 ;
  assign y16193 = ~n35116 ;
  assign y16194 = ~n35120 ;
  assign y16195 = ~1'b0 ;
  assign y16196 = n35123 ;
  assign y16197 = 1'b0 ;
  assign y16198 = n35124 ;
  assign y16199 = ~n35125 ;
  assign y16200 = n35127 ;
  assign y16201 = ~1'b0 ;
  assign y16202 = ~n35129 ;
  assign y16203 = ~1'b0 ;
  assign y16204 = ~n12576 ;
  assign y16205 = ~1'b0 ;
  assign y16206 = n35131 ;
  assign y16207 = ~n35134 ;
  assign y16208 = ~1'b0 ;
  assign y16209 = n35135 ;
  assign y16210 = ~n24559 ;
  assign y16211 = n35141 ;
  assign y16212 = ~1'b0 ;
  assign y16213 = n35142 ;
  assign y16214 = ~n35144 ;
  assign y16215 = n35145 ;
  assign y16216 = n35146 ;
  assign y16217 = n35147 ;
  assign y16218 = ~n35148 ;
  assign y16219 = n35152 ;
  assign y16220 = ~1'b0 ;
  assign y16221 = n10175 ;
  assign y16222 = ~1'b0 ;
  assign y16223 = ~1'b0 ;
  assign y16224 = ~n35158 ;
  assign y16225 = ~n35171 ;
  assign y16226 = ~n25552 ;
  assign y16227 = ~1'b0 ;
  assign y16228 = n35187 ;
  assign y16229 = n35189 ;
  assign y16230 = n35193 ;
  assign y16231 = n35196 ;
  assign y16232 = n35197 ;
  assign y16233 = ~1'b0 ;
  assign y16234 = n35198 ;
  assign y16235 = ~n35204 ;
  assign y16236 = ~1'b0 ;
  assign y16237 = ~1'b0 ;
  assign y16238 = n25343 ;
  assign y16239 = ~n35205 ;
  assign y16240 = ~n35207 ;
  assign y16241 = n35208 ;
  assign y16242 = n35215 ;
  assign y16243 = ~1'b0 ;
  assign y16244 = n35224 ;
  assign y16245 = ~1'b0 ;
  assign y16246 = n35229 ;
  assign y16247 = n35232 ;
  assign y16248 = n35234 ;
  assign y16249 = n35236 ;
  assign y16250 = ~n35239 ;
  assign y16251 = n35240 ;
  assign y16252 = ~1'b0 ;
  assign y16253 = ~1'b0 ;
  assign y16254 = n35242 ;
  assign y16255 = n35243 ;
  assign y16256 = ~n35245 ;
  assign y16257 = ~n35246 ;
  assign y16258 = n35248 ;
  assign y16259 = n35258 ;
  assign y16260 = ~n35260 ;
  assign y16261 = n35261 ;
  assign y16262 = ~n35262 ;
  assign y16263 = n33370 ;
  assign y16264 = n35263 ;
  assign y16265 = ~n35266 ;
  assign y16266 = n35267 ;
  assign y16267 = ~1'b0 ;
  assign y16268 = ~1'b0 ;
  assign y16269 = ~1'b0 ;
  assign y16270 = n35269 ;
  assign y16271 = ~n35272 ;
  assign y16272 = n35279 ;
  assign y16273 = ~1'b0 ;
  assign y16274 = ~n35281 ;
  assign y16275 = ~1'b0 ;
  assign y16276 = ~n35282 ;
  assign y16277 = ~n35290 ;
  assign y16278 = n35291 ;
  assign y16279 = ~n35293 ;
  assign y16280 = ~1'b0 ;
  assign y16281 = ~n35297 ;
  assign y16282 = ~n35298 ;
  assign y16283 = ~n35299 ;
  assign y16284 = ~n35303 ;
  assign y16285 = ~n15239 ;
  assign y16286 = ~n35307 ;
  assign y16287 = ~n35308 ;
  assign y16288 = 1'b0 ;
  assign y16289 = ~1'b0 ;
  assign y16290 = ~n35310 ;
  assign y16291 = ~n35313 ;
  assign y16292 = ~n7481 ;
  assign y16293 = ~n35315 ;
  assign y16294 = ~n35317 ;
  assign y16295 = ~1'b0 ;
  assign y16296 = ~n35319 ;
  assign y16297 = ~n35322 ;
  assign y16298 = ~n35327 ;
  assign y16299 = ~1'b0 ;
  assign y16300 = ~n35329 ;
  assign y16301 = n35334 ;
  assign y16302 = ~1'b0 ;
  assign y16303 = n18842 ;
  assign y16304 = ~n35335 ;
  assign y16305 = ~n35336 ;
  assign y16306 = ~n35338 ;
  assign y16307 = n35340 ;
  assign y16308 = ~n35342 ;
  assign y16309 = ~1'b0 ;
  assign y16310 = ~1'b0 ;
  assign y16311 = ~n35348 ;
  assign y16312 = ~n19695 ;
  assign y16313 = n35349 ;
  assign y16314 = n35352 ;
  assign y16315 = n35353 ;
  assign y16316 = ~n35354 ;
  assign y16317 = ~1'b0 ;
  assign y16318 = ~n35356 ;
  assign y16319 = ~1'b0 ;
  assign y16320 = ~n35358 ;
  assign y16321 = ~n35361 ;
  assign y16322 = ~n35362 ;
  assign y16323 = ~n35365 ;
  assign y16324 = ~1'b0 ;
  assign y16325 = n35367 ;
  assign y16326 = n35370 ;
  assign y16327 = ~n35373 ;
  assign y16328 = 1'b0 ;
  assign y16329 = ~n30260 ;
  assign y16330 = n35376 ;
  assign y16331 = ~n35377 ;
  assign y16332 = ~1'b0 ;
  assign y16333 = ~1'b0 ;
  assign y16334 = n35389 ;
  assign y16335 = ~n35393 ;
  assign y16336 = ~n35396 ;
  assign y16337 = ~n35397 ;
  assign y16338 = ~n35399 ;
  assign y16339 = n35403 ;
  assign y16340 = ~1'b0 ;
  assign y16341 = n35408 ;
  assign y16342 = n8501 ;
  assign y16343 = ~1'b0 ;
  assign y16344 = n35412 ;
  assign y16345 = n35413 ;
  assign y16346 = ~n35415 ;
  assign y16347 = ~n35420 ;
  assign y16348 = ~1'b0 ;
  assign y16349 = n35422 ;
  assign y16350 = n35425 ;
  assign y16351 = n35426 ;
  assign y16352 = ~1'b0 ;
  assign y16353 = 1'b0 ;
  assign y16354 = ~n35430 ;
  assign y16355 = n35431 ;
  assign y16356 = ~1'b0 ;
  assign y16357 = n35436 ;
  assign y16358 = n35437 ;
  assign y16359 = n35438 ;
  assign y16360 = ~n35439 ;
  assign y16361 = n35440 ;
  assign y16362 = n35443 ;
  assign y16363 = ~n3359 ;
  assign y16364 = ~1'b0 ;
  assign y16365 = n35457 ;
  assign y16366 = n35458 ;
  assign y16367 = ~1'b0 ;
  assign y16368 = n35459 ;
  assign y16369 = n35460 ;
  assign y16370 = ~n35461 ;
  assign y16371 = ~1'b0 ;
  assign y16372 = n35465 ;
  assign y16373 = ~1'b0 ;
  assign y16374 = ~1'b0 ;
  assign y16375 = ~n35466 ;
  assign y16376 = n35470 ;
  assign y16377 = n35472 ;
  assign y16378 = n35474 ;
  assign y16379 = n35478 ;
  assign y16380 = ~n35481 ;
  assign y16381 = ~n35482 ;
  assign y16382 = n15005 ;
  assign y16383 = ~n35483 ;
  assign y16384 = ~1'b0 ;
  assign y16385 = ~1'b0 ;
  assign y16386 = n35487 ;
  assign y16387 = n19287 ;
  assign y16388 = ~1'b0 ;
  assign y16389 = n35492 ;
  assign y16390 = n35493 ;
  assign y16391 = ~n35496 ;
  assign y16392 = ~1'b0 ;
  assign y16393 = ~n35498 ;
  assign y16394 = n35500 ;
  assign y16395 = ~1'b0 ;
  assign y16396 = ~n35505 ;
  assign y16397 = ~n35509 ;
  assign y16398 = ~n35513 ;
  assign y16399 = ~1'b0 ;
  assign y16400 = n35515 ;
  assign y16401 = n35520 ;
  assign y16402 = ~n35521 ;
  assign y16403 = ~n35522 ;
  assign y16404 = ~n35524 ;
  assign y16405 = ~n13054 ;
  assign y16406 = n35526 ;
  assign y16407 = n35528 ;
  assign y16408 = ~n35529 ;
  assign y16409 = ~1'b0 ;
  assign y16410 = ~1'b0 ;
  assign y16411 = ~n35533 ;
  assign y16412 = n35534 ;
  assign y16413 = ~n35535 ;
  assign y16414 = ~n4073 ;
  assign y16415 = n35537 ;
  assign y16416 = ~1'b0 ;
  assign y16417 = ~1'b0 ;
  assign y16418 = ~1'b0 ;
  assign y16419 = ~1'b0 ;
  assign y16420 = ~n35539 ;
  assign y16421 = ~n35541 ;
  assign y16422 = ~1'b0 ;
  assign y16423 = ~1'b0 ;
  assign y16424 = n35546 ;
  assign y16425 = ~1'b0 ;
  assign y16426 = ~n16419 ;
  assign y16427 = 1'b0 ;
  assign y16428 = 1'b0 ;
  assign y16429 = n3104 ;
  assign y16430 = ~n35547 ;
  assign y16431 = ~1'b0 ;
  assign y16432 = n35549 ;
  assign y16433 = ~1'b0 ;
  assign y16434 = ~1'b0 ;
  assign y16435 = n35550 ;
  assign y16436 = n35553 ;
  assign y16437 = ~n35555 ;
  assign y16438 = n35558 ;
  assign y16439 = n35559 ;
  assign y16440 = 1'b0 ;
  assign y16441 = ~n35561 ;
  assign y16442 = ~1'b0 ;
  assign y16443 = ~n35566 ;
  assign y16444 = n35567 ;
  assign y16445 = ~n35568 ;
  assign y16446 = n35570 ;
  assign y16447 = n35573 ;
  assign y16448 = ~1'b0 ;
  assign y16449 = ~n35576 ;
  assign y16450 = n35579 ;
  assign y16451 = n35585 ;
  assign y16452 = ~1'b0 ;
  assign y16453 = n35589 ;
  assign y16454 = ~n35592 ;
  assign y16455 = ~n35593 ;
  assign y16456 = ~n35595 ;
  assign y16457 = ~n35596 ;
  assign y16458 = ~n35599 ;
  assign y16459 = n35601 ;
  assign y16460 = n35605 ;
  assign y16461 = n35607 ;
  assign y16462 = n35608 ;
  assign y16463 = n9056 ;
  assign y16464 = n35609 ;
  assign y16465 = ~n35610 ;
  assign y16466 = ~n35614 ;
  assign y16467 = ~n10560 ;
  assign y16468 = ~1'b0 ;
  assign y16469 = ~n35616 ;
  assign y16470 = n35618 ;
  assign y16471 = n35620 ;
  assign y16472 = ~n35623 ;
  assign y16473 = 1'b0 ;
  assign y16474 = ~1'b0 ;
  assign y16475 = ~1'b0 ;
  assign y16476 = ~n1805 ;
  assign y16477 = n35628 ;
  assign y16478 = ~1'b0 ;
  assign y16479 = n35630 ;
  assign y16480 = ~1'b0 ;
  assign y16481 = ~n35631 ;
  assign y16482 = ~n35632 ;
  assign y16483 = ~1'b0 ;
  assign y16484 = n35634 ;
  assign y16485 = 1'b0 ;
  assign y16486 = ~1'b0 ;
  assign y16487 = n35639 ;
  assign y16488 = n35640 ;
  assign y16489 = n35641 ;
  assign y16490 = ~1'b0 ;
  assign y16491 = ~n18399 ;
  assign y16492 = ~n35643 ;
  assign y16493 = ~1'b0 ;
  assign y16494 = 1'b0 ;
  assign y16495 = n35646 ;
  assign y16496 = ~n35647 ;
  assign y16497 = n24097 ;
  assign y16498 = ~n35648 ;
  assign y16499 = n35652 ;
  assign y16500 = ~n35654 ;
  assign y16501 = ~n35656 ;
  assign y16502 = ~n35657 ;
  assign y16503 = n12355 ;
  assign y16504 = ~1'b0 ;
  assign y16505 = ~n35659 ;
  assign y16506 = ~n35660 ;
  assign y16507 = ~1'b0 ;
  assign y16508 = ~1'b0 ;
  assign y16509 = ~n35661 ;
  assign y16510 = ~1'b0 ;
  assign y16511 = ~n35663 ;
  assign y16512 = ~n35664 ;
  assign y16513 = n35665 ;
  assign y16514 = n19157 ;
  assign y16515 = n35668 ;
  assign y16516 = n35672 ;
  assign y16517 = ~n22256 ;
  assign y16518 = ~1'b0 ;
  assign y16519 = ~n35675 ;
  assign y16520 = ~1'b0 ;
  assign y16521 = ~n35680 ;
  assign y16522 = ~1'b0 ;
  assign y16523 = ~n35683 ;
  assign y16524 = ~n35684 ;
  assign y16525 = n35686 ;
  assign y16526 = n9501 ;
  assign y16527 = ~1'b0 ;
  assign y16528 = n35691 ;
  assign y16529 = n35693 ;
  assign y16530 = n35695 ;
  assign y16531 = ~n35696 ;
  assign y16532 = ~n35697 ;
  assign y16533 = ~n35700 ;
  assign y16534 = ~n35701 ;
  assign y16535 = ~n3540 ;
  assign y16536 = ~n35706 ;
  assign y16537 = n35710 ;
  assign y16538 = n35711 ;
  assign y16539 = ~1'b0 ;
  assign y16540 = ~1'b0 ;
  assign y16541 = ~1'b0 ;
  assign y16542 = ~1'b0 ;
  assign y16543 = n35713 ;
  assign y16544 = n35714 ;
  assign y16545 = ~n35715 ;
  assign y16546 = ~n35718 ;
  assign y16547 = ~1'b0 ;
  assign y16548 = ~1'b0 ;
  assign y16549 = ~n35720 ;
  assign y16550 = ~n35721 ;
  assign y16551 = n35722 ;
  assign y16552 = ~n35726 ;
  assign y16553 = ~n35730 ;
  assign y16554 = n16082 ;
  assign y16555 = n3148 ;
  assign y16556 = n35731 ;
  assign y16557 = ~n35736 ;
  assign y16558 = ~n35740 ;
  assign y16559 = n35742 ;
  assign y16560 = n35743 ;
  assign y16561 = n35747 ;
  assign y16562 = ~n35749 ;
  assign y16563 = ~n35752 ;
  assign y16564 = n35755 ;
  assign y16565 = n35756 ;
  assign y16566 = n35757 ;
  assign y16567 = ~1'b0 ;
  assign y16568 = n35760 ;
  assign y16569 = ~1'b0 ;
  assign y16570 = ~n35764 ;
  assign y16571 = n35766 ;
  assign y16572 = n35767 ;
  assign y16573 = n35768 ;
  assign y16574 = n35771 ;
  assign y16575 = ~n35774 ;
  assign y16576 = ~n18218 ;
  assign y16577 = n35776 ;
  assign y16578 = n35777 ;
  assign y16579 = n35778 ;
  assign y16580 = ~n35780 ;
  assign y16581 = ~n35784 ;
  assign y16582 = n35786 ;
  assign y16583 = ~1'b0 ;
  assign y16584 = ~n35787 ;
  assign y16585 = n35788 ;
  assign y16586 = ~n35793 ;
  assign y16587 = n35795 ;
  assign y16588 = ~n35796 ;
  assign y16589 = ~1'b0 ;
  assign y16590 = ~1'b0 ;
  assign y16591 = n35798 ;
  assign y16592 = ~n35800 ;
  assign y16593 = n35802 ;
  assign y16594 = n35803 ;
  assign y16595 = n35805 ;
  assign y16596 = ~n35807 ;
  assign y16597 = ~n35809 ;
  assign y16598 = ~n35811 ;
  assign y16599 = ~n35812 ;
  assign y16600 = ~n35813 ;
  assign y16601 = ~n35814 ;
  assign y16602 = n35817 ;
  assign y16603 = ~n35818 ;
  assign y16604 = ~n35821 ;
  assign y16605 = ~n35825 ;
  assign y16606 = ~1'b0 ;
  assign y16607 = 1'b0 ;
  assign y16608 = n35828 ;
  assign y16609 = ~n35829 ;
  assign y16610 = ~1'b0 ;
  assign y16611 = ~n35832 ;
  assign y16612 = n35833 ;
  assign y16613 = ~1'b0 ;
  assign y16614 = ~n35835 ;
  assign y16615 = n781 ;
  assign y16616 = ~1'b0 ;
  assign y16617 = ~1'b0 ;
  assign y16618 = ~1'b0 ;
  assign y16619 = ~n35837 ;
  assign y16620 = ~n35839 ;
  assign y16621 = n25440 ;
  assign y16622 = ~n35842 ;
  assign y16623 = ~n35844 ;
  assign y16624 = ~n35849 ;
  assign y16625 = ~1'b0 ;
  assign y16626 = ~n35850 ;
  assign y16627 = n35856 ;
  assign y16628 = n35859 ;
  assign y16629 = ~1'b0 ;
  assign y16630 = 1'b0 ;
  assign y16631 = n35861 ;
  assign y16632 = ~n35862 ;
  assign y16633 = ~1'b0 ;
  assign y16634 = ~n12571 ;
  assign y16635 = ~1'b0 ;
  assign y16636 = n35863 ;
  assign y16637 = ~n12191 ;
  assign y16638 = 1'b0 ;
  assign y16639 = n35868 ;
  assign y16640 = ~1'b0 ;
  assign y16641 = ~n35871 ;
  assign y16642 = ~n35876 ;
  assign y16643 = n35879 ;
  assign y16644 = ~1'b0 ;
  assign y16645 = ~1'b0 ;
  assign y16646 = n35880 ;
  assign y16647 = 1'b0 ;
  assign y16648 = n35882 ;
  assign y16649 = ~n35884 ;
  assign y16650 = n35885 ;
  assign y16651 = n35886 ;
  assign y16652 = ~1'b0 ;
  assign y16653 = ~1'b0 ;
  assign y16654 = n5375 ;
  assign y16655 = ~n35892 ;
  assign y16656 = ~n35897 ;
  assign y16657 = ~n35898 ;
  assign y16658 = ~n35899 ;
  assign y16659 = ~n7992 ;
  assign y16660 = ~1'b0 ;
  assign y16661 = ~n35903 ;
  assign y16662 = ~n35904 ;
  assign y16663 = ~1'b0 ;
  assign y16664 = ~n35906 ;
  assign y16665 = ~n35907 ;
  assign y16666 = n35911 ;
  assign y16667 = ~n35913 ;
  assign y16668 = ~1'b0 ;
  assign y16669 = ~1'b0 ;
  assign y16670 = ~n35915 ;
  assign y16671 = ~n35917 ;
  assign y16672 = ~1'b0 ;
  assign y16673 = ~n35925 ;
  assign y16674 = n35928 ;
  assign y16675 = n35931 ;
  assign y16676 = n35936 ;
  assign y16677 = ~1'b0 ;
  assign y16678 = n35938 ;
  assign y16679 = n15388 ;
  assign y16680 = ~1'b0 ;
  assign y16681 = n35939 ;
  assign y16682 = ~n35941 ;
  assign y16683 = n35942 ;
  assign y16684 = n35946 ;
  assign y16685 = ~n35948 ;
  assign y16686 = n35950 ;
  assign y16687 = ~n8632 ;
  assign y16688 = ~1'b0 ;
  assign y16689 = ~1'b0 ;
  assign y16690 = ~n35951 ;
  assign y16691 = n35953 ;
  assign y16692 = ~n35955 ;
  assign y16693 = ~1'b0 ;
  assign y16694 = ~n35957 ;
  assign y16695 = n35958 ;
  assign y16696 = n16823 ;
  assign y16697 = n35964 ;
  assign y16698 = ~n35967 ;
  assign y16699 = n35971 ;
  assign y16700 = ~n35977 ;
  assign y16701 = ~n35979 ;
  assign y16702 = ~n35981 ;
  assign y16703 = ~n35983 ;
  assign y16704 = n35984 ;
  assign y16705 = ~1'b0 ;
  assign y16706 = n35985 ;
  assign y16707 = ~n35986 ;
  assign y16708 = ~n35989 ;
  assign y16709 = n35991 ;
  assign y16710 = ~n35994 ;
  assign y16711 = ~1'b0 ;
  assign y16712 = ~n36001 ;
  assign y16713 = ~1'b0 ;
  assign y16714 = ~1'b0 ;
  assign y16715 = ~n36004 ;
  assign y16716 = n36006 ;
  assign y16717 = ~1'b0 ;
  assign y16718 = n36007 ;
  assign y16719 = n36010 ;
  assign y16720 = ~1'b0 ;
  assign y16721 = ~1'b0 ;
  assign y16722 = ~n36013 ;
  assign y16723 = ~n36017 ;
  assign y16724 = n36021 ;
  assign y16725 = ~n36024 ;
  assign y16726 = n36026 ;
  assign y16727 = n36029 ;
  assign y16728 = ~n36032 ;
  assign y16729 = n36034 ;
  assign y16730 = ~n36036 ;
  assign y16731 = n36044 ;
  assign y16732 = ~n36045 ;
  assign y16733 = n36046 ;
  assign y16734 = n36049 ;
  assign y16735 = ~n36051 ;
  assign y16736 = ~n36054 ;
  assign y16737 = n36057 ;
  assign y16738 = ~1'b0 ;
  assign y16739 = ~n36058 ;
  assign y16740 = 1'b0 ;
  assign y16741 = ~n36061 ;
  assign y16742 = n36064 ;
  assign y16743 = ~n36065 ;
  assign y16744 = ~n36068 ;
  assign y16745 = ~n36069 ;
  assign y16746 = ~1'b0 ;
  assign y16747 = n30878 ;
  assign y16748 = ~n36070 ;
  assign y16749 = n36073 ;
  assign y16750 = n36074 ;
  assign y16751 = ~n36075 ;
  assign y16752 = ~1'b0 ;
  assign y16753 = ~n36084 ;
  assign y16754 = ~n36087 ;
  assign y16755 = ~n583 ;
  assign y16756 = ~1'b0 ;
  assign y16757 = ~1'b0 ;
  assign y16758 = ~n36088 ;
  assign y16759 = ~n36089 ;
  assign y16760 = ~n36091 ;
  assign y16761 = ~n25953 ;
  assign y16762 = n36092 ;
  assign y16763 = ~1'b0 ;
  assign y16764 = ~1'b0 ;
  assign y16765 = ~n36093 ;
  assign y16766 = n36096 ;
  assign y16767 = ~1'b0 ;
  assign y16768 = ~n36098 ;
  assign y16769 = ~n36100 ;
  assign y16770 = ~1'b0 ;
  assign y16771 = n36101 ;
  assign y16772 = ~1'b0 ;
  assign y16773 = n36102 ;
  assign y16774 = n36104 ;
  assign y16775 = ~n36109 ;
  assign y16776 = ~n36111 ;
  assign y16777 = ~n36114 ;
  assign y16778 = ~1'b0 ;
  assign y16779 = ~1'b0 ;
  assign y16780 = ~1'b0 ;
  assign y16781 = ~n2380 ;
  assign y16782 = ~1'b0 ;
  assign y16783 = ~n36116 ;
  assign y16784 = ~n36117 ;
  assign y16785 = n36120 ;
  assign y16786 = ~1'b0 ;
  assign y16787 = ~n36126 ;
  assign y16788 = ~1'b0 ;
  assign y16789 = ~1'b0 ;
  assign y16790 = n36129 ;
  assign y16791 = n36133 ;
  assign y16792 = ~1'b0 ;
  assign y16793 = ~n36134 ;
  assign y16794 = ~n36135 ;
  assign y16795 = ~n36138 ;
  assign y16796 = ~n9304 ;
  assign y16797 = ~1'b0 ;
  assign y16798 = ~n36143 ;
  assign y16799 = n28927 ;
  assign y16800 = ~n36145 ;
  assign y16801 = ~n36147 ;
  assign y16802 = n36149 ;
  assign y16803 = ~n36152 ;
  assign y16804 = ~n36156 ;
  assign y16805 = ~n36158 ;
  assign y16806 = n36160 ;
  assign y16807 = n36161 ;
  assign y16808 = n36163 ;
  assign y16809 = ~n36166 ;
  assign y16810 = n36173 ;
  assign y16811 = ~1'b0 ;
  assign y16812 = n36174 ;
  assign y16813 = ~n32738 ;
  assign y16814 = ~n36175 ;
  assign y16815 = ~n36179 ;
  assign y16816 = n36182 ;
  assign y16817 = n36184 ;
  assign y16818 = ~n36193 ;
  assign y16819 = ~1'b0 ;
  assign y16820 = ~n36194 ;
  assign y16821 = ~n36195 ;
  assign y16822 = ~1'b0 ;
  assign y16823 = n36197 ;
  assign y16824 = n1506 ;
  assign y16825 = ~1'b0 ;
  assign y16826 = ~n36198 ;
  assign y16827 = n36200 ;
  assign y16828 = ~n36203 ;
  assign y16829 = ~n36205 ;
  assign y16830 = ~1'b0 ;
  assign y16831 = n36209 ;
  assign y16832 = n36210 ;
  assign y16833 = ~n36213 ;
  assign y16834 = n36214 ;
  assign y16835 = n36216 ;
  assign y16836 = ~n36217 ;
  assign y16837 = ~1'b0 ;
  assign y16838 = ~n36219 ;
  assign y16839 = ~n36220 ;
  assign y16840 = n36221 ;
  assign y16841 = n36222 ;
  assign y16842 = ~1'b0 ;
  assign y16843 = n36224 ;
  assign y16844 = n36226 ;
  assign y16845 = n36228 ;
  assign y16846 = ~1'b0 ;
  assign y16847 = n36233 ;
  assign y16848 = 1'b0 ;
  assign y16849 = n36234 ;
  assign y16850 = ~1'b0 ;
  assign y16851 = ~n36236 ;
  assign y16852 = ~n36243 ;
  assign y16853 = n36244 ;
  assign y16854 = n36246 ;
  assign y16855 = ~1'b0 ;
  assign y16856 = ~n36253 ;
  assign y16857 = n36263 ;
  assign y16858 = ~n36264 ;
  assign y16859 = n36267 ;
  assign y16860 = ~n36271 ;
  assign y16861 = n36276 ;
  assign y16862 = ~1'b0 ;
  assign y16863 = n36277 ;
  assign y16864 = n36279 ;
  assign y16865 = n36280 ;
  assign y16866 = ~n36284 ;
  assign y16867 = n36285 ;
  assign y16868 = n16077 ;
  assign y16869 = n36286 ;
  assign y16870 = ~1'b0 ;
  assign y16871 = n36290 ;
  assign y16872 = n36293 ;
  assign y16873 = ~1'b0 ;
  assign y16874 = ~n36295 ;
  assign y16875 = n36300 ;
  assign y16876 = ~n36301 ;
  assign y16877 = n36302 ;
  assign y16878 = n36303 ;
  assign y16879 = ~n36307 ;
  assign y16880 = ~1'b0 ;
  assign y16881 = ~n36308 ;
  assign y16882 = ~n36310 ;
  assign y16883 = x124 ;
  assign y16884 = ~n36314 ;
  assign y16885 = ~n36317 ;
  assign y16886 = n36322 ;
  assign y16887 = n36324 ;
  assign y16888 = n36326 ;
  assign y16889 = ~1'b0 ;
  assign y16890 = n36327 ;
  assign y16891 = n36331 ;
  assign y16892 = n36332 ;
  assign y16893 = ~n36334 ;
  assign y16894 = ~n36339 ;
  assign y16895 = ~n36342 ;
  assign y16896 = n36345 ;
  assign y16897 = n36346 ;
  assign y16898 = n5963 ;
  assign y16899 = ~n36350 ;
  assign y16900 = n36351 ;
  assign y16901 = n36353 ;
  assign y16902 = ~1'b0 ;
  assign y16903 = ~n36356 ;
  assign y16904 = n296 ;
  assign y16905 = n36357 ;
  assign y16906 = n36358 ;
  assign y16907 = n36362 ;
  assign y16908 = 1'b0 ;
  assign y16909 = n36364 ;
  assign y16910 = n36365 ;
  assign y16911 = ~1'b0 ;
  assign y16912 = n36366 ;
  assign y16913 = ~n36367 ;
  assign y16914 = ~n36368 ;
  assign y16915 = n36370 ;
  assign y16916 = ~1'b0 ;
  assign y16917 = ~n36372 ;
  assign y16918 = n36373 ;
  assign y16919 = ~n36374 ;
  assign y16920 = ~n36375 ;
  assign y16921 = ~n36378 ;
  assign y16922 = n36379 ;
  assign y16923 = ~1'b0 ;
  assign y16924 = n36383 ;
  assign y16925 = ~1'b0 ;
  assign y16926 = n36384 ;
  assign y16927 = n36386 ;
  assign y16928 = n36387 ;
  assign y16929 = ~n36388 ;
  assign y16930 = n36391 ;
  assign y16931 = n36392 ;
  assign y16932 = ~n15014 ;
  assign y16933 = ~1'b0 ;
  assign y16934 = ~n36396 ;
  assign y16935 = ~n36402 ;
  assign y16936 = ~1'b0 ;
  assign y16937 = ~1'b0 ;
  assign y16938 = ~1'b0 ;
  assign y16939 = ~n36404 ;
  assign y16940 = n36405 ;
  assign y16941 = ~n36407 ;
  assign y16942 = n36413 ;
  assign y16943 = n36414 ;
  assign y16944 = n36415 ;
  assign y16945 = ~1'b0 ;
  assign y16946 = ~n36419 ;
  assign y16947 = n36421 ;
  assign y16948 = n36422 ;
  assign y16949 = ~n36426 ;
  assign y16950 = ~n36427 ;
  assign y16951 = n36431 ;
  assign y16952 = n36435 ;
  assign y16953 = n36436 ;
  assign y16954 = ~1'b0 ;
  assign y16955 = n17669 ;
  assign y16956 = ~n36437 ;
  assign y16957 = n36440 ;
  assign y16958 = ~1'b0 ;
  assign y16959 = ~n36442 ;
  assign y16960 = ~n36445 ;
  assign y16961 = ~n36452 ;
  assign y16962 = ~n36453 ;
  assign y16963 = ~n36455 ;
  assign y16964 = n36456 ;
  assign y16965 = n36457 ;
  assign y16966 = 1'b0 ;
  assign y16967 = n36458 ;
  assign y16968 = n36459 ;
  assign y16969 = ~n36461 ;
  assign y16970 = ~1'b0 ;
  assign y16971 = ~n36462 ;
  assign y16972 = 1'b0 ;
  assign y16973 = n36464 ;
  assign y16974 = ~n36465 ;
  assign y16975 = n36466 ;
  assign y16976 = n36467 ;
  assign y16977 = ~1'b0 ;
  assign y16978 = n36474 ;
  assign y16979 = n36475 ;
  assign y16980 = n36479 ;
  assign y16981 = ~1'b0 ;
  assign y16982 = ~1'b0 ;
  assign y16983 = ~n36483 ;
  assign y16984 = ~n36486 ;
  assign y16985 = ~n36487 ;
  assign y16986 = n36490 ;
  assign y16987 = ~1'b0 ;
  assign y16988 = ~n36491 ;
  assign y16989 = n36496 ;
  assign y16990 = n36500 ;
  assign y16991 = 1'b0 ;
  assign y16992 = n36501 ;
  assign y16993 = ~1'b0 ;
  assign y16994 = n36503 ;
  assign y16995 = n36505 ;
  assign y16996 = ~n36509 ;
  assign y16997 = ~n36510 ;
  assign y16998 = n36512 ;
  assign y16999 = ~1'b0 ;
  assign y17000 = ~n35908 ;
  assign y17001 = ~n36515 ;
  assign y17002 = ~1'b0 ;
  assign y17003 = ~n36517 ;
  assign y17004 = n36519 ;
  assign y17005 = n36522 ;
  assign y17006 = ~n36525 ;
  assign y17007 = ~1'b0 ;
  assign y17008 = ~n36529 ;
  assign y17009 = ~n36531 ;
  assign y17010 = n36534 ;
  assign y17011 = n36535 ;
  assign y17012 = n36536 ;
  assign y17013 = ~n36538 ;
  assign y17014 = n36540 ;
  assign y17015 = n36542 ;
  assign y17016 = n36544 ;
  assign y17017 = n36545 ;
  assign y17018 = ~n36547 ;
  assign y17019 = n36552 ;
  assign y17020 = ~1'b0 ;
  assign y17021 = ~n36554 ;
  assign y17022 = n36557 ;
  assign y17023 = n17063 ;
  assign y17024 = n36560 ;
  assign y17025 = ~1'b0 ;
  assign y17026 = n36561 ;
  assign y17027 = n36562 ;
  assign y17028 = n36566 ;
  assign y17029 = n36569 ;
  assign y17030 = n36573 ;
  assign y17031 = ~n36577 ;
  assign y17032 = ~n36579 ;
  assign y17033 = n36581 ;
  assign y17034 = n36582 ;
  assign y17035 = ~1'b0 ;
  assign y17036 = ~n36583 ;
  assign y17037 = n36586 ;
  assign y17038 = ~n36589 ;
  assign y17039 = n36592 ;
  assign y17040 = n36593 ;
  assign y17041 = ~n36595 ;
  assign y17042 = ~1'b0 ;
  assign y17043 = ~1'b0 ;
  assign y17044 = ~1'b0 ;
  assign y17045 = ~1'b0 ;
  assign y17046 = n36596 ;
  assign y17047 = n36598 ;
  assign y17048 = n36601 ;
  assign y17049 = ~1'b0 ;
  assign y17050 = ~1'b0 ;
  assign y17051 = ~1'b0 ;
  assign y17052 = n36602 ;
  assign y17053 = n36604 ;
  assign y17054 = n36605 ;
  assign y17055 = n36606 ;
  assign y17056 = ~n36610 ;
  assign y17057 = ~1'b0 ;
  assign y17058 = ~n36612 ;
  assign y17059 = ~1'b0 ;
  assign y17060 = ~n36613 ;
  assign y17061 = ~n36614 ;
  assign y17062 = ~n36616 ;
  assign y17063 = ~n36618 ;
  assign y17064 = n36620 ;
  assign y17065 = ~1'b0 ;
  assign y17066 = ~1'b0 ;
  assign y17067 = n36621 ;
  assign y17068 = ~n36624 ;
  assign y17069 = n36625 ;
  assign y17070 = n36626 ;
  assign y17071 = ~n36627 ;
  assign y17072 = ~1'b0 ;
  assign y17073 = ~1'b0 ;
  assign y17074 = n36630 ;
  assign y17075 = ~n36634 ;
  assign y17076 = ~1'b0 ;
  assign y17077 = n36635 ;
  assign y17078 = ~1'b0 ;
  assign y17079 = n36638 ;
  assign y17080 = ~n36643 ;
  assign y17081 = ~n36647 ;
  assign y17082 = n36648 ;
  assign y17083 = ~1'b0 ;
  assign y17084 = ~n36649 ;
  assign y17085 = ~n36653 ;
  assign y17086 = n31119 ;
  assign y17087 = ~n36656 ;
  assign y17088 = n16310 ;
  assign y17089 = n36661 ;
  assign y17090 = n36669 ;
  assign y17091 = ~n36671 ;
  assign y17092 = n36673 ;
  assign y17093 = n36675 ;
  assign y17094 = ~n36677 ;
  assign y17095 = ~1'b0 ;
  assign y17096 = ~n327 ;
  assign y17097 = n7817 ;
  assign y17098 = ~n36681 ;
  assign y17099 = ~1'b0 ;
  assign y17100 = n36684 ;
  assign y17101 = n36687 ;
  assign y17102 = n36689 ;
  assign y17103 = n36691 ;
  assign y17104 = ~n36693 ;
  assign y17105 = ~n36696 ;
  assign y17106 = ~n36698 ;
  assign y17107 = ~n36699 ;
  assign y17108 = ~1'b0 ;
  assign y17109 = ~n36701 ;
  assign y17110 = ~1'b0 ;
  assign y17111 = ~1'b0 ;
  assign y17112 = ~1'b0 ;
  assign y17113 = ~1'b0 ;
  assign y17114 = ~n36702 ;
  assign y17115 = ~n36703 ;
  assign y17116 = n36704 ;
  assign y17117 = ~n36707 ;
  assign y17118 = n36708 ;
  assign y17119 = n36711 ;
  assign y17120 = ~1'b0 ;
  assign y17121 = n36718 ;
  assign y17122 = ~n36719 ;
  assign y17123 = ~1'b0 ;
  assign y17124 = ~n36723 ;
  assign y17125 = ~1'b0 ;
  assign y17126 = ~n36724 ;
  assign y17127 = ~1'b0 ;
  assign y17128 = n36725 ;
  assign y17129 = n36727 ;
  assign y17130 = n36729 ;
  assign y17131 = ~n36733 ;
  assign y17132 = ~n36738 ;
  assign y17133 = ~n36746 ;
  assign y17134 = ~n5689 ;
  assign y17135 = ~1'b0 ;
  assign y17136 = n36747 ;
  assign y17137 = 1'b0 ;
  assign y17138 = n36750 ;
  assign y17139 = ~n36753 ;
  assign y17140 = ~n36755 ;
  assign y17141 = ~1'b0 ;
  assign y17142 = ~n36761 ;
  assign y17143 = n36762 ;
  assign y17144 = n36768 ;
  assign y17145 = ~1'b0 ;
  assign y17146 = ~1'b0 ;
  assign y17147 = 1'b0 ;
  assign y17148 = ~n36771 ;
  assign y17149 = n36773 ;
  assign y17150 = n36775 ;
  assign y17151 = n36776 ;
  assign y17152 = ~n36777 ;
  assign y17153 = n36778 ;
  assign y17154 = ~n36782 ;
  assign y17155 = ~1'b0 ;
  assign y17156 = ~n36784 ;
  assign y17157 = n36786 ;
  assign y17158 = ~n36787 ;
  assign y17159 = ~1'b0 ;
  assign y17160 = n36791 ;
  assign y17161 = ~n36793 ;
  assign y17162 = ~n24737 ;
  assign y17163 = n36796 ;
  assign y17164 = ~n36798 ;
  assign y17165 = ~n36799 ;
  assign y17166 = ~n36800 ;
  assign y17167 = ~1'b0 ;
  assign y17168 = n36804 ;
  assign y17169 = n36810 ;
  assign y17170 = n36814 ;
  assign y17171 = ~1'b0 ;
  assign y17172 = n36816 ;
  assign y17173 = ~n9783 ;
  assign y17174 = ~1'b0 ;
  assign y17175 = n36820 ;
  assign y17176 = ~n36822 ;
  assign y17177 = n36823 ;
  assign y17178 = n36824 ;
  assign y17179 = ~1'b0 ;
  assign y17180 = n36826 ;
  assign y17181 = 1'b0 ;
  assign y17182 = ~1'b0 ;
  assign y17183 = n36833 ;
  assign y17184 = ~1'b0 ;
  assign y17185 = n16642 ;
  assign y17186 = n36835 ;
  assign y17187 = ~1'b0 ;
  assign y17188 = ~n36839 ;
  assign y17189 = ~n36843 ;
  assign y17190 = ~n36845 ;
  assign y17191 = n36846 ;
  assign y17192 = ~1'b0 ;
  assign y17193 = ~n36848 ;
  assign y17194 = ~n36849 ;
  assign y17195 = n36852 ;
  assign y17196 = 1'b0 ;
  assign y17197 = n36853 ;
  assign y17198 = ~n36855 ;
  assign y17199 = ~n36857 ;
  assign y17200 = ~n36859 ;
  assign y17201 = ~n36860 ;
  assign y17202 = ~n11237 ;
  assign y17203 = n36861 ;
  assign y17204 = ~1'b0 ;
  assign y17205 = ~n36865 ;
  assign y17206 = n36870 ;
  assign y17207 = n36872 ;
  assign y17208 = n36873 ;
  assign y17209 = n36875 ;
  assign y17210 = ~n36883 ;
  assign y17211 = ~n36884 ;
  assign y17212 = n36885 ;
  assign y17213 = n34404 ;
  assign y17214 = 1'b0 ;
  assign y17215 = ~1'b0 ;
  assign y17216 = ~1'b0 ;
  assign y17217 = ~1'b0 ;
  assign y17218 = n36886 ;
  assign y17219 = ~n20098 ;
  assign y17220 = ~n36894 ;
  assign y17221 = ~n36895 ;
  assign y17222 = n36900 ;
  assign y17223 = ~1'b0 ;
  assign y17224 = n36902 ;
  assign y17225 = ~1'b0 ;
  assign y17226 = ~1'b0 ;
  assign y17227 = ~n36906 ;
  assign y17228 = ~1'b0 ;
  assign y17229 = ~1'b0 ;
  assign y17230 = n36911 ;
  assign y17231 = ~1'b0 ;
  assign y17232 = 1'b0 ;
  assign y17233 = n36915 ;
  assign y17234 = ~1'b0 ;
  assign y17235 = ~1'b0 ;
  assign y17236 = ~n36919 ;
  assign y17237 = n36921 ;
  assign y17238 = n36922 ;
  assign y17239 = n36928 ;
  assign y17240 = ~1'b0 ;
  assign y17241 = ~1'b0 ;
  assign y17242 = ~n36929 ;
  assign y17243 = n36932 ;
  assign y17244 = 1'b0 ;
  assign y17245 = ~1'b0 ;
  assign y17246 = ~1'b0 ;
  assign y17247 = n36933 ;
  assign y17248 = ~1'b0 ;
  assign y17249 = ~n10329 ;
  assign y17250 = ~1'b0 ;
  assign y17251 = n36935 ;
  assign y17252 = ~1'b0 ;
  assign y17253 = ~1'b0 ;
  assign y17254 = ~n36936 ;
  assign y17255 = n36938 ;
  assign y17256 = ~n36940 ;
  assign y17257 = ~n36941 ;
  assign y17258 = ~n36943 ;
  assign y17259 = ~n36944 ;
  assign y17260 = ~1'b0 ;
  assign y17261 = n36947 ;
  assign y17262 = 1'b0 ;
  assign y17263 = ~n36951 ;
  assign y17264 = ~1'b0 ;
  assign y17265 = ~1'b0 ;
  assign y17266 = ~n36952 ;
  assign y17267 = ~1'b0 ;
  assign y17268 = ~1'b0 ;
  assign y17269 = ~1'b0 ;
  assign y17270 = n36954 ;
  assign y17271 = ~n36955 ;
  assign y17272 = ~n36956 ;
  assign y17273 = ~1'b0 ;
  assign y17274 = ~1'b0 ;
  assign y17275 = ~1'b0 ;
  assign y17276 = ~n36957 ;
  assign y17277 = ~n35504 ;
  assign y17278 = 1'b0 ;
  assign y17279 = n36958 ;
  assign y17280 = ~n36959 ;
  assign y17281 = ~1'b0 ;
  assign y17282 = ~n36963 ;
  assign y17283 = ~n36965 ;
  assign y17284 = n36966 ;
  assign y17285 = n36970 ;
  assign y17286 = ~n36976 ;
  assign y17287 = n36977 ;
  assign y17288 = ~n36980 ;
  assign y17289 = ~1'b0 ;
  assign y17290 = n36984 ;
  assign y17291 = ~n36986 ;
  assign y17292 = n36987 ;
  assign y17293 = ~n11033 ;
  assign y17294 = n36991 ;
  assign y17295 = n36993 ;
  assign y17296 = ~1'b0 ;
  assign y17297 = ~1'b0 ;
  assign y17298 = n36995 ;
  assign y17299 = n36997 ;
  assign y17300 = n36999 ;
  assign y17301 = n37001 ;
  assign y17302 = ~n37002 ;
  assign y17303 = ~1'b0 ;
  assign y17304 = n37003 ;
  assign y17305 = ~n37004 ;
  assign y17306 = ~1'b0 ;
  assign y17307 = ~n37007 ;
  assign y17308 = ~n32419 ;
  assign y17309 = ~1'b0 ;
  assign y17310 = n37009 ;
  assign y17311 = ~n37014 ;
  assign y17312 = n37015 ;
  assign y17313 = ~1'b0 ;
  assign y17314 = ~1'b0 ;
  assign y17315 = ~n37017 ;
  assign y17316 = n37019 ;
  assign y17317 = ~1'b0 ;
  assign y17318 = ~1'b0 ;
  assign y17319 = ~1'b0 ;
  assign y17320 = n37022 ;
  assign y17321 = ~1'b0 ;
  assign y17322 = ~n37023 ;
  assign y17323 = ~1'b0 ;
  assign y17324 = ~n37025 ;
  assign y17325 = ~n37033 ;
  assign y17326 = n37035 ;
  assign y17327 = ~n37039 ;
  assign y17328 = n37041 ;
  assign y17329 = n37047 ;
  assign y17330 = ~n37048 ;
  assign y17331 = ~n37051 ;
  assign y17332 = n37061 ;
  assign y17333 = ~1'b0 ;
  assign y17334 = ~n37064 ;
  assign y17335 = n37066 ;
  assign y17336 = ~n37070 ;
  assign y17337 = ~n37071 ;
  assign y17338 = ~1'b0 ;
  assign y17339 = 1'b0 ;
  assign y17340 = ~n37073 ;
  assign y17341 = n37079 ;
  assign y17342 = n37080 ;
  assign y17343 = ~1'b0 ;
  assign y17344 = n37084 ;
  assign y17345 = ~n37085 ;
  assign y17346 = ~1'b0 ;
  assign y17347 = ~n37086 ;
  assign y17348 = n37090 ;
  assign y17349 = ~n37093 ;
  assign y17350 = ~1'b0 ;
  assign y17351 = ~1'b0 ;
  assign y17352 = n37096 ;
  assign y17353 = n37097 ;
  assign y17354 = ~n37098 ;
  assign y17355 = ~n37100 ;
  assign y17356 = n37104 ;
  assign y17357 = ~1'b0 ;
  assign y17358 = ~1'b0 ;
  assign y17359 = n37110 ;
  assign y17360 = ~1'b0 ;
  assign y17361 = n37111 ;
  assign y17362 = ~n37114 ;
  assign y17363 = n37118 ;
  assign y17364 = ~n37120 ;
  assign y17365 = ~n37124 ;
  assign y17366 = ~1'b0 ;
  assign y17367 = ~1'b0 ;
  assign y17368 = ~1'b0 ;
  assign y17369 = ~n37126 ;
  assign y17370 = ~n37128 ;
  assign y17371 = ~1'b0 ;
  assign y17372 = n37129 ;
  assign y17373 = n37131 ;
  assign y17374 = ~1'b0 ;
  assign y17375 = ~1'b0 ;
  assign y17376 = ~n37132 ;
  assign y17377 = ~1'b0 ;
  assign y17378 = n37134 ;
  assign y17379 = n37138 ;
  assign y17380 = ~n37139 ;
  assign y17381 = n37141 ;
  assign y17382 = ~1'b0 ;
  assign y17383 = ~n37145 ;
  assign y17384 = ~n37146 ;
  assign y17385 = ~1'b0 ;
  assign y17386 = ~n37147 ;
  assign y17387 = n37150 ;
  assign y17388 = ~1'b0 ;
  assign y17389 = ~1'b0 ;
  assign y17390 = ~n37154 ;
  assign y17391 = n37155 ;
  assign y17392 = n37158 ;
  assign y17393 = n37160 ;
  assign y17394 = ~1'b0 ;
  assign y17395 = ~1'b0 ;
  assign y17396 = n37161 ;
  assign y17397 = ~1'b0 ;
  assign y17398 = n37163 ;
  assign y17399 = ~n37165 ;
  assign y17400 = ~n37169 ;
  assign y17401 = n37170 ;
  assign y17402 = n37174 ;
  assign y17403 = ~n37179 ;
  assign y17404 = ~n37184 ;
  assign y17405 = n37186 ;
  assign y17406 = ~n37188 ;
  assign y17407 = n37189 ;
  assign y17408 = ~n37190 ;
  assign y17409 = n37192 ;
  assign y17410 = ~n37197 ;
  assign y17411 = ~n37201 ;
  assign y17412 = n37203 ;
  assign y17413 = n37214 ;
  assign y17414 = n37217 ;
  assign y17415 = n37218 ;
  assign y17416 = n37219 ;
  assign y17417 = 1'b0 ;
  assign y17418 = n37223 ;
  assign y17419 = ~1'b0 ;
  assign y17420 = ~n37224 ;
  assign y17421 = ~1'b0 ;
  assign y17422 = ~1'b0 ;
  assign y17423 = ~n16228 ;
  assign y17424 = ~n37226 ;
  assign y17425 = n37230 ;
  assign y17426 = n37232 ;
  assign y17427 = ~1'b0 ;
  assign y17428 = ~n32273 ;
  assign y17429 = ~1'b0 ;
  assign y17430 = n37233 ;
  assign y17431 = n37235 ;
  assign y17432 = n37236 ;
  assign y17433 = n37238 ;
  assign y17434 = n37240 ;
  assign y17435 = n37243 ;
  assign y17436 = ~1'b0 ;
  assign y17437 = n37244 ;
  assign y17438 = ~1'b0 ;
  assign y17439 = ~n37247 ;
  assign y17440 = ~1'b0 ;
  assign y17441 = n37249 ;
  assign y17442 = n37250 ;
  assign y17443 = n37251 ;
  assign y17444 = n37253 ;
  assign y17445 = ~1'b0 ;
  assign y17446 = ~n37255 ;
  assign y17447 = ~1'b0 ;
  assign y17448 = ~1'b0 ;
  assign y17449 = ~n37257 ;
  assign y17450 = ~n37261 ;
  assign y17451 = n37262 ;
  assign y17452 = ~n37263 ;
  assign y17453 = ~n37266 ;
  assign y17454 = n37267 ;
  assign y17455 = n37269 ;
  assign y17456 = n37273 ;
  assign y17457 = n37275 ;
  assign y17458 = ~1'b0 ;
  assign y17459 = n3543 ;
  assign y17460 = n37277 ;
  assign y17461 = ~n37280 ;
  assign y17462 = ~1'b0 ;
  assign y17463 = ~n8533 ;
  assign y17464 = ~1'b0 ;
  assign y17465 = ~1'b0 ;
  assign y17466 = n37282 ;
  assign y17467 = ~n37284 ;
  assign y17468 = n37285 ;
  assign y17469 = n37290 ;
  assign y17470 = n37291 ;
  assign y17471 = ~1'b0 ;
  assign y17472 = ~n37294 ;
  assign y17473 = n37298 ;
  assign y17474 = n37301 ;
  assign y17475 = ~1'b0 ;
  assign y17476 = ~n37302 ;
  assign y17477 = n1201 ;
  assign y17478 = n37307 ;
  assign y17479 = ~n37309 ;
  assign y17480 = ~n37311 ;
  assign y17481 = n37313 ;
  assign y17482 = n37314 ;
  assign y17483 = n37319 ;
  assign y17484 = n37320 ;
  assign y17485 = n37322 ;
  assign y17486 = ~n37329 ;
  assign y17487 = ~n37332 ;
  assign y17488 = ~n37333 ;
  assign y17489 = n37334 ;
  assign y17490 = n37337 ;
  assign y17491 = ~1'b0 ;
  assign y17492 = ~1'b0 ;
  assign y17493 = ~1'b0 ;
  assign y17494 = ~n37339 ;
  assign y17495 = ~1'b0 ;
  assign y17496 = n37340 ;
  assign y17497 = n37341 ;
  assign y17498 = ~n37348 ;
  assign y17499 = ~1'b0 ;
  assign y17500 = ~n15562 ;
  assign y17501 = ~1'b0 ;
  assign y17502 = ~1'b0 ;
  assign y17503 = ~n37350 ;
  assign y17504 = ~1'b0 ;
  assign y17505 = ~1'b0 ;
  assign y17506 = 1'b0 ;
  assign y17507 = ~n37351 ;
  assign y17508 = ~n37354 ;
  assign y17509 = ~n341 ;
  assign y17510 = ~n37361 ;
  assign y17511 = ~n37364 ;
  assign y17512 = n37365 ;
  assign y17513 = n37369 ;
  assign y17514 = ~1'b0 ;
  assign y17515 = ~n37371 ;
  assign y17516 = ~n37375 ;
  assign y17517 = n37376 ;
  assign y17518 = ~1'b0 ;
  assign y17519 = ~n37377 ;
  assign y17520 = ~n37378 ;
  assign y17521 = ~n37384 ;
  assign y17522 = n37386 ;
  assign y17523 = n37388 ;
  assign y17524 = ~n37389 ;
  assign y17525 = ~n37397 ;
  assign y17526 = ~n37400 ;
  assign y17527 = ~1'b0 ;
  assign y17528 = n37402 ;
  assign y17529 = ~n37405 ;
  assign y17530 = ~n37408 ;
  assign y17531 = n37410 ;
  assign y17532 = ~1'b0 ;
  assign y17533 = n37411 ;
  assign y17534 = n37413 ;
  assign y17535 = ~n37414 ;
  assign y17536 = ~1'b0 ;
  assign y17537 = n37418 ;
  assign y17538 = n4514 ;
  assign y17539 = ~n37421 ;
  assign y17540 = n37423 ;
  assign y17541 = ~n37426 ;
  assign y17542 = ~1'b0 ;
  assign y17543 = n37432 ;
  assign y17544 = ~n37433 ;
  assign y17545 = ~n37436 ;
  assign y17546 = ~n12255 ;
  assign y17547 = n37442 ;
  assign y17548 = n3926 ;
  assign y17549 = n37443 ;
  assign y17550 = ~n25718 ;
  assign y17551 = ~1'b0 ;
  assign y17552 = ~1'b0 ;
  assign y17553 = n37444 ;
  assign y17554 = ~1'b0 ;
  assign y17555 = n37446 ;
  assign y17556 = n37447 ;
  assign y17557 = ~1'b0 ;
  assign y17558 = ~1'b0 ;
  assign y17559 = ~1'b0 ;
  assign y17560 = ~n37449 ;
  assign y17561 = ~n37454 ;
  assign y17562 = n37456 ;
  assign y17563 = ~n37460 ;
  assign y17564 = n37464 ;
  assign y17565 = ~n37465 ;
  assign y17566 = ~n37467 ;
  assign y17567 = ~1'b0 ;
  assign y17568 = n37468 ;
  assign y17569 = ~n37379 ;
  assign y17570 = n37469 ;
  assign y17571 = n37471 ;
  assign y17572 = ~n37478 ;
  assign y17573 = ~n37479 ;
  assign y17574 = ~n37480 ;
  assign y17575 = ~n37484 ;
  assign y17576 = ~1'b0 ;
  assign y17577 = n37487 ;
  assign y17578 = n37488 ;
  assign y17579 = ~n37490 ;
  assign y17580 = ~n37494 ;
  assign y17581 = n37495 ;
  assign y17582 = n37496 ;
  assign y17583 = ~n37498 ;
  assign y17584 = ~n8328 ;
  assign y17585 = ~1'b0 ;
  assign y17586 = ~1'b0 ;
  assign y17587 = n37499 ;
  assign y17588 = ~n37500 ;
  assign y17589 = n37505 ;
  assign y17590 = ~1'b0 ;
  assign y17591 = ~n37506 ;
  assign y17592 = ~n37508 ;
  assign y17593 = ~1'b0 ;
  assign y17594 = ~n37511 ;
  assign y17595 = ~n37512 ;
  assign y17596 = ~1'b0 ;
  assign y17597 = ~n37513 ;
  assign y17598 = ~n37515 ;
  assign y17599 = n11221 ;
  assign y17600 = n8328 ;
  assign y17601 = ~n37518 ;
  assign y17602 = n37519 ;
  assign y17603 = ~1'b0 ;
  assign y17604 = ~n37524 ;
  assign y17605 = n37526 ;
  assign y17606 = ~n37527 ;
  assign y17607 = ~n37528 ;
  assign y17608 = ~n37531 ;
  assign y17609 = ~n37533 ;
  assign y17610 = n37540 ;
  assign y17611 = n37542 ;
  assign y17612 = ~n37544 ;
  assign y17613 = ~n37547 ;
  assign y17614 = ~n37550 ;
  assign y17615 = n37554 ;
  assign y17616 = ~n37559 ;
  assign y17617 = n37561 ;
  assign y17618 = ~1'b0 ;
  assign y17619 = ~1'b0 ;
  assign y17620 = ~n37563 ;
  assign y17621 = n37564 ;
  assign y17622 = ~n37565 ;
  assign y17623 = ~n37568 ;
  assign y17624 = ~1'b0 ;
  assign y17625 = ~1'b0 ;
  assign y17626 = n37569 ;
  assign y17627 = ~n37570 ;
  assign y17628 = ~n37576 ;
  assign y17629 = ~n1168 ;
  assign y17630 = n37577 ;
  assign y17631 = ~n37579 ;
  assign y17632 = n37585 ;
  assign y17633 = n37588 ;
  assign y17634 = n11634 ;
  assign y17635 = n37589 ;
  assign y17636 = ~n37591 ;
  assign y17637 = ~n37594 ;
  assign y17638 = n37596 ;
  assign y17639 = ~n37597 ;
  assign y17640 = n37601 ;
  assign y17641 = ~n19971 ;
  assign y17642 = n37602 ;
  assign y17643 = n37603 ;
  assign y17644 = ~1'b0 ;
  assign y17645 = ~n37604 ;
  assign y17646 = n37605 ;
  assign y17647 = n37613 ;
  assign y17648 = ~1'b0 ;
  assign y17649 = n37620 ;
  assign y17650 = ~1'b0 ;
  assign y17651 = n37630 ;
  assign y17652 = ~n37631 ;
  assign y17653 = n37634 ;
  assign y17654 = ~1'b0 ;
  assign y17655 = n37635 ;
  assign y17656 = ~n37636 ;
  assign y17657 = n37638 ;
  assign y17658 = ~n35627 ;
  assign y17659 = n37639 ;
  assign y17660 = ~1'b0 ;
  assign y17661 = ~n3633 ;
  assign y17662 = n37640 ;
  assign y17663 = ~n37641 ;
  assign y17664 = n3844 ;
  assign y17665 = n5589 ;
  assign y17666 = ~1'b0 ;
  assign y17667 = ~1'b0 ;
  assign y17668 = ~1'b0 ;
  assign y17669 = n37643 ;
  assign y17670 = n37644 ;
  assign y17671 = ~n37651 ;
  assign y17672 = ~n37654 ;
  assign y17673 = ~n37656 ;
  assign y17674 = n37658 ;
  assign y17675 = n37664 ;
  assign y17676 = n37666 ;
  assign y17677 = ~n37669 ;
  assign y17678 = n37670 ;
  assign y17679 = ~1'b0 ;
  assign y17680 = ~n29549 ;
  assign y17681 = n37674 ;
  assign y17682 = ~n37681 ;
  assign y17683 = n37686 ;
  assign y17684 = ~n20041 ;
  assign y17685 = n37692 ;
  assign y17686 = n18868 ;
  assign y17687 = 1'b0 ;
  assign y17688 = n37693 ;
  assign y17689 = 1'b0 ;
  assign y17690 = ~n37694 ;
  assign y17691 = ~1'b0 ;
  assign y17692 = ~n37697 ;
  assign y17693 = ~n37698 ;
  assign y17694 = n37700 ;
  assign y17695 = ~1'b0 ;
  assign y17696 = ~1'b0 ;
  assign y17697 = ~n37702 ;
  assign y17698 = n37703 ;
  assign y17699 = ~1'b0 ;
  assign y17700 = ~n37706 ;
  assign y17701 = ~n37708 ;
  assign y17702 = n37709 ;
  assign y17703 = ~1'b0 ;
  assign y17704 = ~n26332 ;
  assign y17705 = n37711 ;
  assign y17706 = ~n37712 ;
  assign y17707 = n37716 ;
  assign y17708 = n37723 ;
  assign y17709 = ~1'b0 ;
  assign y17710 = ~1'b0 ;
  assign y17711 = ~n37724 ;
  assign y17712 = ~n37726 ;
  assign y17713 = ~n37728 ;
  assign y17714 = ~n37730 ;
  assign y17715 = ~1'b0 ;
  assign y17716 = ~n37734 ;
  assign y17717 = ~1'b0 ;
  assign y17718 = ~n37736 ;
  assign y17719 = ~n27747 ;
  assign y17720 = ~n37737 ;
  assign y17721 = ~n37743 ;
  assign y17722 = n37744 ;
  assign y17723 = n37745 ;
  assign y17724 = ~1'b0 ;
  assign y17725 = ~1'b0 ;
  assign y17726 = ~n37750 ;
  assign y17727 = ~1'b0 ;
  assign y17728 = n37754 ;
  assign y17729 = n37758 ;
  assign y17730 = ~n37760 ;
  assign y17731 = n37763 ;
  assign y17732 = n37764 ;
  assign y17733 = ~1'b0 ;
  assign y17734 = ~n37766 ;
  assign y17735 = ~1'b0 ;
  assign y17736 = ~1'b0 ;
  assign y17737 = ~n37769 ;
  assign y17738 = ~n37771 ;
  assign y17739 = ~n37772 ;
  assign y17740 = n37778 ;
  assign y17741 = ~n37780 ;
  assign y17742 = n37781 ;
  assign y17743 = ~n37782 ;
  assign y17744 = ~n37785 ;
  assign y17745 = ~n37786 ;
  assign y17746 = ~1'b0 ;
  assign y17747 = ~1'b0 ;
  assign y17748 = ~n37787 ;
  assign y17749 = ~1'b0 ;
  assign y17750 = ~n37790 ;
  assign y17751 = n37791 ;
  assign y17752 = ~n37792 ;
  assign y17753 = n37796 ;
  assign y17754 = n37799 ;
  assign y17755 = ~1'b0 ;
  assign y17756 = ~n37801 ;
  assign y17757 = ~1'b0 ;
  assign y17758 = ~n37803 ;
  assign y17759 = ~1'b0 ;
  assign y17760 = n37804 ;
  assign y17761 = ~n37073 ;
  assign y17762 = ~1'b0 ;
  assign y17763 = n25655 ;
  assign y17764 = n37810 ;
  assign y17765 = ~n37813 ;
  assign y17766 = ~n37814 ;
  assign y17767 = ~n37815 ;
  assign y17768 = n37817 ;
  assign y17769 = n37819 ;
  assign y17770 = ~1'b0 ;
  assign y17771 = n37820 ;
  assign y17772 = n37824 ;
  assign y17773 = ~1'b0 ;
  assign y17774 = n37831 ;
  assign y17775 = ~n37832 ;
  assign y17776 = n37835 ;
  assign y17777 = n10588 ;
  assign y17778 = ~n37838 ;
  assign y17779 = ~1'b0 ;
  assign y17780 = ~1'b0 ;
  assign y17781 = n37840 ;
  assign y17782 = ~n37847 ;
  assign y17783 = n37851 ;
  assign y17784 = ~n37852 ;
  assign y17785 = n37853 ;
  assign y17786 = n37857 ;
  assign y17787 = ~n37859 ;
  assign y17788 = n37861 ;
  assign y17789 = n27390 ;
  assign y17790 = ~1'b0 ;
  assign y17791 = ~1'b0 ;
  assign y17792 = n16435 ;
  assign y17793 = ~n37865 ;
  assign y17794 = n37866 ;
  assign y17795 = ~1'b0 ;
  assign y17796 = n37868 ;
  assign y17797 = ~1'b0 ;
  assign y17798 = ~n37869 ;
  assign y17799 = n37876 ;
  assign y17800 = ~n4029 ;
  assign y17801 = ~1'b0 ;
  assign y17802 = ~n37877 ;
  assign y17803 = ~n37880 ;
  assign y17804 = n37883 ;
  assign y17805 = n37885 ;
  assign y17806 = ~1'b0 ;
  assign y17807 = n37888 ;
  assign y17808 = ~1'b0 ;
  assign y17809 = ~1'b0 ;
  assign y17810 = ~1'b0 ;
  assign y17811 = ~n37889 ;
  assign y17812 = n37894 ;
  assign y17813 = ~n37895 ;
  assign y17814 = n37896 ;
  assign y17815 = ~1'b0 ;
  assign y17816 = ~n37899 ;
  assign y17817 = ~1'b0 ;
  assign y17818 = ~n34835 ;
  assign y17819 = ~n37902 ;
  assign y17820 = ~n37903 ;
  assign y17821 = n37905 ;
  assign y17822 = ~1'b0 ;
  assign y17823 = n37910 ;
  assign y17824 = ~n37911 ;
  assign y17825 = ~n37912 ;
  assign y17826 = ~n37915 ;
  assign y17827 = ~1'b0 ;
  assign y17828 = n37918 ;
  assign y17829 = ~1'b0 ;
  assign y17830 = ~n37919 ;
  assign y17831 = ~n37921 ;
  assign y17832 = ~n37925 ;
  assign y17833 = n37926 ;
  assign y17834 = ~1'b0 ;
  assign y17835 = ~n37933 ;
  assign y17836 = ~n37935 ;
  assign y17837 = n37936 ;
  assign y17838 = n37939 ;
  assign y17839 = ~n37940 ;
  assign y17840 = ~1'b0 ;
  assign y17841 = 1'b0 ;
  assign y17842 = ~n37947 ;
  assign y17843 = n9375 ;
  assign y17844 = ~n37953 ;
  assign y17845 = n37955 ;
  assign y17846 = ~n37957 ;
  assign y17847 = ~1'b0 ;
  assign y17848 = 1'b0 ;
  assign y17849 = ~n37960 ;
  assign y17850 = n37964 ;
  assign y17851 = ~n37966 ;
  assign y17852 = n37967 ;
  assign y17853 = ~1'b0 ;
  assign y17854 = ~n37976 ;
  assign y17855 = ~n24734 ;
  assign y17856 = n37977 ;
  assign y17857 = ~n37979 ;
  assign y17858 = ~1'b0 ;
  assign y17859 = ~1'b0 ;
  assign y17860 = ~1'b0 ;
  assign y17861 = n5754 ;
  assign y17862 = n37980 ;
  assign y17863 = ~n37981 ;
  assign y17864 = ~1'b0 ;
  assign y17865 = n37982 ;
  assign y17866 = ~n37983 ;
  assign y17867 = 1'b0 ;
  assign y17868 = ~n37984 ;
  assign y17869 = ~n37985 ;
  assign y17870 = ~1'b0 ;
  assign y17871 = ~n37988 ;
  assign y17872 = n37989 ;
  assign y17873 = ~n37990 ;
  assign y17874 = ~n37992 ;
  assign y17875 = ~n37998 ;
  assign y17876 = n37999 ;
  assign y17877 = ~n29597 ;
  assign y17878 = n38002 ;
  assign y17879 = ~1'b0 ;
  assign y17880 = ~1'b0 ;
  assign y17881 = ~1'b0 ;
  assign y17882 = ~n38004 ;
  assign y17883 = n29490 ;
  assign y17884 = ~n38007 ;
  assign y17885 = n38009 ;
  assign y17886 = ~1'b0 ;
  assign y17887 = ~n38011 ;
  assign y17888 = n38012 ;
  assign y17889 = ~n38013 ;
  assign y17890 = ~1'b0 ;
  assign y17891 = n38017 ;
  assign y17892 = ~n38018 ;
  assign y17893 = ~n38021 ;
  assign y17894 = ~n38023 ;
  assign y17895 = ~n38025 ;
  assign y17896 = ~n38027 ;
  assign y17897 = ~n38028 ;
  assign y17898 = ~n38030 ;
  assign y17899 = n38032 ;
  assign y17900 = ~n38035 ;
  assign y17901 = n38036 ;
  assign y17902 = ~n38040 ;
  assign y17903 = ~n38045 ;
  assign y17904 = n38047 ;
  assign y17905 = ~1'b0 ;
  assign y17906 = n38048 ;
  assign y17907 = ~1'b0 ;
  assign y17908 = ~1'b0 ;
  assign y17909 = ~n38050 ;
  assign y17910 = ~n38051 ;
  assign y17911 = ~1'b0 ;
  assign y17912 = ~n38052 ;
  assign y17913 = ~n38057 ;
  assign y17914 = ~n18559 ;
  assign y17915 = ~n38059 ;
  assign y17916 = n38066 ;
  assign y17917 = n10289 ;
  assign y17918 = n38070 ;
  assign y17919 = n38076 ;
  assign y17920 = ~n30097 ;
  assign y17921 = ~n38077 ;
  assign y17922 = ~1'b0 ;
  assign y17923 = ~n38079 ;
  assign y17924 = ~n38083 ;
  assign y17925 = n38086 ;
  assign y17926 = n38090 ;
  assign y17927 = ~1'b0 ;
  assign y17928 = n38092 ;
  assign y17929 = ~n38094 ;
  assign y17930 = n30080 ;
  assign y17931 = n38099 ;
  assign y17932 = ~1'b0 ;
  assign y17933 = n38100 ;
  assign y17934 = 1'b0 ;
  assign y17935 = ~1'b0 ;
  assign y17936 = ~n38105 ;
  assign y17937 = ~n38106 ;
  assign y17938 = ~n38108 ;
  assign y17939 = ~n38114 ;
  assign y17940 = ~1'b0 ;
  assign y17941 = ~n38115 ;
  assign y17942 = ~n38118 ;
  assign y17943 = n38119 ;
  assign y17944 = ~1'b0 ;
  assign y17945 = ~1'b0 ;
  assign y17946 = n38120 ;
  assign y17947 = ~n38122 ;
  assign y17948 = n38123 ;
  assign y17949 = n38124 ;
  assign y17950 = n38125 ;
  assign y17951 = ~1'b0 ;
  assign y17952 = ~1'b0 ;
  assign y17953 = ~1'b0 ;
  assign y17954 = 1'b0 ;
  assign y17955 = ~1'b0 ;
  assign y17956 = n38126 ;
  assign y17957 = n4241 ;
  assign y17958 = ~n38127 ;
  assign y17959 = ~1'b0 ;
  assign y17960 = ~n38130 ;
  assign y17961 = n38133 ;
  assign y17962 = n38138 ;
  assign y17963 = n38139 ;
  assign y17964 = n38142 ;
  assign y17965 = ~1'b0 ;
  assign y17966 = ~n38144 ;
  assign y17967 = ~n38147 ;
  assign y17968 = ~n38148 ;
  assign y17969 = ~1'b0 ;
  assign y17970 = ~n38149 ;
  assign y17971 = ~1'b0 ;
  assign y17972 = n38151 ;
  assign y17973 = ~1'b0 ;
  assign y17974 = n38154 ;
  assign y17975 = ~1'b0 ;
  assign y17976 = n38155 ;
  assign y17977 = n38156 ;
  assign y17978 = n38160 ;
  assign y17979 = n38161 ;
  assign y17980 = n38164 ;
  assign y17981 = ~1'b0 ;
  assign y17982 = ~1'b0 ;
  assign y17983 = n38168 ;
  assign y17984 = ~n38172 ;
  assign y17985 = ~n38175 ;
  assign y17986 = ~n38176 ;
  assign y17987 = ~n38178 ;
  assign y17988 = ~n38180 ;
  assign y17989 = ~n38186 ;
  assign y17990 = ~n18479 ;
  assign y17991 = ~1'b0 ;
  assign y17992 = ~1'b0 ;
  assign y17993 = ~n38189 ;
  assign y17994 = ~n38193 ;
  assign y17995 = ~n38195 ;
  assign y17996 = ~1'b0 ;
  assign y17997 = ~1'b0 ;
  assign y17998 = n38198 ;
  assign y17999 = ~n38201 ;
  assign y18000 = ~1'b0 ;
  assign y18001 = ~n38204 ;
  assign y18002 = ~1'b0 ;
  assign y18003 = n38205 ;
  assign y18004 = n38206 ;
  assign y18005 = ~n38207 ;
  assign y18006 = ~n7457 ;
  assign y18007 = n22995 ;
  assign y18008 = n38208 ;
  assign y18009 = n38213 ;
  assign y18010 = n38218 ;
  assign y18011 = ~n38224 ;
  assign y18012 = ~n38225 ;
  assign y18013 = ~n38228 ;
  assign y18014 = n38231 ;
  assign y18015 = ~n38233 ;
  assign y18016 = ~1'b0 ;
  assign y18017 = ~1'b0 ;
  assign y18018 = ~1'b0 ;
  assign y18019 = ~n38235 ;
  assign y18020 = n38237 ;
  assign y18021 = ~1'b0 ;
  assign y18022 = ~n38239 ;
  assign y18023 = ~n38158 ;
  assign y18024 = n38240 ;
  assign y18025 = ~n38242 ;
  assign y18026 = ~1'b0 ;
  assign y18027 = ~n24035 ;
  assign y18028 = ~n20722 ;
  assign y18029 = ~1'b0 ;
  assign y18030 = n10348 ;
  assign y18031 = n7154 ;
  assign y18032 = ~n38245 ;
  assign y18033 = ~1'b0 ;
  assign y18034 = n38246 ;
  assign y18035 = n38247 ;
  assign y18036 = ~1'b0 ;
  assign y18037 = n38248 ;
  assign y18038 = ~n38259 ;
  assign y18039 = n38261 ;
  assign y18040 = ~n38263 ;
  assign y18041 = n38264 ;
  assign y18042 = ~1'b0 ;
  assign y18043 = n38265 ;
  assign y18044 = ~n38269 ;
  assign y18045 = n38270 ;
  assign y18046 = n38271 ;
  assign y18047 = n38272 ;
  assign y18048 = ~n38274 ;
  assign y18049 = n38275 ;
  assign y18050 = n38277 ;
  assign y18051 = ~n38280 ;
  assign y18052 = n38282 ;
  assign y18053 = ~1'b0 ;
  assign y18054 = ~n38286 ;
  assign y18055 = n38287 ;
  assign y18056 = ~n38290 ;
  assign y18057 = ~n38293 ;
  assign y18058 = ~n38294 ;
  assign y18059 = ~1'b0 ;
  assign y18060 = n38296 ;
  assign y18061 = ~n38298 ;
  assign y18062 = ~n38304 ;
  assign y18063 = n9962 ;
  assign y18064 = ~n38305 ;
  assign y18065 = ~n38309 ;
  assign y18066 = n38311 ;
  assign y18067 = ~1'b0 ;
  assign y18068 = n38312 ;
  assign y18069 = n38315 ;
  assign y18070 = n38318 ;
  assign y18071 = n38320 ;
  assign y18072 = n38322 ;
  assign y18073 = ~n38325 ;
  assign y18074 = n38326 ;
  assign y18075 = ~n38333 ;
  assign y18076 = ~1'b0 ;
  assign y18077 = ~1'b0 ;
  assign y18078 = ~1'b0 ;
  assign y18079 = ~n38336 ;
  assign y18080 = ~n38338 ;
  assign y18081 = ~n38343 ;
  assign y18082 = ~1'b0 ;
  assign y18083 = ~n38347 ;
  assign y18084 = n38349 ;
  assign y18085 = n38351 ;
  assign y18086 = n38353 ;
  assign y18087 = ~1'b0 ;
  assign y18088 = n38354 ;
  assign y18089 = ~1'b0 ;
  assign y18090 = ~1'b0 ;
  assign y18091 = n38356 ;
  assign y18092 = ~n38357 ;
  assign y18093 = n38366 ;
  assign y18094 = n38367 ;
  assign y18095 = ~n38368 ;
  assign y18096 = ~n38371 ;
  assign y18097 = n38373 ;
  assign y18098 = n38374 ;
  assign y18099 = ~1'b0 ;
  assign y18100 = ~1'b0 ;
  assign y18101 = n38377 ;
  assign y18102 = n38379 ;
  assign y18103 = n38381 ;
  assign y18104 = n38384 ;
  assign y18105 = ~n38386 ;
  assign y18106 = n38387 ;
  assign y18107 = ~n38389 ;
  assign y18108 = n38392 ;
  assign y18109 = ~n38396 ;
  assign y18110 = n35845 ;
  assign y18111 = n38397 ;
  assign y18112 = ~n11249 ;
  assign y18113 = n38399 ;
  assign y18114 = ~1'b0 ;
  assign y18115 = ~n33097 ;
  assign y18116 = n38401 ;
  assign y18117 = ~n38403 ;
  assign y18118 = ~1'b0 ;
  assign y18119 = ~n38405 ;
  assign y18120 = ~n38406 ;
  assign y18121 = n38411 ;
  assign y18122 = n38413 ;
  assign y18123 = n17811 ;
  assign y18124 = ~n38420 ;
  assign y18125 = n38424 ;
  assign y18126 = ~1'b0 ;
  assign y18127 = ~1'b0 ;
  assign y18128 = 1'b0 ;
  assign y18129 = n38429 ;
  assign y18130 = ~1'b0 ;
  assign y18131 = n38430 ;
  assign y18132 = n38431 ;
  assign y18133 = ~1'b0 ;
  assign y18134 = ~1'b0 ;
  assign y18135 = ~1'b0 ;
  assign y18136 = ~1'b0 ;
  assign y18137 = n38432 ;
  assign y18138 = n38435 ;
  assign y18139 = ~n38437 ;
  assign y18140 = ~n38448 ;
  assign y18141 = n38450 ;
  assign y18142 = ~1'b0 ;
  assign y18143 = ~n38452 ;
  assign y18144 = ~n38457 ;
  assign y18145 = n38460 ;
  assign y18146 = n38464 ;
  assign y18147 = n38465 ;
  assign y18148 = ~n38466 ;
  assign y18149 = ~n38467 ;
  assign y18150 = ~n38469 ;
  assign y18151 = n38470 ;
  assign y18152 = ~n38476 ;
  assign y18153 = ~1'b0 ;
  assign y18154 = ~n38477 ;
  assign y18155 = n38481 ;
  assign y18156 = n38486 ;
  assign y18157 = ~n38493 ;
  assign y18158 = n38494 ;
  assign y18159 = n38495 ;
  assign y18160 = n38496 ;
  assign y18161 = ~n38498 ;
  assign y18162 = ~n38501 ;
  assign y18163 = ~n38508 ;
  assign y18164 = ~n38510 ;
  assign y18165 = n23471 ;
  assign y18166 = ~n38511 ;
  assign y18167 = n38512 ;
  assign y18168 = ~n38513 ;
  assign y18169 = ~n38514 ;
  assign y18170 = n38515 ;
  assign y18171 = ~n34778 ;
  assign y18172 = n38516 ;
  assign y18173 = ~1'b0 ;
  assign y18174 = n38517 ;
  assign y18175 = n38518 ;
  assign y18176 = ~1'b0 ;
  assign y18177 = n38520 ;
  assign y18178 = n20550 ;
  assign y18179 = ~n38523 ;
  assign y18180 = ~1'b0 ;
  assign y18181 = ~n38524 ;
  assign y18182 = ~n38526 ;
  assign y18183 = n38528 ;
  assign y18184 = n38529 ;
  assign y18185 = n38535 ;
  assign y18186 = n38537 ;
  assign y18187 = n38539 ;
  assign y18188 = n38541 ;
  assign y18189 = ~n38542 ;
  assign y18190 = ~n38544 ;
  assign y18191 = ~1'b0 ;
  assign y18192 = n38545 ;
  assign y18193 = n38548 ;
  assign y18194 = ~n38550 ;
  assign y18195 = n38551 ;
  assign y18196 = ~n38554 ;
  assign y18197 = ~1'b0 ;
  assign y18198 = n38555 ;
  assign y18199 = n38556 ;
  assign y18200 = ~n38560 ;
  assign y18201 = n38561 ;
  assign y18202 = ~n38563 ;
  assign y18203 = ~1'b0 ;
  assign y18204 = n38568 ;
  assign y18205 = n38571 ;
  assign y18206 = ~1'b0 ;
  assign y18207 = n38573 ;
  assign y18208 = n38575 ;
  assign y18209 = ~n30080 ;
  assign y18210 = ~n38577 ;
  assign y18211 = n38580 ;
  assign y18212 = ~1'b0 ;
  assign y18213 = n38583 ;
  assign y18214 = n38585 ;
  assign y18215 = ~n38586 ;
  assign y18216 = n38587 ;
  assign y18217 = ~n38588 ;
  assign y18218 = ~n38590 ;
  assign y18219 = ~n38594 ;
  assign y18220 = n38595 ;
  assign y18221 = ~n38597 ;
  assign y18222 = ~1'b0 ;
  assign y18223 = n38600 ;
  assign y18224 = n38601 ;
  assign y18225 = n38603 ;
  assign y18226 = ~n38604 ;
  assign y18227 = ~1'b0 ;
  assign y18228 = ~n38608 ;
  assign y18229 = ~1'b0 ;
  assign y18230 = ~n38610 ;
  assign y18231 = ~1'b0 ;
  assign y18232 = ~n38611 ;
  assign y18233 = n38616 ;
  assign y18234 = n38618 ;
  assign y18235 = ~n38619 ;
  assign y18236 = n38621 ;
  assign y18237 = n38622 ;
  assign y18238 = ~n38624 ;
  assign y18239 = ~n8041 ;
  assign y18240 = ~n38631 ;
  assign y18241 = ~n38633 ;
  assign y18242 = n38637 ;
  assign y18243 = n38638 ;
  assign y18244 = ~n38639 ;
  assign y18245 = n38641 ;
  assign y18246 = ~n38642 ;
  assign y18247 = ~n38646 ;
  assign y18248 = ~1'b0 ;
  assign y18249 = n38648 ;
  assign y18250 = n12197 ;
  assign y18251 = ~1'b0 ;
  assign y18252 = ~n38651 ;
  assign y18253 = n38655 ;
  assign y18254 = n38658 ;
  assign y18255 = ~n38663 ;
  assign y18256 = ~1'b0 ;
  assign y18257 = ~1'b0 ;
  assign y18258 = n38664 ;
  assign y18259 = n38666 ;
  assign y18260 = ~1'b0 ;
  assign y18261 = ~n38668 ;
  assign y18262 = ~n38675 ;
  assign y18263 = n2442 ;
  assign y18264 = ~1'b0 ;
  assign y18265 = ~n38676 ;
  assign y18266 = n38677 ;
  assign y18267 = ~1'b0 ;
  assign y18268 = 1'b0 ;
  assign y18269 = ~n38680 ;
  assign y18270 = ~1'b0 ;
  assign y18271 = n38681 ;
  assign y18272 = n38682 ;
  assign y18273 = ~n38687 ;
  assign y18274 = ~n38688 ;
  assign y18275 = ~1'b0 ;
  assign y18276 = n38690 ;
  assign y18277 = n38691 ;
  assign y18278 = ~1'b0 ;
  assign y18279 = ~1'b0 ;
  assign y18280 = ~n38694 ;
  assign y18281 = n38699 ;
  assign y18282 = ~1'b0 ;
  assign y18283 = ~n38702 ;
  assign y18284 = n34645 ;
  assign y18285 = n38705 ;
  assign y18286 = n38706 ;
  assign y18287 = ~n38713 ;
  assign y18288 = ~1'b0 ;
  assign y18289 = ~n38714 ;
  assign y18290 = ~n38715 ;
  assign y18291 = ~1'b0 ;
  assign y18292 = n35122 ;
  assign y18293 = ~n38716 ;
  assign y18294 = n38717 ;
  assign y18295 = n38718 ;
  assign y18296 = ~1'b0 ;
  assign y18297 = n38719 ;
  assign y18298 = ~n38720 ;
  assign y18299 = ~1'b0 ;
  assign y18300 = n38723 ;
  assign y18301 = n38729 ;
  assign y18302 = n4016 ;
  assign y18303 = ~n38730 ;
  assign y18304 = ~1'b0 ;
  assign y18305 = ~1'b0 ;
  assign y18306 = ~1'b0 ;
  assign y18307 = ~n38731 ;
  assign y18308 = n27138 ;
  assign y18309 = n38732 ;
  assign y18310 = ~n38733 ;
  assign y18311 = ~n38735 ;
  assign y18312 = ~1'b0 ;
  assign y18313 = ~n38739 ;
  assign y18314 = n38745 ;
  assign y18315 = ~1'b0 ;
  assign y18316 = ~1'b0 ;
  assign y18317 = n38746 ;
  assign y18318 = n38748 ;
  assign y18319 = n38750 ;
  assign y18320 = ~n38753 ;
  assign y18321 = n38754 ;
  assign y18322 = n38756 ;
  assign y18323 = ~1'b0 ;
  assign y18324 = n38757 ;
  assign y18325 = ~1'b0 ;
  assign y18326 = ~n38762 ;
  assign y18327 = ~n38765 ;
  assign y18328 = ~n38766 ;
  assign y18329 = ~n38769 ;
  assign y18330 = 1'b0 ;
  assign y18331 = n38771 ;
  assign y18332 = n38772 ;
  assign y18333 = n38773 ;
  assign y18334 = n38777 ;
  assign y18335 = n38779 ;
  assign y18336 = ~n38781 ;
  assign y18337 = ~1'b0 ;
  assign y18338 = ~n38788 ;
  assign y18339 = n38792 ;
  assign y18340 = ~n38796 ;
  assign y18341 = ~1'b0 ;
  assign y18342 = ~1'b0 ;
  assign y18343 = n38797 ;
  assign y18344 = ~n38801 ;
  assign y18345 = n38803 ;
  assign y18346 = ~1'b0 ;
  assign y18347 = ~1'b0 ;
  assign y18348 = n38805 ;
  assign y18349 = ~1'b0 ;
  assign y18350 = ~1'b0 ;
  assign y18351 = n38807 ;
  assign y18352 = n9435 ;
  assign y18353 = n38808 ;
  assign y18354 = n38809 ;
  assign y18355 = n38811 ;
  assign y18356 = n38813 ;
  assign y18357 = ~1'b0 ;
  assign y18358 = n38814 ;
  assign y18359 = ~1'b0 ;
  assign y18360 = n38818 ;
  assign y18361 = ~n38819 ;
  assign y18362 = ~n38821 ;
  assign y18363 = n38824 ;
  assign y18364 = n38826 ;
  assign y18365 = ~n38827 ;
  assign y18366 = ~1'b0 ;
  assign y18367 = ~n38830 ;
  assign y18368 = ~n38836 ;
  assign y18369 = ~n38838 ;
  assign y18370 = ~n12031 ;
  assign y18371 = n38839 ;
  assign y18372 = ~n27181 ;
  assign y18373 = n38841 ;
  assign y18374 = n38851 ;
  assign y18375 = n38856 ;
  assign y18376 = ~1'b0 ;
  assign y18377 = ~1'b0 ;
  assign y18378 = n38857 ;
  assign y18379 = n19941 ;
  assign y18380 = n38859 ;
  assign y18381 = ~1'b0 ;
  assign y18382 = ~1'b0 ;
  assign y18383 = ~1'b0 ;
  assign y18384 = ~n38861 ;
  assign y18385 = ~n38863 ;
  assign y18386 = ~1'b0 ;
  assign y18387 = ~1'b0 ;
  assign y18388 = n38866 ;
  assign y18389 = n38872 ;
  assign y18390 = ~n38874 ;
  assign y18391 = n38876 ;
  assign y18392 = ~1'b0 ;
  assign y18393 = ~n38880 ;
  assign y18394 = n38883 ;
  assign y18395 = n38887 ;
  assign y18396 = ~1'b0 ;
  assign y18397 = n38889 ;
  assign y18398 = n38890 ;
  assign y18399 = n38891 ;
  assign y18400 = n38900 ;
  assign y18401 = n38905 ;
  assign y18402 = ~1'b0 ;
  assign y18403 = ~1'b0 ;
  assign y18404 = ~n38907 ;
  assign y18405 = ~1'b0 ;
  assign y18406 = n38909 ;
  assign y18407 = ~n38910 ;
  assign y18408 = n38920 ;
  assign y18409 = n38921 ;
  assign y18410 = n38924 ;
  assign y18411 = ~n38928 ;
  assign y18412 = n38929 ;
  assign y18413 = ~1'b0 ;
  assign y18414 = ~n38933 ;
  assign y18415 = n38938 ;
  assign y18416 = n38943 ;
  assign y18417 = ~n38944 ;
  assign y18418 = ~n38945 ;
  assign y18419 = ~n38949 ;
  assign y18420 = ~1'b0 ;
  assign y18421 = ~1'b0 ;
  assign y18422 = ~n38951 ;
  assign y18423 = n38952 ;
  assign y18424 = ~1'b0 ;
  assign y18425 = ~n38963 ;
  assign y18426 = ~n38970 ;
  assign y18427 = n38971 ;
  assign y18428 = n38972 ;
  assign y18429 = n38974 ;
  assign y18430 = n38975 ;
  assign y18431 = n38978 ;
  assign y18432 = ~n38983 ;
  assign y18433 = ~n38986 ;
  assign y18434 = ~n38988 ;
  assign y18435 = n38992 ;
  assign y18436 = ~n38996 ;
  assign y18437 = ~n16539 ;
  assign y18438 = ~n38997 ;
  assign y18439 = ~n39002 ;
  assign y18440 = ~n39003 ;
  assign y18441 = ~n39005 ;
  assign y18442 = ~1'b0 ;
  assign y18443 = ~n39006 ;
  assign y18444 = ~1'b0 ;
  assign y18445 = ~n39007 ;
  assign y18446 = ~n39008 ;
  assign y18447 = n39010 ;
  assign y18448 = ~1'b0 ;
  assign y18449 = ~n39012 ;
  assign y18450 = n39017 ;
  assign y18451 = ~1'b0 ;
  assign y18452 = ~n39024 ;
  assign y18453 = n39028 ;
  assign y18454 = ~1'b0 ;
  assign y18455 = ~n39029 ;
  assign y18456 = ~n39033 ;
  assign y18457 = n39034 ;
  assign y18458 = ~n39038 ;
  assign y18459 = n39039 ;
  assign y18460 = ~n39042 ;
  assign y18461 = ~1'b0 ;
  assign y18462 = ~n39043 ;
  assign y18463 = n39045 ;
  assign y18464 = ~1'b0 ;
  assign y18465 = n39046 ;
  assign y18466 = ~1'b0 ;
  assign y18467 = ~n39047 ;
  assign y18468 = ~n39048 ;
  assign y18469 = ~1'b0 ;
  assign y18470 = ~1'b0 ;
  assign y18471 = ~n39051 ;
  assign y18472 = ~n39058 ;
  assign y18473 = ~1'b0 ;
  assign y18474 = n39060 ;
  assign y18475 = ~n39061 ;
  assign y18476 = n39064 ;
  assign y18477 = ~n16515 ;
  assign y18478 = ~n39071 ;
  assign y18479 = ~n39075 ;
  assign y18480 = n39077 ;
  assign y18481 = ~1'b0 ;
  assign y18482 = ~1'b0 ;
  assign y18483 = n39078 ;
  assign y18484 = n39079 ;
  assign y18485 = n39080 ;
  assign y18486 = n39083 ;
  assign y18487 = n39085 ;
  assign y18488 = ~n39087 ;
  assign y18489 = ~1'b0 ;
  assign y18490 = ~1'b0 ;
  assign y18491 = ~n39089 ;
  assign y18492 = ~1'b0 ;
  assign y18493 = n6907 ;
  assign y18494 = n39090 ;
  assign y18495 = ~n39094 ;
  assign y18496 = ~1'b0 ;
  assign y18497 = ~n39095 ;
  assign y18498 = ~n39098 ;
  assign y18499 = ~1'b0 ;
  assign y18500 = n39101 ;
  assign y18501 = n39102 ;
  assign y18502 = ~n39105 ;
  assign y18503 = n39107 ;
  assign y18504 = n39109 ;
  assign y18505 = n39111 ;
  assign y18506 = ~1'b0 ;
  assign y18507 = ~1'b0 ;
  assign y18508 = n28291 ;
  assign y18509 = ~n22814 ;
  assign y18510 = ~n6232 ;
  assign y18511 = n39112 ;
  assign y18512 = ~n39113 ;
  assign y18513 = ~n39115 ;
  assign y18514 = ~n39118 ;
  assign y18515 = ~n39119 ;
  assign y18516 = ~1'b0 ;
  assign y18517 = ~n39120 ;
  assign y18518 = ~n39122 ;
  assign y18519 = ~n39123 ;
  assign y18520 = ~1'b0 ;
  assign y18521 = ~n39128 ;
  assign y18522 = ~n39131 ;
  assign y18523 = n39133 ;
  assign y18524 = ~1'b0 ;
  assign y18525 = ~1'b0 ;
  assign y18526 = n39140 ;
  assign y18527 = ~1'b0 ;
  assign y18528 = n39146 ;
  assign y18529 = ~1'b0 ;
  assign y18530 = ~1'b0 ;
  assign y18531 = ~n39147 ;
  assign y18532 = n39151 ;
  assign y18533 = ~n39155 ;
  assign y18534 = n39158 ;
  assign y18535 = ~1'b0 ;
  assign y18536 = ~n39160 ;
  assign y18537 = ~1'b0 ;
  assign y18538 = 1'b0 ;
  assign y18539 = ~1'b0 ;
  assign y18540 = n39161 ;
  assign y18541 = ~n39163 ;
  assign y18542 = ~n39165 ;
  assign y18543 = n1223 ;
  assign y18544 = n39167 ;
  assign y18545 = ~n39169 ;
  assign y18546 = ~1'b0 ;
  assign y18547 = n39171 ;
  assign y18548 = ~n39181 ;
  assign y18549 = ~n39184 ;
  assign y18550 = ~n39190 ;
  assign y18551 = ~n39193 ;
  assign y18552 = ~1'b0 ;
  assign y18553 = ~n39194 ;
  assign y18554 = ~1'b0 ;
  assign y18555 = ~n39196 ;
  assign y18556 = ~n39199 ;
  assign y18557 = ~n39204 ;
  assign y18558 = n39205 ;
  assign y18559 = ~n39207 ;
  assign y18560 = ~n39209 ;
  assign y18561 = ~n39210 ;
  assign y18562 = n39213 ;
  assign y18563 = ~1'b0 ;
  assign y18564 = ~n39215 ;
  assign y18565 = n23253 ;
  assign y18566 = ~1'b0 ;
  assign y18567 = ~n39222 ;
  assign y18568 = ~n39223 ;
  assign y18569 = ~n39224 ;
  assign y18570 = ~n39228 ;
  assign y18571 = ~n39233 ;
  assign y18572 = ~n39235 ;
  assign y18573 = n39237 ;
  assign y18574 = ~n39239 ;
  assign y18575 = ~1'b0 ;
  assign y18576 = n39241 ;
  assign y18577 = ~n39242 ;
  assign y18578 = n39245 ;
  assign y18579 = n39248 ;
  assign y18580 = ~1'b0 ;
  assign y18581 = ~1'b0 ;
  assign y18582 = ~1'b0 ;
  assign y18583 = n39250 ;
  assign y18584 = n39253 ;
  assign y18585 = ~1'b0 ;
  assign y18586 = n39254 ;
  assign y18587 = 1'b0 ;
  assign y18588 = 1'b0 ;
  assign y18589 = ~n39256 ;
  assign y18590 = ~1'b0 ;
  assign y18591 = n39259 ;
  assign y18592 = ~1'b0 ;
  assign y18593 = ~1'b0 ;
  assign y18594 = ~n39261 ;
  assign y18595 = ~n39262 ;
  assign y18596 = ~1'b0 ;
  assign y18597 = n39265 ;
  assign y18598 = n39270 ;
  assign y18599 = n39271 ;
  assign y18600 = n39272 ;
  assign y18601 = n39273 ;
  assign y18602 = ~1'b0 ;
  assign y18603 = ~n1703 ;
  assign y18604 = ~1'b0 ;
  assign y18605 = n39276 ;
  assign y18606 = n39279 ;
  assign y18607 = n39283 ;
  assign y18608 = n39285 ;
  assign y18609 = ~n39286 ;
  assign y18610 = n39288 ;
  assign y18611 = ~1'b0 ;
  assign y18612 = ~n39291 ;
  assign y18613 = n39292 ;
  assign y18614 = n39294 ;
  assign y18615 = ~1'b0 ;
  assign y18616 = n39295 ;
  assign y18617 = ~1'b0 ;
  assign y18618 = n39296 ;
  assign y18619 = ~n39298 ;
  assign y18620 = ~1'b0 ;
  assign y18621 = n39305 ;
  assign y18622 = ~n39312 ;
  assign y18623 = n39313 ;
  assign y18624 = ~1'b0 ;
  assign y18625 = ~1'b0 ;
  assign y18626 = n39314 ;
  assign y18627 = n39316 ;
  assign y18628 = n39318 ;
  assign y18629 = ~n39319 ;
  assign y18630 = ~n39328 ;
  assign y18631 = ~1'b0 ;
  assign y18632 = ~n39329 ;
  assign y18633 = n39331 ;
  assign y18634 = ~1'b0 ;
  assign y18635 = n39333 ;
  assign y18636 = ~n39335 ;
  assign y18637 = n39336 ;
  assign y18638 = 1'b0 ;
  assign y18639 = ~n39337 ;
  assign y18640 = n39341 ;
  assign y18641 = ~1'b0 ;
  assign y18642 = n39342 ;
  assign y18643 = n24348 ;
  assign y18644 = ~1'b0 ;
  assign y18645 = ~1'b0 ;
  assign y18646 = n39343 ;
  assign y18647 = n39347 ;
  assign y18648 = n39353 ;
  assign y18649 = ~1'b0 ;
  assign y18650 = ~1'b0 ;
  assign y18651 = n39355 ;
  assign y18652 = ~1'b0 ;
  assign y18653 = ~n39356 ;
  assign y18654 = n39359 ;
  assign y18655 = ~n39360 ;
  assign y18656 = ~n17233 ;
  assign y18657 = n39367 ;
  assign y18658 = n39370 ;
  assign y18659 = n39372 ;
  assign y18660 = ~1'b0 ;
  assign y18661 = ~1'b0 ;
  assign y18662 = n39374 ;
  assign y18663 = ~n39375 ;
  assign y18664 = ~n39377 ;
  assign y18665 = n21784 ;
  assign y18666 = ~1'b0 ;
  assign y18667 = n39379 ;
  assign y18668 = ~1'b0 ;
  assign y18669 = ~1'b0 ;
  assign y18670 = ~n39386 ;
  assign y18671 = ~n39388 ;
  assign y18672 = n39391 ;
  assign y18673 = ~n39392 ;
  assign y18674 = ~1'b0 ;
  assign y18675 = ~n39396 ;
  assign y18676 = ~n39397 ;
  assign y18677 = n6429 ;
  assign y18678 = ~n39404 ;
  assign y18679 = ~n39410 ;
  assign y18680 = n39415 ;
  assign y18681 = n39418 ;
  assign y18682 = n39420 ;
  assign y18683 = n39428 ;
  assign y18684 = n26588 ;
  assign y18685 = ~1'b0 ;
  assign y18686 = n39430 ;
  assign y18687 = ~n39432 ;
  assign y18688 = ~n39434 ;
  assign y18689 = ~n39436 ;
  assign y18690 = ~n39441 ;
  assign y18691 = ~n39448 ;
  assign y18692 = ~n30208 ;
  assign y18693 = ~n26120 ;
  assign y18694 = ~1'b0 ;
  assign y18695 = ~1'b0 ;
  assign y18696 = ~1'b0 ;
  assign y18697 = ~n39449 ;
  assign y18698 = ~n39450 ;
  assign y18699 = n39451 ;
  assign y18700 = n39456 ;
  assign y18701 = n39458 ;
  assign y18702 = ~1'b0 ;
  assign y18703 = ~n39461 ;
  assign y18704 = n39466 ;
  assign y18705 = ~n39467 ;
  assign y18706 = ~n39470 ;
  assign y18707 = ~1'b0 ;
  assign y18708 = n39472 ;
  assign y18709 = n36185 ;
  assign y18710 = ~n39474 ;
  assign y18711 = n39476 ;
  assign y18712 = ~n39479 ;
  assign y18713 = n23094 ;
  assign y18714 = ~n39481 ;
  assign y18715 = ~1'b0 ;
  assign y18716 = ~1'b0 ;
  assign y18717 = ~1'b0 ;
  assign y18718 = ~n39483 ;
  assign y18719 = ~1'b0 ;
  assign y18720 = ~n39486 ;
  assign y18721 = 1'b0 ;
  assign y18722 = n39488 ;
  assign y18723 = n39490 ;
  assign y18724 = n39495 ;
  assign y18725 = ~n39500 ;
  assign y18726 = ~1'b0 ;
  assign y18727 = ~1'b0 ;
  assign y18728 = ~n39504 ;
  assign y18729 = ~n39505 ;
  assign y18730 = n39506 ;
  assign y18731 = ~n39509 ;
  assign y18732 = n39512 ;
  assign y18733 = ~n39515 ;
  assign y18734 = n39519 ;
  assign y18735 = n39520 ;
  assign y18736 = ~n39522 ;
  assign y18737 = n39523 ;
  assign y18738 = ~1'b0 ;
  assign y18739 = ~1'b0 ;
  assign y18740 = ~1'b0 ;
  assign y18741 = n39531 ;
  assign y18742 = ~n39533 ;
  assign y18743 = n39534 ;
  assign y18744 = ~n39540 ;
  assign y18745 = n39544 ;
  assign y18746 = ~1'b0 ;
  assign y18747 = ~1'b0 ;
  assign y18748 = ~1'b0 ;
  assign y18749 = ~1'b0 ;
  assign y18750 = ~1'b0 ;
  assign y18751 = ~1'b0 ;
  assign y18752 = ~1'b0 ;
  assign y18753 = n39545 ;
  assign y18754 = ~n39546 ;
  assign y18755 = n39548 ;
  assign y18756 = n39550 ;
  assign y18757 = ~1'b0 ;
  assign y18758 = 1'b0 ;
  assign y18759 = ~n3630 ;
  assign y18760 = ~n39554 ;
  assign y18761 = ~n39556 ;
  assign y18762 = ~n39560 ;
  assign y18763 = n39568 ;
  assign y18764 = ~1'b0 ;
  assign y18765 = n39573 ;
  assign y18766 = ~1'b0 ;
  assign y18767 = n39580 ;
  assign y18768 = n37800 ;
  assign y18769 = ~1'b0 ;
  assign y18770 = ~n39582 ;
  assign y18771 = ~n39586 ;
  assign y18772 = n39587 ;
  assign y18773 = ~n39588 ;
  assign y18774 = ~n39590 ;
  assign y18775 = n39591 ;
  assign y18776 = ~1'b0 ;
  assign y18777 = ~1'b0 ;
  assign y18778 = n21326 ;
  assign y18779 = ~n39593 ;
  assign y18780 = n39594 ;
  assign y18781 = ~n39595 ;
  assign y18782 = n39596 ;
  assign y18783 = ~n39598 ;
  assign y18784 = n39599 ;
  assign y18785 = n39600 ;
  assign y18786 = ~1'b0 ;
  assign y18787 = ~n39601 ;
  assign y18788 = ~n39607 ;
  assign y18789 = n39608 ;
  assign y18790 = n39610 ;
  assign y18791 = n39611 ;
  assign y18792 = n39612 ;
  assign y18793 = n39616 ;
  assign y18794 = ~n39617 ;
  assign y18795 = n39620 ;
  assign y18796 = ~n39621 ;
  assign y18797 = ~n39624 ;
  assign y18798 = ~n12341 ;
  assign y18799 = n39625 ;
  assign y18800 = ~n39628 ;
  assign y18801 = n36817 ;
  assign y18802 = ~1'b0 ;
  assign y18803 = 1'b0 ;
  assign y18804 = ~n39630 ;
  assign y18805 = n39635 ;
  assign y18806 = n39636 ;
  assign y18807 = n39640 ;
  assign y18808 = ~1'b0 ;
  assign y18809 = n39641 ;
  assign y18810 = ~n39645 ;
  assign y18811 = n39647 ;
  assign y18812 = ~n39652 ;
  assign y18813 = n39658 ;
  assign y18814 = ~1'b0 ;
  assign y18815 = ~1'b0 ;
  assign y18816 = n39659 ;
  assign y18817 = n39660 ;
  assign y18818 = ~n39667 ;
  assign y18819 = ~n39671 ;
  assign y18820 = ~1'b0 ;
  assign y18821 = n39694 ;
  assign y18822 = n39698 ;
  assign y18823 = ~n39699 ;
  assign y18824 = ~n39701 ;
  assign y18825 = ~n11667 ;
  assign y18826 = ~1'b0 ;
  assign y18827 = ~n39707 ;
  assign y18828 = n39708 ;
  assign y18829 = n19863 ;
  assign y18830 = n39710 ;
  assign y18831 = ~n39714 ;
  assign y18832 = n39717 ;
  assign y18833 = ~n39721 ;
  assign y18834 = ~n39725 ;
  assign y18835 = n39727 ;
  assign y18836 = ~1'b0 ;
  assign y18837 = n39729 ;
  assign y18838 = ~n39731 ;
  assign y18839 = ~n1440 ;
  assign y18840 = n39732 ;
  assign y18841 = n39736 ;
  assign y18842 = n39738 ;
  assign y18843 = ~1'b0 ;
  assign y18844 = n39739 ;
  assign y18845 = ~1'b0 ;
  assign y18846 = n39741 ;
  assign y18847 = ~n39744 ;
  assign y18848 = n39747 ;
  assign y18849 = ~n39753 ;
  assign y18850 = n39755 ;
  assign y18851 = n39757 ;
  assign y18852 = n39763 ;
  assign y18853 = ~1'b0 ;
  assign y18854 = n39765 ;
  assign y18855 = ~1'b0 ;
  assign y18856 = ~n39766 ;
  assign y18857 = ~1'b0 ;
  assign y18858 = n39767 ;
  assign y18859 = n39770 ;
  assign y18860 = ~1'b0 ;
  assign y18861 = ~1'b0 ;
  assign y18862 = 1'b0 ;
  assign y18863 = ~n39773 ;
  assign y18864 = n34196 ;
  assign y18865 = ~1'b0 ;
  assign y18866 = n39774 ;
  assign y18867 = n39775 ;
  assign y18868 = n39779 ;
  assign y18869 = ~1'b0 ;
  assign y18870 = n39781 ;
  assign y18871 = n39782 ;
  assign y18872 = ~n39783 ;
  assign y18873 = ~1'b0 ;
  assign y18874 = ~n39785 ;
  assign y18875 = n39789 ;
  assign y18876 = ~n39790 ;
  assign y18877 = n39792 ;
  assign y18878 = n39797 ;
  assign y18879 = n39799 ;
  assign y18880 = ~n39801 ;
  assign y18881 = ~n39802 ;
  assign y18882 = ~1'b0 ;
  assign y18883 = ~n39804 ;
  assign y18884 = n39806 ;
  assign y18885 = n39809 ;
  assign y18886 = n39815 ;
  assign y18887 = n30821 ;
  assign y18888 = ~1'b0 ;
  assign y18889 = n16602 ;
  assign y18890 = ~1'b0 ;
  assign y18891 = 1'b0 ;
  assign y18892 = ~n4509 ;
  assign y18893 = n39816 ;
  assign y18894 = ~n39818 ;
  assign y18895 = ~n39821 ;
  assign y18896 = ~n39823 ;
  assign y18897 = ~1'b0 ;
  assign y18898 = n39824 ;
  assign y18899 = n39826 ;
  assign y18900 = n39827 ;
  assign y18901 = n39829 ;
  assign y18902 = n39832 ;
  assign y18903 = n39838 ;
  assign y18904 = n39839 ;
  assign y18905 = n39840 ;
  assign y18906 = n39846 ;
  assign y18907 = ~1'b0 ;
  assign y18908 = n39851 ;
  assign y18909 = ~n39852 ;
  assign y18910 = n39855 ;
  assign y18911 = n39857 ;
  assign y18912 = ~n39859 ;
  assign y18913 = ~n39862 ;
  assign y18914 = ~1'b0 ;
  assign y18915 = ~n39863 ;
  assign y18916 = ~1'b0 ;
  assign y18917 = n39870 ;
  assign y18918 = n39872 ;
  assign y18919 = n39874 ;
  assign y18920 = n39876 ;
  assign y18921 = ~n7559 ;
  assign y18922 = ~n39877 ;
  assign y18923 = n10697 ;
  assign y18924 = ~n39883 ;
  assign y18925 = ~1'b0 ;
  assign y18926 = ~n39884 ;
  assign y18927 = n39890 ;
  assign y18928 = ~1'b0 ;
  assign y18929 = 1'b0 ;
  assign y18930 = ~n39891 ;
  assign y18931 = ~n39892 ;
  assign y18932 = ~n39894 ;
  assign y18933 = ~1'b0 ;
  assign y18934 = ~1'b0 ;
  assign y18935 = ~1'b0 ;
  assign y18936 = n39895 ;
  assign y18937 = n39897 ;
  assign y18938 = n39898 ;
  assign y18939 = n39901 ;
  assign y18940 = ~1'b0 ;
  assign y18941 = ~n39904 ;
  assign y18942 = ~1'b0 ;
  assign y18943 = ~n39906 ;
  assign y18944 = n39907 ;
  assign y18945 = ~1'b0 ;
  assign y18946 = n39908 ;
  assign y18947 = n31412 ;
  assign y18948 = ~n39912 ;
  assign y18949 = ~n39913 ;
  assign y18950 = ~1'b0 ;
  assign y18951 = ~n39917 ;
  assign y18952 = ~n39919 ;
  assign y18953 = ~1'b0 ;
  assign y18954 = ~n39921 ;
  assign y18955 = n39927 ;
  assign y18956 = ~1'b0 ;
  assign y18957 = ~n39929 ;
  assign y18958 = n39931 ;
  assign y18959 = ~n39932 ;
  assign y18960 = n39934 ;
  assign y18961 = n39935 ;
  assign y18962 = n39938 ;
  assign y18963 = n39943 ;
  assign y18964 = ~1'b0 ;
  assign y18965 = ~1'b0 ;
  assign y18966 = n39944 ;
  assign y18967 = ~n39945 ;
  assign y18968 = n39946 ;
  assign y18969 = ~1'b0 ;
  assign y18970 = n39951 ;
  assign y18971 = ~n39954 ;
  assign y18972 = 1'b0 ;
  assign y18973 = ~1'b0 ;
  assign y18974 = n39956 ;
  assign y18975 = ~1'b0 ;
  assign y18976 = ~n11772 ;
  assign y18977 = n39958 ;
  assign y18978 = ~n39960 ;
  assign y18979 = n39964 ;
  assign y18980 = n39965 ;
  assign y18981 = ~n39967 ;
  assign y18982 = ~n39972 ;
  assign y18983 = ~n39974 ;
  assign y18984 = ~n39976 ;
  assign y18985 = n39982 ;
  assign y18986 = ~1'b0 ;
  assign y18987 = ~n39986 ;
  assign y18988 = ~n39988 ;
  assign y18989 = n39990 ;
  assign y18990 = ~1'b0 ;
  assign y18991 = ~1'b0 ;
  assign y18992 = ~1'b0 ;
  assign y18993 = ~n39994 ;
  assign y18994 = ~n39995 ;
  assign y18995 = n39997 ;
  assign y18996 = ~n21608 ;
  assign y18997 = ~n40000 ;
  assign y18998 = ~1'b0 ;
  assign y18999 = ~n40004 ;
  assign y19000 = ~1'b0 ;
  assign y19001 = ~n40006 ;
  assign y19002 = n40009 ;
  assign y19003 = n40011 ;
  assign y19004 = ~1'b0 ;
  assign y19005 = n40015 ;
  assign y19006 = ~n40016 ;
  assign y19007 = n40020 ;
  assign y19008 = ~n40025 ;
  assign y19009 = ~1'b0 ;
  assign y19010 = n40028 ;
  assign y19011 = ~1'b0 ;
  assign y19012 = ~n40031 ;
  assign y19013 = ~1'b0 ;
  assign y19014 = n40032 ;
  assign y19015 = ~n40036 ;
  assign y19016 = n40039 ;
  assign y19017 = ~n40040 ;
  assign y19018 = n40041 ;
  assign y19019 = 1'b0 ;
  assign y19020 = ~n40042 ;
  assign y19021 = ~n40043 ;
  assign y19022 = ~n40046 ;
  assign y19023 = ~n40047 ;
  assign y19024 = ~n19916 ;
  assign y19025 = ~n40049 ;
  assign y19026 = ~n40053 ;
  assign y19027 = n40054 ;
  assign y19028 = ~n40060 ;
  assign y19029 = ~n10707 ;
  assign y19030 = ~n40063 ;
  assign y19031 = ~n40064 ;
  assign y19032 = ~n40065 ;
  assign y19033 = n40067 ;
  assign y19034 = n40068 ;
  assign y19035 = ~n40070 ;
  assign y19036 = n40077 ;
  assign y19037 = ~n40080 ;
  assign y19038 = n40081 ;
  assign y19039 = n40082 ;
  assign y19040 = ~1'b0 ;
  assign y19041 = ~n40085 ;
  assign y19042 = ~1'b0 ;
  assign y19043 = ~n40086 ;
  assign y19044 = n40088 ;
  assign y19045 = ~n40089 ;
  assign y19046 = n40093 ;
  assign y19047 = n40095 ;
  assign y19048 = ~n40097 ;
  assign y19049 = ~n40098 ;
  assign y19050 = 1'b0 ;
  assign y19051 = ~1'b0 ;
  assign y19052 = ~1'b0 ;
  assign y19053 = n40100 ;
  assign y19054 = n40102 ;
  assign y19055 = ~n40106 ;
  assign y19056 = n40111 ;
  assign y19057 = ~1'b0 ;
  assign y19058 = ~n40112 ;
  assign y19059 = n40114 ;
  assign y19060 = ~1'b0 ;
  assign y19061 = n40117 ;
  assign y19062 = ~1'b0 ;
  assign y19063 = ~1'b0 ;
  assign y19064 = n40119 ;
  assign y19065 = 1'b0 ;
  assign y19066 = ~n40123 ;
  assign y19067 = ~n40124 ;
  assign y19068 = n40127 ;
  assign y19069 = n40128 ;
  assign y19070 = n40132 ;
  assign y19071 = n40137 ;
  assign y19072 = ~n40139 ;
  assign y19073 = ~n40144 ;
  assign y19074 = n40150 ;
  assign y19075 = ~n40152 ;
  assign y19076 = ~n40156 ;
  assign y19077 = n24253 ;
  assign y19078 = ~n40158 ;
  assign y19079 = ~n40163 ;
  assign y19080 = ~n40165 ;
  assign y19081 = n40167 ;
  assign y19082 = ~n40168 ;
  assign y19083 = ~n40171 ;
  assign y19084 = n40172 ;
  assign y19085 = n40175 ;
  assign y19086 = n40176 ;
  assign y19087 = n40178 ;
  assign y19088 = n40181 ;
  assign y19089 = ~n40185 ;
  assign y19090 = ~n40188 ;
  assign y19091 = ~n40189 ;
  assign y19092 = ~n40190 ;
  assign y19093 = n40192 ;
  assign y19094 = n585 ;
  assign y19095 = ~n40194 ;
  assign y19096 = ~1'b0 ;
  assign y19097 = 1'b0 ;
  assign y19098 = ~n40195 ;
  assign y19099 = ~1'b0 ;
  assign y19100 = ~n40196 ;
  assign y19101 = n40202 ;
  assign y19102 = n40204 ;
  assign y19103 = n7485 ;
  assign y19104 = ~1'b0 ;
  assign y19105 = n40205 ;
  assign y19106 = ~n40208 ;
  assign y19107 = ~1'b0 ;
  assign y19108 = ~1'b0 ;
  assign y19109 = n40209 ;
  assign y19110 = ~n40212 ;
  assign y19111 = ~1'b0 ;
  assign y19112 = ~1'b0 ;
  assign y19113 = ~1'b0 ;
  assign y19114 = ~1'b0 ;
  assign y19115 = ~1'b0 ;
  assign y19116 = ~1'b0 ;
  assign y19117 = ~n40219 ;
  assign y19118 = 1'b0 ;
  assign y19119 = ~n40222 ;
  assign y19120 = ~n40227 ;
  assign y19121 = ~n30701 ;
  assign y19122 = ~n40228 ;
  assign y19123 = ~1'b0 ;
  assign y19124 = n40232 ;
  assign y19125 = ~n40236 ;
  assign y19126 = ~n40237 ;
  assign y19127 = ~1'b0 ;
  assign y19128 = ~n40238 ;
  assign y19129 = ~1'b0 ;
  assign y19130 = ~n40240 ;
  assign y19131 = n40242 ;
  assign y19132 = ~n40244 ;
  assign y19133 = ~n40246 ;
  assign y19134 = ~n40247 ;
  assign y19135 = n40254 ;
  assign y19136 = ~n40255 ;
  assign y19137 = n40256 ;
  assign y19138 = ~1'b0 ;
  assign y19139 = ~n40257 ;
  assign y19140 = ~n40259 ;
  assign y19141 = ~n40261 ;
  assign y19142 = ~1'b0 ;
  assign y19143 = ~1'b0 ;
  assign y19144 = ~n40267 ;
  assign y19145 = n40268 ;
  assign y19146 = ~1'b0 ;
  assign y19147 = n40270 ;
  assign y19148 = ~n40272 ;
  assign y19149 = ~1'b0 ;
  assign y19150 = ~n40276 ;
  assign y19151 = n40278 ;
  assign y19152 = ~n40279 ;
  assign y19153 = n40281 ;
  assign y19154 = ~n40282 ;
  assign y19155 = ~n40285 ;
  assign y19156 = n40288 ;
  assign y19157 = ~1'b0 ;
  assign y19158 = ~n40289 ;
  assign y19159 = ~1'b0 ;
  assign y19160 = n40290 ;
  assign y19161 = ~n40292 ;
  assign y19162 = n40293 ;
  assign y19163 = n40295 ;
  assign y19164 = ~n40296 ;
  assign y19165 = ~n40297 ;
  assign y19166 = ~n40300 ;
  assign y19167 = 1'b0 ;
  assign y19168 = ~1'b0 ;
  assign y19169 = n40301 ;
  assign y19170 = n40302 ;
  assign y19171 = n40304 ;
  assign y19172 = ~1'b0 ;
  assign y19173 = n40305 ;
  assign y19174 = ~1'b0 ;
  assign y19175 = n40306 ;
  assign y19176 = ~n40310 ;
  assign y19177 = ~n40312 ;
  assign y19178 = n13700 ;
  assign y19179 = ~n40314 ;
  assign y19180 = ~n19467 ;
  assign y19181 = ~1'b0 ;
  assign y19182 = n40316 ;
  assign y19183 = ~n40319 ;
  assign y19184 = n40325 ;
  assign y19185 = ~1'b0 ;
  assign y19186 = ~1'b0 ;
  assign y19187 = ~1'b0 ;
  assign y19188 = n40327 ;
  assign y19189 = ~n40328 ;
  assign y19190 = ~n40329 ;
  assign y19191 = ~1'b0 ;
  assign y19192 = ~n40330 ;
  assign y19193 = n40332 ;
  assign y19194 = ~n40333 ;
  assign y19195 = ~1'b0 ;
  assign y19196 = ~1'b0 ;
  assign y19197 = n40336 ;
  assign y19198 = n40337 ;
  assign y19199 = ~1'b0 ;
  assign y19200 = n40343 ;
  assign y19201 = ~n40344 ;
  assign y19202 = ~n40345 ;
  assign y19203 = ~1'b0 ;
  assign y19204 = n16130 ;
  assign y19205 = ~n15717 ;
  assign y19206 = ~n40346 ;
  assign y19207 = ~1'b0 ;
  assign y19208 = ~n40351 ;
  assign y19209 = ~n40355 ;
  assign y19210 = ~n34579 ;
  assign y19211 = ~1'b0 ;
  assign y19212 = ~1'b0 ;
  assign y19213 = n40356 ;
  assign y19214 = ~n40360 ;
  assign y19215 = n40362 ;
  assign y19216 = ~1'b0 ;
  assign y19217 = n40365 ;
  assign y19218 = ~n40367 ;
  assign y19219 = ~n40369 ;
  assign y19220 = n40371 ;
  assign y19221 = ~1'b0 ;
  assign y19222 = ~n40374 ;
  assign y19223 = ~1'b0 ;
  assign y19224 = ~n40378 ;
  assign y19225 = ~n40379 ;
  assign y19226 = n40380 ;
  assign y19227 = ~n40383 ;
  assign y19228 = ~1'b0 ;
  assign y19229 = n40387 ;
  assign y19230 = 1'b0 ;
  assign y19231 = 1'b0 ;
  assign y19232 = ~n40392 ;
  assign y19233 = n40394 ;
  assign y19234 = ~n40399 ;
  assign y19235 = ~n40400 ;
  assign y19236 = n40402 ;
  assign y19237 = ~1'b0 ;
  assign y19238 = n40405 ;
  assign y19239 = ~1'b0 ;
  assign y19240 = ~n40408 ;
  assign y19241 = n40411 ;
  assign y19242 = ~1'b0 ;
  assign y19243 = n40412 ;
  assign y19244 = ~n40413 ;
  assign y19245 = ~n40415 ;
  assign y19246 = n40417 ;
  assign y19247 = n40418 ;
  assign y19248 = n40422 ;
  assign y19249 = n40425 ;
  assign y19250 = ~n40426 ;
  assign y19251 = ~1'b0 ;
  assign y19252 = n40429 ;
  assign y19253 = ~1'b0 ;
  assign y19254 = n40433 ;
  assign y19255 = ~1'b0 ;
  assign y19256 = n9822 ;
  assign y19257 = n40434 ;
  assign y19258 = n40437 ;
  assign y19259 = ~n34980 ;
  assign y19260 = ~1'b0 ;
  assign y19261 = ~1'b0 ;
  assign y19262 = ~1'b0 ;
  assign y19263 = ~n40439 ;
  assign y19264 = ~n40444 ;
  assign y19265 = ~n40446 ;
  assign y19266 = ~n40447 ;
  assign y19267 = n40448 ;
  assign y19268 = ~n28270 ;
  assign y19269 = ~n40450 ;
  assign y19270 = n40453 ;
  assign y19271 = ~n40455 ;
  assign y19272 = ~1'b0 ;
  assign y19273 = ~n40457 ;
  assign y19274 = n40460 ;
  assign y19275 = n40461 ;
  assign y19276 = n40465 ;
  assign y19277 = ~1'b0 ;
  assign y19278 = ~n31478 ;
  assign y19279 = ~n40466 ;
  assign y19280 = n40467 ;
  assign y19281 = ~n40471 ;
  assign y19282 = ~n40478 ;
  assign y19283 = ~n40479 ;
  assign y19284 = n31972 ;
  assign y19285 = n40486 ;
  assign y19286 = ~1'b0 ;
  assign y19287 = n40490 ;
  assign y19288 = n1913 ;
  assign y19289 = n40493 ;
  assign y19290 = n40494 ;
  assign y19291 = ~n40495 ;
  assign y19292 = ~1'b0 ;
  assign y19293 = ~1'b0 ;
  assign y19294 = n40496 ;
  assign y19295 = ~1'b0 ;
  assign y19296 = n40500 ;
  assign y19297 = ~n40502 ;
  assign y19298 = ~n40503 ;
  assign y19299 = n40505 ;
  assign y19300 = ~n40507 ;
  assign y19301 = ~1'b0 ;
  assign y19302 = ~1'b0 ;
  assign y19303 = ~n40512 ;
  assign y19304 = ~1'b0 ;
  assign y19305 = n31832 ;
  assign y19306 = ~1'b0 ;
  assign y19307 = n40514 ;
  assign y19308 = ~n40515 ;
  assign y19309 = ~n40516 ;
  assign y19310 = ~1'b0 ;
  assign y19311 = ~n40520 ;
  assign y19312 = ~n40521 ;
  assign y19313 = ~n40522 ;
  assign y19314 = n40525 ;
  assign y19315 = ~n40527 ;
  assign y19316 = ~1'b0 ;
  assign y19317 = n40531 ;
  assign y19318 = n40534 ;
  assign y19319 = ~n40535 ;
  assign y19320 = n23614 ;
  assign y19321 = ~1'b0 ;
  assign y19322 = ~n40536 ;
  assign y19323 = ~1'b0 ;
  assign y19324 = ~1'b0 ;
  assign y19325 = n40541 ;
  assign y19326 = ~n40544 ;
  assign y19327 = ~n40545 ;
  assign y19328 = n40546 ;
  assign y19329 = n31669 ;
  assign y19330 = n40549 ;
  assign y19331 = n40550 ;
  assign y19332 = ~n40554 ;
  assign y19333 = ~1'b0 ;
  assign y19334 = ~n40560 ;
  assign y19335 = ~n40563 ;
  assign y19336 = n19225 ;
  assign y19337 = n40564 ;
  assign y19338 = ~1'b0 ;
  assign y19339 = n40566 ;
  assign y19340 = n33339 ;
  assign y19341 = ~n40567 ;
  assign y19342 = n40568 ;
  assign y19343 = ~1'b0 ;
  assign y19344 = ~n40570 ;
  assign y19345 = ~1'b0 ;
  assign y19346 = ~n40571 ;
  assign y19347 = ~n40572 ;
  assign y19348 = n40579 ;
  assign y19349 = ~1'b0 ;
  assign y19350 = ~n40581 ;
  assign y19351 = n40589 ;
  assign y19352 = ~n40595 ;
  assign y19353 = ~1'b0 ;
  assign y19354 = ~1'b0 ;
  assign y19355 = ~1'b0 ;
  assign y19356 = ~1'b0 ;
  assign y19357 = n40596 ;
  assign y19358 = n40597 ;
  assign y19359 = ~n13754 ;
  assign y19360 = ~n40601 ;
  assign y19361 = ~n40607 ;
  assign y19362 = n40610 ;
  assign y19363 = ~n40612 ;
  assign y19364 = ~n40614 ;
  assign y19365 = n40615 ;
  assign y19366 = n40617 ;
  assign y19367 = n40618 ;
  assign y19368 = ~1'b0 ;
  assign y19369 = ~1'b0 ;
  assign y19370 = ~n40619 ;
  assign y19371 = n40625 ;
  assign y19372 = ~n4024 ;
  assign y19373 = ~n40626 ;
  assign y19374 = ~n40628 ;
  assign y19375 = n40630 ;
  assign y19376 = n40631 ;
  assign y19377 = n40633 ;
  assign y19378 = ~1'b0 ;
  assign y19379 = ~n40635 ;
  assign y19380 = ~1'b0 ;
  assign y19381 = ~1'b0 ;
  assign y19382 = n40638 ;
  assign y19383 = ~1'b0 ;
  assign y19384 = ~n40641 ;
  assign y19385 = n40642 ;
  assign y19386 = ~n40643 ;
  assign y19387 = n40647 ;
  assign y19388 = ~n40652 ;
  assign y19389 = n40658 ;
  assign y19390 = ~1'b0 ;
  assign y19391 = ~1'b0 ;
  assign y19392 = ~n40660 ;
  assign y19393 = ~1'b0 ;
  assign y19394 = ~n15867 ;
  assign y19395 = n40662 ;
  assign y19396 = ~n40663 ;
  assign y19397 = ~n40667 ;
  assign y19398 = ~1'b0 ;
  assign y19399 = ~n40671 ;
  assign y19400 = ~n40675 ;
  assign y19401 = ~n40679 ;
  assign y19402 = ~1'b0 ;
  assign y19403 = ~n40685 ;
  assign y19404 = ~n40688 ;
  assign y19405 = n40691 ;
  assign y19406 = n40692 ;
  assign y19407 = ~n40693 ;
  assign y19408 = n40695 ;
  assign y19409 = ~1'b0 ;
  assign y19410 = ~n40697 ;
  assign y19411 = ~1'b0 ;
  assign y19412 = n34847 ;
  assign y19413 = n40698 ;
  assign y19414 = ~n40700 ;
  assign y19415 = ~n40701 ;
  assign y19416 = ~n7839 ;
  assign y19417 = n40702 ;
  assign y19418 = n40704 ;
  assign y19419 = n40708 ;
  assign y19420 = ~1'b0 ;
  assign y19421 = n40709 ;
  assign y19422 = ~n40713 ;
  assign y19423 = ~1'b0 ;
  assign y19424 = ~1'b0 ;
  assign y19425 = ~n40717 ;
  assign y19426 = ~n40718 ;
  assign y19427 = x184 ;
  assign y19428 = n40719 ;
  assign y19429 = ~1'b0 ;
  assign y19430 = n40721 ;
  assign y19431 = ~1'b0 ;
  assign y19432 = ~n40723 ;
  assign y19433 = ~1'b0 ;
  assign y19434 = ~n40726 ;
  assign y19435 = ~n40733 ;
  assign y19436 = ~1'b0 ;
  assign y19437 = n40734 ;
  assign y19438 = n40737 ;
  assign y19439 = ~n19671 ;
  assign y19440 = ~1'b0 ;
  assign y19441 = n40738 ;
  assign y19442 = n40740 ;
  assign y19443 = n40743 ;
  assign y19444 = n40745 ;
  assign y19445 = n40749 ;
  assign y19446 = ~n40750 ;
  assign y19447 = ~1'b0 ;
  assign y19448 = ~1'b0 ;
  assign y19449 = n40752 ;
  assign y19450 = n15712 ;
  assign y19451 = ~1'b0 ;
  assign y19452 = ~n40757 ;
  assign y19453 = n40758 ;
  assign y19454 = 1'b0 ;
  assign y19455 = ~n40761 ;
  assign y19456 = 1'b0 ;
  assign y19457 = ~1'b0 ;
  assign y19458 = ~1'b0 ;
  assign y19459 = ~1'b0 ;
  assign y19460 = ~n40762 ;
  assign y19461 = ~n40765 ;
  assign y19462 = ~n40767 ;
  assign y19463 = n40769 ;
  assign y19464 = ~n40770 ;
  assign y19465 = n40772 ;
  assign y19466 = ~1'b0 ;
  assign y19467 = n40773 ;
  assign y19468 = n40776 ;
  assign y19469 = n40777 ;
  assign y19470 = n40778 ;
  assign y19471 = ~n40779 ;
  assign y19472 = n40783 ;
  assign y19473 = ~1'b0 ;
  assign y19474 = n21652 ;
  assign y19475 = ~1'b0 ;
  assign y19476 = n40785 ;
  assign y19477 = n40787 ;
  assign y19478 = n40789 ;
  assign y19479 = ~n40790 ;
  assign y19480 = ~n40792 ;
  assign y19481 = ~n40793 ;
  assign y19482 = ~n40794 ;
  assign y19483 = ~1'b0 ;
  assign y19484 = n40797 ;
  assign y19485 = ~1'b0 ;
  assign y19486 = n40799 ;
  assign y19487 = ~n40801 ;
  assign y19488 = n40806 ;
  assign y19489 = n40808 ;
  assign y19490 = ~n40809 ;
  assign y19491 = ~n40810 ;
  assign y19492 = ~n40813 ;
  assign y19493 = ~1'b0 ;
  assign y19494 = ~n40815 ;
  assign y19495 = ~1'b0 ;
  assign y19496 = ~1'b0 ;
  assign y19497 = ~n3430 ;
  assign y19498 = ~n40816 ;
  assign y19499 = ~n40818 ;
  assign y19500 = ~1'b0 ;
  assign y19501 = ~1'b0 ;
  assign y19502 = ~1'b0 ;
  assign y19503 = ~1'b0 ;
  assign y19504 = 1'b0 ;
  assign y19505 = ~n40826 ;
  assign y19506 = ~n40829 ;
  assign y19507 = ~n40833 ;
  assign y19508 = n40839 ;
  assign y19509 = ~n40840 ;
  assign y19510 = ~1'b0 ;
  assign y19511 = ~n40842 ;
  assign y19512 = ~n40843 ;
  assign y19513 = ~n40844 ;
  assign y19514 = ~1'b0 ;
  assign y19515 = ~1'b0 ;
  assign y19516 = ~1'b0 ;
  assign y19517 = ~n40845 ;
  assign y19518 = ~n40846 ;
  assign y19519 = n25755 ;
  assign y19520 = ~n40849 ;
  assign y19521 = n40850 ;
  assign y19522 = ~1'b0 ;
  assign y19523 = ~1'b0 ;
  assign y19524 = ~1'b0 ;
  assign y19525 = ~1'b0 ;
  assign y19526 = ~1'b0 ;
  assign y19527 = n40851 ;
  assign y19528 = n5433 ;
  assign y19529 = ~n40852 ;
  assign y19530 = ~n40854 ;
  assign y19531 = ~1'b0 ;
  assign y19532 = n40855 ;
  assign y19533 = ~n40857 ;
  assign y19534 = n1768 ;
  assign y19535 = ~1'b0 ;
  assign y19536 = n40858 ;
  assign y19537 = ~n40860 ;
  assign y19538 = n40861 ;
  assign y19539 = ~n40862 ;
  assign y19540 = n40869 ;
  assign y19541 = n40870 ;
  assign y19542 = ~n40872 ;
  assign y19543 = ~n40876 ;
  assign y19544 = n40878 ;
  assign y19545 = ~n40880 ;
  assign y19546 = ~n40882 ;
  assign y19547 = ~1'b0 ;
  assign y19548 = ~n40886 ;
  assign y19549 = ~n29837 ;
  assign y19550 = n40887 ;
  assign y19551 = ~1'b0 ;
  assign y19552 = n40888 ;
  assign y19553 = n40890 ;
  assign y19554 = ~1'b0 ;
  assign y19555 = ~1'b0 ;
  assign y19556 = ~n40892 ;
  assign y19557 = ~1'b0 ;
  assign y19558 = n40893 ;
  assign y19559 = ~n40895 ;
  assign y19560 = n40896 ;
  assign y19561 = ~1'b0 ;
  assign y19562 = n40897 ;
  assign y19563 = ~n40899 ;
  assign y19564 = ~n40901 ;
  assign y19565 = ~n40902 ;
  assign y19566 = ~n31893 ;
  assign y19567 = n40903 ;
  assign y19568 = ~n40907 ;
  assign y19569 = n40909 ;
  assign y19570 = n40910 ;
  assign y19571 = ~1'b0 ;
  assign y19572 = ~n40913 ;
  assign y19573 = ~1'b0 ;
  assign y19574 = n40915 ;
  assign y19575 = ~1'b0 ;
  assign y19576 = n40916 ;
  assign y19577 = n40917 ;
  assign y19578 = n40920 ;
  assign y19579 = ~n40922 ;
  assign y19580 = ~n40926 ;
  assign y19581 = n1187 ;
  assign y19582 = n40928 ;
  assign y19583 = ~n40931 ;
  assign y19584 = ~n40935 ;
  assign y19585 = n40939 ;
  assign y19586 = ~1'b0 ;
  assign y19587 = ~n40941 ;
  assign y19588 = ~n40942 ;
  assign y19589 = ~1'b0 ;
  assign y19590 = ~1'b0 ;
  assign y19591 = ~1'b0 ;
  assign y19592 = n40944 ;
  assign y19593 = n40945 ;
  assign y19594 = ~n40947 ;
  assign y19595 = n35776 ;
  assign y19596 = ~1'b0 ;
  assign y19597 = n40948 ;
  assign y19598 = ~n40949 ;
  assign y19599 = ~1'b0 ;
  assign y19600 = ~n40956 ;
  assign y19601 = n40957 ;
  assign y19602 = n12885 ;
  assign y19603 = ~1'b0 ;
  assign y19604 = ~n40958 ;
  assign y19605 = n40961 ;
  assign y19606 = n40962 ;
  assign y19607 = ~1'b0 ;
  assign y19608 = ~1'b0 ;
  assign y19609 = ~n40967 ;
  assign y19610 = ~1'b0 ;
  assign y19611 = ~n40969 ;
  assign y19612 = ~1'b0 ;
  assign y19613 = n40971 ;
  assign y19614 = n40975 ;
  assign y19615 = ~n40976 ;
  assign y19616 = ~n40977 ;
  assign y19617 = ~1'b0 ;
  assign y19618 = ~n40979 ;
  assign y19619 = n40981 ;
  assign y19620 = ~1'b0 ;
  assign y19621 = n795 ;
  assign y19622 = ~n40983 ;
  assign y19623 = ~n40984 ;
  assign y19624 = ~1'b0 ;
  assign y19625 = ~n40985 ;
  assign y19626 = ~n40986 ;
  assign y19627 = n40987 ;
  assign y19628 = ~n40990 ;
  assign y19629 = ~1'b0 ;
  assign y19630 = ~1'b0 ;
  assign y19631 = ~n40991 ;
  assign y19632 = n40992 ;
  assign y19633 = n40995 ;
  assign y19634 = ~1'b0 ;
  assign y19635 = ~1'b0 ;
  assign y19636 = n40999 ;
  assign y19637 = n11301 ;
  assign y19638 = ~1'b0 ;
  assign y19639 = ~1'b0 ;
  assign y19640 = ~1'b0 ;
  assign y19641 = n41004 ;
  assign y19642 = n41005 ;
  assign y19643 = ~n41009 ;
  assign y19644 = ~n41011 ;
  assign y19645 = ~1'b0 ;
  assign y19646 = n41013 ;
  assign y19647 = n41014 ;
  assign y19648 = ~n41016 ;
  assign y19649 = ~n41022 ;
  assign y19650 = n41025 ;
  assign y19651 = ~n41028 ;
  assign y19652 = ~n41029 ;
  assign y19653 = ~1'b0 ;
  assign y19654 = ~n41030 ;
  assign y19655 = ~n41031 ;
  assign y19656 = ~n41036 ;
  assign y19657 = 1'b0 ;
  assign y19658 = n25602 ;
  assign y19659 = n41037 ;
  assign y19660 = ~n41041 ;
  assign y19661 = n41044 ;
  assign y19662 = n41046 ;
  assign y19663 = n41048 ;
  assign y19664 = ~n41050 ;
  assign y19665 = n41055 ;
  assign y19666 = ~n41057 ;
  assign y19667 = ~n41058 ;
  assign y19668 = ~n41061 ;
  assign y19669 = n41062 ;
  assign y19670 = ~1'b0 ;
  assign y19671 = ~n41063 ;
  assign y19672 = ~1'b0 ;
  assign y19673 = ~1'b0 ;
  assign y19674 = n41065 ;
  assign y19675 = n41071 ;
  assign y19676 = ~n41074 ;
  assign y19677 = n5228 ;
  assign y19678 = ~n41077 ;
  assign y19679 = ~n41078 ;
  assign y19680 = n41080 ;
  assign y19681 = ~1'b0 ;
  assign y19682 = ~n41082 ;
  assign y19683 = ~n41084 ;
  assign y19684 = ~1'b0 ;
  assign y19685 = ~1'b0 ;
  assign y19686 = ~1'b0 ;
  assign y19687 = ~n31404 ;
  assign y19688 = ~n41087 ;
  assign y19689 = ~n41088 ;
  assign y19690 = ~n30444 ;
  assign y19691 = ~1'b0 ;
  assign y19692 = ~n41090 ;
  assign y19693 = ~n41092 ;
  assign y19694 = ~n41096 ;
  assign y19695 = n41098 ;
  assign y19696 = ~n41099 ;
  assign y19697 = ~n41102 ;
  assign y19698 = ~1'b0 ;
  assign y19699 = n41104 ;
  assign y19700 = ~1'b0 ;
  assign y19701 = n41106 ;
  assign y19702 = ~n41111 ;
  assign y19703 = ~1'b0 ;
  assign y19704 = n41112 ;
  assign y19705 = ~n41114 ;
  assign y19706 = ~n22877 ;
  assign y19707 = n41115 ;
  assign y19708 = n41120 ;
  assign y19709 = n41122 ;
  assign y19710 = ~n29751 ;
  assign y19711 = 1'b0 ;
  assign y19712 = n41123 ;
  assign y19713 = ~n41129 ;
  assign y19714 = ~n41130 ;
  assign y19715 = ~1'b0 ;
  assign y19716 = n41133 ;
  assign y19717 = ~n41135 ;
  assign y19718 = ~n41136 ;
  assign y19719 = ~n41137 ;
  assign y19720 = ~1'b0 ;
  assign y19721 = ~1'b0 ;
  assign y19722 = n41140 ;
  assign y19723 = ~n41142 ;
  assign y19724 = n41143 ;
  assign y19725 = n41144 ;
  assign y19726 = n41146 ;
  assign y19727 = n41147 ;
  assign y19728 = ~1'b0 ;
  assign y19729 = ~1'b0 ;
  assign y19730 = ~n41148 ;
  assign y19731 = ~1'b0 ;
  assign y19732 = ~n41152 ;
  assign y19733 = n41154 ;
  assign y19734 = ~n41155 ;
  assign y19735 = n41163 ;
  assign y19736 = ~n41165 ;
  assign y19737 = n41172 ;
  assign y19738 = n41173 ;
  assign y19739 = ~n41175 ;
  assign y19740 = ~1'b0 ;
  assign y19741 = ~1'b0 ;
  assign y19742 = ~n41176 ;
  assign y19743 = n41177 ;
  assign y19744 = ~n41178 ;
  assign y19745 = n41180 ;
  assign y19746 = ~n41185 ;
  assign y19747 = ~n41187 ;
  assign y19748 = ~1'b0 ;
  assign y19749 = ~1'b0 ;
  assign y19750 = ~n20783 ;
  assign y19751 = ~n41193 ;
  assign y19752 = ~n32350 ;
  assign y19753 = ~n41195 ;
  assign y19754 = n41199 ;
  assign y19755 = n41200 ;
  assign y19756 = n16233 ;
  assign y19757 = ~1'b0 ;
  assign y19758 = n41204 ;
  assign y19759 = n41205 ;
  assign y19760 = ~1'b0 ;
  assign y19761 = ~1'b0 ;
  assign y19762 = ~n41206 ;
  assign y19763 = ~1'b0 ;
  assign y19764 = ~1'b0 ;
  assign y19765 = n41207 ;
  assign y19766 = n41210 ;
  assign y19767 = n41215 ;
  assign y19768 = ~1'b0 ;
  assign y19769 = ~1'b0 ;
  assign y19770 = n41216 ;
  assign y19771 = n41217 ;
  assign y19772 = ~n41219 ;
  assign y19773 = ~1'b0 ;
  assign y19774 = ~n41220 ;
  assign y19775 = n11219 ;
  assign y19776 = ~n41222 ;
  assign y19777 = ~n41226 ;
  assign y19778 = n41227 ;
  assign y19779 = n41232 ;
  assign y19780 = ~n41233 ;
  assign y19781 = n41236 ;
  assign y19782 = n41238 ;
  assign y19783 = ~1'b0 ;
  assign y19784 = ~n41240 ;
  assign y19785 = ~n41242 ;
  assign y19786 = ~n41243 ;
  assign y19787 = ~n41244 ;
  assign y19788 = ~1'b0 ;
  assign y19789 = n41245 ;
  assign y19790 = n41247 ;
  assign y19791 = n41249 ;
  assign y19792 = n41250 ;
  assign y19793 = ~1'b0 ;
  assign y19794 = ~n41252 ;
  assign y19795 = n41255 ;
  assign y19796 = ~n41258 ;
  assign y19797 = n41259 ;
  assign y19798 = n41261 ;
  assign y19799 = ~n41263 ;
  assign y19800 = n41264 ;
  assign y19801 = ~1'b0 ;
  assign y19802 = ~1'b0 ;
  assign y19803 = ~n41266 ;
  assign y19804 = ~n41271 ;
  assign y19805 = ~n41272 ;
  assign y19806 = ~n41273 ;
  assign y19807 = n41278 ;
  assign y19808 = n41285 ;
  assign y19809 = ~n41288 ;
  assign y19810 = ~1'b0 ;
  assign y19811 = n41289 ;
  assign y19812 = ~1'b0 ;
  assign y19813 = ~n41291 ;
  assign y19814 = ~n41292 ;
  assign y19815 = n41295 ;
  assign y19816 = ~n41296 ;
  assign y19817 = ~1'b0 ;
  assign y19818 = n41299 ;
  assign y19819 = ~n41303 ;
  assign y19820 = n41304 ;
  assign y19821 = n41306 ;
  assign y19822 = ~n41307 ;
  assign y19823 = n41311 ;
  assign y19824 = ~1'b0 ;
  assign y19825 = ~n41312 ;
  assign y19826 = ~1'b0 ;
  assign y19827 = ~n16480 ;
  assign y19828 = ~1'b0 ;
  assign y19829 = ~n41314 ;
  assign y19830 = n41316 ;
  assign y19831 = ~n41317 ;
  assign y19832 = ~n41318 ;
  assign y19833 = ~n17148 ;
  assign y19834 = ~1'b0 ;
  assign y19835 = n41323 ;
  assign y19836 = ~1'b0 ;
  assign y19837 = n41327 ;
  assign y19838 = n41328 ;
  assign y19839 = n41329 ;
  assign y19840 = n41334 ;
  assign y19841 = ~n41342 ;
  assign y19842 = n41343 ;
  assign y19843 = ~n41346 ;
  assign y19844 = n41347 ;
  assign y19845 = 1'b0 ;
  assign y19846 = ~n41349 ;
  assign y19847 = ~1'b0 ;
  assign y19848 = n41350 ;
  assign y19849 = 1'b0 ;
  assign y19850 = ~n41352 ;
  assign y19851 = ~1'b0 ;
  assign y19852 = ~n41353 ;
  assign y19853 = n34505 ;
  assign y19854 = ~n41355 ;
  assign y19855 = ~1'b0 ;
  assign y19856 = ~1'b0 ;
  assign y19857 = n41357 ;
  assign y19858 = n41358 ;
  assign y19859 = ~n41359 ;
  assign y19860 = n41361 ;
  assign y19861 = ~1'b0 ;
  assign y19862 = ~1'b0 ;
  assign y19863 = ~n41364 ;
  assign y19864 = ~1'b0 ;
  assign y19865 = ~n41365 ;
  assign y19866 = n41366 ;
  assign y19867 = ~n41367 ;
  assign y19868 = ~n41368 ;
  assign y19869 = ~1'b0 ;
  assign y19870 = n41370 ;
  assign y19871 = ~1'b0 ;
  assign y19872 = ~n41381 ;
  assign y19873 = ~1'b0 ;
  assign y19874 = ~n15227 ;
  assign y19875 = ~1'b0 ;
  assign y19876 = ~n41382 ;
  assign y19877 = n41389 ;
  assign y19878 = ~n41390 ;
  assign y19879 = ~1'b0 ;
  assign y19880 = n41391 ;
  assign y19881 = n41393 ;
  assign y19882 = ~n41394 ;
  assign y19883 = ~1'b0 ;
  assign y19884 = ~n41395 ;
  assign y19885 = ~n41396 ;
  assign y19886 = n18899 ;
  assign y19887 = n41399 ;
  assign y19888 = ~n41402 ;
  assign y19889 = ~n41406 ;
  assign y19890 = ~n41410 ;
  assign y19891 = ~1'b0 ;
  assign y19892 = n41413 ;
  assign y19893 = n41415 ;
  assign y19894 = ~1'b0 ;
  assign y19895 = n41419 ;
  assign y19896 = n41420 ;
  assign y19897 = n26986 ;
  assign y19898 = n41424 ;
  assign y19899 = ~1'b0 ;
  assign y19900 = n41427 ;
  assign y19901 = ~n41428 ;
  assign y19902 = n41429 ;
  assign y19903 = ~n41431 ;
  assign y19904 = ~1'b0 ;
  assign y19905 = n41433 ;
  assign y19906 = ~n41436 ;
  assign y19907 = n41437 ;
  assign y19908 = ~1'b0 ;
  assign y19909 = ~1'b0 ;
  assign y19910 = ~1'b0 ;
  assign y19911 = n41438 ;
  assign y19912 = ~n41444 ;
  assign y19913 = ~n41445 ;
  assign y19914 = n41447 ;
  assign y19915 = ~n41449 ;
  assign y19916 = n41456 ;
  assign y19917 = ~1'b0 ;
  assign y19918 = ~n41458 ;
  assign y19919 = ~1'b0 ;
  assign y19920 = n41459 ;
  assign y19921 = n41470 ;
  assign y19922 = n26463 ;
  assign y19923 = ~n41476 ;
  assign y19924 = n41483 ;
  assign y19925 = ~1'b0 ;
  assign y19926 = ~1'b0 ;
  assign y19927 = ~1'b0 ;
  assign y19928 = ~n41491 ;
  assign y19929 = ~1'b0 ;
  assign y19930 = ~n41493 ;
  assign y19931 = ~1'b0 ;
  assign y19932 = x210 ;
  assign y19933 = n41495 ;
  assign y19934 = n41497 ;
  assign y19935 = ~1'b0 ;
  assign y19936 = 1'b0 ;
  assign y19937 = ~n41498 ;
  assign y19938 = n41499 ;
  assign y19939 = n41500 ;
  assign y19940 = n41504 ;
  assign y19941 = n18888 ;
  assign y19942 = ~n41506 ;
  assign y19943 = ~n41507 ;
  assign y19944 = ~1'b0 ;
  assign y19945 = ~n41509 ;
  assign y19946 = ~n41511 ;
  assign y19947 = ~n41512 ;
  assign y19948 = ~n30427 ;
  assign y19949 = ~n41516 ;
  assign y19950 = ~n41520 ;
  assign y19951 = n41524 ;
  assign y19952 = ~1'b0 ;
  assign y19953 = ~1'b0 ;
  assign y19954 = ~n41525 ;
  assign y19955 = ~n41526 ;
  assign y19956 = ~n41529 ;
  assign y19957 = n41532 ;
  assign y19958 = ~n41533 ;
  assign y19959 = n41535 ;
  assign y19960 = ~n41537 ;
  assign y19961 = ~n41539 ;
  assign y19962 = ~n41541 ;
  assign y19963 = ~1'b0 ;
  assign y19964 = ~n41542 ;
  assign y19965 = ~n41543 ;
  assign y19966 = ~n41545 ;
  assign y19967 = ~n41546 ;
  assign y19968 = n36740 ;
  assign y19969 = ~n41550 ;
  assign y19970 = n41554 ;
  assign y19971 = ~1'b0 ;
  assign y19972 = ~n16129 ;
  assign y19973 = n41556 ;
  assign y19974 = ~1'b0 ;
  assign y19975 = n41558 ;
  assign y19976 = n41559 ;
  assign y19977 = ~n41560 ;
  assign y19978 = ~n41565 ;
  assign y19979 = n41566 ;
  assign y19980 = n24904 ;
  assign y19981 = n41568 ;
  assign y19982 = ~n41569 ;
  assign y19983 = ~1'b0 ;
  assign y19984 = ~1'b0 ;
  assign y19985 = ~n41572 ;
  assign y19986 = n23855 ;
  assign y19987 = ~1'b0 ;
  assign y19988 = n41574 ;
  assign y19989 = ~n41576 ;
  assign y19990 = n41579 ;
  assign y19991 = ~n41580 ;
  assign y19992 = ~1'b0 ;
  assign y19993 = ~1'b0 ;
  assign y19994 = ~n41582 ;
  assign y19995 = ~1'b0 ;
  assign y19996 = n41585 ;
  assign y19997 = n41589 ;
  assign y19998 = ~n41592 ;
  assign y19999 = ~1'b0 ;
  assign y20000 = ~1'b0 ;
  assign y20001 = ~1'b0 ;
  assign y20002 = n41594 ;
  assign y20003 = ~n41596 ;
  assign y20004 = n41597 ;
  assign y20005 = ~n41600 ;
  assign y20006 = ~1'b0 ;
  assign y20007 = ~n41601 ;
  assign y20008 = ~n41603 ;
  assign y20009 = ~n41604 ;
  assign y20010 = ~n41605 ;
  assign y20011 = 1'b0 ;
  assign y20012 = n41608 ;
  assign y20013 = n41611 ;
  assign y20014 = ~1'b0 ;
  assign y20015 = n41616 ;
  assign y20016 = n41624 ;
  assign y20017 = ~n41626 ;
  assign y20018 = n41627 ;
  assign y20019 = ~n41628 ;
  assign y20020 = ~n41630 ;
  assign y20021 = n41632 ;
  assign y20022 = ~1'b0 ;
  assign y20023 = n41634 ;
  assign y20024 = n29577 ;
  assign y20025 = ~1'b0 ;
  assign y20026 = ~1'b0 ;
  assign y20027 = ~n41635 ;
  assign y20028 = ~n41636 ;
  assign y20029 = ~n41637 ;
  assign y20030 = ~n41643 ;
  assign y20031 = ~n10218 ;
  assign y20032 = ~n41644 ;
  assign y20033 = n41647 ;
  assign y20034 = ~n41648 ;
  assign y20035 = n41653 ;
  assign y20036 = ~1'b0 ;
  assign y20037 = ~1'b0 ;
  assign y20038 = ~n41654 ;
  assign y20039 = n41656 ;
  assign y20040 = n41657 ;
  assign y20041 = n41661 ;
  assign y20042 = ~n41662 ;
  assign y20043 = ~n41666 ;
  assign y20044 = 1'b0 ;
  assign y20045 = n41668 ;
  assign y20046 = ~n41672 ;
  assign y20047 = ~n41673 ;
  assign y20048 = ~n41674 ;
  assign y20049 = n41675 ;
  assign y20050 = n9582 ;
  assign y20051 = ~n41676 ;
  assign y20052 = ~n41680 ;
  assign y20053 = n41681 ;
  assign y20054 = 1'b0 ;
  assign y20055 = ~n41682 ;
  assign y20056 = ~n41684 ;
  assign y20057 = n41686 ;
  assign y20058 = n41688 ;
  assign y20059 = ~n41690 ;
  assign y20060 = ~n41691 ;
  assign y20061 = n41695 ;
  assign y20062 = ~n41696 ;
  assign y20063 = n41697 ;
  assign y20064 = n41699 ;
  assign y20065 = ~1'b0 ;
  assign y20066 = ~1'b0 ;
  assign y20067 = ~n41705 ;
  assign y20068 = ~n41713 ;
  assign y20069 = ~n41715 ;
  assign y20070 = ~n41718 ;
  assign y20071 = ~n41720 ;
  assign y20072 = ~1'b0 ;
  assign y20073 = ~n41723 ;
  assign y20074 = ~n41724 ;
  assign y20075 = n41725 ;
  assign y20076 = ~n41728 ;
  assign y20077 = n41729 ;
  assign y20078 = n22081 ;
  assign y20079 = n41737 ;
  assign y20080 = ~n41738 ;
  assign y20081 = ~n8080 ;
  assign y20082 = ~1'b0 ;
  assign y20083 = ~n20996 ;
  assign y20084 = ~n36023 ;
  assign y20085 = ~n41740 ;
  assign y20086 = n41746 ;
  assign y20087 = ~n41747 ;
  assign y20088 = ~n41748 ;
  assign y20089 = ~n41750 ;
  assign y20090 = n41753 ;
  assign y20091 = ~n41755 ;
  assign y20092 = ~1'b0 ;
  assign y20093 = ~n41758 ;
  assign y20094 = n41764 ;
  assign y20095 = ~n41768 ;
  assign y20096 = n41769 ;
  assign y20097 = n41770 ;
  assign y20098 = n41771 ;
  assign y20099 = ~n41772 ;
  assign y20100 = n41775 ;
  assign y20101 = n41778 ;
  assign y20102 = n41781 ;
  assign y20103 = ~n41783 ;
  assign y20104 = ~1'b0 ;
  assign y20105 = ~n41785 ;
  assign y20106 = ~1'b0 ;
  assign y20107 = n41786 ;
  assign y20108 = ~n41790 ;
  assign y20109 = ~n41791 ;
  assign y20110 = n41792 ;
  assign y20111 = ~n41795 ;
  assign y20112 = ~n41800 ;
  assign y20113 = n41802 ;
  assign y20114 = ~n41807 ;
  assign y20115 = ~n41809 ;
  assign y20116 = ~1'b0 ;
  assign y20117 = ~n41814 ;
  assign y20118 = n41819 ;
  assign y20119 = n41822 ;
  assign y20120 = ~n41829 ;
  assign y20121 = n41831 ;
  assign y20122 = n41838 ;
  assign y20123 = ~1'b0 ;
  assign y20124 = ~1'b0 ;
  assign y20125 = ~1'b0 ;
  assign y20126 = ~n41841 ;
  assign y20127 = ~n41842 ;
  assign y20128 = n41844 ;
  assign y20129 = ~n41845 ;
  assign y20130 = n41848 ;
  assign y20131 = ~n41851 ;
  assign y20132 = ~n41853 ;
  assign y20133 = ~n41855 ;
  assign y20134 = n41858 ;
  assign y20135 = n41859 ;
  assign y20136 = ~n41860 ;
  assign y20137 = n41861 ;
  assign y20138 = n41862 ;
  assign y20139 = n10743 ;
  assign y20140 = n41863 ;
  assign y20141 = n41865 ;
  assign y20142 = ~n41869 ;
  assign y20143 = ~n6851 ;
  assign y20144 = ~n41877 ;
  assign y20145 = n41878 ;
  assign y20146 = ~n41879 ;
  assign y20147 = ~n41883 ;
  assign y20148 = ~1'b0 ;
  assign y20149 = ~n41885 ;
  assign y20150 = ~n41886 ;
  assign y20151 = ~1'b0 ;
  assign y20152 = ~n41888 ;
  assign y20153 = ~1'b0 ;
  assign y20154 = n41890 ;
  assign y20155 = ~n41892 ;
  assign y20156 = n41895 ;
  assign y20157 = ~n41897 ;
  assign y20158 = ~n41899 ;
  assign y20159 = n41900 ;
  assign y20160 = n41901 ;
  assign y20161 = n41908 ;
  assign y20162 = ~n41911 ;
  assign y20163 = ~n41913 ;
  assign y20164 = ~1'b0 ;
  assign y20165 = n41914 ;
  assign y20166 = ~n41917 ;
  assign y20167 = n41919 ;
  assign y20168 = ~n41921 ;
  assign y20169 = n41922 ;
  assign y20170 = ~1'b0 ;
  assign y20171 = ~n18449 ;
  assign y20172 = ~1'b0 ;
  assign y20173 = n41926 ;
  assign y20174 = ~n41927 ;
  assign y20175 = n41930 ;
  assign y20176 = ~1'b0 ;
  assign y20177 = n41936 ;
  assign y20178 = ~n41937 ;
  assign y20179 = ~n41938 ;
  assign y20180 = ~n41939 ;
  assign y20181 = ~1'b0 ;
  assign y20182 = ~n41940 ;
  assign y20183 = n5217 ;
  assign y20184 = n41942 ;
  assign y20185 = ~n41946 ;
  assign y20186 = ~1'b0 ;
  assign y20187 = ~1'b0 ;
  assign y20188 = ~n41949 ;
  assign y20189 = ~n41950 ;
  assign y20190 = ~n41954 ;
  assign y20191 = ~n41955 ;
  assign y20192 = ~n41962 ;
  assign y20193 = n41963 ;
  assign y20194 = ~1'b0 ;
  assign y20195 = n41965 ;
  assign y20196 = ~n3000 ;
  assign y20197 = ~1'b0 ;
  assign y20198 = ~n41968 ;
  assign y20199 = ~1'b0 ;
  assign y20200 = ~n4902 ;
  assign y20201 = ~n41971 ;
  assign y20202 = ~1'b0 ;
  assign y20203 = ~n41973 ;
  assign y20204 = ~1'b0 ;
  assign y20205 = ~1'b0 ;
  assign y20206 = ~n41974 ;
  assign y20207 = n41979 ;
  assign y20208 = ~n41981 ;
  assign y20209 = ~n41982 ;
  assign y20210 = n41986 ;
  assign y20211 = ~n41992 ;
  assign y20212 = ~n41995 ;
  assign y20213 = n41998 ;
  assign y20214 = 1'b0 ;
  assign y20215 = ~1'b0 ;
  assign y20216 = ~n42000 ;
  assign y20217 = n42004 ;
  assign y20218 = n42008 ;
  assign y20219 = n42010 ;
  assign y20220 = n42013 ;
  assign y20221 = ~n42014 ;
  assign y20222 = ~n42015 ;
  assign y20223 = n42016 ;
  assign y20224 = ~n42019 ;
  assign y20225 = ~n42021 ;
  assign y20226 = ~1'b0 ;
  assign y20227 = n42022 ;
  assign y20228 = ~n42023 ;
  assign y20229 = ~1'b0 ;
  assign y20230 = ~n42030 ;
  assign y20231 = n42031 ;
  assign y20232 = n42032 ;
  assign y20233 = ~n42038 ;
  assign y20234 = n42040 ;
  assign y20235 = n5452 ;
  assign y20236 = ~1'b0 ;
  assign y20237 = n42041 ;
  assign y20238 = n42045 ;
  assign y20239 = 1'b0 ;
  assign y20240 = ~n42047 ;
  assign y20241 = ~n42048 ;
  assign y20242 = n42051 ;
  assign y20243 = n42055 ;
  assign y20244 = ~n42056 ;
  assign y20245 = ~1'b0 ;
  assign y20246 = n42057 ;
  assign y20247 = ~1'b0 ;
  assign y20248 = ~1'b0 ;
  assign y20249 = n42058 ;
  assign y20250 = ~n42063 ;
  assign y20251 = ~n42064 ;
  assign y20252 = ~n42066 ;
  assign y20253 = ~n42069 ;
  assign y20254 = ~1'b0 ;
  assign y20255 = ~1'b0 ;
  assign y20256 = ~n42072 ;
  assign y20257 = ~n42074 ;
  assign y20258 = ~n42078 ;
  assign y20259 = ~n42079 ;
  assign y20260 = ~n42082 ;
  assign y20261 = n42084 ;
  assign y20262 = ~1'b0 ;
  assign y20263 = ~n42088 ;
  assign y20264 = n42089 ;
  assign y20265 = ~n42091 ;
  assign y20266 = n42093 ;
  assign y20267 = ~n42096 ;
  assign y20268 = ~1'b0 ;
  assign y20269 = ~1'b0 ;
  assign y20270 = ~n42098 ;
  assign y20271 = 1'b0 ;
  assign y20272 = ~n42100 ;
  assign y20273 = ~n42102 ;
  assign y20274 = n42104 ;
  assign y20275 = ~n42109 ;
  assign y20276 = ~n42111 ;
  assign y20277 = ~1'b0 ;
  assign y20278 = ~n42113 ;
  assign y20279 = ~n42120 ;
  assign y20280 = ~n42122 ;
  assign y20281 = ~n42126 ;
  assign y20282 = ~n32418 ;
  assign y20283 = ~n42132 ;
  assign y20284 = ~n42134 ;
  assign y20285 = ~n2155 ;
  assign y20286 = ~1'b0 ;
  assign y20287 = ~1'b0 ;
  assign y20288 = ~1'b0 ;
  assign y20289 = ~1'b0 ;
  assign y20290 = ~n42141 ;
  assign y20291 = ~n42142 ;
  assign y20292 = ~n42145 ;
  assign y20293 = n42146 ;
  assign y20294 = ~n42150 ;
  assign y20295 = n42152 ;
  assign y20296 = ~n42156 ;
  assign y20297 = 1'b0 ;
  assign y20298 = ~n42158 ;
  assign y20299 = n42159 ;
  assign y20300 = ~1'b0 ;
  assign y20301 = ~n42161 ;
  assign y20302 = n42163 ;
  assign y20303 = ~n21394 ;
  assign y20304 = ~n42164 ;
  assign y20305 = n42166 ;
  assign y20306 = ~n42168 ;
  assign y20307 = n42172 ;
  assign y20308 = ~n42175 ;
  assign y20309 = ~n42177 ;
  assign y20310 = ~1'b0 ;
  assign y20311 = n42179 ;
  assign y20312 = n42180 ;
  assign y20313 = n42185 ;
  assign y20314 = ~n42186 ;
  assign y20315 = ~n42187 ;
  assign y20316 = n42192 ;
  assign y20317 = ~1'b0 ;
  assign y20318 = n42195 ;
  assign y20319 = n42196 ;
  assign y20320 = ~1'b0 ;
  assign y20321 = n42198 ;
  assign y20322 = n42204 ;
  assign y20323 = n42205 ;
  assign y20324 = n42206 ;
  assign y20325 = ~n20509 ;
  assign y20326 = ~n42207 ;
  assign y20327 = n42211 ;
  assign y20328 = ~1'b0 ;
  assign y20329 = ~n42213 ;
  assign y20330 = ~n42215 ;
  assign y20331 = ~1'b0 ;
  assign y20332 = ~1'b0 ;
  assign y20333 = ~n42216 ;
  assign y20334 = n42218 ;
  assign y20335 = n42220 ;
  assign y20336 = ~1'b0 ;
  assign y20337 = ~n42222 ;
  assign y20338 = ~n42226 ;
  assign y20339 = ~n42227 ;
  assign y20340 = n42229 ;
  assign y20341 = n42235 ;
  assign y20342 = n42240 ;
  assign y20343 = ~1'b0 ;
  assign y20344 = ~n42241 ;
  assign y20345 = n42243 ;
  assign y20346 = n42246 ;
  assign y20347 = n42248 ;
  assign y20348 = ~n42254 ;
  assign y20349 = ~1'b0 ;
  assign y20350 = ~n42255 ;
  assign y20351 = n42270 ;
  assign y20352 = n34530 ;
  assign y20353 = ~1'b0 ;
  assign y20354 = n42271 ;
  assign y20355 = ~n42275 ;
  assign y20356 = n42279 ;
  assign y20357 = ~n42280 ;
  assign y20358 = ~n42284 ;
  assign y20359 = n42285 ;
  assign y20360 = n42287 ;
  assign y20361 = ~1'b0 ;
  assign y20362 = ~1'b0 ;
  assign y20363 = ~1'b0 ;
  assign y20364 = n42291 ;
  assign y20365 = n42298 ;
  assign y20366 = ~n42301 ;
  assign y20367 = ~n42305 ;
  assign y20368 = ~1'b0 ;
  assign y20369 = ~n42310 ;
  assign y20370 = ~n42312 ;
  assign y20371 = n42316 ;
  assign y20372 = ~n42319 ;
  assign y20373 = ~1'b0 ;
  assign y20374 = n15284 ;
  assign y20375 = n42326 ;
  assign y20376 = n42327 ;
  assign y20377 = ~1'b0 ;
  assign y20378 = ~n42330 ;
  assign y20379 = ~n42334 ;
  assign y20380 = n42336 ;
  assign y20381 = n42339 ;
  assign y20382 = ~1'b0 ;
  assign y20383 = ~n42341 ;
  assign y20384 = n42343 ;
  assign y20385 = n42344 ;
  assign y20386 = ~n42346 ;
  assign y20387 = ~n42349 ;
  assign y20388 = ~1'b0 ;
  assign y20389 = n42351 ;
  assign y20390 = ~n42353 ;
  assign y20391 = ~n42358 ;
  assign y20392 = ~1'b0 ;
  assign y20393 = ~1'b0 ;
  assign y20394 = n42359 ;
  assign y20395 = ~n42364 ;
  assign y20396 = ~n42365 ;
  assign y20397 = ~1'b0 ;
  assign y20398 = ~n42369 ;
  assign y20399 = ~1'b0 ;
  assign y20400 = ~n42371 ;
  assign y20401 = n42373 ;
  assign y20402 = ~n42378 ;
  assign y20403 = n42380 ;
  assign y20404 = ~n42382 ;
  assign y20405 = n42383 ;
  assign y20406 = ~n42385 ;
  assign y20407 = ~n42387 ;
  assign y20408 = ~n42388 ;
  assign y20409 = ~1'b0 ;
  assign y20410 = ~n42389 ;
  assign y20411 = ~n42392 ;
  assign y20412 = ~1'b0 ;
  assign y20413 = ~1'b0 ;
  assign y20414 = ~n42393 ;
  assign y20415 = n42398 ;
  assign y20416 = ~n42399 ;
  assign y20417 = ~n42400 ;
  assign y20418 = ~n42402 ;
  assign y20419 = ~n42405 ;
  assign y20420 = ~1'b0 ;
  assign y20421 = n42408 ;
  assign y20422 = ~1'b0 ;
  assign y20423 = n42409 ;
  assign y20424 = n42410 ;
  assign y20425 = n42411 ;
  assign y20426 = ~n42414 ;
  assign y20427 = ~n42415 ;
  assign y20428 = ~1'b0 ;
  assign y20429 = n42416 ;
  assign y20430 = ~1'b0 ;
  assign y20431 = ~1'b0 ;
  assign y20432 = n42419 ;
  assign y20433 = n42422 ;
  assign y20434 = n42424 ;
  assign y20435 = ~n42427 ;
  assign y20436 = ~1'b0 ;
  assign y20437 = ~n42429 ;
  assign y20438 = ~1'b0 ;
  assign y20439 = ~1'b0 ;
  assign y20440 = n42431 ;
  assign y20441 = ~n42434 ;
  assign y20442 = n793 ;
  assign y20443 = ~n42436 ;
  assign y20444 = n42438 ;
  assign y20445 = n30261 ;
  assign y20446 = n42440 ;
  assign y20447 = ~n42442 ;
  assign y20448 = ~1'b0 ;
  assign y20449 = n22268 ;
  assign y20450 = ~n42443 ;
  assign y20451 = 1'b0 ;
  assign y20452 = ~n42444 ;
  assign y20453 = ~n42445 ;
  assign y20454 = n42446 ;
  assign y20455 = ~n42452 ;
  assign y20456 = ~1'b0 ;
  assign y20457 = ~n2012 ;
  assign y20458 = ~n42454 ;
  assign y20459 = ~1'b0 ;
  assign y20460 = n11653 ;
  assign y20461 = n42455 ;
  assign y20462 = n42460 ;
  assign y20463 = ~n42463 ;
  assign y20464 = n42476 ;
  assign y20465 = ~n19429 ;
  assign y20466 = ~n42480 ;
  assign y20467 = ~1'b0 ;
  assign y20468 = ~1'b0 ;
  assign y20469 = ~n42482 ;
  assign y20470 = ~n42484 ;
  assign y20471 = ~1'b0 ;
  assign y20472 = n42485 ;
  assign y20473 = ~n42486 ;
  assign y20474 = ~n14574 ;
  assign y20475 = n42487 ;
  assign y20476 = ~n12118 ;
  assign y20477 = 1'b0 ;
  assign y20478 = ~1'b0 ;
  assign y20479 = n32185 ;
  assign y20480 = ~n42491 ;
  assign y20481 = ~n42494 ;
  assign y20482 = n42495 ;
  assign y20483 = n42499 ;
  assign y20484 = ~n42503 ;
  assign y20485 = ~n42504 ;
  assign y20486 = ~1'b0 ;
  assign y20487 = ~n42505 ;
  assign y20488 = ~n42510 ;
  assign y20489 = n42513 ;
  assign y20490 = n42517 ;
  assign y20491 = n42518 ;
  assign y20492 = ~n42519 ;
  assign y20493 = ~1'b0 ;
  assign y20494 = n42524 ;
  assign y20495 = n42532 ;
  assign y20496 = 1'b0 ;
  assign y20497 = ~n42535 ;
  assign y20498 = ~1'b0 ;
  assign y20499 = ~1'b0 ;
  assign y20500 = ~n42537 ;
  assign y20501 = ~n42538 ;
  assign y20502 = n652 ;
  assign y20503 = ~n42542 ;
  assign y20504 = ~1'b0 ;
  assign y20505 = ~1'b0 ;
  assign y20506 = ~1'b0 ;
  assign y20507 = n42547 ;
  assign y20508 = ~n42551 ;
  assign y20509 = n42557 ;
  assign y20510 = n42558 ;
  assign y20511 = ~n42560 ;
  assign y20512 = ~1'b0 ;
  assign y20513 = ~1'b0 ;
  assign y20514 = ~1'b0 ;
  assign y20515 = ~1'b0 ;
  assign y20516 = ~1'b0 ;
  assign y20517 = ~1'b0 ;
  assign y20518 = n42561 ;
  assign y20519 = ~n26404 ;
  assign y20520 = ~1'b0 ;
  assign y20521 = ~1'b0 ;
  assign y20522 = n42563 ;
  assign y20523 = n42567 ;
  assign y20524 = ~n42573 ;
  assign y20525 = n9715 ;
  assign y20526 = n42578 ;
  assign y20527 = ~n42579 ;
  assign y20528 = ~n42580 ;
  assign y20529 = ~n42581 ;
  assign y20530 = ~n42582 ;
  assign y20531 = ~1'b0 ;
  assign y20532 = ~1'b0 ;
  assign y20533 = n42583 ;
  assign y20534 = ~1'b0 ;
  assign y20535 = ~1'b0 ;
  assign y20536 = ~1'b0 ;
  assign y20537 = ~n42586 ;
  assign y20538 = ~n42587 ;
  assign y20539 = ~n42588 ;
  assign y20540 = ~n42590 ;
  assign y20541 = ~n42591 ;
  assign y20542 = ~n42595 ;
  assign y20543 = ~n10592 ;
  assign y20544 = n42597 ;
  assign y20545 = ~n42599 ;
  assign y20546 = ~1'b0 ;
  assign y20547 = ~n42601 ;
  assign y20548 = ~n42603 ;
  assign y20549 = ~n42606 ;
  assign y20550 = ~n42607 ;
  assign y20551 = ~1'b0 ;
  assign y20552 = ~n42609 ;
  assign y20553 = ~n42611 ;
  assign y20554 = n42614 ;
  assign y20555 = ~1'b0 ;
  assign y20556 = ~n8363 ;
  assign y20557 = n42616 ;
  assign y20558 = ~n42618 ;
  assign y20559 = n42620 ;
  assign y20560 = ~1'b0 ;
  assign y20561 = ~1'b0 ;
  assign y20562 = n42625 ;
  assign y20563 = ~n42626 ;
  assign y20564 = ~1'b0 ;
  assign y20565 = n42633 ;
  assign y20566 = n42635 ;
  assign y20567 = ~n42638 ;
  assign y20568 = ~n42640 ;
  assign y20569 = ~1'b0 ;
  assign y20570 = ~n42643 ;
  assign y20571 = ~1'b0 ;
  assign y20572 = ~1'b0 ;
  assign y20573 = 1'b0 ;
  assign y20574 = ~1'b0 ;
  assign y20575 = ~n42651 ;
  assign y20576 = ~n42652 ;
  assign y20577 = ~n42654 ;
  assign y20578 = ~1'b0 ;
  assign y20579 = ~1'b0 ;
  assign y20580 = n42656 ;
  assign y20581 = ~n8526 ;
  assign y20582 = 1'b0 ;
  assign y20583 = ~1'b0 ;
  assign y20584 = n42658 ;
  assign y20585 = n42659 ;
  assign y20586 = n42661 ;
  assign y20587 = ~n42663 ;
  assign y20588 = n42664 ;
  assign y20589 = ~1'b0 ;
  assign y20590 = n9952 ;
  assign y20591 = n42669 ;
  assign y20592 = ~n42670 ;
  assign y20593 = ~1'b0 ;
  assign y20594 = n42671 ;
  assign y20595 = n42675 ;
  assign y20596 = n42678 ;
  assign y20597 = n42684 ;
  assign y20598 = ~n42685 ;
  assign y20599 = ~n42687 ;
  assign y20600 = n42688 ;
  assign y20601 = ~n3558 ;
  assign y20602 = ~n42690 ;
  assign y20603 = ~1'b0 ;
  assign y20604 = ~1'b0 ;
  assign y20605 = 1'b0 ;
  assign y20606 = n35168 ;
  assign y20607 = ~n42696 ;
  assign y20608 = ~n42699 ;
  assign y20609 = n42702 ;
  assign y20610 = ~1'b0 ;
  assign y20611 = n42704 ;
  assign y20612 = ~1'b0 ;
  assign y20613 = n42707 ;
  assign y20614 = ~1'b0 ;
  assign y20615 = ~1'b0 ;
  assign y20616 = ~1'b0 ;
  assign y20617 = n42710 ;
  assign y20618 = ~n42712 ;
  assign y20619 = n42713 ;
  assign y20620 = ~n42714 ;
  assign y20621 = ~1'b0 ;
  assign y20622 = n42715 ;
  assign y20623 = ~n42716 ;
  assign y20624 = ~1'b0 ;
  assign y20625 = ~1'b0 ;
  assign y20626 = n467 ;
  assign y20627 = ~n42717 ;
  assign y20628 = n38530 ;
  assign y20629 = n42720 ;
  assign y20630 = n42727 ;
  assign y20631 = n42732 ;
  assign y20632 = ~1'b0 ;
  assign y20633 = ~1'b0 ;
  assign y20634 = ~n42735 ;
  assign y20635 = n42736 ;
  assign y20636 = ~n42737 ;
  assign y20637 = n42741 ;
  assign y20638 = ~1'b0 ;
  assign y20639 = ~n42743 ;
  assign y20640 = ~n42745 ;
  assign y20641 = ~n42750 ;
  assign y20642 = ~n42753 ;
  assign y20643 = ~n42756 ;
  assign y20644 = ~n42757 ;
  assign y20645 = ~n42759 ;
  assign y20646 = ~1'b0 ;
  assign y20647 = ~1'b0 ;
  assign y20648 = n30330 ;
  assign y20649 = n42763 ;
  assign y20650 = ~n42764 ;
  assign y20651 = ~n42765 ;
  assign y20652 = ~1'b0 ;
  assign y20653 = ~1'b0 ;
  assign y20654 = ~n42769 ;
  assign y20655 = n42771 ;
  assign y20656 = n42773 ;
  assign y20657 = ~1'b0 ;
  assign y20658 = n42775 ;
  assign y20659 = ~n42776 ;
  assign y20660 = ~n42782 ;
  assign y20661 = ~n42783 ;
  assign y20662 = ~n38355 ;
  assign y20663 = ~1'b0 ;
  assign y20664 = ~n42786 ;
  assign y20665 = ~n42788 ;
  assign y20666 = ~n42789 ;
  assign y20667 = ~1'b0 ;
  assign y20668 = ~1'b0 ;
  assign y20669 = ~n42790 ;
  assign y20670 = n42793 ;
  assign y20671 = ~n42794 ;
  assign y20672 = ~n42795 ;
  assign y20673 = ~n42797 ;
  assign y20674 = ~1'b0 ;
  assign y20675 = ~1'b0 ;
  assign y20676 = ~n42803 ;
  assign y20677 = ~n42805 ;
  assign y20678 = n42806 ;
  assign y20679 = ~n42811 ;
  assign y20680 = ~n42812 ;
  assign y20681 = ~n42814 ;
  assign y20682 = 1'b0 ;
  assign y20683 = ~1'b0 ;
  assign y20684 = ~1'b0 ;
  assign y20685 = ~n42819 ;
  assign y20686 = ~1'b0 ;
  assign y20687 = n42821 ;
  assign y20688 = ~n42822 ;
  assign y20689 = n42823 ;
  assign y20690 = n42825 ;
  assign y20691 = n42826 ;
  assign y20692 = ~1'b0 ;
  assign y20693 = ~n42830 ;
  assign y20694 = ~n42831 ;
  assign y20695 = ~1'b0 ;
  assign y20696 = n42837 ;
  assign y20697 = n42839 ;
  assign y20698 = ~n42843 ;
  assign y20699 = n42844 ;
  assign y20700 = n42846 ;
  assign y20701 = ~1'b0 ;
  assign y20702 = ~n42848 ;
  assign y20703 = ~n42850 ;
  assign y20704 = n42851 ;
  assign y20705 = n42852 ;
  assign y20706 = ~1'b0 ;
  assign y20707 = ~1'b0 ;
  assign y20708 = ~1'b0 ;
  assign y20709 = ~n42853 ;
  assign y20710 = n42855 ;
  assign y20711 = n42858 ;
  assign y20712 = n42859 ;
  assign y20713 = n42861 ;
  assign y20714 = n2801 ;
  assign y20715 = ~1'b0 ;
  assign y20716 = ~1'b0 ;
  assign y20717 = ~1'b0 ;
  assign y20718 = ~n42864 ;
  assign y20719 = n42865 ;
  assign y20720 = ~n42867 ;
  assign y20721 = n42869 ;
  assign y20722 = n42873 ;
  assign y20723 = ~1'b0 ;
  assign y20724 = n42877 ;
  assign y20725 = n42878 ;
  assign y20726 = ~n16362 ;
  assign y20727 = ~1'b0 ;
  assign y20728 = ~n42879 ;
  assign y20729 = n42884 ;
  assign y20730 = ~n42887 ;
  assign y20731 = n42888 ;
  assign y20732 = ~n42890 ;
  assign y20733 = ~1'b0 ;
  assign y20734 = n42891 ;
  assign y20735 = n42893 ;
  assign y20736 = ~1'b0 ;
  assign y20737 = n42895 ;
  assign y20738 = ~n42899 ;
  assign y20739 = ~n42902 ;
  assign y20740 = n42903 ;
  assign y20741 = n42905 ;
  assign y20742 = ~n42908 ;
  assign y20743 = n42913 ;
  assign y20744 = n42915 ;
  assign y20745 = ~n42919 ;
  assign y20746 = ~1'b0 ;
  assign y20747 = ~n42922 ;
  assign y20748 = 1'b0 ;
  assign y20749 = ~1'b0 ;
  assign y20750 = ~n28378 ;
  assign y20751 = n42926 ;
  assign y20752 = ~n42927 ;
  assign y20753 = ~n42929 ;
  assign y20754 = ~1'b0 ;
  assign y20755 = n42932 ;
  assign y20756 = ~n7710 ;
  assign y20757 = ~n42934 ;
  assign y20758 = n42936 ;
  assign y20759 = ~1'b0 ;
  assign y20760 = ~n42937 ;
  assign y20761 = ~n42940 ;
  assign y20762 = n42941 ;
  assign y20763 = ~n42943 ;
  assign y20764 = ~1'b0 ;
  assign y20765 = ~n42945 ;
  assign y20766 = n42952 ;
  assign y20767 = ~1'b0 ;
  assign y20768 = n42953 ;
  assign y20769 = 1'b0 ;
  assign y20770 = ~n42957 ;
  assign y20771 = n42958 ;
  assign y20772 = n25766 ;
  assign y20773 = n42959 ;
  assign y20774 = n42960 ;
  assign y20775 = ~n42963 ;
  assign y20776 = n42964 ;
  assign y20777 = n42965 ;
  assign y20778 = ~n42969 ;
  assign y20779 = n42970 ;
  assign y20780 = n42973 ;
  assign y20781 = ~n42975 ;
  assign y20782 = n42978 ;
  assign y20783 = ~1'b0 ;
  assign y20784 = ~n19393 ;
  assign y20785 = n42982 ;
  assign y20786 = ~n42985 ;
  assign y20787 = ~n42989 ;
  assign y20788 = n42990 ;
  assign y20789 = ~n29322 ;
  assign y20790 = n42994 ;
  assign y20791 = ~n42996 ;
  assign y20792 = ~1'b0 ;
  assign y20793 = n42997 ;
  assign y20794 = n19069 ;
  assign y20795 = ~1'b0 ;
  assign y20796 = ~n42998 ;
  assign y20797 = ~1'b0 ;
  assign y20798 = ~n42999 ;
  assign y20799 = n43000 ;
  assign y20800 = ~n43002 ;
  assign y20801 = ~n43004 ;
  assign y20802 = ~n43007 ;
  assign y20803 = n15320 ;
  assign y20804 = ~n43008 ;
  assign y20805 = n43011 ;
  assign y20806 = n43015 ;
  assign y20807 = ~1'b0 ;
  assign y20808 = n43017 ;
  assign y20809 = n43019 ;
  assign y20810 = ~n43023 ;
  assign y20811 = ~1'b0 ;
  assign y20812 = ~1'b0 ;
  assign y20813 = ~1'b0 ;
  assign y20814 = n43024 ;
  assign y20815 = n43026 ;
  assign y20816 = n43028 ;
  assign y20817 = n43029 ;
  assign y20818 = n43031 ;
  assign y20819 = n17228 ;
  assign y20820 = ~1'b0 ;
  assign y20821 = n43034 ;
  assign y20822 = ~n43037 ;
  assign y20823 = ~n43038 ;
  assign y20824 = ~n43040 ;
  assign y20825 = ~1'b0 ;
  assign y20826 = ~n43041 ;
  assign y20827 = ~n43042 ;
  assign y20828 = ~n43048 ;
  assign y20829 = n43054 ;
  assign y20830 = ~1'b0 ;
  assign y20831 = ~1'b0 ;
  assign y20832 = ~1'b0 ;
  assign y20833 = ~1'b0 ;
  assign y20834 = ~1'b0 ;
  assign y20835 = n43057 ;
  assign y20836 = ~1'b0 ;
  assign y20837 = ~n43061 ;
  assign y20838 = ~n43068 ;
  assign y20839 = n43070 ;
  assign y20840 = n43072 ;
  assign y20841 = n43073 ;
  assign y20842 = ~1'b0 ;
  assign y20843 = n43075 ;
  assign y20844 = ~1'b0 ;
  assign y20845 = ~n43077 ;
  assign y20846 = ~1'b0 ;
  assign y20847 = n43079 ;
  assign y20848 = ~n43081 ;
  assign y20849 = ~n29375 ;
  assign y20850 = ~n43084 ;
  assign y20851 = n43087 ;
  assign y20852 = ~1'b0 ;
  assign y20853 = n43090 ;
  assign y20854 = n43093 ;
  assign y20855 = ~n43094 ;
  assign y20856 = ~n43095 ;
  assign y20857 = ~1'b0 ;
  assign y20858 = n43097 ;
  assign y20859 = ~n43098 ;
  assign y20860 = ~n43099 ;
  assign y20861 = n26973 ;
  assign y20862 = n43100 ;
  assign y20863 = n43101 ;
  assign y20864 = n43102 ;
  assign y20865 = n43104 ;
  assign y20866 = ~n43106 ;
  assign y20867 = ~n43107 ;
  assign y20868 = n43109 ;
  assign y20869 = ~n43110 ;
  assign y20870 = n43111 ;
  assign y20871 = ~n43115 ;
  assign y20872 = ~1'b0 ;
  assign y20873 = n43116 ;
  assign y20874 = n43117 ;
  assign y20875 = ~n43118 ;
  assign y20876 = ~1'b0 ;
  assign y20877 = n43120 ;
  assign y20878 = n43121 ;
  assign y20879 = n43124 ;
  assign y20880 = ~n43127 ;
  assign y20881 = n43131 ;
  assign y20882 = ~1'b0 ;
  assign y20883 = ~n43134 ;
  assign y20884 = ~1'b0 ;
  assign y20885 = ~n43135 ;
  assign y20886 = ~1'b0 ;
  assign y20887 = ~n43138 ;
  assign y20888 = ~n43140 ;
  assign y20889 = n43144 ;
  assign y20890 = ~n36700 ;
  assign y20891 = ~1'b0 ;
  assign y20892 = ~n20631 ;
  assign y20893 = n43147 ;
  assign y20894 = ~n43148 ;
  assign y20895 = ~1'b0 ;
  assign y20896 = ~1'b0 ;
  assign y20897 = ~n43152 ;
  assign y20898 = n43155 ;
  assign y20899 = ~n43158 ;
  assign y20900 = n43159 ;
  assign y20901 = ~n43163 ;
  assign y20902 = 1'b0 ;
  assign y20903 = n43166 ;
  assign y20904 = n43168 ;
  assign y20905 = ~n43170 ;
  assign y20906 = ~1'b0 ;
  assign y20907 = n43175 ;
  assign y20908 = ~n43176 ;
  assign y20909 = n43177 ;
  assign y20910 = ~n43179 ;
  assign y20911 = ~n43180 ;
  assign y20912 = n43185 ;
  assign y20913 = ~n43189 ;
  assign y20914 = n14079 ;
  assign y20915 = ~n43191 ;
  assign y20916 = n43194 ;
  assign y20917 = ~n43196 ;
  assign y20918 = ~n43200 ;
  assign y20919 = ~n41601 ;
  assign y20920 = n43201 ;
  assign y20921 = n43206 ;
  assign y20922 = ~n43208 ;
  assign y20923 = ~1'b0 ;
  assign y20924 = ~1'b0 ;
  assign y20925 = ~1'b0 ;
  assign y20926 = n43209 ;
  assign y20927 = ~n43210 ;
  assign y20928 = ~1'b0 ;
  assign y20929 = n43211 ;
  assign y20930 = ~1'b0 ;
  assign y20931 = ~n43212 ;
  assign y20932 = ~n43213 ;
  assign y20933 = n43218 ;
  assign y20934 = n43219 ;
  assign y20935 = n31078 ;
  assign y20936 = ~n43220 ;
  assign y20937 = n43221 ;
  assign y20938 = ~1'b0 ;
  assign y20939 = ~n43223 ;
  assign y20940 = ~n43224 ;
  assign y20941 = ~n43226 ;
  assign y20942 = ~n3752 ;
  assign y20943 = n43229 ;
  assign y20944 = n43230 ;
  assign y20945 = ~1'b0 ;
  assign y20946 = ~n43236 ;
  assign y20947 = ~n43239 ;
  assign y20948 = ~n43245 ;
  assign y20949 = n43247 ;
  assign y20950 = ~1'b0 ;
  assign y20951 = ~n43248 ;
  assign y20952 = ~n43249 ;
  assign y20953 = ~n43251 ;
  assign y20954 = n43252 ;
  assign y20955 = ~n43255 ;
  assign y20956 = n43256 ;
  assign y20957 = n43258 ;
  assign y20958 = n43260 ;
  assign y20959 = ~n43262 ;
  assign y20960 = ~1'b0 ;
  assign y20961 = ~1'b0 ;
  assign y20962 = ~n43263 ;
  assign y20963 = n43271 ;
  assign y20964 = ~n43277 ;
  assign y20965 = ~n43283 ;
  assign y20966 = n43285 ;
  assign y20967 = ~n43287 ;
  assign y20968 = ~n43288 ;
  assign y20969 = n43289 ;
  assign y20970 = n43290 ;
  assign y20971 = ~n43293 ;
  assign y20972 = ~n43294 ;
  assign y20973 = ~n43295 ;
  assign y20974 = ~n43296 ;
  assign y20975 = n43297 ;
  assign y20976 = ~n43298 ;
  assign y20977 = ~1'b0 ;
  assign y20978 = n28691 ;
  assign y20979 = ~n43300 ;
  assign y20980 = ~n43302 ;
  assign y20981 = n43304 ;
  assign y20982 = ~n43308 ;
  assign y20983 = ~n43309 ;
  assign y20984 = ~n43312 ;
  assign y20985 = ~1'b0 ;
  assign y20986 = ~1'b0 ;
  assign y20987 = ~1'b0 ;
  assign y20988 = ~n21151 ;
  assign y20989 = ~1'b0 ;
  assign y20990 = n43314 ;
  assign y20991 = ~n20397 ;
  assign y20992 = ~n43315 ;
  assign y20993 = ~1'b0 ;
  assign y20994 = ~1'b0 ;
  assign y20995 = ~1'b0 ;
  assign y20996 = n43317 ;
  assign y20997 = ~n43318 ;
  assign y20998 = ~n43321 ;
  assign y20999 = ~1'b0 ;
  assign y21000 = ~n43325 ;
  assign y21001 = n43328 ;
  assign y21002 = n43339 ;
  assign y21003 = n43340 ;
  assign y21004 = ~n8194 ;
  assign y21005 = n43346 ;
  assign y21006 = ~n43348 ;
  assign y21007 = n43357 ;
  assign y21008 = n43359 ;
  assign y21009 = ~1'b0 ;
  assign y21010 = ~1'b0 ;
  assign y21011 = ~n43360 ;
  assign y21012 = ~n43361 ;
  assign y21013 = ~n43364 ;
  assign y21014 = 1'b0 ;
  assign y21015 = ~n43366 ;
  assign y21016 = ~n43369 ;
  assign y21017 = ~n43371 ;
  assign y21018 = n24007 ;
  assign y21019 = ~n636 ;
  assign y21020 = 1'b0 ;
  assign y21021 = ~1'b0 ;
  assign y21022 = n43374 ;
  assign y21023 = n43375 ;
  assign y21024 = n43376 ;
  assign y21025 = n22694 ;
  assign y21026 = ~n43377 ;
  assign y21027 = ~1'b0 ;
  assign y21028 = n43381 ;
  assign y21029 = n43382 ;
  assign y21030 = ~1'b0 ;
  assign y21031 = ~n43384 ;
  assign y21032 = ~n43385 ;
  assign y21033 = ~1'b0 ;
  assign y21034 = n43393 ;
  assign y21035 = ~n43395 ;
  assign y21036 = n43399 ;
  assign y21037 = n43401 ;
  assign y21038 = ~1'b0 ;
  assign y21039 = ~1'b0 ;
  assign y21040 = ~n43404 ;
  assign y21041 = ~n43407 ;
  assign y21042 = n43408 ;
  assign y21043 = n43410 ;
  assign y21044 = n43412 ;
  assign y21045 = n43413 ;
  assign y21046 = 1'b0 ;
  assign y21047 = ~1'b0 ;
  assign y21048 = ~n43414 ;
  assign y21049 = ~n43420 ;
  assign y21050 = n43421 ;
  assign y21051 = ~1'b0 ;
  assign y21052 = n43422 ;
  assign y21053 = ~1'b0 ;
  assign y21054 = ~n43423 ;
  assign y21055 = n43425 ;
  assign y21056 = ~n43428 ;
  assign y21057 = n41055 ;
  assign y21058 = n43430 ;
  assign y21059 = ~n43431 ;
  assign y21060 = ~n43434 ;
  assign y21061 = n43436 ;
  assign y21062 = n43438 ;
  assign y21063 = n43440 ;
  assign y21064 = ~n43442 ;
  assign y21065 = n43445 ;
  assign y21066 = n43447 ;
  assign y21067 = n43448 ;
  assign y21068 = n43450 ;
  assign y21069 = n43451 ;
  assign y21070 = n43452 ;
  assign y21071 = n43454 ;
  assign y21072 = n43455 ;
  assign y21073 = ~1'b0 ;
  assign y21074 = n43457 ;
  assign y21075 = ~n43458 ;
  assign y21076 = n43460 ;
  assign y21077 = ~n43462 ;
  assign y21078 = ~n43463 ;
  assign y21079 = ~n43465 ;
  assign y21080 = ~n43470 ;
  assign y21081 = ~n43472 ;
  assign y21082 = ~1'b0 ;
  assign y21083 = ~n43474 ;
  assign y21084 = 1'b0 ;
  assign y21085 = ~n43475 ;
  assign y21086 = n43476 ;
  assign y21087 = n11274 ;
  assign y21088 = n43478 ;
  assign y21089 = n43479 ;
  assign y21090 = ~1'b0 ;
  assign y21091 = ~1'b0 ;
  assign y21092 = ~1'b0 ;
  assign y21093 = ~1'b0 ;
  assign y21094 = n43481 ;
  assign y21095 = n43485 ;
  assign y21096 = ~n43489 ;
  assign y21097 = n43490 ;
  assign y21098 = n43492 ;
  assign y21099 = ~n43498 ;
  assign y21100 = n43500 ;
  assign y21101 = n36188 ;
  assign y21102 = n43502 ;
  assign y21103 = ~1'b0 ;
  assign y21104 = ~n43507 ;
  assign y21105 = ~1'b0 ;
  assign y21106 = ~1'b0 ;
  assign y21107 = ~n43508 ;
  assign y21108 = ~n20651 ;
  assign y21109 = ~n43509 ;
  assign y21110 = ~n43512 ;
  assign y21111 = n43514 ;
  assign y21112 = ~n43516 ;
  assign y21113 = ~n43517 ;
  assign y21114 = ~n43522 ;
  assign y21115 = ~n43525 ;
  assign y21116 = ~n43527 ;
  assign y21117 = ~n43531 ;
  assign y21118 = n43533 ;
  assign y21119 = n43534 ;
  assign y21120 = ~n43535 ;
  assign y21121 = n43536 ;
  assign y21122 = ~1'b0 ;
  assign y21123 = ~1'b0 ;
  assign y21124 = ~n43542 ;
  assign y21125 = ~n43544 ;
  assign y21126 = ~n14380 ;
  assign y21127 = ~n43546 ;
  assign y21128 = n43548 ;
  assign y21129 = ~x241 ;
  assign y21130 = n43549 ;
  assign y21131 = n43552 ;
  assign y21132 = ~n43554 ;
  assign y21133 = n43556 ;
  assign y21134 = ~1'b0 ;
  assign y21135 = ~n43557 ;
  assign y21136 = ~n43561 ;
  assign y21137 = ~n43563 ;
  assign y21138 = ~1'b0 ;
  assign y21139 = ~n43564 ;
  assign y21140 = ~n43565 ;
  assign y21141 = n43566 ;
  assign y21142 = n42506 ;
  assign y21143 = 1'b0 ;
  assign y21144 = n43571 ;
  assign y21145 = ~n43573 ;
  assign y21146 = ~1'b0 ;
  assign y21147 = ~n43575 ;
  assign y21148 = n43576 ;
  assign y21149 = n43577 ;
  assign y21150 = ~n43580 ;
  assign y21151 = ~n43583 ;
  assign y21152 = n43593 ;
  assign y21153 = n43594 ;
  assign y21154 = ~1'b0 ;
  assign y21155 = ~n43598 ;
  assign y21156 = ~1'b0 ;
  assign y21157 = ~1'b0 ;
  assign y21158 = n43602 ;
  assign y21159 = ~n43603 ;
  assign y21160 = ~n43605 ;
  assign y21161 = n43606 ;
  assign y21162 = n43609 ;
  assign y21163 = n43611 ;
  assign y21164 = ~n43613 ;
  assign y21165 = ~n43617 ;
  assign y21166 = ~1'b0 ;
  assign y21167 = ~n43620 ;
  assign y21168 = ~n43623 ;
  assign y21169 = ~n33397 ;
  assign y21170 = n43628 ;
  assign y21171 = n43630 ;
  assign y21172 = ~n43631 ;
  assign y21173 = ~n43633 ;
  assign y21174 = ~n43637 ;
  assign y21175 = n43641 ;
  assign y21176 = ~n43643 ;
  assign y21177 = n7607 ;
  assign y21178 = ~n43647 ;
  assign y21179 = n43648 ;
  assign y21180 = n43649 ;
  assign y21181 = ~n43650 ;
  assign y21182 = ~1'b0 ;
  assign y21183 = ~n43653 ;
  assign y21184 = n23786 ;
  assign y21185 = ~n43654 ;
  assign y21186 = ~1'b0 ;
  assign y21187 = ~1'b0 ;
  assign y21188 = ~n43655 ;
  assign y21189 = n43657 ;
  assign y21190 = ~n43660 ;
  assign y21191 = n43667 ;
  assign y21192 = ~1'b0 ;
  assign y21193 = ~n43669 ;
  assign y21194 = n43672 ;
  assign y21195 = ~n43674 ;
  assign y21196 = n43681 ;
  assign y21197 = ~n43682 ;
  assign y21198 = n43683 ;
  assign y21199 = n43684 ;
  assign y21200 = n43688 ;
  assign y21201 = n43692 ;
  assign y21202 = ~1'b0 ;
  assign y21203 = ~1'b0 ;
  assign y21204 = n43694 ;
  assign y21205 = n43696 ;
  assign y21206 = ~n43698 ;
  assign y21207 = ~n43701 ;
  assign y21208 = ~n43702 ;
  assign y21209 = ~1'b0 ;
  assign y21210 = ~1'b0 ;
  assign y21211 = n43703 ;
  assign y21212 = n43704 ;
  assign y21213 = n43708 ;
  assign y21214 = ~1'b0 ;
  assign y21215 = ~1'b0 ;
  assign y21216 = ~1'b0 ;
  assign y21217 = n43710 ;
  assign y21218 = ~n28088 ;
  assign y21219 = n43712 ;
  assign y21220 = ~n43713 ;
  assign y21221 = ~n43715 ;
  assign y21222 = n43717 ;
  assign y21223 = ~n43719 ;
  assign y21224 = ~1'b0 ;
  assign y21225 = n43721 ;
  assign y21226 = n43724 ;
  assign y21227 = ~n17094 ;
  assign y21228 = ~n43725 ;
  assign y21229 = n43727 ;
  assign y21230 = ~1'b0 ;
  assign y21231 = ~1'b0 ;
  assign y21232 = ~n43730 ;
  assign y21233 = n43735 ;
  assign y21234 = ~1'b0 ;
  assign y21235 = n43738 ;
  assign y21236 = ~1'b0 ;
  assign y21237 = n43739 ;
  assign y21238 = ~n43740 ;
  assign y21239 = ~n43741 ;
  assign y21240 = ~1'b0 ;
  assign y21241 = ~n43744 ;
  assign y21242 = 1'b0 ;
  assign y21243 = ~1'b0 ;
  assign y21244 = ~1'b0 ;
  assign y21245 = ~n43745 ;
  assign y21246 = ~1'b0 ;
  assign y21247 = ~1'b0 ;
  assign y21248 = ~n43747 ;
  assign y21249 = ~n43748 ;
  assign y21250 = ~n43749 ;
  assign y21251 = ~n1409 ;
  assign y21252 = ~1'b0 ;
  assign y21253 = ~n43751 ;
  assign y21254 = ~1'b0 ;
  assign y21255 = ~1'b0 ;
  assign y21256 = ~n9327 ;
  assign y21257 = ~n43755 ;
  assign y21258 = ~n43757 ;
  assign y21259 = n43762 ;
  assign y21260 = n43763 ;
  assign y21261 = ~1'b0 ;
  assign y21262 = ~n43768 ;
  assign y21263 = ~n43771 ;
  assign y21264 = ~n43772 ;
  assign y21265 = n43773 ;
  assign y21266 = ~1'b0 ;
  assign y21267 = n43778 ;
  assign y21268 = n43779 ;
  assign y21269 = n43781 ;
  assign y21270 = ~n43787 ;
  assign y21271 = ~n43788 ;
  assign y21272 = n43791 ;
  assign y21273 = n21176 ;
  assign y21274 = ~1'b0 ;
  assign y21275 = ~1'b0 ;
  assign y21276 = ~1'b0 ;
  assign y21277 = ~1'b0 ;
  assign y21278 = n43795 ;
  assign y21279 = ~n43798 ;
  assign y21280 = ~n12227 ;
  assign y21281 = n43801 ;
  assign y21282 = ~n43805 ;
  assign y21283 = ~n43806 ;
  assign y21284 = ~1'b0 ;
  assign y21285 = n43807 ;
  assign y21286 = 1'b0 ;
  assign y21287 = ~1'b0 ;
  assign y21288 = n43808 ;
  assign y21289 = n43812 ;
  assign y21290 = ~n26046 ;
  assign y21291 = ~n43818 ;
  assign y21292 = n43819 ;
  assign y21293 = ~1'b0 ;
  assign y21294 = n43821 ;
  assign y21295 = ~n43822 ;
  assign y21296 = n43824 ;
  assign y21297 = n43826 ;
  assign y21298 = ~1'b0 ;
  assign y21299 = ~1'b0 ;
  assign y21300 = ~1'b0 ;
  assign y21301 = ~n43829 ;
  assign y21302 = ~n43833 ;
  assign y21303 = ~n43834 ;
  assign y21304 = n43836 ;
  assign y21305 = ~n43840 ;
  assign y21306 = n43843 ;
  assign y21307 = ~1'b0 ;
  assign y21308 = ~1'b0 ;
  assign y21309 = n43845 ;
  assign y21310 = 1'b0 ;
  assign y21311 = n43846 ;
  assign y21312 = n43847 ;
  assign y21313 = n43849 ;
  assign y21314 = ~n43852 ;
  assign y21315 = ~n43854 ;
  assign y21316 = n43856 ;
  assign y21317 = ~n43857 ;
  assign y21318 = n43860 ;
  assign y21319 = ~n43861 ;
  assign y21320 = n43863 ;
  assign y21321 = ~1'b0 ;
  assign y21322 = ~n34353 ;
  assign y21323 = n43866 ;
  assign y21324 = ~n43869 ;
  assign y21325 = n43873 ;
  assign y21326 = ~n43874 ;
  assign y21327 = ~n43875 ;
  assign y21328 = ~n21851 ;
  assign y21329 = ~1'b0 ;
  assign y21330 = ~1'b0 ;
  assign y21331 = ~n43876 ;
  assign y21332 = ~n43881 ;
  assign y21333 = ~n43882 ;
  assign y21334 = ~n43883 ;
  assign y21335 = n43888 ;
  assign y21336 = n43890 ;
  assign y21337 = ~1'b0 ;
  assign y21338 = ~1'b0 ;
  assign y21339 = ~1'b0 ;
  assign y21340 = n43892 ;
  assign y21341 = ~1'b0 ;
  assign y21342 = n43897 ;
  assign y21343 = n43898 ;
  assign y21344 = ~n43900 ;
  assign y21345 = ~1'b0 ;
  assign y21346 = ~n43902 ;
  assign y21347 = n43903 ;
  assign y21348 = ~n43907 ;
  assign y21349 = ~n43908 ;
  assign y21350 = ~n791 ;
  assign y21351 = n43909 ;
  assign y21352 = n43914 ;
  assign y21353 = n43916 ;
  assign y21354 = n43924 ;
  assign y21355 = ~n43927 ;
  assign y21356 = ~n43930 ;
  assign y21357 = n43932 ;
  assign y21358 = n43934 ;
  assign y21359 = ~1'b0 ;
  assign y21360 = ~1'b0 ;
  assign y21361 = n43935 ;
  assign y21362 = n43938 ;
  assign y21363 = n43942 ;
  assign y21364 = ~n43943 ;
  assign y21365 = ~n43947 ;
  assign y21366 = ~n43955 ;
  assign y21367 = ~n25748 ;
  assign y21368 = ~n22724 ;
  assign y21369 = ~n43957 ;
  assign y21370 = ~n43958 ;
  assign y21371 = n43960 ;
  assign y21372 = ~n43961 ;
  assign y21373 = ~1'b0 ;
  assign y21374 = n43964 ;
  assign y21375 = n43967 ;
  assign y21376 = ~n43969 ;
  assign y21377 = ~n43972 ;
  assign y21378 = ~1'b0 ;
  assign y21379 = ~1'b0 ;
  assign y21380 = n43975 ;
  assign y21381 = ~n43979 ;
  assign y21382 = n43980 ;
  assign y21383 = ~n43981 ;
  assign y21384 = ~n43982 ;
  assign y21385 = ~n43985 ;
  assign y21386 = ~n43986 ;
  assign y21387 = ~n43991 ;
  assign y21388 = ~n43993 ;
  assign y21389 = ~n43994 ;
  assign y21390 = ~1'b0 ;
  assign y21391 = ~n43997 ;
  assign y21392 = ~n44000 ;
  assign y21393 = ~1'b0 ;
  assign y21394 = ~n18387 ;
  assign y21395 = ~n44002 ;
  assign y21396 = n44003 ;
  assign y21397 = n44008 ;
  assign y21398 = ~1'b0 ;
  assign y21399 = n44010 ;
  assign y21400 = ~1'b0 ;
  assign y21401 = ~1'b0 ;
  assign y21402 = ~n44011 ;
  assign y21403 = ~n44012 ;
  assign y21404 = ~n44014 ;
  assign y21405 = n44019 ;
  assign y21406 = ~n44020 ;
  assign y21407 = ~n44023 ;
  assign y21408 = n44025 ;
  assign y21409 = ~n44026 ;
  assign y21410 = 1'b0 ;
  assign y21411 = ~n44028 ;
  assign y21412 = n44031 ;
  assign y21413 = ~1'b0 ;
  assign y21414 = ~1'b0 ;
  assign y21415 = ~n44032 ;
  assign y21416 = 1'b0 ;
  assign y21417 = n44035 ;
  assign y21418 = ~n44040 ;
  assign y21419 = ~n44042 ;
  assign y21420 = 1'b0 ;
  assign y21421 = n44046 ;
  assign y21422 = ~n44047 ;
  assign y21423 = ~1'b0 ;
  assign y21424 = ~1'b0 ;
  assign y21425 = n44048 ;
  assign y21426 = ~n44051 ;
  assign y21427 = 1'b0 ;
  assign y21428 = ~1'b0 ;
  assign y21429 = n44052 ;
  assign y21430 = ~1'b0 ;
  assign y21431 = 1'b0 ;
  assign y21432 = ~1'b0 ;
  assign y21433 = ~n44054 ;
  assign y21434 = ~n44058 ;
  assign y21435 = ~n44060 ;
  assign y21436 = ~n44062 ;
  assign y21437 = ~n44067 ;
  assign y21438 = ~n44070 ;
  assign y21439 = ~n44073 ;
  assign y21440 = ~n44075 ;
  assign y21441 = ~1'b0 ;
  assign y21442 = 1'b0 ;
  assign y21443 = n44076 ;
  assign y21444 = ~n44082 ;
  assign y21445 = ~n44085 ;
  assign y21446 = ~n33339 ;
  assign y21447 = n29415 ;
  assign y21448 = ~n44089 ;
  assign y21449 = ~n44092 ;
  assign y21450 = n44094 ;
  assign y21451 = ~n44101 ;
  assign y21452 = ~1'b0 ;
  assign y21453 = ~n44103 ;
  assign y21454 = n44105 ;
  assign y21455 = n44110 ;
  assign y21456 = n44117 ;
  assign y21457 = ~n44118 ;
  assign y21458 = n44119 ;
  assign y21459 = n44120 ;
  assign y21460 = ~n44121 ;
  assign y21461 = ~1'b0 ;
  assign y21462 = ~1'b0 ;
  assign y21463 = n44125 ;
  assign y21464 = ~n44126 ;
  assign y21465 = ~n44130 ;
  assign y21466 = ~1'b0 ;
  assign y21467 = n32545 ;
  assign y21468 = n44131 ;
  assign y21469 = n44132 ;
  assign y21470 = ~n44134 ;
  assign y21471 = ~n44135 ;
  assign y21472 = n44140 ;
  assign y21473 = ~n44142 ;
  assign y21474 = ~n44143 ;
  assign y21475 = ~n24594 ;
  assign y21476 = ~1'b0 ;
  assign y21477 = n44145 ;
  assign y21478 = ~n44146 ;
  assign y21479 = ~n44147 ;
  assign y21480 = ~n44150 ;
  assign y21481 = ~1'b0 ;
  assign y21482 = n44151 ;
  assign y21483 = n44154 ;
  assign y21484 = ~n4175 ;
  assign y21485 = ~1'b0 ;
  assign y21486 = n44157 ;
  assign y21487 = n44158 ;
  assign y21488 = ~1'b0 ;
  assign y21489 = ~n44162 ;
  assign y21490 = ~n44163 ;
  assign y21491 = ~n44164 ;
  assign y21492 = ~1'b0 ;
  assign y21493 = ~1'b0 ;
  assign y21494 = ~1'b0 ;
  assign y21495 = ~n44165 ;
  assign y21496 = n44168 ;
  assign y21497 = ~n44171 ;
  assign y21498 = n44173 ;
  assign y21499 = n44176 ;
  assign y21500 = ~n44179 ;
  assign y21501 = ~n44183 ;
  assign y21502 = ~n44190 ;
  assign y21503 = n44192 ;
  assign y21504 = ~1'b0 ;
  assign y21505 = ~1'b0 ;
  assign y21506 = ~1'b0 ;
  assign y21507 = n44193 ;
  assign y21508 = n44198 ;
  assign y21509 = ~1'b0 ;
  assign y21510 = ~1'b0 ;
  assign y21511 = ~1'b0 ;
  assign y21512 = n44199 ;
  assign y21513 = ~n44200 ;
  assign y21514 = ~1'b0 ;
  assign y21515 = n44201 ;
  assign y21516 = n44203 ;
  assign y21517 = n44204 ;
  assign y21518 = ~n44205 ;
  assign y21519 = ~1'b0 ;
  assign y21520 = ~1'b0 ;
  assign y21521 = n44207 ;
  assign y21522 = n44208 ;
  assign y21523 = n15922 ;
  assign y21524 = ~1'b0 ;
  assign y21525 = ~1'b0 ;
  assign y21526 = n44211 ;
  assign y21527 = ~n44213 ;
  assign y21528 = ~n44214 ;
  assign y21529 = ~1'b0 ;
  assign y21530 = n44216 ;
  assign y21531 = n44218 ;
  assign y21532 = ~n44219 ;
  assign y21533 = n44220 ;
  assign y21534 = ~1'b0 ;
  assign y21535 = n44221 ;
  assign y21536 = ~1'b0 ;
  assign y21537 = ~n44222 ;
  assign y21538 = ~n44224 ;
  assign y21539 = n44225 ;
  assign y21540 = ~1'b0 ;
  assign y21541 = n44229 ;
  assign y21542 = ~n44230 ;
  assign y21543 = ~n44231 ;
  assign y21544 = n44232 ;
  assign y21545 = ~1'b0 ;
  assign y21546 = n44233 ;
  assign y21547 = n44234 ;
  assign y21548 = ~1'b0 ;
  assign y21549 = ~n44239 ;
  assign y21550 = ~1'b0 ;
  assign y21551 = ~n44241 ;
  assign y21552 = ~n44243 ;
  assign y21553 = n44244 ;
  assign y21554 = n44248 ;
  assign y21555 = n44252 ;
  assign y21556 = ~1'b0 ;
  assign y21557 = n44253 ;
  assign y21558 = ~n44255 ;
  assign y21559 = ~1'b0 ;
  assign y21560 = n44257 ;
  assign y21561 = ~n44259 ;
  assign y21562 = ~1'b0 ;
  assign y21563 = n44260 ;
  assign y21564 = n44263 ;
  assign y21565 = n44264 ;
  assign y21566 = ~n44266 ;
  assign y21567 = ~1'b0 ;
  assign y21568 = ~1'b0 ;
  assign y21569 = ~n44268 ;
  assign y21570 = ~1'b0 ;
  assign y21571 = ~n44272 ;
  assign y21572 = ~1'b0 ;
  assign y21573 = ~1'b0 ;
  assign y21574 = ~1'b0 ;
  assign y21575 = ~n44273 ;
  assign y21576 = ~n44274 ;
  assign y21577 = ~n465 ;
  assign y21578 = ~n44276 ;
  assign y21579 = ~1'b0 ;
  assign y21580 = ~n44278 ;
  assign y21581 = ~1'b0 ;
  assign y21582 = ~1'b0 ;
  assign y21583 = ~n44281 ;
  assign y21584 = ~n44283 ;
  assign y21585 = ~n44285 ;
  assign y21586 = n44286 ;
  assign y21587 = n44290 ;
  assign y21588 = ~n44292 ;
  assign y21589 = ~n44295 ;
  assign y21590 = ~n44296 ;
  assign y21591 = ~1'b0 ;
  assign y21592 = ~1'b0 ;
  assign y21593 = ~1'b0 ;
  assign y21594 = n44301 ;
  assign y21595 = n44304 ;
  assign y21596 = ~1'b0 ;
  assign y21597 = ~n44306 ;
  assign y21598 = n44309 ;
  assign y21599 = ~n19305 ;
  assign y21600 = n44311 ;
  assign y21601 = ~1'b0 ;
  assign y21602 = ~n44313 ;
  assign y21603 = ~n44314 ;
  assign y21604 = ~n44315 ;
  assign y21605 = ~n44321 ;
  assign y21606 = ~1'b0 ;
  assign y21607 = ~1'b0 ;
  assign y21608 = ~n24342 ;
  assign y21609 = n44323 ;
  assign y21610 = ~n44325 ;
  assign y21611 = n44327 ;
  assign y21612 = ~1'b0 ;
  assign y21613 = ~n44332 ;
  assign y21614 = n44333 ;
  assign y21615 = n44334 ;
  assign y21616 = ~n44335 ;
  assign y21617 = n44336 ;
  assign y21618 = n44340 ;
  assign y21619 = ~n44344 ;
  assign y21620 = ~1'b0 ;
  assign y21621 = ~1'b0 ;
  assign y21622 = ~1'b0 ;
  assign y21623 = n44348 ;
  assign y21624 = ~1'b0 ;
  assign y21625 = ~n44351 ;
  assign y21626 = n44355 ;
  assign y21627 = n44359 ;
  assign y21628 = ~1'b0 ;
  assign y21629 = n44361 ;
  assign y21630 = 1'b0 ;
  assign y21631 = 1'b0 ;
  assign y21632 = ~1'b0 ;
  assign y21633 = n44363 ;
  assign y21634 = ~n44364 ;
  assign y21635 = ~n44369 ;
  assign y21636 = n44370 ;
  assign y21637 = ~n44371 ;
  assign y21638 = n44372 ;
  assign y21639 = n44375 ;
  assign y21640 = ~1'b0 ;
  assign y21641 = n44377 ;
  assign y21642 = n44378 ;
  assign y21643 = n44379 ;
  assign y21644 = ~1'b0 ;
  assign y21645 = n44381 ;
  assign y21646 = n23653 ;
  assign y21647 = n44382 ;
  assign y21648 = n44383 ;
  assign y21649 = ~1'b0 ;
  assign y21650 = n44386 ;
  assign y21651 = n44388 ;
  assign y21652 = ~1'b0 ;
  assign y21653 = n44389 ;
  assign y21654 = n44391 ;
  assign y21655 = ~n44392 ;
  assign y21656 = ~n44395 ;
  assign y21657 = ~n44397 ;
  assign y21658 = ~n44398 ;
  assign y21659 = n44399 ;
  assign y21660 = ~n30683 ;
  assign y21661 = ~1'b0 ;
  assign y21662 = n44405 ;
  assign y21663 = ~1'b0 ;
  assign y21664 = ~n44407 ;
  assign y21665 = ~n44409 ;
  assign y21666 = ~n44412 ;
  assign y21667 = ~n44413 ;
  assign y21668 = n44417 ;
  assign y21669 = n44418 ;
  assign y21670 = ~1'b0 ;
  assign y21671 = n44420 ;
  assign y21672 = ~1'b0 ;
  assign y21673 = ~n44422 ;
  assign y21674 = ~1'b0 ;
  assign y21675 = n44425 ;
  assign y21676 = n44426 ;
  assign y21677 = ~n44429 ;
  assign y21678 = n44430 ;
  assign y21679 = n44433 ;
  assign y21680 = ~1'b0 ;
  assign y21681 = ~n44434 ;
  assign y21682 = ~n44435 ;
  assign y21683 = ~1'b0 ;
  assign y21684 = ~1'b0 ;
  assign y21685 = n44436 ;
  assign y21686 = ~1'b0 ;
  assign y21687 = n44439 ;
  assign y21688 = ~n44441 ;
  assign y21689 = ~n44444 ;
  assign y21690 = n44447 ;
  assign y21691 = n44453 ;
  assign y21692 = ~n44454 ;
  assign y21693 = ~1'b0 ;
  assign y21694 = n44455 ;
  assign y21695 = ~1'b0 ;
  assign y21696 = n44458 ;
  assign y21697 = ~n44459 ;
  assign y21698 = n44462 ;
  assign y21699 = n44465 ;
  assign y21700 = n44467 ;
  assign y21701 = ~n44468 ;
  assign y21702 = ~1'b0 ;
  assign y21703 = ~n44469 ;
  assign y21704 = n44470 ;
  assign y21705 = ~1'b0 ;
  assign y21706 = n44472 ;
  assign y21707 = ~n13156 ;
  assign y21708 = n44475 ;
  assign y21709 = n44477 ;
  assign y21710 = n44478 ;
  assign y21711 = ~1'b0 ;
  assign y21712 = n44480 ;
  assign y21713 = ~1'b0 ;
  assign y21714 = ~1'b0 ;
  assign y21715 = n44488 ;
  assign y21716 = n26251 ;
  assign y21717 = n44490 ;
  assign y21718 = n44491 ;
  assign y21719 = n44495 ;
  assign y21720 = ~n44498 ;
  assign y21721 = ~n44504 ;
  assign y21722 = n44508 ;
  assign y21723 = n44514 ;
  assign y21724 = ~1'b0 ;
  assign y21725 = ~1'b0 ;
  assign y21726 = n44515 ;
  assign y21727 = ~1'b0 ;
  assign y21728 = n44516 ;
  assign y21729 = n44517 ;
  assign y21730 = n44518 ;
  assign y21731 = ~n44521 ;
  assign y21732 = ~n44522 ;
  assign y21733 = ~n44524 ;
  assign y21734 = ~1'b0 ;
  assign y21735 = ~1'b0 ;
  assign y21736 = n44527 ;
  assign y21737 = ~n44531 ;
  assign y21738 = ~n44536 ;
  assign y21739 = n44538 ;
  assign y21740 = ~n44539 ;
  assign y21741 = ~n44543 ;
  assign y21742 = n44544 ;
  assign y21743 = ~n44545 ;
  assign y21744 = ~1'b0 ;
  assign y21745 = n44546 ;
  assign y21746 = ~n44550 ;
  assign y21747 = n44553 ;
  assign y21748 = ~1'b0 ;
  assign y21749 = ~n44554 ;
  assign y21750 = ~n8354 ;
  assign y21751 = ~n44556 ;
  assign y21752 = ~n44557 ;
  assign y21753 = n44558 ;
  assign y21754 = ~n44559 ;
  assign y21755 = n44561 ;
  assign y21756 = ~n40826 ;
  assign y21757 = ~1'b0 ;
  assign y21758 = ~1'b0 ;
  assign y21759 = n44562 ;
  assign y21760 = n44564 ;
  assign y21761 = n44568 ;
  assign y21762 = n44569 ;
  assign y21763 = ~n44571 ;
  assign y21764 = ~1'b0 ;
  assign y21765 = ~n44573 ;
  assign y21766 = ~n44576 ;
  assign y21767 = ~1'b0 ;
  assign y21768 = ~n44579 ;
  assign y21769 = ~n44581 ;
  assign y21770 = ~n44585 ;
  assign y21771 = ~1'b0 ;
  assign y21772 = ~n44586 ;
  assign y21773 = ~n44587 ;
  assign y21774 = n26398 ;
  assign y21775 = ~1'b0 ;
  assign y21776 = n44588 ;
  assign y21777 = ~n38624 ;
  assign y21778 = ~n44590 ;
  assign y21779 = ~1'b0 ;
  assign y21780 = ~1'b0 ;
  assign y21781 = ~n44592 ;
  assign y21782 = n44593 ;
  assign y21783 = ~n44595 ;
  assign y21784 = ~n44598 ;
  assign y21785 = n9644 ;
  assign y21786 = ~n44600 ;
  assign y21787 = ~1'b0 ;
  assign y21788 = ~n44605 ;
  assign y21789 = n44606 ;
  assign y21790 = ~1'b0 ;
  assign y21791 = n44607 ;
  assign y21792 = ~n22438 ;
  assign y21793 = n44609 ;
  assign y21794 = n44612 ;
  assign y21795 = n44614 ;
  assign y21796 = n44620 ;
  assign y21797 = n44623 ;
  assign y21798 = ~1'b0 ;
  assign y21799 = n8377 ;
  assign y21800 = ~1'b0 ;
  assign y21801 = ~n44624 ;
  assign y21802 = n44626 ;
  assign y21803 = ~1'b0 ;
  assign y21804 = n44627 ;
  assign y21805 = ~1'b0 ;
  assign y21806 = n44630 ;
  assign y21807 = ~1'b0 ;
  assign y21808 = n44631 ;
  assign y21809 = ~n44633 ;
  assign y21810 = ~1'b0 ;
  assign y21811 = ~n44635 ;
  assign y21812 = n44636 ;
  assign y21813 = ~n44637 ;
  assign y21814 = ~n44640 ;
  assign y21815 = ~n44642 ;
  assign y21816 = ~1'b0 ;
  assign y21817 = ~n44644 ;
  assign y21818 = ~n44645 ;
  assign y21819 = ~n2286 ;
  assign y21820 = n44649 ;
  assign y21821 = ~1'b0 ;
  assign y21822 = 1'b0 ;
  assign y21823 = ~n44651 ;
  assign y21824 = ~n44657 ;
  assign y21825 = ~n44660 ;
  assign y21826 = ~n44664 ;
  assign y21827 = ~1'b0 ;
  assign y21828 = ~n44665 ;
  assign y21829 = n44667 ;
  assign y21830 = ~n44669 ;
  assign y21831 = n44672 ;
  assign y21832 = ~n26102 ;
  assign y21833 = n44674 ;
  assign y21834 = n44676 ;
  assign y21835 = n44679 ;
  assign y21836 = n44683 ;
  assign y21837 = ~1'b0 ;
  assign y21838 = ~1'b0 ;
  assign y21839 = ~1'b0 ;
  assign y21840 = n44686 ;
  assign y21841 = n44687 ;
  assign y21842 = ~1'b0 ;
  assign y21843 = n20544 ;
  assign y21844 = ~n44690 ;
  assign y21845 = ~n44691 ;
  assign y21846 = ~n44692 ;
  assign y21847 = ~1'b0 ;
  assign y21848 = n44693 ;
  assign y21849 = ~1'b0 ;
  assign y21850 = n44696 ;
  assign y21851 = ~n44700 ;
  assign y21852 = n44702 ;
  assign y21853 = n44703 ;
  assign y21854 = n44706 ;
  assign y21855 = ~n44708 ;
  assign y21856 = ~n44709 ;
  assign y21857 = n44711 ;
  assign y21858 = ~1'b0 ;
  assign y21859 = ~n44714 ;
  assign y21860 = n44717 ;
  assign y21861 = ~1'b0 ;
  assign y21862 = n44719 ;
  assign y21863 = ~n44721 ;
  assign y21864 = n44722 ;
  assign y21865 = ~n25818 ;
  assign y21866 = ~n23240 ;
  assign y21867 = n44723 ;
  assign y21868 = ~n44725 ;
  assign y21869 = ~1'b0 ;
  assign y21870 = ~n44727 ;
  assign y21871 = ~n44728 ;
  assign y21872 = ~n44729 ;
  assign y21873 = n44735 ;
  assign y21874 = n44737 ;
  assign y21875 = n44741 ;
  assign y21876 = ~n44742 ;
  assign y21877 = ~n44743 ;
  assign y21878 = ~n44751 ;
  assign y21879 = ~n44754 ;
  assign y21880 = n44755 ;
  assign y21881 = ~1'b0 ;
  assign y21882 = n44757 ;
  assign y21883 = ~n44759 ;
  assign y21884 = ~n44766 ;
  assign y21885 = ~n44767 ;
  assign y21886 = ~1'b0 ;
  assign y21887 = ~n44770 ;
  assign y21888 = ~n44771 ;
  assign y21889 = n44772 ;
  assign y21890 = ~n44774 ;
  assign y21891 = ~n44775 ;
  assign y21892 = ~1'b0 ;
  assign y21893 = n44779 ;
  assign y21894 = ~1'b0 ;
  assign y21895 = n44782 ;
  assign y21896 = n44783 ;
  assign y21897 = ~n6262 ;
  assign y21898 = n44787 ;
  assign y21899 = n44791 ;
  assign y21900 = ~1'b0 ;
  assign y21901 = ~1'b0 ;
  assign y21902 = ~1'b0 ;
  assign y21903 = ~1'b0 ;
  assign y21904 = n44792 ;
  assign y21905 = n44798 ;
  assign y21906 = ~1'b0 ;
  assign y21907 = ~n33594 ;
  assign y21908 = ~n44800 ;
  assign y21909 = ~n44803 ;
  assign y21910 = n44807 ;
  assign y21911 = ~n44810 ;
  assign y21912 = n44812 ;
  assign y21913 = ~n44818 ;
  assign y21914 = ~1'b0 ;
  assign y21915 = n44820 ;
  assign y21916 = ~n44823 ;
  assign y21917 = 1'b0 ;
  assign y21918 = ~n44824 ;
  assign y21919 = n44825 ;
  assign y21920 = n44827 ;
  assign y21921 = n44828 ;
  assign y21922 = n44830 ;
  assign y21923 = ~n44832 ;
  assign y21924 = ~n44834 ;
  assign y21925 = n44836 ;
  assign y21926 = ~1'b0 ;
  assign y21927 = ~1'b0 ;
  assign y21928 = n44838 ;
  assign y21929 = ~n44840 ;
  assign y21930 = ~n44841 ;
  assign y21931 = ~n44844 ;
  assign y21932 = n44846 ;
  assign y21933 = ~1'b0 ;
  assign y21934 = ~n44849 ;
  assign y21935 = ~n44852 ;
  assign y21936 = ~n44855 ;
  assign y21937 = ~1'b0 ;
  assign y21938 = n44861 ;
  assign y21939 = ~n44862 ;
  assign y21940 = ~n44863 ;
  assign y21941 = 1'b0 ;
  assign y21942 = ~n44865 ;
  assign y21943 = ~n44866 ;
  assign y21944 = n44867 ;
  assign y21945 = ~n44877 ;
  assign y21946 = n44881 ;
  assign y21947 = n44883 ;
  assign y21948 = ~n44889 ;
  assign y21949 = n44891 ;
  assign y21950 = ~1'b0 ;
  assign y21951 = ~n44893 ;
  assign y21952 = ~n44896 ;
  assign y21953 = ~n44897 ;
  assign y21954 = ~1'b0 ;
  assign y21955 = ~1'b0 ;
  assign y21956 = n22969 ;
  assign y21957 = n44899 ;
  assign y21958 = ~n44902 ;
  assign y21959 = ~n44904 ;
  assign y21960 = n44906 ;
  assign y21961 = n44907 ;
  assign y21962 = ~n44908 ;
  assign y21963 = ~n44909 ;
  assign y21964 = n44911 ;
  assign y21965 = ~n44912 ;
  assign y21966 = ~n44913 ;
  assign y21967 = ~1'b0 ;
  assign y21968 = n44914 ;
  assign y21969 = 1'b0 ;
  assign y21970 = ~1'b0 ;
  assign y21971 = n44918 ;
  assign y21972 = ~n44919 ;
  assign y21973 = n44921 ;
  assign y21974 = ~1'b0 ;
  assign y21975 = ~1'b0 ;
  assign y21976 = n44923 ;
  assign y21977 = n44927 ;
  assign y21978 = ~n44929 ;
  assign y21979 = n44932 ;
  assign y21980 = ~1'b0 ;
  assign y21981 = n44933 ;
  assign y21982 = ~n44943 ;
  assign y21983 = ~n44946 ;
  assign y21984 = n44949 ;
  assign y21985 = ~n44954 ;
  assign y21986 = ~n44955 ;
  assign y21987 = ~n44959 ;
  assign y21988 = n44962 ;
  assign y21989 = ~1'b0 ;
  assign y21990 = ~1'b0 ;
  assign y21991 = ~n44971 ;
  assign y21992 = ~n44972 ;
  assign y21993 = ~n44973 ;
  assign y21994 = n44974 ;
  assign y21995 = n44975 ;
  assign y21996 = ~n44978 ;
  assign y21997 = ~n44982 ;
  assign y21998 = ~1'b0 ;
  assign y21999 = ~1'b0 ;
  assign y22000 = n44985 ;
  assign y22001 = n44986 ;
  assign y22002 = ~n44987 ;
  assign y22003 = n44990 ;
  assign y22004 = ~1'b0 ;
  assign y22005 = n17146 ;
  assign y22006 = ~n44991 ;
  assign y22007 = n44402 ;
  assign y22008 = ~n44996 ;
  assign y22009 = ~n44997 ;
  assign y22010 = ~1'b0 ;
  assign y22011 = n45002 ;
  assign y22012 = n45004 ;
  assign y22013 = ~n45006 ;
  assign y22014 = ~1'b0 ;
  assign y22015 = ~1'b0 ;
  assign y22016 = n45007 ;
  assign y22017 = ~n4380 ;
  assign y22018 = n45014 ;
  assign y22019 = n45018 ;
  assign y22020 = ~n45019 ;
  assign y22021 = ~1'b0 ;
  assign y22022 = ~1'b0 ;
  assign y22023 = n45020 ;
  assign y22024 = ~n45022 ;
  assign y22025 = ~1'b0 ;
  assign y22026 = ~x182 ;
  assign y22027 = ~1'b0 ;
  assign y22028 = ~n45025 ;
  assign y22029 = ~n45026 ;
  assign y22030 = ~1'b0 ;
  assign y22031 = ~1'b0 ;
  assign y22032 = ~n45029 ;
  assign y22033 = ~n45030 ;
  assign y22034 = n45033 ;
  assign y22035 = n45035 ;
  assign y22036 = n45038 ;
  assign y22037 = n45044 ;
  assign y22038 = ~n45050 ;
  assign y22039 = n45053 ;
  assign y22040 = n852 ;
  assign y22041 = n45055 ;
  assign y22042 = ~1'b0 ;
  assign y22043 = n45057 ;
  assign y22044 = ~n45058 ;
  assign y22045 = ~n45061 ;
  assign y22046 = ~n45063 ;
  assign y22047 = ~n45064 ;
  assign y22048 = n45065 ;
  assign y22049 = ~n14422 ;
  assign y22050 = ~n45067 ;
  assign y22051 = ~n45071 ;
  assign y22052 = 1'b0 ;
  assign y22053 = n45072 ;
  assign y22054 = ~1'b0 ;
  assign y22055 = ~1'b0 ;
  assign y22056 = ~n45077 ;
  assign y22057 = ~n45081 ;
  assign y22058 = ~n45082 ;
  assign y22059 = ~1'b0 ;
  assign y22060 = n45083 ;
  assign y22061 = ~n45086 ;
  assign y22062 = n45087 ;
  assign y22063 = ~n45092 ;
  assign y22064 = ~1'b0 ;
  assign y22065 = ~n45093 ;
  assign y22066 = ~n45095 ;
  assign y22067 = ~n45098 ;
  assign y22068 = ~n45101 ;
  assign y22069 = ~n45102 ;
  assign y22070 = ~1'b0 ;
  assign y22071 = ~n36837 ;
  assign y22072 = n26438 ;
  assign y22073 = ~n45104 ;
  assign y22074 = ~n45106 ;
  assign y22075 = ~n45108 ;
  assign y22076 = 1'b0 ;
  assign y22077 = n45111 ;
  assign y22078 = ~n45116 ;
  assign y22079 = ~1'b0 ;
  assign y22080 = n45119 ;
  assign y22081 = ~n45121 ;
  assign y22082 = ~1'b0 ;
  assign y22083 = ~n45125 ;
  assign y22084 = ~n45127 ;
  assign y22085 = ~n45129 ;
  assign y22086 = ~1'b0 ;
  assign y22087 = n45130 ;
  assign y22088 = 1'b0 ;
  assign y22089 = ~n45133 ;
  assign y22090 = ~n45134 ;
  assign y22091 = n45135 ;
  assign y22092 = ~n45137 ;
  assign y22093 = ~1'b0 ;
  assign y22094 = n45139 ;
  assign y22095 = ~1'b0 ;
  assign y22096 = ~n45144 ;
  assign y22097 = ~n45148 ;
  assign y22098 = n45152 ;
  assign y22099 = ~n45154 ;
  assign y22100 = n45155 ;
  assign y22101 = ~n45156 ;
  assign y22102 = ~1'b0 ;
  assign y22103 = ~1'b0 ;
  assign y22104 = ~n45159 ;
  assign y22105 = ~n23232 ;
  assign y22106 = ~n45161 ;
  assign y22107 = ~1'b0 ;
  assign y22108 = ~1'b0 ;
  assign y22109 = n45162 ;
  assign y22110 = n45163 ;
  assign y22111 = ~n45168 ;
  assign y22112 = ~n45176 ;
  assign y22113 = 1'b0 ;
  assign y22114 = ~1'b0 ;
  assign y22115 = ~1'b0 ;
  assign y22116 = ~1'b0 ;
  assign y22117 = ~1'b0 ;
  assign y22118 = ~1'b0 ;
  assign y22119 = ~1'b0 ;
  assign y22120 = 1'b0 ;
  assign y22121 = n45180 ;
  assign y22122 = ~n45185 ;
  assign y22123 = n45195 ;
  assign y22124 = n45199 ;
  assign y22125 = ~1'b0 ;
  assign y22126 = ~1'b0 ;
  assign y22127 = n45200 ;
  assign y22128 = ~n42906 ;
  assign y22129 = ~n45201 ;
  assign y22130 = n45202 ;
  assign y22131 = ~n45203 ;
  assign y22132 = n45206 ;
  assign y22133 = ~n10717 ;
  assign y22134 = ~1'b0 ;
  assign y22135 = ~1'b0 ;
  assign y22136 = ~1'b0 ;
  assign y22137 = n45208 ;
  assign y22138 = ~1'b0 ;
  assign y22139 = ~n45209 ;
  assign y22140 = ~n45215 ;
  assign y22141 = n45217 ;
  assign y22142 = n45226 ;
  assign y22143 = n45229 ;
  assign y22144 = ~n45230 ;
  assign y22145 = ~n45231 ;
  assign y22146 = n45234 ;
  assign y22147 = ~1'b0 ;
  assign y22148 = ~n45237 ;
  assign y22149 = n45239 ;
  assign y22150 = ~1'b0 ;
  assign y22151 = ~n45240 ;
  assign y22152 = ~n45241 ;
  assign y22153 = n45242 ;
  assign y22154 = n45243 ;
  assign y22155 = ~n45245 ;
  assign y22156 = ~1'b0 ;
  assign y22157 = n45249 ;
  assign y22158 = ~1'b0 ;
  assign y22159 = ~1'b0 ;
  assign y22160 = ~n45252 ;
  assign y22161 = ~1'b0 ;
  assign y22162 = ~n45254 ;
  assign y22163 = ~n45255 ;
  assign y22164 = ~n45258 ;
  assign y22165 = n45260 ;
  assign y22166 = n45261 ;
  assign y22167 = n45264 ;
  assign y22168 = ~1'b0 ;
  assign y22169 = ~1'b0 ;
  assign y22170 = ~1'b0 ;
  assign y22171 = ~n35000 ;
  assign y22172 = n45266 ;
  assign y22173 = n45267 ;
  assign y22174 = n45272 ;
  assign y22175 = ~n45273 ;
  assign y22176 = ~n45274 ;
  assign y22177 = 1'b0 ;
  assign y22178 = ~1'b0 ;
  assign y22179 = n45276 ;
  assign y22180 = ~1'b0 ;
  assign y22181 = ~1'b0 ;
  assign y22182 = n45277 ;
  assign y22183 = ~1'b0 ;
  assign y22184 = n45280 ;
  assign y22185 = ~n45281 ;
  assign y22186 = ~n45282 ;
  assign y22187 = ~1'b0 ;
  assign y22188 = ~1'b0 ;
  assign y22189 = ~1'b0 ;
  assign y22190 = ~n45284 ;
  assign y22191 = ~n45288 ;
  assign y22192 = ~n45290 ;
  assign y22193 = n45292 ;
  assign y22194 = ~1'b0 ;
  assign y22195 = ~n45294 ;
  assign y22196 = ~n45297 ;
  assign y22197 = ~n45298 ;
  assign y22198 = ~1'b0 ;
  assign y22199 = n45299 ;
  assign y22200 = ~1'b0 ;
  assign y22201 = ~n45303 ;
  assign y22202 = n45306 ;
  assign y22203 = ~1'b0 ;
  assign y22204 = ~n45310 ;
  assign y22205 = n45312 ;
  assign y22206 = ~n45318 ;
  assign y22207 = ~n45323 ;
  assign y22208 = ~n1987 ;
  assign y22209 = ~1'b0 ;
  assign y22210 = ~1'b0 ;
  assign y22211 = ~n45329 ;
  assign y22212 = ~n45330 ;
  assign y22213 = ~n45332 ;
  assign y22214 = ~n45333 ;
  assign y22215 = n45335 ;
  assign y22216 = ~1'b0 ;
  assign y22217 = ~n9032 ;
  assign y22218 = ~n45336 ;
  assign y22219 = ~n45339 ;
  assign y22220 = n45340 ;
  assign y22221 = n45342 ;
  assign y22222 = n45345 ;
  assign y22223 = n45346 ;
  assign y22224 = ~n28166 ;
  assign y22225 = ~1'b0 ;
  assign y22226 = n45349 ;
  assign y22227 = 1'b0 ;
  assign y22228 = n45352 ;
  assign y22229 = n45354 ;
  assign y22230 = ~n45356 ;
  assign y22231 = ~1'b0 ;
  assign y22232 = ~1'b0 ;
  assign y22233 = ~1'b0 ;
  assign y22234 = n45362 ;
  assign y22235 = n45364 ;
  assign y22236 = n29216 ;
  assign y22237 = ~n45365 ;
  assign y22238 = n45367 ;
  assign y22239 = n45369 ;
  assign y22240 = ~n45370 ;
  assign y22241 = ~n45371 ;
  assign y22242 = ~n45372 ;
  assign y22243 = ~n45374 ;
  assign y22244 = n45379 ;
  assign y22245 = ~1'b0 ;
  assign y22246 = n45381 ;
  assign y22247 = n45383 ;
  assign y22248 = n45385 ;
  assign y22249 = ~n45386 ;
  assign y22250 = ~n45387 ;
  assign y22251 = ~n45391 ;
  assign y22252 = n1304 ;
  assign y22253 = n45399 ;
  assign y22254 = n45401 ;
  assign y22255 = n45404 ;
  assign y22256 = ~1'b0 ;
  assign y22257 = ~n45406 ;
  assign y22258 = n17240 ;
  assign y22259 = n45409 ;
  assign y22260 = ~n45410 ;
  assign y22261 = n45411 ;
  assign y22262 = ~1'b0 ;
  assign y22263 = n45414 ;
  assign y22264 = ~n45418 ;
  assign y22265 = ~n45422 ;
  assign y22266 = ~n17045 ;
  assign y22267 = ~n39710 ;
  assign y22268 = ~1'b0 ;
  assign y22269 = n45426 ;
  assign y22270 = n45433 ;
  assign y22271 = n45434 ;
  assign y22272 = ~n45435 ;
  assign y22273 = n45438 ;
  assign y22274 = ~1'b0 ;
  assign y22275 = n45439 ;
  assign y22276 = n45440 ;
  assign y22277 = n45441 ;
  assign y22278 = n45443 ;
  assign y22279 = ~n45446 ;
  assign y22280 = n45450 ;
  assign y22281 = n45451 ;
  assign y22282 = n45452 ;
  assign y22283 = ~1'b0 ;
  assign y22284 = n45453 ;
  assign y22285 = ~n45458 ;
  assign y22286 = n45463 ;
  assign y22287 = n45464 ;
  assign y22288 = ~1'b0 ;
  assign y22289 = ~1'b0 ;
  assign y22290 = ~n45466 ;
  assign y22291 = ~n45468 ;
  assign y22292 = ~1'b0 ;
  assign y22293 = ~n45470 ;
  assign y22294 = ~n45473 ;
  assign y22295 = ~n45476 ;
  assign y22296 = n45478 ;
  assign y22297 = ~1'b0 ;
  assign y22298 = ~1'b0 ;
  assign y22299 = ~n45480 ;
  assign y22300 = ~1'b0 ;
  assign y22301 = ~n45481 ;
  assign y22302 = ~1'b0 ;
  assign y22303 = ~n45483 ;
  assign y22304 = ~n45485 ;
  assign y22305 = n15276 ;
  assign y22306 = n13880 ;
  assign y22307 = 1'b0 ;
  assign y22308 = ~n45489 ;
  assign y22309 = n45493 ;
  assign y22310 = ~1'b0 ;
  assign y22311 = n45499 ;
  assign y22312 = ~n45505 ;
  assign y22313 = n45506 ;
  assign y22314 = n45509 ;
  assign y22315 = n45512 ;
  assign y22316 = n45513 ;
  assign y22317 = ~n45516 ;
  assign y22318 = n45518 ;
  assign y22319 = n45520 ;
  assign y22320 = ~n45522 ;
  assign y22321 = ~n45523 ;
  assign y22322 = ~1'b0 ;
  assign y22323 = n4542 ;
  assign y22324 = n45524 ;
  assign y22325 = n45526 ;
  assign y22326 = n45529 ;
  assign y22327 = n45531 ;
  assign y22328 = ~1'b0 ;
  assign y22329 = ~1'b0 ;
  assign y22330 = ~n45533 ;
  assign y22331 = ~1'b0 ;
  assign y22332 = n45534 ;
  assign y22333 = n45539 ;
  assign y22334 = ~n45545 ;
  assign y22335 = ~n31768 ;
  assign y22336 = n45548 ;
  assign y22337 = n45549 ;
  assign y22338 = ~1'b0 ;
  assign y22339 = n45554 ;
  assign y22340 = n45555 ;
  assign y22341 = ~n45556 ;
  assign y22342 = n45557 ;
  assign y22343 = n45559 ;
  assign y22344 = ~n45560 ;
  assign y22345 = ~n45563 ;
  assign y22346 = n45566 ;
  assign y22347 = ~n45567 ;
  assign y22348 = n45569 ;
  assign y22349 = ~n37413 ;
  assign y22350 = n45570 ;
  assign y22351 = ~1'b0 ;
  assign y22352 = ~n45573 ;
  assign y22353 = ~n45574 ;
  assign y22354 = ~1'b0 ;
  assign y22355 = ~n45576 ;
  assign y22356 = ~n45577 ;
  assign y22357 = ~n45578 ;
  assign y22358 = n3376 ;
  assign y22359 = n45579 ;
  assign y22360 = ~1'b0 ;
  assign y22361 = ~1'b0 ;
  assign y22362 = ~n45586 ;
  assign y22363 = ~n45587 ;
  assign y22364 = n45589 ;
  assign y22365 = ~n23249 ;
  assign y22366 = n45592 ;
  assign y22367 = n45593 ;
  assign y22368 = ~n20756 ;
  assign y22369 = ~n45597 ;
  assign y22370 = ~n45598 ;
  assign y22371 = ~n45599 ;
  assign y22372 = ~1'b0 ;
  assign y22373 = n45603 ;
  assign y22374 = ~1'b0 ;
  assign y22375 = ~n45604 ;
  assign y22376 = ~n45606 ;
  assign y22377 = ~n45608 ;
  assign y22378 = n45611 ;
  assign y22379 = n45612 ;
  assign y22380 = n45613 ;
  assign y22381 = ~n45614 ;
  assign y22382 = ~n45616 ;
  assign y22383 = n813 ;
  assign y22384 = ~n45617 ;
  assign y22385 = ~n45618 ;
  assign y22386 = ~n45619 ;
  assign y22387 = n45620 ;
  assign y22388 = n45622 ;
  assign y22389 = n45625 ;
  assign y22390 = n45628 ;
  assign y22391 = n45630 ;
  assign y22392 = n45632 ;
  assign y22393 = ~n45635 ;
  assign y22394 = n9318 ;
  assign y22395 = ~n45639 ;
  assign y22396 = ~1'b0 ;
  assign y22397 = n45641 ;
  assign y22398 = ~1'b0 ;
  assign y22399 = n13364 ;
  assign y22400 = ~n45643 ;
  assign y22401 = ~n45647 ;
  assign y22402 = n45651 ;
  assign y22403 = n45652 ;
  assign y22404 = ~n27264 ;
  assign y22405 = ~1'b0 ;
  assign y22406 = ~n31336 ;
  assign y22407 = n45655 ;
  assign y22408 = ~1'b0 ;
  assign y22409 = ~n45658 ;
  assign y22410 = n45660 ;
  assign y22411 = ~1'b0 ;
  assign y22412 = ~n45667 ;
  assign y22413 = n45670 ;
  assign y22414 = ~n45672 ;
  assign y22415 = ~1'b0 ;
  assign y22416 = n45673 ;
  assign y22417 = 1'b0 ;
  assign y22418 = ~n45675 ;
  assign y22419 = ~n45677 ;
  assign y22420 = n45679 ;
  assign y22421 = ~1'b0 ;
  assign y22422 = ~1'b0 ;
  assign y22423 = ~n45682 ;
  assign y22424 = ~n45685 ;
  assign y22425 = ~n45686 ;
  assign y22426 = ~n45688 ;
  assign y22427 = n45690 ;
  assign y22428 = ~n45692 ;
  assign y22429 = n45695 ;
  assign y22430 = n45697 ;
  assign y22431 = ~1'b0 ;
  assign y22432 = n45700 ;
  assign y22433 = ~1'b0 ;
  assign y22434 = ~n45701 ;
  assign y22435 = ~n45703 ;
  assign y22436 = ~n45708 ;
  assign y22437 = n45709 ;
  assign y22438 = n4860 ;
  assign y22439 = ~n45710 ;
  assign y22440 = ~1'b0 ;
  assign y22441 = ~n45714 ;
  assign y22442 = ~1'b0 ;
  assign y22443 = ~n45717 ;
  assign y22444 = ~1'b0 ;
  assign y22445 = n45718 ;
  assign y22446 = ~n45719 ;
  assign y22447 = ~n45720 ;
  assign y22448 = ~1'b0 ;
  assign y22449 = ~n45721 ;
  assign y22450 = n45722 ;
  assign y22451 = n45723 ;
  assign y22452 = n45727 ;
  assign y22453 = ~n45732 ;
  assign y22454 = n15410 ;
  assign y22455 = ~n45734 ;
  assign y22456 = ~n45739 ;
  assign y22457 = ~n45740 ;
  assign y22458 = ~1'b0 ;
  assign y22459 = ~1'b0 ;
  assign y22460 = n45743 ;
  assign y22461 = ~1'b0 ;
  assign y22462 = ~1'b0 ;
  assign y22463 = ~n45753 ;
  assign y22464 = ~n45754 ;
  assign y22465 = ~1'b0 ;
  assign y22466 = n45755 ;
  assign y22467 = n45758 ;
  assign y22468 = ~n45759 ;
  assign y22469 = ~1'b0 ;
  assign y22470 = ~n45760 ;
  assign y22471 = ~1'b0 ;
  assign y22472 = ~n45763 ;
  assign y22473 = ~1'b0 ;
  assign y22474 = 1'b0 ;
  assign y22475 = n45765 ;
  assign y22476 = ~n45766 ;
  assign y22477 = n45768 ;
  assign y22478 = ~n45769 ;
  assign y22479 = n45770 ;
  assign y22480 = n26692 ;
  assign y22481 = n45772 ;
  assign y22482 = n45776 ;
  assign y22483 = ~1'b0 ;
  assign y22484 = ~1'b0 ;
  assign y22485 = ~n45777 ;
  assign y22486 = ~n45779 ;
  assign y22487 = ~n45780 ;
  assign y22488 = n45784 ;
  assign y22489 = ~1'b0 ;
  assign y22490 = ~n45785 ;
  assign y22491 = ~n45791 ;
  assign y22492 = n45793 ;
  assign y22493 = ~1'b0 ;
  assign y22494 = ~n45798 ;
  assign y22495 = ~1'b0 ;
  assign y22496 = n45803 ;
  assign y22497 = n45804 ;
  assign y22498 = n45809 ;
  assign y22499 = ~n45812 ;
  assign y22500 = n45813 ;
  assign y22501 = ~1'b0 ;
  assign y22502 = ~1'b0 ;
  assign y22503 = ~n45814 ;
  assign y22504 = n45815 ;
  assign y22505 = ~1'b0 ;
  assign y22506 = ~1'b0 ;
  assign y22507 = ~1'b0 ;
  assign y22508 = ~1'b0 ;
  assign y22509 = ~n45817 ;
  assign y22510 = n45818 ;
  assign y22511 = n45819 ;
  assign y22512 = ~n31294 ;
  assign y22513 = ~1'b0 ;
  assign y22514 = ~1'b0 ;
  assign y22515 = ~1'b0 ;
  assign y22516 = ~n45820 ;
  assign y22517 = ~1'b0 ;
  assign y22518 = ~1'b0 ;
  assign y22519 = n45821 ;
  assign y22520 = n45826 ;
  assign y22521 = n45827 ;
  assign y22522 = ~1'b0 ;
  assign y22523 = ~n45829 ;
  assign y22524 = ~n45832 ;
  assign y22525 = ~1'b0 ;
  assign y22526 = ~1'b0 ;
  assign y22527 = n45834 ;
  assign y22528 = n45835 ;
  assign y22529 = ~n45836 ;
  assign y22530 = ~n45838 ;
  assign y22531 = n45841 ;
  assign y22532 = ~n45842 ;
  assign y22533 = ~n45846 ;
  assign y22534 = ~n45848 ;
  assign y22535 = n45849 ;
  assign y22536 = ~n45858 ;
  assign y22537 = n45859 ;
  assign y22538 = ~1'b0 ;
  assign y22539 = ~1'b0 ;
  assign y22540 = 1'b0 ;
  assign y22541 = ~n45862 ;
  assign y22542 = n45863 ;
  assign y22543 = n45864 ;
  assign y22544 = ~1'b0 ;
  assign y22545 = ~n45866 ;
  assign y22546 = ~1'b0 ;
  assign y22547 = ~n45870 ;
  assign y22548 = ~1'b0 ;
  assign y22549 = ~n45879 ;
  assign y22550 = n45881 ;
  assign y22551 = ~n45882 ;
  assign y22552 = n45883 ;
  assign y22553 = n45885 ;
  assign y22554 = ~n45892 ;
  assign y22555 = n45894 ;
  assign y22556 = n45899 ;
  assign y22557 = n45909 ;
  assign y22558 = ~n45912 ;
  assign y22559 = ~1'b0 ;
  assign y22560 = ~1'b0 ;
  assign y22561 = ~n45914 ;
  assign y22562 = ~1'b0 ;
  assign y22563 = ~n45915 ;
  assign y22564 = n44318 ;
  assign y22565 = ~n45916 ;
  assign y22566 = n45918 ;
  assign y22567 = n45922 ;
  assign y22568 = ~1'b0 ;
  assign y22569 = ~n45925 ;
  assign y22570 = ~n45927 ;
  assign y22571 = n45930 ;
  assign y22572 = ~n45931 ;
  assign y22573 = n45932 ;
  assign y22574 = ~n45933 ;
  assign y22575 = n45935 ;
  assign y22576 = n45936 ;
  assign y22577 = n45937 ;
  assign y22578 = ~n45938 ;
  assign y22579 = ~n45942 ;
  assign y22580 = n5356 ;
  assign y22581 = n45944 ;
  assign y22582 = ~n26207 ;
  assign y22583 = ~n45948 ;
  assign y22584 = n45950 ;
  assign y22585 = n45951 ;
  assign y22586 = n45954 ;
  assign y22587 = ~n45958 ;
  assign y22588 = n45960 ;
  assign y22589 = n28099 ;
  assign y22590 = ~1'b0 ;
  assign y22591 = n45963 ;
  assign y22592 = ~n45965 ;
  assign y22593 = n45970 ;
  assign y22594 = ~n45972 ;
  assign y22595 = ~1'b0 ;
  assign y22596 = ~n45973 ;
  assign y22597 = ~n45974 ;
  assign y22598 = n45975 ;
  assign y22599 = ~n45977 ;
  assign y22600 = ~n45979 ;
  assign y22601 = ~1'b0 ;
  assign y22602 = n3007 ;
  assign y22603 = ~1'b0 ;
  assign y22604 = ~n45981 ;
  assign y22605 = n45982 ;
  assign y22606 = n45984 ;
  assign y22607 = ~n45990 ;
  assign y22608 = n45999 ;
  assign y22609 = n46006 ;
  assign y22610 = ~1'b0 ;
  assign y22611 = n46008 ;
  assign y22612 = ~1'b0 ;
  assign y22613 = ~n46011 ;
  assign y22614 = ~n46012 ;
  assign y22615 = ~1'b0 ;
  assign y22616 = n46013 ;
  assign y22617 = ~1'b0 ;
  assign y22618 = n46015 ;
  assign y22619 = ~n46016 ;
  assign y22620 = n46018 ;
  assign y22621 = ~1'b0 ;
  assign y22622 = ~1'b0 ;
  assign y22623 = n46019 ;
  assign y22624 = ~1'b0 ;
  assign y22625 = n46020 ;
  assign y22626 = ~n46021 ;
  assign y22627 = ~n46023 ;
  assign y22628 = ~n46024 ;
  assign y22629 = ~n46025 ;
  assign y22630 = ~n46026 ;
  assign y22631 = n46027 ;
  assign y22632 = ~n46028 ;
  assign y22633 = ~1'b0 ;
  assign y22634 = n46030 ;
  assign y22635 = ~n46032 ;
  assign y22636 = n46034 ;
  assign y22637 = ~n46036 ;
  assign y22638 = n46038 ;
  assign y22639 = ~1'b0 ;
  assign y22640 = ~n46039 ;
  assign y22641 = n46040 ;
  assign y22642 = n46044 ;
  assign y22643 = n46046 ;
  assign y22644 = ~n46049 ;
  assign y22645 = 1'b0 ;
  assign y22646 = n46053 ;
  assign y22647 = n46056 ;
  assign y22648 = n46057 ;
  assign y22649 = ~1'b0 ;
  assign y22650 = n46059 ;
  assign y22651 = n46062 ;
  assign y22652 = ~n46063 ;
  assign y22653 = n46069 ;
  assign y22654 = n46071 ;
  assign y22655 = ~1'b0 ;
  assign y22656 = ~1'b0 ;
  assign y22657 = ~1'b0 ;
  assign y22658 = ~n46074 ;
  assign y22659 = n46075 ;
  assign y22660 = n46076 ;
  assign y22661 = n46077 ;
  assign y22662 = ~n46078 ;
  assign y22663 = ~n46080 ;
  assign y22664 = ~n46081 ;
  assign y22665 = ~n46083 ;
  assign y22666 = ~n46085 ;
  assign y22667 = n46087 ;
  assign y22668 = n46088 ;
  assign y22669 = ~1'b0 ;
  assign y22670 = ~n46090 ;
  assign y22671 = n46092 ;
  assign y22672 = ~1'b0 ;
  assign y22673 = n46095 ;
  assign y22674 = n46098 ;
  assign y22675 = n46101 ;
  assign y22676 = ~1'b0 ;
  assign y22677 = ~n46108 ;
  assign y22678 = n46111 ;
  assign y22679 = ~n46112 ;
  assign y22680 = ~1'b0 ;
  assign y22681 = ~1'b0 ;
  assign y22682 = n46113 ;
  assign y22683 = n46116 ;
  assign y22684 = n46117 ;
  assign y22685 = ~1'b0 ;
  assign y22686 = n46118 ;
  assign y22687 = n46122 ;
  assign y22688 = ~n46128 ;
  assign y22689 = ~n46130 ;
  assign y22690 = ~n46132 ;
  assign y22691 = ~n46134 ;
  assign y22692 = n33898 ;
  assign y22693 = ~1'b0 ;
  assign y22694 = ~1'b0 ;
  assign y22695 = ~1'b0 ;
  assign y22696 = n46136 ;
  assign y22697 = n46137 ;
  assign y22698 = ~1'b0 ;
  assign y22699 = ~1'b0 ;
  assign y22700 = ~n46138 ;
  assign y22701 = ~n46139 ;
  assign y22702 = ~n46141 ;
  assign y22703 = ~1'b0 ;
  assign y22704 = ~n46143 ;
  assign y22705 = ~n46146 ;
  assign y22706 = ~n46148 ;
  assign y22707 = ~n46150 ;
  assign y22708 = ~n34439 ;
  assign y22709 = n46152 ;
  assign y22710 = ~n46153 ;
  assign y22711 = ~n46156 ;
  assign y22712 = ~n46158 ;
  assign y22713 = n46160 ;
  assign y22714 = ~n46162 ;
  assign y22715 = n46163 ;
  assign y22716 = ~n46165 ;
  assign y22717 = ~n46171 ;
  assign y22718 = ~n46172 ;
  assign y22719 = n46173 ;
  assign y22720 = ~n46174 ;
  assign y22721 = n46178 ;
  assign y22722 = ~n46179 ;
  assign y22723 = ~n46180 ;
  assign y22724 = n46184 ;
  assign y22725 = ~1'b0 ;
  assign y22726 = n46186 ;
  assign y22727 = 1'b0 ;
  assign y22728 = n46187 ;
  assign y22729 = ~n46190 ;
  assign y22730 = ~n46194 ;
  assign y22731 = ~1'b0 ;
  assign y22732 = ~n46196 ;
  assign y22733 = n407 ;
  assign y22734 = ~1'b0 ;
  assign y22735 = ~1'b0 ;
  assign y22736 = ~n9439 ;
  assign y22737 = ~1'b0 ;
  assign y22738 = ~1'b0 ;
  assign y22739 = ~n46201 ;
  assign y22740 = ~n46208 ;
  assign y22741 = ~n46213 ;
  assign y22742 = n46217 ;
  assign y22743 = n46219 ;
  assign y22744 = ~1'b0 ;
  assign y22745 = ~n46221 ;
  assign y22746 = n46223 ;
endmodule
