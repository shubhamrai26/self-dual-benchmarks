module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 ;
  assign n129 = x106 ^ x93 ^ x27 ;
  assign n130 = x23 & x125 ;
  assign n131 = ~x75 & n130 ;
  assign n132 = x97 ^ x83 ^ 1'b0 ;
  assign n133 = x36 & x112 ;
  assign n134 = n133 ^ x46 ^ 1'b0 ;
  assign n135 = x79 & ~x103 ;
  assign n136 = x105 ^ x3 ^ 1'b0 ;
  assign n137 = x31 & n136 ;
  assign n138 = x103 & x125 ;
  assign n139 = ~x127 & n138 ;
  assign n140 = x107 ^ x11 ^ 1'b0 ;
  assign n141 = ~n139 & n140 ;
  assign n142 = n141 ^ x126 ^ 1'b0 ;
  assign n143 = x65 & n142 ;
  assign n144 = x118 ^ x113 ^ x70 ;
  assign n145 = x96 & x99 ;
  assign n146 = n145 ^ x82 ^ 1'b0 ;
  assign n147 = x100 & ~n146 ;
  assign n148 = n147 ^ x98 ^ 1'b0 ;
  assign n149 = n139 ^ x12 ^ 1'b0 ;
  assign n150 = x46 & ~n149 ;
  assign n151 = x103 ^ x79 ^ 1'b0 ;
  assign n152 = x26 & n151 ;
  assign n153 = x93 ^ x6 ^ x1 ;
  assign n154 = x99 & ~n153 ;
  assign n155 = ~x46 & n154 ;
  assign n156 = ( ~x31 & x38 ) | ( ~x31 & x44 ) | ( x38 & x44 ) ;
  assign n157 = x89 ^ x66 ^ 1'b0 ;
  assign n158 = x62 & n157 ;
  assign n159 = x25 & x65 ;
  assign n162 = x118 ^ x30 ^ 1'b0 ;
  assign n163 = x20 & n162 ;
  assign n160 = x124 ^ x48 ^ 1'b0 ;
  assign n161 = x89 & n160 ;
  assign n164 = n163 ^ n161 ^ 1'b0 ;
  assign n165 = ( x7 & x16 ) | ( x7 & ~x36 ) | ( x16 & ~x36 ) ;
  assign n166 = n146 ^ x52 ^ 1'b0 ;
  assign n167 = x108 & ~n166 ;
  assign n168 = x18 & x91 ;
  assign n169 = ~n167 & n168 ;
  assign n170 = n165 & ~n169 ;
  assign n171 = n170 ^ x18 ^ 1'b0 ;
  assign n172 = x98 ^ x62 ^ 1'b0 ;
  assign n173 = x68 & n172 ;
  assign n174 = x68 & n163 ;
  assign n175 = n174 ^ x58 ^ 1'b0 ;
  assign n176 = n173 & ~n175 ;
  assign n177 = n176 ^ x30 ^ 1'b0 ;
  assign n178 = x122 ^ x104 ^ 1'b0 ;
  assign n179 = x5 & n178 ;
  assign n180 = x10 ^ x4 ^ 1'b0 ;
  assign n181 = n179 & n180 ;
  assign n182 = x37 & x104 ;
  assign n183 = ~x73 & n182 ;
  assign n184 = x0 & x113 ;
  assign n185 = ~n141 & n184 ;
  assign n187 = x16 ^ x2 ^ 1'b0 ;
  assign n188 = x7 & n187 ;
  assign n186 = x82 & x83 ;
  assign n189 = n188 ^ n186 ^ 1'b0 ;
  assign n190 = ~x9 & x58 ;
  assign n191 = x15 & x116 ;
  assign n192 = n191 ^ n143 ^ 1'b0 ;
  assign n194 = ~x24 & x40 ;
  assign n195 = n139 & n194 ;
  assign n193 = x97 & x121 ;
  assign n196 = n195 ^ n193 ^ 1'b0 ;
  assign n202 = x63 & x78 ;
  assign n203 = n202 ^ n131 ^ 1'b0 ;
  assign n197 = x59 & x118 ;
  assign n198 = n197 ^ x102 ^ 1'b0 ;
  assign n199 = x79 & ~n198 ;
  assign n200 = n199 ^ x71 ^ 1'b0 ;
  assign n201 = n200 ^ n194 ^ x58 ;
  assign n204 = n203 ^ n201 ^ 1'b0 ;
  assign n205 = x45 & n204 ;
  assign n206 = x42 & x91 ;
  assign n207 = ~x44 & n206 ;
  assign n208 = ( x19 & n164 ) | ( x19 & n207 ) | ( n164 & n207 ) ;
  assign n209 = x95 ^ x2 ^ 1'b0 ;
  assign n210 = x74 & n209 ;
  assign n211 = ~x2 & n210 ;
  assign n212 = x67 ^ x59 ^ 1'b0 ;
  assign n213 = x70 & n212 ;
  assign n214 = ~n129 & n213 ;
  assign n215 = ~x29 & n214 ;
  assign n216 = x110 | n215 ;
  assign n217 = n165 | n171 ;
  assign n218 = x0 & x13 ;
  assign n219 = n218 ^ x9 ^ 1'b0 ;
  assign n220 = n219 ^ x125 ^ x47 ;
  assign n221 = x49 & x112 ;
  assign n222 = x54 ^ x24 ^ x13 ;
  assign n223 = n219 | n222 ;
  assign n224 = n223 ^ x4 ^ 1'b0 ;
  assign n225 = x108 & ~n224 ;
  assign n228 = x99 ^ x83 ^ 1'b0 ;
  assign n229 = x7 & n228 ;
  assign n232 = n229 ^ x39 ^ 1'b0 ;
  assign n233 = x114 & n232 ;
  assign n226 = x3 & x30 ;
  assign n227 = ~x18 & n226 ;
  assign n230 = n229 ^ n175 ^ 1'b0 ;
  assign n231 = ( x76 & n227 ) | ( x76 & n230 ) | ( n227 & n230 ) ;
  assign n234 = n233 ^ n231 ^ 1'b0 ;
  assign n235 = x50 & n234 ;
  assign n236 = x72 & n203 ;
  assign n237 = n236 ^ n139 ^ 1'b0 ;
  assign n238 = ~x5 & x69 ;
  assign n239 = x29 ^ x4 ^ 1'b0 ;
  assign n240 = x121 & n239 ;
  assign n241 = x57 ^ x42 ^ 1'b0 ;
  assign n242 = x31 & n241 ;
  assign n243 = ~n240 & n242 ;
  assign n244 = n167 & n233 ;
  assign n245 = n244 ^ n179 ^ 1'b0 ;
  assign n246 = x59 & ~n245 ;
  assign n247 = n246 ^ n135 ^ 1'b0 ;
  assign n248 = n179 & n247 ;
  assign n249 = x51 & x82 ;
  assign n250 = n249 ^ n165 ^ 1'b0 ;
  assign n251 = x53 | n250 ;
  assign n252 = ( x52 & x56 ) | ( x52 & ~n242 ) | ( x56 & ~n242 ) ;
  assign n253 = x82 & x106 ;
  assign n254 = n129 & n253 ;
  assign n255 = n254 ^ x108 ^ 1'b0 ;
  assign n256 = n252 & ~n255 ;
  assign n257 = x24 & n256 ;
  assign n258 = n257 ^ n158 ^ 1'b0 ;
  assign n259 = ( ~x50 & n181 ) | ( ~x50 & n238 ) | ( n181 & n238 ) ;
  assign n267 = n158 ^ x1 ^ 1'b0 ;
  assign n260 = x2 & x87 ;
  assign n261 = ~x67 & n260 ;
  assign n262 = x127 ^ x27 ^ x9 ;
  assign n263 = n262 ^ n159 ^ 1'b0 ;
  assign n264 = n135 & ~n263 ;
  assign n265 = n264 ^ x2 ^ 1'b0 ;
  assign n266 = ~n261 & n265 ;
  assign n268 = n267 ^ n266 ^ 1'b0 ;
  assign n269 = n268 ^ n169 ^ 1'b0 ;
  assign n270 = x100 & n269 ;
  assign n271 = x43 & x102 ;
  assign n272 = n271 ^ x37 ^ 1'b0 ;
  assign n273 = n272 ^ n163 ^ 1'b0 ;
  assign n275 = x71 & x98 ;
  assign n276 = n275 ^ x16 ^ 1'b0 ;
  assign n274 = x39 & x121 ;
  assign n277 = n276 ^ n274 ^ 1'b0 ;
  assign n278 = n256 & n277 ;
  assign n279 = ~x69 & n278 ;
  assign n280 = x6 & ~n279 ;
  assign n281 = n280 ^ n219 ^ 1'b0 ;
  assign n282 = x122 ^ x23 ^ 1'b0 ;
  assign n283 = x14 & n282 ;
  assign n284 = x111 & n283 ;
  assign n285 = n208 & n284 ;
  assign n286 = n281 & ~n285 ;
  assign n287 = ~x14 & n286 ;
  assign n288 = n261 ^ x91 ^ 1'b0 ;
  assign n289 = n288 ^ n243 ^ 1'b0 ;
  assign n290 = x88 & ~x109 ;
  assign n291 = n179 & n246 ;
  assign n292 = ~n290 & n291 ;
  assign n293 = ~x49 & x56 ;
  assign n294 = x86 ^ x55 ^ 1'b0 ;
  assign n295 = x84 & ~n175 ;
  assign n296 = n295 ^ x81 ^ 1'b0 ;
  assign n297 = n141 & n296 ;
  assign n298 = x29 & n163 ;
  assign n299 = ~n290 & n298 ;
  assign n300 = x66 & n299 ;
  assign n301 = n250 ^ n181 ^ 1'b0 ;
  assign n302 = n300 | n301 ;
  assign n303 = x53 & n242 ;
  assign n304 = n303 ^ n134 ^ 1'b0 ;
  assign n306 = x90 & x114 ;
  assign n307 = n306 ^ x20 ^ 1'b0 ;
  assign n305 = x58 & ~n248 ;
  assign n308 = n307 ^ n305 ^ 1'b0 ;
  assign n309 = n211 ^ x13 ^ 1'b0 ;
  assign n310 = n276 | n309 ;
  assign n311 = ~n238 & n310 ;
  assign n313 = n238 | n287 ;
  assign n314 = n248 | n313 ;
  assign n312 = x38 & ~n245 ;
  assign n315 = n314 ^ n312 ^ 1'b0 ;
  assign n316 = ( x8 & ~x97 ) | ( x8 & n264 ) | ( ~x97 & n264 ) ;
  assign n317 = ~n175 & n316 ;
  assign n318 = n317 ^ n224 ^ 1'b0 ;
  assign n319 = x74 ^ x31 ^ 1'b0 ;
  assign n320 = x69 & n319 ;
  assign n321 = x31 & n177 ;
  assign n322 = ~n288 & n321 ;
  assign n323 = n322 ^ x111 ^ 1'b0 ;
  assign n324 = n159 | n323 ;
  assign n325 = n270 ^ x48 ^ 1'b0 ;
  assign n326 = x34 & n314 ;
  assign n327 = n213 & ~n292 ;
  assign n328 = n146 & n327 ;
  assign n329 = n139 | n222 ;
  assign n330 = n329 ^ x9 ^ 1'b0 ;
  assign n331 = n179 ^ x51 ^ 1'b0 ;
  assign n332 = n330 & n331 ;
  assign n333 = ~x35 & n332 ;
  assign n334 = n135 ^ x107 ^ 1'b0 ;
  assign n335 = ~n259 & n334 ;
  assign n336 = n208 ^ x25 ^ 1'b0 ;
  assign n337 = n141 & n240 ;
  assign n338 = n337 ^ n229 ^ 1'b0 ;
  assign n339 = n338 ^ n252 ^ 1'b0 ;
  assign n340 = n326 ^ x19 ^ 1'b0 ;
  assign n341 = x61 & n314 ;
  assign n342 = n341 ^ n339 ^ 1'b0 ;
  assign n343 = ~x79 & x95 ;
  assign n344 = ( x73 & ~x74 ) | ( x73 & n129 ) | ( ~x74 & n129 ) ;
  assign n345 = x16 & n325 ;
  assign n346 = n345 ^ x112 ^ 1'b0 ;
  assign n356 = n194 ^ n175 ^ n144 ;
  assign n357 = n330 & ~n356 ;
  assign n358 = n357 ^ x53 ^ 1'b0 ;
  assign n348 = x49 ^ x33 ^ 1'b0 ;
  assign n349 = n173 & n348 ;
  assign n350 = x75 & x125 ;
  assign n351 = n350 ^ n167 ^ 1'b0 ;
  assign n352 = n349 & ~n351 ;
  assign n353 = ~x64 & n352 ;
  assign n354 = x82 & ~n353 ;
  assign n355 = ~x107 & n354 ;
  assign n359 = n358 ^ n355 ^ n246 ;
  assign n347 = x82 & x99 ;
  assign n360 = n359 ^ n347 ^ 1'b0 ;
  assign n361 = x64 | n360 ;
  assign n362 = n283 ^ x32 ^ 1'b0 ;
  assign n363 = n229 & n362 ;
  assign n364 = n363 ^ n353 ^ 1'b0 ;
  assign n365 = x44 & ~n364 ;
  assign n366 = ~n134 & n195 ;
  assign n367 = ~x51 & n366 ;
  assign n368 = n315 | n367 ;
  assign n369 = n216 & ~n368 ;
  assign n370 = x53 ^ x26 ^ 1'b0 ;
  assign n371 = ~n169 & n370 ;
  assign n372 = x81 & n159 ;
  assign n373 = n164 & n372 ;
  assign n374 = n371 & ~n373 ;
  assign n375 = n374 ^ n181 ^ 1'b0 ;
  assign n376 = x7 & ~x114 ;
  assign n377 = x33 & x112 ;
  assign n378 = ~n143 & n377 ;
  assign n379 = x68 & x113 ;
  assign n380 = ~x125 & n379 ;
  assign n381 = x10 & n380 ;
  assign n382 = ~n378 & n381 ;
  assign n383 = n382 ^ n221 ^ 1'b0 ;
  assign n384 = x117 & ~n383 ;
  assign n385 = n376 & n384 ;
  assign n386 = n353 ^ x89 ^ 1'b0 ;
  assign n387 = x66 & ~n386 ;
  assign n388 = n163 & ~n268 ;
  assign n389 = ~x127 & n388 ;
  assign n390 = n314 ^ x59 ^ 1'b0 ;
  assign n391 = x21 | n297 ;
  assign n392 = x98 ^ x8 ^ 1'b0 ;
  assign n393 = n259 | n392 ;
  assign n394 = n393 ^ n248 ^ 1'b0 ;
  assign n395 = x46 & n217 ;
  assign n396 = n395 ^ n281 ^ 1'b0 ;
  assign n397 = x94 & ~n220 ;
  assign n398 = n396 | n397 ;
  assign n399 = n273 & ~n398 ;
  assign n400 = ( x8 & ~x53 ) | ( x8 & n141 ) | ( ~x53 & n141 ) ;
  assign n401 = n283 ^ x19 ^ 1'b0 ;
  assign n402 = x99 & n401 ;
  assign n403 = n161 & n402 ;
  assign n404 = n403 ^ n167 ^ 1'b0 ;
  assign n405 = x55 & ~n404 ;
  assign n406 = n405 ^ x105 ^ 1'b0 ;
  assign n407 = n404 ^ n201 ^ 1'b0 ;
  assign n408 = x35 ^ x8 ^ 1'b0 ;
  assign n409 = ~n164 & n408 ;
  assign n410 = x31 & ~n402 ;
  assign n411 = x97 & x115 ;
  assign n412 = ~n201 & n411 ;
  assign n413 = n285 ^ x12 ^ 1'b0 ;
  assign n414 = ( x37 & ~x122 ) | ( x37 & n233 ) | ( ~x122 & n233 ) ;
  assign n415 = n373 | n414 ;
  assign n416 = x96 & n415 ;
  assign n417 = n318 & n416 ;
  assign n418 = ~x53 & x115 ;
  assign n419 = n207 ^ x45 ^ 1'b0 ;
  assign n420 = n201 & ~n419 ;
  assign n421 = n420 ^ x11 ^ 1'b0 ;
  assign n422 = x20 & n421 ;
  assign n423 = n252 ^ x44 ^ 1'b0 ;
  assign n424 = x57 & n423 ;
  assign n425 = ( ~x68 & x93 ) | ( ~x68 & x108 ) | ( x93 & x108 ) ;
  assign n426 = ~n219 & n425 ;
  assign n427 = n426 ^ x117 ^ 1'b0 ;
  assign n428 = x57 & n287 ;
  assign n429 = n396 ^ n167 ^ 1'b0 ;
  assign n430 = n428 | n429 ;
  assign n431 = x81 & ~n367 ;
  assign n432 = ~x87 & n431 ;
  assign n433 = n304 ^ n231 ^ 1'b0 ;
  assign n434 = x45 & ~n433 ;
  assign n435 = ~n432 & n434 ;
  assign n436 = x85 | n250 ;
  assign n437 = n425 ^ n141 ^ 1'b0 ;
  assign n438 = ~n146 & n437 ;
  assign n439 = n438 ^ n242 ^ n229 ;
  assign n440 = x15 & n150 ;
  assign n441 = ~x119 & n440 ;
  assign n442 = ~n287 & n371 ;
  assign n443 = x43 & n156 ;
  assign n444 = n443 ^ x33 ^ 1'b0 ;
  assign n445 = n296 & ~n378 ;
  assign n446 = ~n299 & n445 ;
  assign n447 = x60 & ~n446 ;
  assign n448 = n447 ^ n216 ^ 1'b0 ;
  assign n449 = x63 & n205 ;
  assign n450 = n449 ^ n296 ^ 1'b0 ;
  assign n451 = n450 ^ n400 ^ n285 ;
  assign n452 = x14 & n451 ;
  assign n453 = ~n448 & n452 ;
  assign n454 = x11 & x112 ;
  assign n455 = ~x101 & n454 ;
  assign n456 = n455 ^ x23 ^ 1'b0 ;
  assign n457 = ~n177 & n189 ;
  assign n458 = n188 & ~n375 ;
  assign n459 = n457 & n458 ;
  assign n460 = n316 ^ x69 ^ 1'b0 ;
  assign n461 = ~n459 & n460 ;
  assign n462 = n150 ^ x65 ^ 1'b0 ;
  assign n463 = ~n432 & n462 ;
  assign n464 = x74 & ~n463 ;
  assign n465 = n308 & ~n444 ;
  assign n466 = ~n270 & n465 ;
  assign n467 = n466 ^ n279 ^ 1'b0 ;
  assign n468 = ~n173 & n446 ;
  assign n469 = ~x85 & x115 ;
  assign n470 = n324 | n469 ;
  assign n471 = n287 & ~n470 ;
  assign n472 = x94 & ~n469 ;
  assign n473 = n472 ^ n137 ^ 1'b0 ;
  assign n474 = x118 & n473 ;
  assign n475 = ( ~x31 & x119 ) | ( ~x31 & n304 ) | ( x119 & n304 ) ;
  assign n476 = n475 ^ x67 ^ 1'b0 ;
  assign n477 = x40 & n476 ;
  assign n478 = x50 & ~n477 ;
  assign n479 = n262 | n432 ;
  assign n480 = n171 & ~n479 ;
  assign n481 = n439 & ~n480 ;
  assign n482 = n481 ^ n208 ^ 1'b0 ;
  assign n483 = n159 & n356 ;
  assign n484 = ( ~x37 & n353 ) | ( ~x37 & n483 ) | ( n353 & n483 ) ;
  assign n485 = x46 ^ x23 ^ 1'b0 ;
  assign n486 = n485 ^ n404 ^ 1'b0 ;
  assign n487 = ~n404 & n486 ;
  assign n488 = n179 & ~n328 ;
  assign n489 = n488 ^ n333 ^ 1'b0 ;
  assign n490 = n194 & n330 ;
  assign n491 = n489 & n490 ;
  assign n492 = n324 & ~n344 ;
  assign n493 = n316 ^ x97 ^ 1'b0 ;
  assign n494 = n493 ^ x126 ^ x77 ;
  assign n495 = x5 & n167 ;
  assign n496 = ~x125 & n495 ;
  assign n497 = ~x39 & x40 ;
  assign n498 = n497 ^ x81 ^ 1'b0 ;
  assign n499 = n131 | n498 ;
  assign n500 = n463 ^ x106 ^ 1'b0 ;
  assign n501 = n499 | n500 ;
  assign n502 = n392 & ~n501 ;
  assign n503 = n365 & ~n502 ;
  assign n504 = n289 ^ x61 ^ 1'b0 ;
  assign n505 = ~n501 & n504 ;
  assign n506 = n505 ^ n354 ^ 1'b0 ;
  assign n507 = n171 ^ x55 ^ x32 ;
  assign n508 = n323 & n507 ;
  assign n509 = x42 & n242 ;
  assign n510 = n509 ^ n321 ^ 1'b0 ;
  assign n511 = n461 & n467 ;
  assign n512 = n510 & n511 ;
  assign n513 = x60 & x73 ;
  assign n514 = n513 ^ x114 ^ 1'b0 ;
  assign n515 = n514 ^ x9 ^ 1'b0 ;
  assign n516 = x92 & ~n515 ;
  assign n517 = x54 & n516 ;
  assign n518 = n517 ^ n242 ^ 1'b0 ;
  assign n519 = n281 ^ x52 ^ 1'b0 ;
  assign n520 = n519 ^ n299 ^ 1'b0 ;
  assign n521 = n261 | n474 ;
  assign n522 = n521 ^ n453 ^ 1'b0 ;
  assign n523 = n201 & ~n338 ;
  assign n524 = n523 ^ n466 ^ 1'b0 ;
  assign n525 = n445 ^ x124 ^ 1'b0 ;
  assign n526 = n504 & ~n525 ;
  assign n527 = n277 ^ n210 ^ 1'b0 ;
  assign n528 = n526 & n527 ;
  assign n529 = n528 ^ n134 ^ 1'b0 ;
  assign n530 = n529 ^ x15 ^ 1'b0 ;
  assign n531 = n522 ^ x24 ^ x9 ;
  assign n532 = x21 ^ x20 ^ 1'b0 ;
  assign n533 = x109 & n532 ;
  assign n535 = n196 ^ n135 ^ 1'b0 ;
  assign n536 = x56 & n535 ;
  assign n537 = n536 ^ x6 ^ 1'b0 ;
  assign n538 = n336 ^ n287 ^ 1'b0 ;
  assign n539 = ( ~n320 & n537 ) | ( ~n320 & n538 ) | ( n537 & n538 ) ;
  assign n534 = x5 & x45 ;
  assign n540 = n539 ^ n534 ^ 1'b0 ;
  assign n541 = n215 | n261 ;
  assign n542 = n541 ^ x21 ^ 1'b0 ;
  assign n543 = x105 & n320 ;
  assign n544 = n543 ^ x9 ^ 1'b0 ;
  assign n545 = n542 & n544 ;
  assign n546 = n545 ^ x96 ^ 1'b0 ;
  assign n547 = n467 & n546 ;
  assign n548 = n135 & n230 ;
  assign n549 = n432 & n491 ;
  assign n550 = ~x26 & n477 ;
  assign n551 = x42 & ~n380 ;
  assign n552 = n155 & n551 ;
  assign n553 = n336 ^ n129 ^ 1'b0 ;
  assign n554 = ~n323 & n553 ;
  assign n555 = ~n354 & n554 ;
  assign n556 = x73 & ~n555 ;
  assign n557 = n556 ^ x9 ^ 1'b0 ;
  assign n558 = n552 & ~n557 ;
  assign n559 = ~n189 & n270 ;
  assign n560 = ~x7 & n559 ;
  assign n561 = n297 | n560 ;
  assign n562 = x99 | n561 ;
  assign n563 = x123 & n349 ;
  assign n564 = n563 ^ n413 ^ 1'b0 ;
  assign n565 = ~n279 & n333 ;
  assign n566 = n565 ^ n188 ^ 1'b0 ;
  assign n567 = n510 ^ n139 ^ 1'b0 ;
  assign n568 = ( ~n196 & n459 ) | ( ~n196 & n567 ) | ( n459 & n567 ) ;
  assign n569 = x77 & n267 ;
  assign n570 = ~x94 & n569 ;
  assign n571 = n336 | n570 ;
  assign n572 = n164 & n400 ;
  assign n573 = n432 | n572 ;
  assign n574 = n373 & ~n573 ;
  assign n575 = n451 ^ n222 ^ n148 ;
  assign n576 = n560 ^ x9 ^ 1'b0 ;
  assign n577 = n420 ^ x116 ^ x53 ;
  assign n578 = x58 & ~n445 ;
  assign n579 = n134 & n578 ;
  assign n580 = n335 & ~n358 ;
  assign n581 = n385 & n580 ;
  assign n582 = x94 & ~x126 ;
  assign n583 = x11 & ~n582 ;
  assign n584 = n349 & ~n583 ;
  assign n587 = x1 & n152 ;
  assign n588 = n587 ^ n277 ^ 1'b0 ;
  assign n585 = n173 ^ x45 ^ 1'b0 ;
  assign n586 = ~n148 & n585 ;
  assign n589 = n588 ^ n586 ^ 1'b0 ;
  assign n590 = n391 | n589 ;
  assign n591 = n333 ^ x15 ^ 1'b0 ;
  assign n592 = x71 & x112 ;
  assign n593 = ~n229 & n592 ;
  assign n594 = ~n591 & n593 ;
  assign n595 = x18 & x76 ;
  assign n596 = n595 ^ n444 ^ 1'b0 ;
  assign n597 = n409 & ~n596 ;
  assign n599 = x119 & ~n153 ;
  assign n600 = n599 ^ x0 ^ 1'b0 ;
  assign n598 = x78 & x94 ;
  assign n601 = n600 ^ n598 ^ 1'b0 ;
  assign n602 = n190 ^ x127 ^ 1'b0 ;
  assign n603 = ~n296 & n602 ;
  assign n604 = n603 ^ x107 ^ 1'b0 ;
  assign n605 = n604 ^ n292 ^ 1'b0 ;
  assign n606 = n169 | n605 ;
  assign n607 = n601 | n606 ;
  assign n608 = n375 & n607 ;
  assign n609 = ~n153 & n293 ;
  assign n610 = n609 ^ x60 ^ 1'b0 ;
  assign n611 = n593 ^ n501 ^ 1'b0 ;
  assign n612 = n576 & n611 ;
  assign n613 = x85 | n439 ;
  assign n622 = n425 ^ x106 ^ 1'b0 ;
  assign n623 = n179 & n622 ;
  assign n614 = n256 ^ x54 ^ 1'b0 ;
  assign n615 = n194 & ~n614 ;
  assign n616 = n615 ^ n216 ^ 1'b0 ;
  assign n617 = n376 ^ x122 ^ 1'b0 ;
  assign n618 = x44 & ~n617 ;
  assign n619 = n616 & n618 ;
  assign n620 = n619 ^ n471 ^ 1'b0 ;
  assign n621 = x103 & n620 ;
  assign n624 = n623 ^ n621 ^ 1'b0 ;
  assign n625 = n210 ^ x94 ^ x60 ;
  assign n626 = n625 ^ n318 ^ 1'b0 ;
  assign n627 = n194 & n626 ;
  assign n628 = n627 ^ x111 ^ 1'b0 ;
  assign n629 = n475 & n628 ;
  assign n630 = x103 ^ x68 ^ 1'b0 ;
  assign n631 = n373 | n514 ;
  assign n632 = x59 | n631 ;
  assign n633 = n632 ^ x15 ^ 1'b0 ;
  assign n634 = x17 & n520 ;
  assign n635 = x69 & n181 ;
  assign n636 = n146 & n635 ;
  assign n637 = x59 & n290 ;
  assign n638 = ~n163 & n637 ;
  assign n639 = n603 & ~n638 ;
  assign n640 = ~n607 & n639 ;
  assign n644 = n235 & n475 ;
  assign n645 = n644 ^ n369 ^ 1'b0 ;
  assign n641 = x0 & n242 ;
  assign n642 = ~x68 & n641 ;
  assign n643 = x92 & ~n642 ;
  assign n646 = n645 ^ n643 ^ 1'b0 ;
  assign n647 = x5 & n646 ;
  assign n654 = x12 & ~n287 ;
  assign n655 = n654 ^ n638 ^ 1'b0 ;
  assign n649 = n381 & ~n392 ;
  assign n650 = ~x106 & n649 ;
  assign n648 = ~x26 & n252 ;
  assign n651 = n650 ^ n648 ^ 1'b0 ;
  assign n652 = n354 & n651 ;
  assign n653 = x13 & n652 ;
  assign n656 = n655 ^ n653 ^ 1'b0 ;
  assign n661 = x54 & n475 ;
  assign n662 = ~x100 & n661 ;
  assign n657 = n553 ^ n383 ^ 1'b0 ;
  assign n658 = x11 & ~n657 ;
  assign n659 = x8 & n658 ;
  assign n660 = n659 ^ n407 ^ 1'b0 ;
  assign n663 = n662 ^ n660 ^ 1'b0 ;
  assign n664 = n333 ^ x55 ^ 1'b0 ;
  assign n665 = n550 & n664 ;
  assign n666 = n353 ^ n196 ^ 1'b0 ;
  assign n667 = ~n402 & n647 ;
  assign n668 = n201 & n230 ;
  assign n669 = n668 ^ x17 ^ 1'b0 ;
  assign n670 = n669 ^ n487 ^ 1'b0 ;
  assign n671 = x3 & n670 ;
  assign n672 = n528 ^ x73 ^ x35 ;
  assign n673 = n672 ^ n288 ^ 1'b0 ;
  assign n674 = n321 & ~n673 ;
  assign n675 = n674 ^ x124 ^ 1'b0 ;
  assign n676 = x66 & x74 ;
  assign n677 = n614 & n676 ;
  assign n678 = n457 ^ n355 ^ 1'b0 ;
  assign n679 = ~n171 & n678 ;
  assign n680 = n677 & n679 ;
  assign n681 = n243 & ~n680 ;
  assign n682 = n614 ^ x126 ^ 1'b0 ;
  assign n683 = n169 | n682 ;
  assign n684 = n683 ^ x3 ^ 1'b0 ;
  assign n685 = x91 & ~n684 ;
  assign n686 = ~x60 & n685 ;
  assign n687 = n189 & n509 ;
  assign n688 = n528 & n687 ;
  assign n689 = n688 ^ n512 ^ 1'b0 ;
  assign n690 = ~n406 & n689 ;
  assign n691 = ~n378 & n408 ;
  assign n692 = ~n504 & n691 ;
  assign n693 = n200 ^ x12 ^ 1'b0 ;
  assign n694 = n656 ^ n213 ^ 1'b0 ;
  assign n695 = ~n258 & n557 ;
  assign n696 = n624 ^ n381 ^ 1'b0 ;
  assign n697 = n316 ^ n153 ^ 1'b0 ;
  assign n698 = x84 & ~n697 ;
  assign n700 = n356 ^ x12 ^ 1'b0 ;
  assign n699 = x91 & ~n339 ;
  assign n701 = n700 ^ n699 ^ 1'b0 ;
  assign n702 = n652 ^ n494 ^ 1'b0 ;
  assign n703 = n535 ^ n281 ^ 1'b0 ;
  assign n704 = n390 & ~n638 ;
  assign n705 = x101 & n433 ;
  assign n706 = n507 ^ n281 ^ 1'b0 ;
  assign n707 = ~n216 & n706 ;
  assign n708 = n707 ^ n497 ^ 1'b0 ;
  assign n709 = n438 ^ x64 ^ x12 ;
  assign n710 = x25 & ~n709 ;
  assign n711 = n710 ^ x63 ^ 1'b0 ;
  assign n712 = n627 & ~n711 ;
  assign n713 = n708 & n712 ;
  assign n714 = n200 ^ n134 ^ 1'b0 ;
  assign n715 = ~n131 & n714 ;
  assign n716 = n715 ^ n512 ^ 1'b0 ;
  assign n717 = x35 ^ x21 ^ 1'b0 ;
  assign n718 = n717 ^ n205 ^ 1'b0 ;
  assign n719 = n718 ^ n281 ^ 1'b0 ;
  assign n720 = n529 | n719 ;
  assign n721 = x42 ^ x30 ^ 1'b0 ;
  assign n722 = ( n153 & n254 ) | ( n153 & ~n721 ) | ( n254 & ~n721 ) ;
  assign n723 = n230 & ~n297 ;
  assign n724 = n723 ^ n537 ^ 1'b0 ;
  assign n725 = ( n173 & ~n483 ) | ( n173 & n724 ) | ( ~n483 & n724 ) ;
  assign n726 = n725 ^ x72 ^ 1'b0 ;
  assign n727 = n220 & n726 ;
  assign n728 = x90 & ~x118 ;
  assign n729 = n221 | n704 ;
  assign n730 = n555 ^ n225 ^ 1'b0 ;
  assign n731 = x104 & n730 ;
  assign n732 = n647 ^ x105 ^ 1'b0 ;
  assign n733 = ~n300 & n732 ;
  assign n734 = ~n200 & n733 ;
  assign n735 = n432 & n734 ;
  assign n740 = n243 & ~n514 ;
  assign n741 = n740 ^ n207 ^ 1'b0 ;
  assign n736 = n158 & n237 ;
  assign n737 = n736 ^ x10 ^ 1'b0 ;
  assign n738 = n705 ^ n616 ^ 1'b0 ;
  assign n739 = ~n737 & n738 ;
  assign n742 = n741 ^ n739 ^ n351 ;
  assign n743 = x70 & n456 ;
  assign n744 = n614 & n743 ;
  assign n745 = n330 ^ n144 ^ 1'b0 ;
  assign n746 = n333 & ~n737 ;
  assign n747 = ~n224 & n746 ;
  assign n748 = n422 & ~n747 ;
  assign n749 = n406 & n748 ;
  assign n750 = x26 & x106 ;
  assign n752 = n185 | n225 ;
  assign n753 = n752 ^ n183 ^ 1'b0 ;
  assign n754 = x106 ^ x35 ^ 1'b0 ;
  assign n755 = n754 ^ x75 ^ 1'b0 ;
  assign n756 = n753 & ~n755 ;
  assign n751 = x76 & ~n740 ;
  assign n757 = n756 ^ n751 ^ 1'b0 ;
  assign n758 = n264 & ~n514 ;
  assign n759 = ~x68 & n758 ;
  assign n760 = n759 ^ x120 ^ 1'b0 ;
  assign n761 = n367 | n760 ;
  assign n762 = n328 ^ x48 ^ 1'b0 ;
  assign n763 = n224 & ~n762 ;
  assign n764 = ( n336 & n442 ) | ( n336 & ~n450 ) | ( n442 & ~n450 ) ;
  assign n765 = x91 & ~n155 ;
  assign n766 = ~x10 & n765 ;
  assign n767 = n173 | n250 ;
  assign n768 = n320 | n767 ;
  assign n769 = ~n766 & n768 ;
  assign n770 = n769 ^ x105 ^ 1'b0 ;
  assign n771 = x5 & ~n338 ;
  assign n772 = ~n439 & n771 ;
  assign n773 = n772 ^ x37 ^ 1'b0 ;
  assign n774 = n311 & ~n773 ;
  assign n775 = n774 ^ n367 ^ 1'b0 ;
  assign n776 = n351 ^ x8 ^ 1'b0 ;
  assign n777 = n687 ^ n250 ^ 1'b0 ;
  assign n778 = n776 | n777 ;
  assign n780 = ~n300 & n639 ;
  assign n781 = ~n538 & n780 ;
  assign n779 = n252 & n409 ;
  assign n782 = n781 ^ n779 ^ 1'b0 ;
  assign n783 = x15 & ~x81 ;
  assign n784 = x119 & ~n267 ;
  assign n785 = n783 | n784 ;
  assign n786 = n290 | n373 ;
  assign n787 = n786 ^ n200 ^ 1'b0 ;
  assign n788 = ~n614 & n787 ;
  assign n791 = n233 ^ x104 ^ 1'b0 ;
  assign n792 = x48 & n791 ;
  assign n789 = n165 ^ x69 ^ 1'b0 ;
  assign n790 = x99 & n789 ;
  assign n793 = n792 ^ n790 ^ 1'b0 ;
  assign n794 = n415 ^ x75 ^ 1'b0 ;
  assign n799 = ~n413 & n489 ;
  assign n800 = n799 ^ n408 ^ n264 ;
  assign n795 = x55 & n544 ;
  assign n796 = n795 ^ x23 ^ 1'b0 ;
  assign n797 = n796 ^ n566 ^ 1'b0 ;
  assign n798 = x98 & n797 ;
  assign n801 = n800 ^ n798 ^ 1'b0 ;
  assign n802 = x42 & ~n645 ;
  assign n803 = x31 & ~n571 ;
  assign n804 = ~n359 & n803 ;
  assign n805 = ~n245 & n804 ;
  assign n806 = n340 & ~n600 ;
  assign n807 = x96 ^ x11 ^ 1'b0 ;
  assign n808 = ~n761 & n807 ;
  assign n809 = ~n717 & n753 ;
  assign n810 = n167 | n788 ;
  assign n811 = n477 ^ x40 ^ 1'b0 ;
  assign n812 = x124 & n811 ;
  assign n813 = n812 ^ n692 ^ x61 ;
  assign n814 = n224 & n801 ;
  assign n816 = n173 & n325 ;
  assign n817 = n216 & n816 ;
  assign n818 = n205 & ~n817 ;
  assign n819 = n818 ^ x47 ^ 1'b0 ;
  assign n820 = n819 ^ x46 ^ 1'b0 ;
  assign n821 = n579 | n820 ;
  assign n822 = n821 ^ x74 ^ 1'b0 ;
  assign n823 = ( n361 & ~n603 ) | ( n361 & n822 ) | ( ~n603 & n822 ) ;
  assign n815 = n564 & n813 ;
  assign n824 = n823 ^ n815 ^ 1'b0 ;
  assign n825 = n540 | n624 ;
  assign n826 = n739 ^ n459 ^ 1'b0 ;
  assign n827 = ~n245 & n289 ;
  assign n828 = n827 ^ x110 ^ 1'b0 ;
  assign n829 = n828 ^ n363 ^ 1'b0 ;
  assign n830 = n340 | n829 ;
  assign n831 = n830 ^ n645 ^ 1'b0 ;
  assign n832 = n831 ^ n721 ^ 1'b0 ;
  assign n833 = n832 ^ n155 ^ 1'b0 ;
  assign n834 = ( n351 & ~n516 ) | ( n351 & n547 ) | ( ~n516 & n547 ) ;
  assign n835 = n242 | n834 ;
  assign n836 = ~x18 & n835 ;
  assign n837 = n586 & ~n810 ;
  assign n838 = n296 ^ n240 ^ 1'b0 ;
  assign n839 = n200 | n838 ;
  assign n840 = n839 ^ n332 ^ 1'b0 ;
  assign n841 = n595 & ~n840 ;
  assign n842 = ~n163 & n642 ;
  assign n843 = n360 ^ n194 ^ 1'b0 ;
  assign n844 = ~x12 & n843 ;
  assign n845 = n542 | n740 ;
  assign n846 = n817 ^ n396 ^ 1'b0 ;
  assign n849 = x0 & ~x67 ;
  assign n850 = ~n134 & n849 ;
  assign n851 = ~n667 & n850 ;
  assign n852 = x55 | n851 ;
  assign n847 = n417 ^ x85 ^ 1'b0 ;
  assign n848 = ~n747 & n847 ;
  assign n853 = n852 ^ n848 ^ 1'b0 ;
  assign n854 = n240 ^ n205 ^ x91 ;
  assign n855 = x70 & x90 ;
  assign n856 = n220 & n235 ;
  assign n857 = ~n316 & n856 ;
  assign n858 = ~n297 & n857 ;
  assign n859 = n415 ^ n281 ^ 1'b0 ;
  assign n860 = n853 ^ n553 ^ 1'b0 ;
  assign n861 = n859 & ~n860 ;
  assign n864 = n139 | n175 ;
  assign n865 = n514 & ~n864 ;
  assign n862 = n709 ^ n438 ^ 1'b0 ;
  assign n863 = n862 ^ n491 ^ 1'b0 ;
  assign n866 = n865 ^ n863 ^ n439 ;
  assign n867 = ~n198 & n731 ;
  assign n868 = n481 ^ n144 ^ 1'b0 ;
  assign n869 = x65 & n753 ;
  assign n870 = n181 | n552 ;
  assign n871 = x41 & n158 ;
  assign n872 = n871 ^ x103 ^ 1'b0 ;
  assign n873 = n297 ^ x70 ^ 1'b0 ;
  assign n874 = x6 & n873 ;
  assign n875 = n872 | n874 ;
  assign n876 = n875 ^ x77 ^ 1'b0 ;
  assign n877 = n161 ^ x73 ^ 1'b0 ;
  assign n878 = x106 & n220 ;
  assign n879 = ~n425 & n878 ;
  assign n880 = n512 ^ n442 ^ 1'b0 ;
  assign n881 = n281 ^ n229 ^ 1'b0 ;
  assign n882 = x91 & n881 ;
  assign n883 = n455 ^ x118 ^ 1'b0 ;
  assign n884 = n882 & ~n883 ;
  assign n885 = n656 & n884 ;
  assign n886 = n211 & n363 ;
  assign n887 = n731 ^ n544 ^ 1'b0 ;
  assign n888 = ~n886 & n887 ;
  assign n889 = ~n507 & n645 ;
  assign n890 = n164 ^ x96 ^ 1'b0 ;
  assign n891 = n776 ^ n369 ^ 1'b0 ;
  assign n892 = ~x108 & n845 ;
  assign n893 = n227 & ~n744 ;
  assign n894 = x12 & ~n496 ;
  assign n895 = n473 & ~n555 ;
  assign n896 = ( n169 & n499 ) | ( n169 & ~n895 ) | ( n499 & ~n895 ) ;
  assign n897 = n248 ^ x110 ^ 1'b0 ;
  assign n898 = x97 & n593 ;
  assign n899 = x112 & n849 ;
  assign n900 = ~n432 & n899 ;
  assign n901 = n900 ^ n756 ^ 1'b0 ;
  assign n902 = n898 | n901 ;
  assign n903 = n230 & n849 ;
  assign n904 = ~n277 & n903 ;
  assign n905 = n904 ^ n230 ^ 1'b0 ;
  assign n907 = n314 & ~n461 ;
  assign n906 = x17 & ~n686 ;
  assign n908 = n907 ^ n906 ^ 1'b0 ;
  assign n909 = n667 ^ n153 ^ 1'b0 ;
  assign n910 = n684 | n909 ;
  assign n911 = x119 | n910 ;
  assign n912 = n823 ^ n418 ^ 1'b0 ;
  assign n913 = x25 & n420 ;
  assign n914 = ~n205 & n913 ;
  assign n915 = n914 ^ x39 ^ 1'b0 ;
  assign n916 = x73 & ~n915 ;
  assign n917 = x57 & n916 ;
  assign n918 = n917 ^ n480 ^ 1'b0 ;
  assign n919 = n508 | n781 ;
  assign n920 = n349 | n919 ;
  assign n921 = ~n918 & n920 ;
  assign n922 = n171 & n414 ;
  assign n923 = n489 ^ x11 ^ 1'b0 ;
  assign n924 = n922 | n923 ;
  assign n925 = n455 | n480 ;
  assign n926 = n623 | n925 ;
  assign n933 = x9 & ~n638 ;
  assign n934 = n412 & n933 ;
  assign n928 = x63 & n144 ;
  assign n929 = x113 & n415 ;
  assign n930 = ~n928 & n929 ;
  assign n931 = ~n708 & n930 ;
  assign n927 = ~n571 & n782 ;
  assign n932 = n931 ^ n927 ^ 1'b0 ;
  assign n935 = n934 ^ n932 ^ 1'b0 ;
  assign n936 = n926 & ~n935 ;
  assign n937 = x29 & ~x37 ;
  assign n938 = n937 ^ n911 ^ 1'b0 ;
  assign n939 = ~n225 & n243 ;
  assign n941 = n753 ^ n135 ^ 1'b0 ;
  assign n942 = x108 & ~n941 ;
  assign n943 = n942 ^ n252 ^ 1'b0 ;
  assign n944 = ~n428 & n943 ;
  assign n940 = ~n481 & n658 ;
  assign n945 = n944 ^ n940 ^ 1'b0 ;
  assign n946 = n731 & ~n800 ;
  assign n947 = x31 & x34 ;
  assign n948 = ~x21 & n947 ;
  assign n949 = n766 | n948 ;
  assign n950 = n846 ^ x47 ^ 1'b0 ;
  assign n951 = n325 & n522 ;
  assign n952 = ~n420 & n951 ;
  assign n953 = n296 | n886 ;
  assign n954 = n953 ^ n408 ^ 1'b0 ;
  assign n955 = n229 & ~n954 ;
  assign n956 = n955 ^ n806 ^ 1'b0 ;
  assign n957 = ~n499 & n823 ;
  assign n958 = n225 & n957 ;
  assign n959 = n153 & n642 ;
  assign n960 = n764 & n959 ;
  assign n961 = ~n143 & n954 ;
  assign n962 = n428 ^ n230 ^ 1'b0 ;
  assign n963 = n962 ^ n321 ^ 1'b0 ;
  assign n964 = n963 ^ n250 ^ 1'b0 ;
  assign n965 = ~n614 & n964 ;
  assign n966 = n143 & n965 ;
  assign n967 = ~n620 & n966 ;
  assign n968 = ~n430 & n876 ;
  assign n969 = n967 & n968 ;
  assign n970 = ~n141 & n795 ;
  assign n971 = n970 ^ n141 ^ 1'b0 ;
  assign n972 = n195 & n376 ;
  assign n973 = ~n971 & n972 ;
  assign n974 = n713 & ~n973 ;
  assign n975 = x102 & ~n485 ;
  assign n976 = x18 & ~n459 ;
  assign n977 = n976 ^ n444 ^ 1'b0 ;
  assign n978 = n254 | n977 ;
  assign n979 = x114 & ~n276 ;
  assign n980 = ~x96 & n979 ;
  assign n981 = ~n302 & n980 ;
  assign n982 = x106 ^ x18 ^ 1'b0 ;
  assign n983 = n369 | n982 ;
  assign n984 = n938 ^ n584 ^ 1'b0 ;
  assign n985 = n245 | n983 ;
  assign n986 = ( n480 & n640 ) | ( n480 & ~n828 ) | ( n640 & ~n828 ) ;
  assign n987 = ~n146 & n381 ;
  assign n988 = ~x70 & n987 ;
  assign n989 = x105 & n222 ;
  assign n990 = n365 & n862 ;
  assign n991 = n990 ^ x32 ^ 1'b0 ;
  assign n993 = n250 | n380 ;
  assign n994 = x81 | n993 ;
  assign n992 = x97 ^ x33 ^ 1'b0 ;
  assign n995 = n994 ^ n992 ^ n360 ;
  assign n996 = n547 ^ n442 ^ 1'b0 ;
  assign n997 = n996 ^ n672 ^ 1'b0 ;
  assign n998 = x74 & ~n997 ;
  assign n999 = n509 ^ x119 ^ 1'b0 ;
  assign n1000 = x92 ^ x70 ^ 1'b0 ;
  assign n1001 = x14 & n1000 ;
  assign n1002 = n438 & ~n695 ;
  assign n1003 = n1001 & ~n1002 ;
  assign n1004 = n999 & n1003 ;
  assign n1005 = x72 | n514 ;
  assign n1006 = x102 & ~n1005 ;
  assign n1007 = n735 | n1006 ;
  assign n1008 = n1007 ^ n681 ^ 1'b0 ;
  assign n1009 = n467 & n553 ;
  assign n1010 = n1009 ^ n210 ^ 1'b0 ;
  assign n1011 = n463 & n570 ;
  assign n1012 = ~n1010 & n1011 ;
  assign n1013 = n630 ^ n238 ^ 1'b0 ;
  assign n1014 = x90 & n325 ;
  assign n1015 = ~n542 & n1014 ;
  assign n1016 = n502 ^ n137 ^ 1'b0 ;
  assign n1017 = n1016 ^ x81 ^ 1'b0 ;
  assign n1018 = n1015 | n1017 ;
  assign n1019 = ~n367 & n448 ;
  assign n1020 = n1019 ^ n210 ^ 1'b0 ;
  assign n1021 = n1020 ^ x16 ^ 1'b0 ;
  assign n1022 = n504 & ~n1021 ;
  assign n1023 = x70 & ~x78 ;
  assign n1024 = n1022 & ~n1023 ;
  assign n1025 = n591 & n1024 ;
  assign n1026 = x26 & ~n642 ;
  assign n1030 = x89 & ~x124 ;
  assign n1027 = ~n482 & n620 ;
  assign n1028 = n1027 ^ n290 ^ 1'b0 ;
  assign n1029 = n754 | n1028 ;
  assign n1031 = n1030 ^ n1029 ^ 1'b0 ;
  assign n1032 = ~n793 & n932 ;
  assign n1033 = n579 & n1032 ;
  assign n1034 = n642 ^ n215 ^ 1'b0 ;
  assign n1035 = x38 | n287 ;
  assign n1036 = n171 ^ x89 ^ 1'b0 ;
  assign n1037 = n1035 & ~n1036 ;
  assign n1038 = ( ~x14 & x78 ) | ( ~x14 & n173 ) | ( x78 & n173 ) ;
  assign n1039 = n1038 ^ n986 ^ 1'b0 ;
  assign n1040 = n1037 & ~n1039 ;
  assign n1041 = n1034 | n1040 ;
  assign n1042 = n189 | n281 ;
  assign n1043 = x125 & n1042 ;
  assign n1044 = n1043 ^ n413 ^ 1'b0 ;
  assign n1045 = n524 ^ n397 ^ 1'b0 ;
  assign n1046 = n1044 & ~n1045 ;
  assign n1047 = n141 & ~n600 ;
  assign n1048 = n1047 ^ x86 ^ 1'b0 ;
  assign n1049 = ~n590 & n1048 ;
  assign n1050 = n1046 & ~n1049 ;
  assign n1051 = n1050 ^ x15 ^ 1'b0 ;
  assign n1052 = ~n529 & n1051 ;
  assign n1054 = ~n404 & n1020 ;
  assign n1055 = n992 | n1054 ;
  assign n1053 = ~n360 & n506 ;
  assign n1056 = n1055 ^ n1053 ^ x32 ;
  assign n1057 = x84 | n380 ;
  assign n1058 = n1057 ^ n595 ^ 1'b0 ;
  assign n1059 = x109 & n1058 ;
  assign n1060 = ~n1010 & n1059 ;
  assign n1061 = n328 | n1060 ;
  assign n1062 = n179 & n1061 ;
  assign n1063 = n1062 ^ n1030 ^ 1'b0 ;
  assign n1064 = n406 ^ n324 ^ 1'b0 ;
  assign n1065 = n1064 ^ n272 ^ 1'b0 ;
  assign n1066 = n190 & ~n1065 ;
  assign n1067 = ~n955 & n1066 ;
  assign n1068 = n394 & ~n630 ;
  assign n1069 = n428 & n1068 ;
  assign n1070 = n509 ^ n487 ^ 1'b0 ;
  assign n1071 = ( n183 & n1069 ) | ( n183 & ~n1070 ) | ( n1069 & ~n1070 ) ;
  assign n1072 = n1071 ^ n478 ^ 1'b0 ;
  assign n1073 = ~n225 & n784 ;
  assign n1074 = n531 & ~n799 ;
  assign n1075 = n1074 ^ n219 ^ 1'b0 ;
  assign n1076 = n1075 ^ n788 ^ 1'b0 ;
  assign n1077 = ( n813 & n1073 ) | ( n813 & ~n1076 ) | ( n1073 & ~n1076 ) ;
  assign n1078 = n276 | n568 ;
  assign n1079 = n1078 ^ n727 ^ 1'b0 ;
  assign n1080 = n333 ^ x107 ^ 1'b0 ;
  assign n1081 = n281 & n1080 ;
  assign n1082 = n1081 ^ n459 ^ 1'b0 ;
  assign n1083 = ~n749 & n870 ;
  assign n1084 = n1083 ^ n243 ^ 1'b0 ;
  assign n1085 = n163 & n562 ;
  assign n1086 = n1085 ^ x68 ^ 1'b0 ;
  assign n1087 = n203 | n1086 ;
  assign n1088 = x94 & n451 ;
  assign n1089 = n1088 ^ x103 ^ 1'b0 ;
  assign n1090 = n640 | n1089 ;
  assign n1091 = n1090 ^ n258 ^ 1'b0 ;
  assign n1092 = n656 | n1091 ;
  assign n1093 = ~x124 & n504 ;
  assign n1097 = x8 & ~n132 ;
  assign n1098 = n1097 ^ x3 ^ 1'b0 ;
  assign n1094 = n571 | n889 ;
  assign n1095 = n1094 ^ x82 ^ 1'b0 ;
  assign n1096 = n188 & n1095 ;
  assign n1099 = n1098 ^ n1096 ^ 1'b0 ;
  assign n1100 = n1099 ^ n555 ^ 1'b0 ;
  assign n1101 = n948 | n1100 ;
  assign n1102 = n273 & ~n391 ;
  assign n1103 = n477 & ~n837 ;
  assign n1104 = n891 & ~n1002 ;
  assign n1105 = n1010 & n1104 ;
  assign n1106 = n952 | n1061 ;
  assign n1107 = n1031 ^ x98 ^ 1'b0 ;
  assign n1108 = n358 | n708 ;
  assign n1109 = n1108 ^ n629 ^ 1'b0 ;
  assign n1110 = n847 ^ n499 ^ 1'b0 ;
  assign n1111 = ~n899 & n1110 ;
  assign n1112 = ~n410 & n1111 ;
  assign n1113 = x74 & ~n1112 ;
  assign n1114 = ~n1109 & n1113 ;
  assign n1115 = ~x4 & x63 ;
  assign n1116 = n1114 | n1115 ;
  assign n1117 = n229 & n438 ;
  assign n1118 = n1117 ^ n844 ^ 1'b0 ;
  assign n1119 = n400 ^ n208 ^ 1'b0 ;
  assign n1120 = x84 & ~n1119 ;
  assign n1121 = n1120 ^ n246 ^ 1'b0 ;
  assign n1122 = ~n1067 & n1121 ;
  assign n1123 = n862 ^ n444 ^ 1'b0 ;
  assign n1124 = ~n759 & n1123 ;
  assign n1125 = ~n958 & n970 ;
  assign n1126 = ~x0 & n1125 ;
  assign n1127 = x10 & n806 ;
  assign n1128 = n717 & n1127 ;
  assign n1129 = n1030 | n1128 ;
  assign n1130 = n165 | n638 ;
  assign n1131 = n1130 ^ n645 ^ n328 ;
  assign n1132 = n485 & ~n506 ;
  assign n1133 = n1131 & ~n1132 ;
  assign n1134 = x0 & ~n358 ;
  assign n1135 = ~x41 & n1134 ;
  assign n1136 = n733 | n1135 ;
  assign n1137 = n766 | n1136 ;
  assign n1138 = n591 ^ n344 ^ 1'b0 ;
  assign n1139 = ~n396 & n1138 ;
  assign n1140 = ~n494 & n845 ;
  assign n1141 = n1140 ^ x16 ^ 1'b0 ;
  assign n1142 = n402 & n764 ;
  assign n1143 = ~n499 & n1142 ;
  assign n1144 = ~n849 & n1143 ;
  assign n1145 = n972 ^ n831 ^ 1'b0 ;
  assign n1146 = ~n538 & n1145 ;
  assign n1147 = n453 | n1146 ;
  assign n1148 = x89 & ~n638 ;
  assign n1149 = ~n229 & n1148 ;
  assign n1150 = n375 & ~n1149 ;
  assign n1151 = ~n884 & n1150 ;
  assign n1152 = n1147 | n1151 ;
  assign n1153 = n701 | n1152 ;
  assign n1154 = n570 & n1153 ;
  assign n1155 = n1154 ^ n1070 ^ 1'b0 ;
  assign n1156 = n652 & ~n1155 ;
  assign n1157 = ( n150 & n246 ) | ( n150 & n625 ) | ( n246 & n625 ) ;
  assign n1158 = n904 | n1157 ;
  assign n1159 = x37 ^ x11 ^ 1'b0 ;
  assign n1160 = n696 & n1159 ;
  assign n1161 = x91 | n375 ;
  assign n1162 = ~n1042 & n1161 ;
  assign n1163 = n1015 ^ n814 ^ 1'b0 ;
  assign n1164 = n825 ^ n150 ^ 1'b0 ;
  assign n1165 = ~n288 & n1164 ;
  assign n1167 = n195 | n215 ;
  assign n1166 = n354 ^ n344 ^ 1'b0 ;
  assign n1168 = n1167 ^ n1166 ^ 1'b0 ;
  assign n1169 = ~n367 & n1168 ;
  assign n1170 = n400 ^ n245 ^ 1'b0 ;
  assign n1171 = n1170 ^ n482 ^ x54 ;
  assign n1172 = n1052 | n1171 ;
  assign n1173 = n1144 ^ n555 ^ 1'b0 ;
  assign n1175 = x68 & ~n134 ;
  assign n1176 = n1175 ^ x26 ^ 1'b0 ;
  assign n1174 = n753 & n1075 ;
  assign n1177 = n1176 ^ n1174 ^ 1'b0 ;
  assign n1178 = n198 & n1177 ;
  assign n1179 = n246 & ~n302 ;
  assign n1180 = ~n872 & n1179 ;
  assign n1181 = n1180 ^ x58 ^ 1'b0 ;
  assign n1182 = x113 & ~n1181 ;
  assign n1183 = ~x39 & n1182 ;
  assign n1184 = n135 & n326 ;
  assign n1185 = n444 & n1184 ;
  assign n1187 = n672 ^ n404 ^ n153 ;
  assign n1186 = n481 | n1115 ;
  assign n1188 = n1187 ^ n1186 ^ 1'b0 ;
  assign n1189 = n967 & ~n1186 ;
  assign n1190 = x114 ^ x82 ^ 1'b0 ;
  assign n1191 = x109 & n1190 ;
  assign n1192 = n1191 ^ n808 ^ 1'b0 ;
  assign n1193 = n742 ^ n487 ^ 1'b0 ;
  assign n1194 = n402 | n1193 ;
  assign n1195 = ( n134 & ~n363 ) | ( n134 & n519 ) | ( ~n363 & n519 ) ;
  assign n1196 = n477 & ~n1106 ;
  assign n1197 = n1196 ^ n991 ^ 1'b0 ;
  assign n1198 = n292 | n1069 ;
  assign n1199 = n1198 ^ n1077 ^ 1'b0 ;
  assign n1200 = n487 | n761 ;
  assign n1201 = n1200 ^ n804 ^ 1'b0 ;
  assign n1202 = n694 ^ n289 ^ 1'b0 ;
  assign n1203 = ~n991 & n1059 ;
  assign n1204 = n795 ^ n574 ^ 1'b0 ;
  assign n1205 = ( n663 & n1109 ) | ( n663 & n1204 ) | ( n1109 & n1204 ) ;
  assign n1206 = x73 | n297 ;
  assign n1207 = x47 & n1206 ;
  assign n1208 = x49 & ~n502 ;
  assign n1209 = n378 ^ x109 ^ x65 ;
  assign n1210 = n1209 ^ n728 ^ 1'b0 ;
  assign n1211 = ~n506 & n1210 ;
  assign n1212 = n442 & n504 ;
  assign n1213 = n770 | n1212 ;
  assign n1214 = n1213 ^ n1156 ^ 1'b0 ;
  assign n1215 = n213 ^ x119 ^ 1'b0 ;
  assign n1216 = n1214 & n1215 ;
  assign n1217 = x119 & ~n394 ;
  assign n1218 = x3 & n1217 ;
  assign n1219 = ~n1216 & n1218 ;
  assign n1220 = n741 ^ x98 ^ 1'b0 ;
  assign n1221 = n834 | n1220 ;
  assign n1222 = n1030 ^ x64 ^ 1'b0 ;
  assign n1223 = n399 | n1222 ;
  assign n1224 = n1223 ^ n747 ^ 1'b0 ;
  assign n1225 = n246 & n753 ;
  assign n1226 = n1224 & n1225 ;
  assign n1227 = n407 ^ n318 ^ 1'b0 ;
  assign n1228 = n420 & n1227 ;
  assign n1229 = n1228 ^ n576 ^ n131 ;
  assign n1230 = ( n399 & n1064 ) | ( n399 & n1179 ) | ( n1064 & n1179 ) ;
  assign n1231 = ~n491 & n618 ;
  assign n1232 = ~n1230 & n1231 ;
  assign n1233 = n399 | n995 ;
  assign n1234 = n1232 & ~n1233 ;
  assign n1235 = n378 & n652 ;
  assign n1236 = n766 & n1031 ;
  assign n1237 = n900 ^ x49 ^ 1'b0 ;
  assign n1238 = n480 | n1237 ;
  assign n1239 = n1238 ^ n418 ^ 1'b0 ;
  assign n1240 = n689 & ~n1239 ;
  assign n1241 = n1240 ^ x90 ^ 1'b0 ;
  assign n1242 = x71 & n938 ;
  assign n1243 = ~n1070 & n1242 ;
  assign n1244 = ( n279 & n373 ) | ( n279 & n643 ) | ( n373 & n643 ) ;
  assign n1245 = n531 ^ n259 ^ 1'b0 ;
  assign n1246 = n1245 ^ n722 ^ 1'b0 ;
  assign n1247 = n289 & n1246 ;
  assign n1248 = n1247 ^ n720 ^ 1'b0 ;
  assign n1249 = n1244 | n1248 ;
  assign n1250 = n669 ^ n497 ^ 1'b0 ;
  assign n1251 = ~n680 & n1250 ;
  assign n1252 = n1251 ^ n300 ^ 1'b0 ;
  assign n1253 = n1030 | n1252 ;
  assign n1254 = n413 ^ x47 ^ 1'b0 ;
  assign n1255 = x15 & n413 ;
  assign n1256 = n1255 ^ n1204 ^ 1'b0 ;
  assign n1257 = n862 ^ n540 ^ 1'b0 ;
  assign n1258 = n1256 | n1257 ;
  assign n1263 = x83 & n332 ;
  assign n1264 = ~n246 & n1263 ;
  assign n1259 = x90 & ~n669 ;
  assign n1260 = n1259 ^ n210 ^ 1'b0 ;
  assign n1261 = n731 ^ x42 ^ 1'b0 ;
  assign n1262 = ~n1260 & n1261 ;
  assign n1265 = n1264 ^ n1262 ^ 1'b0 ;
  assign n1266 = x46 & ~n506 ;
  assign n1267 = n468 & n1266 ;
  assign n1268 = x36 | n1267 ;
  assign n1269 = n845 & ~n1268 ;
  assign n1270 = n616 & n1269 ;
  assign n1271 = x76 & ~x106 ;
  assign n1272 = ~n195 & n1271 ;
  assign n1273 = x27 | n1272 ;
  assign n1274 = n383 | n841 ;
  assign n1275 = n444 | n487 ;
  assign n1276 = ~n1030 & n1275 ;
  assign n1277 = ~n665 & n1276 ;
  assign n1278 = n978 ^ x39 ^ 1'b0 ;
  assign n1279 = n380 | n1278 ;
  assign n1280 = n1016 ^ n800 ^ n360 ;
  assign n1281 = n283 & n576 ;
  assign n1282 = n579 | n851 ;
  assign n1283 = n277 | n1282 ;
  assign n1284 = x99 & n320 ;
  assign n1285 = ~n614 & n1284 ;
  assign n1286 = n1169 & n1285 ;
  assign n1287 = ~n1283 & n1286 ;
  assign n1288 = ~n695 & n1251 ;
  assign n1289 = n1070 & n1288 ;
  assign n1290 = n1289 ^ x70 ^ 1'b0 ;
  assign n1291 = n754 & ~n886 ;
  assign n1292 = n907 | n1291 ;
  assign n1293 = n338 ^ n307 ^ 1'b0 ;
  assign n1294 = n410 & ~n1293 ;
  assign n1295 = n650 & n1294 ;
  assign n1296 = n153 | n1270 ;
  assign n1297 = n567 & ~n1296 ;
  assign n1298 = n1297 ^ n1057 ^ 1'b0 ;
  assign n1299 = x92 & n198 ;
  assign n1300 = n956 | n1144 ;
  assign n1301 = n1300 ^ n433 ^ 1'b0 ;
  assign n1302 = n552 ^ x48 ^ 1'b0 ;
  assign n1303 = n540 & ~n1102 ;
  assign n1304 = n371 ^ x54 ^ 1'b0 ;
  assign n1305 = n1055 ^ n427 ^ 1'b0 ;
  assign n1306 = ~n566 & n1305 ;
  assign n1307 = n1306 ^ n152 ^ 1'b0 ;
  assign n1308 = n1304 & n1307 ;
  assign n1309 = n153 | n328 ;
  assign n1310 = n1309 ^ n396 ^ 1'b0 ;
  assign n1311 = n262 | n1310 ;
  assign n1312 = n516 | n1311 ;
  assign n1313 = ~n251 & n1312 ;
  assign n1314 = n153 & n1313 ;
  assign n1315 = n1245 ^ n731 ^ 1'b0 ;
  assign n1316 = n926 ^ n570 ^ n381 ;
  assign n1317 = n1316 ^ x50 ^ 1'b0 ;
  assign n1318 = x71 & n450 ;
  assign n1319 = ~n1317 & n1318 ;
  assign n1320 = x21 & n701 ;
  assign n1321 = n1320 ^ n439 ^ 1'b0 ;
  assign n1322 = ~n356 & n1321 ;
  assign n1323 = n1322 ^ x127 ^ 1'b0 ;
  assign n1324 = n1173 ^ n1167 ^ x80 ;
  assign n1325 = n625 ^ n217 ^ 1'b0 ;
  assign n1326 = x83 ^ x74 ^ 1'b0 ;
  assign n1327 = ~n660 & n1326 ;
  assign n1328 = n921 | n1062 ;
  assign n1330 = x122 & ~n207 ;
  assign n1331 = n1330 ^ n369 ^ 1'b0 ;
  assign n1329 = n709 ^ n156 ^ 1'b0 ;
  assign n1332 = n1331 ^ n1329 ^ 1'b0 ;
  assign n1333 = ~n1328 & n1332 ;
  assign n1334 = n1327 & n1333 ;
  assign n1335 = n680 | n766 ;
  assign n1336 = n595 & ~n1335 ;
  assign n1337 = n763 & ~n1062 ;
  assign n1338 = ~n1064 & n1337 ;
  assign n1339 = n1336 | n1338 ;
  assign n1340 = n245 & ~n1339 ;
  assign n1342 = x123 & ~n259 ;
  assign n1343 = n687 & n1342 ;
  assign n1344 = n934 & n1343 ;
  assign n1341 = n544 ^ x121 ^ 1'b0 ;
  assign n1345 = n1344 ^ n1341 ^ 1'b0 ;
  assign n1346 = n299 & ~n1345 ;
  assign n1347 = n428 | n1346 ;
  assign n1348 = n487 & ~n1347 ;
  assign n1349 = n259 & ~n272 ;
  assign n1350 = n1035 ^ n909 ^ 1'b0 ;
  assign n1351 = n704 | n1350 ;
  assign n1352 = n684 ^ n363 ^ 1'b0 ;
  assign n1353 = n805 ^ n701 ^ 1'b0 ;
  assign n1354 = n349 & ~n1353 ;
  assign n1355 = n1354 ^ n493 ^ 1'b0 ;
  assign n1356 = n344 & ~n1018 ;
  assign n1357 = n250 ^ x127 ^ 1'b0 ;
  assign n1358 = n288 | n1357 ;
  assign n1359 = n1243 | n1358 ;
  assign n1360 = n1359 ^ n164 ^ 1'b0 ;
  assign n1361 = n296 | n1001 ;
  assign n1362 = x106 & ~n1361 ;
  assign n1363 = ~n775 & n1362 ;
  assign n1364 = n1063 & n1316 ;
  assign n1365 = n221 & ~n1310 ;
  assign n1366 = n1365 ^ n792 ^ 1'b0 ;
  assign n1367 = n1206 & n1366 ;
  assign n1368 = ~n711 & n1367 ;
  assign n1369 = ~n283 & n387 ;
  assign n1370 = x116 & ~n338 ;
  assign n1371 = ~x52 & n1370 ;
  assign n1372 = n1040 & n1371 ;
  assign n1373 = ~n1201 & n1372 ;
  assign n1374 = n491 & n1373 ;
  assign n1375 = x106 ^ x52 ^ 1'b0 ;
  assign n1376 = n741 | n1375 ;
  assign n1377 = x14 & ~n1060 ;
  assign n1378 = n1377 ^ n892 ^ 1'b0 ;
  assign n1379 = n1004 ^ n992 ^ 1'b0 ;
  assign n1380 = n1378 & n1379 ;
  assign n1381 = ~n380 & n594 ;
  assign n1382 = x37 & ~n189 ;
  assign n1383 = n1382 ^ n450 ^ 1'b0 ;
  assign n1384 = n775 & ~n1383 ;
  assign n1385 = n1384 ^ n194 ^ 1'b0 ;
  assign n1386 = n1385 ^ n694 ^ 1'b0 ;
  assign n1387 = n835 & ~n1386 ;
  assign n1388 = n188 & n242 ;
  assign n1389 = n1388 ^ x69 ^ 1'b0 ;
  assign n1390 = n485 ^ x120 ^ 1'b0 ;
  assign n1391 = ~n1389 & n1390 ;
  assign n1392 = n1035 & n1391 ;
  assign n1393 = n315 & n1392 ;
  assign n1394 = n417 & ~n1393 ;
  assign n1395 = n828 ^ n571 ^ 1'b0 ;
  assign n1396 = n311 ^ n240 ^ 1'b0 ;
  assign n1397 = ~n198 & n1396 ;
  assign n1398 = ( n381 & n389 ) | ( n381 & ~n1397 ) | ( n389 & ~n1397 ) ;
  assign n1400 = n308 ^ n240 ^ 1'b0 ;
  assign n1401 = n1400 ^ n189 ^ 1'b0 ;
  assign n1399 = n583 & n857 ;
  assign n1402 = n1401 ^ n1399 ^ 1'b0 ;
  assign n1404 = n1042 ^ n190 ^ 1'b0 ;
  assign n1405 = n407 & n1404 ;
  assign n1406 = x55 & n857 ;
  assign n1407 = ~n1115 & n1406 ;
  assign n1408 = n1407 ^ n969 ^ 1'b0 ;
  assign n1409 = n1405 & ~n1408 ;
  assign n1403 = x114 & ~n238 ;
  assign n1410 = n1409 ^ n1403 ^ 1'b0 ;
  assign n1411 = n451 & ~n896 ;
  assign n1412 = ~n794 & n1411 ;
  assign n1413 = n442 | n1412 ;
  assign n1414 = x23 | n1413 ;
  assign n1415 = ~n481 & n1054 ;
  assign n1416 = ~n916 & n1405 ;
  assign n1417 = ~n828 & n1327 ;
  assign n1418 = ~n516 & n1417 ;
  assign n1419 = n252 | n1418 ;
  assign n1420 = x68 & ~n325 ;
  assign n1421 = n459 | n466 ;
  assign n1422 = x25 | n1421 ;
  assign n1423 = n402 & ~n1422 ;
  assign n1424 = n1423 ^ n1327 ^ 1'b0 ;
  assign n1425 = n1031 & ~n1424 ;
  assign n1426 = n539 | n684 ;
  assign n1427 = n408 | n1426 ;
  assign n1428 = n1427 ^ x91 ^ 1'b0 ;
  assign n1429 = n542 ^ x40 ^ 1'b0 ;
  assign n1430 = x118 & n1429 ;
  assign n1431 = n1430 ^ x88 ^ 1'b0 ;
  assign n1432 = x9 & n1431 ;
  assign n1433 = ~n318 & n1432 ;
  assign n1434 = n1433 ^ n1292 ^ 1'b0 ;
  assign n1435 = n272 | n892 ;
  assign n1436 = n1435 ^ n258 ^ 1'b0 ;
  assign n1437 = n978 ^ n231 ^ 1'b0 ;
  assign n1438 = n400 ^ n190 ^ 1'b0 ;
  assign n1439 = ~n776 & n1438 ;
  assign n1440 = n1439 ^ n390 ^ 1'b0 ;
  assign n1441 = x70 & ~n1440 ;
  assign n1442 = n884 ^ n647 ^ 1'b0 ;
  assign n1443 = ~n749 & n1442 ;
  assign n1444 = n1443 ^ n652 ^ 1'b0 ;
  assign n1445 = n1441 & n1444 ;
  assign n1446 = n1445 ^ x104 ^ 1'b0 ;
  assign n1447 = n487 ^ n230 ^ 1'b0 ;
  assign n1448 = n1447 ^ n258 ^ 1'b0 ;
  assign n1449 = x23 & ~n1448 ;
  assign n1450 = n163 & n1449 ;
  assign n1451 = n950 & n1450 ;
  assign n1452 = n1064 ^ x127 ^ 1'b0 ;
  assign n1453 = n1427 ^ n394 ^ 1'b0 ;
  assign n1454 = n1452 & n1453 ;
  assign n1455 = n1176 & n1454 ;
  assign n1456 = n876 & ~n1446 ;
  assign n1457 = n1291 ^ n698 ^ 1'b0 ;
  assign n1458 = n349 & n375 ;
  assign n1459 = n1458 ^ n1327 ^ 1'b0 ;
  assign n1460 = n932 & ~n1459 ;
  assign n1461 = ~x32 & n1460 ;
  assign n1462 = n237 ^ n173 ^ 1'b0 ;
  assign n1463 = ( n221 & n1051 ) | ( n221 & ~n1462 ) | ( n1051 & ~n1462 ) ;
  assign n1466 = n254 | n261 ;
  assign n1467 = n1466 ^ n321 ^ 1'b0 ;
  assign n1468 = ~x14 & n1467 ;
  assign n1464 = n457 | n461 ;
  assign n1465 = n634 & ~n1464 ;
  assign n1469 = n1468 ^ n1465 ^ 1'b0 ;
  assign n1470 = ~n369 & n852 ;
  assign n1471 = ( ~x53 & n135 ) | ( ~x53 & n724 ) | ( n135 & n724 ) ;
  assign n1472 = n342 & n1471 ;
  assign n1473 = ~n302 & n775 ;
  assign n1474 = ~n852 & n1473 ;
  assign n1475 = n667 & n862 ;
  assign n1476 = n1316 ^ x106 ^ 1'b0 ;
  assign n1477 = n806 | n1476 ;
  assign n1478 = n825 ^ n548 ^ x119 ;
  assign n1479 = n855 ^ n467 ^ 1'b0 ;
  assign n1480 = x77 & ~n1479 ;
  assign n1481 = n288 | n1023 ;
  assign n1482 = n1481 ^ n1243 ^ 1'b0 ;
  assign n1483 = n359 & n858 ;
  assign n1484 = n463 & ~n1483 ;
  assign n1485 = n669 | n793 ;
  assign n1486 = x16 & n173 ;
  assign n1487 = n373 & n1486 ;
  assign n1488 = n1098 ^ x89 ^ 1'b0 ;
  assign n1489 = x116 & ~n1488 ;
  assign n1490 = x21 ^ x5 ^ 1'b0 ;
  assign n1491 = n1489 & n1490 ;
  assign n1492 = ~n773 & n1491 ;
  assign n1493 = n1492 ^ n624 ^ 1'b0 ;
  assign n1494 = x12 | n526 ;
  assign n1495 = n1494 ^ x56 ^ 1'b0 ;
  assign n1496 = x47 | n1468 ;
  assign n1497 = n198 & ~n1258 ;
  assign n1498 = n1056 ^ n457 ^ 1'b0 ;
  assign n1499 = n463 ^ n346 ^ 1'b0 ;
  assign n1500 = x105 & ~n134 ;
  assign n1501 = n1500 ^ n159 ^ 1'b0 ;
  assign n1502 = n1501 ^ n192 ^ 1'b0 ;
  assign n1503 = n972 & ~n1016 ;
  assign n1504 = n1503 ^ n144 ^ 1'b0 ;
  assign n1505 = n387 & n613 ;
  assign n1506 = ~n727 & n1505 ;
  assign n1507 = x54 & x126 ;
  assign n1508 = n1507 ^ n1025 ^ 1'b0 ;
  assign n1509 = ~n1506 & n1508 ;
  assign n1510 = n1509 ^ n378 ^ 1'b0 ;
  assign n1511 = n1504 & n1510 ;
  assign n1512 = n1511 ^ n1202 ^ 1'b0 ;
  assign n1513 = n1512 ^ n1238 ^ 1'b0 ;
  assign n1514 = n568 | n614 ;
  assign n1515 = n1514 ^ n1291 ^ 1'b0 ;
  assign n1516 = ~n131 & n595 ;
  assign n1517 = ~n233 & n1516 ;
  assign n1518 = n1515 & ~n1517 ;
  assign n1519 = ~x104 & n1518 ;
  assign n1520 = n399 ^ n171 ^ 1'b0 ;
  assign n1521 = x81 & n1520 ;
  assign n1522 = ~n344 & n1521 ;
  assign n1523 = n978 & n1522 ;
  assign n1524 = n1519 | n1523 ;
  assign n1525 = n1524 ^ x47 ^ 1'b0 ;
  assign n1526 = n1054 ^ n636 ^ 1'b0 ;
  assign n1527 = n1177 ^ n418 ^ 1'b0 ;
  assign n1528 = n1527 ^ n441 ^ 1'b0 ;
  assign n1529 = x52 & n1528 ;
  assign n1530 = n724 & n1529 ;
  assign n1531 = ~n1526 & n1530 ;
  assign n1532 = ~n450 & n1531 ;
  assign n1533 = n707 & ~n1369 ;
  assign n1534 = n1061 & n1533 ;
  assign n1535 = ~n259 & n267 ;
  assign n1536 = ~n594 & n1535 ;
  assign n1537 = n1180 ^ n144 ^ 1'b0 ;
  assign n1538 = n690 ^ n576 ^ 1'b0 ;
  assign n1539 = ~n285 & n1538 ;
  assign n1540 = ~n733 & n1489 ;
  assign n1541 = ~x109 & x116 ;
  assign n1542 = n1541 ^ n1221 ^ 1'b0 ;
  assign n1543 = n820 ^ n484 ^ 1'b0 ;
  assign n1544 = n311 & ~n464 ;
  assign n1545 = n1258 & n1544 ;
  assign n1546 = n1201 | n1525 ;
  assign n1547 = n1546 ^ n797 ^ 1'b0 ;
  assign n1551 = n739 ^ n708 ^ 1'b0 ;
  assign n1548 = x94 & ~n1098 ;
  assign n1549 = n456 & n1548 ;
  assign n1550 = n1549 ^ x125 ^ 1'b0 ;
  assign n1552 = n1551 ^ n1550 ^ n183 ;
  assign n1553 = n1179 & n1552 ;
  assign n1554 = n675 & n1553 ;
  assign n1555 = n963 ^ n373 ^ 1'b0 ;
  assign n1556 = n235 & n1555 ;
  assign n1557 = x106 & ~n353 ;
  assign n1558 = n1557 ^ n724 ^ 1'b0 ;
  assign n1559 = n1558 ^ n1082 ^ 1'b0 ;
  assign n1560 = n1556 & ~n1559 ;
  assign n1561 = n1560 ^ n394 ^ 1'b0 ;
  assign n1562 = n747 | n1310 ;
  assign n1563 = n900 & ~n1562 ;
  assign n1564 = ~n1115 & n1563 ;
  assign n1565 = n564 ^ n237 ^ 1'b0 ;
  assign n1566 = n483 & n1565 ;
  assign n1567 = n836 | n1049 ;
  assign n1568 = n1567 ^ n381 ^ 1'b0 ;
  assign n1569 = n1568 ^ n292 ^ 1'b0 ;
  assign n1570 = n252 & ~n613 ;
  assign n1571 = n1570 ^ n1070 ^ 1'b0 ;
  assign n1572 = n1060 & ~n1571 ;
  assign n1573 = x100 & ~n346 ;
  assign n1574 = n1573 ^ n570 ^ 1'b0 ;
  assign n1575 = x94 & n586 ;
  assign n1576 = ~n1574 & n1575 ;
  assign n1577 = n1280 & ~n1576 ;
  assign n1578 = ~x6 & n1577 ;
  assign n1579 = n188 | n571 ;
  assign n1580 = ~n825 & n1579 ;
  assign n1581 = n794 & ~n899 ;
  assign n1582 = n155 | n1243 ;
  assign n1583 = n976 | n1582 ;
  assign n1584 = n1260 ^ n464 ^ 1'b0 ;
  assign n1585 = n430 | n1584 ;
  assign n1586 = n692 & ~n1585 ;
  assign n1587 = n916 & ~n1586 ;
  assign n1589 = ~n577 & n826 ;
  assign n1588 = n507 ^ n422 ^ x34 ;
  assign n1590 = n1589 ^ n1588 ^ 1'b0 ;
  assign n1591 = x11 & x117 ;
  assign n1592 = n164 & n1591 ;
  assign n1593 = n781 ^ n230 ^ n139 ;
  assign n1594 = n766 | n1593 ;
  assign n1595 = n1594 ^ n724 ^ 1'b0 ;
  assign n1596 = ( x119 & ~n409 ) | ( x119 & n1268 ) | ( ~n409 & n1268 ) ;
  assign n1597 = n801 & ~n1596 ;
  assign n1598 = n238 | n1597 ;
  assign n1599 = n595 | n1598 ;
  assign n1600 = x127 | n480 ;
  assign n1601 = n1599 | n1600 ;
  assign n1602 = n794 & ~n1601 ;
  assign n1605 = n918 ^ n753 ^ 1'b0 ;
  assign n1606 = ~n287 & n1605 ;
  assign n1603 = n717 | n1383 ;
  assign n1604 = n1406 & ~n1603 ;
  assign n1607 = n1606 ^ n1604 ^ 1'b0 ;
  assign n1608 = n1383 | n1607 ;
  assign n1609 = n797 ^ n315 ^ 1'b0 ;
  assign n1610 = n1609 ^ n1287 ^ x75 ;
  assign n1611 = n811 | n1102 ;
  assign n1612 = n1149 & ~n1611 ;
  assign n1613 = x31 | n904 ;
  assign n1614 = n812 & ~n1054 ;
  assign n1615 = n1609 & n1614 ;
  assign n1616 = n1615 ^ n1316 ^ 1'b0 ;
  assign n1617 = x68 ^ x32 ^ 1'b0 ;
  assign n1618 = n725 & n1617 ;
  assign n1619 = ~n785 & n1618 ;
  assign n1620 = n1619 ^ n1541 ^ 1'b0 ;
  assign n1621 = x9 & n1620 ;
  assign n1622 = n1572 & n1621 ;
  assign n1623 = ~n177 & n397 ;
  assign n1624 = x19 & ~n1623 ;
  assign n1625 = n695 | n1245 ;
  assign n1626 = n1625 ^ n703 ^ 1'b0 ;
  assign n1627 = n958 & ~n1163 ;
  assign n1630 = n722 & ~n796 ;
  assign n1631 = n744 & ~n1630 ;
  assign n1628 = x84 & n572 ;
  assign n1629 = n1628 ^ n1235 ^ 1'b0 ;
  assign n1632 = n1631 ^ n1629 ^ n994 ;
  assign n1633 = n499 | n713 ;
  assign n1634 = n1633 ^ n604 ^ 1'b0 ;
  assign n1635 = ~n886 & n1634 ;
  assign n1636 = n1635 ^ n632 ^ 1'b0 ;
  assign n1637 = ~n836 & n1287 ;
  assign n1638 = n250 ^ x5 ^ 1'b0 ;
  assign n1639 = n1637 & ~n1638 ;
  assign n1640 = n989 | n1395 ;
  assign n1641 = x86 & ~n391 ;
  assign n1642 = n1641 ^ n1380 ^ 1'b0 ;
  assign n1643 = n1640 | n1642 ;
  assign n1644 = n1643 ^ x49 ^ 1'b0 ;
  assign n1645 = n1149 ^ n399 ^ 1'b0 ;
  assign n1646 = n669 ^ n227 ^ 1'b0 ;
  assign n1647 = n484 | n1646 ;
  assign n1648 = n1647 ^ n1558 ^ 1'b0 ;
  assign n1649 = n1114 ^ n584 ^ 1'b0 ;
  assign n1650 = ~n1457 & n1649 ;
  assign n1651 = x17 | n1126 ;
  assign n1652 = n1587 & n1646 ;
  assign n1654 = n841 ^ n451 ^ 1'b0 ;
  assign n1653 = n642 ^ x5 ^ 1'b0 ;
  assign n1655 = n1654 ^ n1653 ^ 1'b0 ;
  assign n1656 = n1655 ^ n1449 ^ 1'b0 ;
  assign n1657 = n795 ^ n538 ^ 1'b0 ;
  assign n1658 = n509 & n1657 ;
  assign n1659 = x102 & n1658 ;
  assign n1660 = ~n373 & n1659 ;
  assign n1661 = ~n826 & n1660 ;
  assign n1662 = ( n544 & n1656 ) | ( n544 & ~n1661 ) | ( n1656 & ~n1661 ) ;
  assign n1663 = n1055 ^ n912 ^ n663 ;
  assign n1664 = ~n851 & n1663 ;
  assign n1665 = x34 & ~n820 ;
  assign n1666 = n826 & ~n1665 ;
  assign n1667 = n1666 ^ n1556 ^ 1'b0 ;
  assign n1668 = n444 & ~n660 ;
  assign n1669 = n177 & ~n1525 ;
  assign n1670 = ~n614 & n1441 ;
  assign n1671 = n1670 ^ n667 ^ 1'b0 ;
  assign n1672 = n1671 ^ n1629 ^ 1'b0 ;
  assign n1673 = n607 & ~n1672 ;
  assign n1674 = n904 ^ n800 ^ 1'b0 ;
  assign n1675 = n568 & n1540 ;
  assign n1676 = ~n718 & n1366 ;
  assign n1677 = n1107 & n1676 ;
  assign n1678 = n288 ^ x19 ^ 1'b0 ;
  assign n1679 = n240 | n1678 ;
  assign n1680 = ~n320 & n1679 ;
  assign n1681 = ~n336 & n796 ;
  assign n1682 = n901 ^ x89 ^ 1'b0 ;
  assign n1683 = x71 & ~n1682 ;
  assign n1684 = n715 & n1683 ;
  assign n1685 = n1684 ^ n778 ^ 1'b0 ;
  assign n1686 = n916 & n1130 ;
  assign n1687 = n158 & n1686 ;
  assign n1688 = ~n775 & n1687 ;
  assign n1689 = n445 | n606 ;
  assign n1690 = n1689 ^ n1012 ^ 1'b0 ;
  assign n1691 = n1037 & ~n1690 ;
  assign n1692 = ~n1191 & n1691 ;
  assign n1693 = ~n781 & n1031 ;
  assign n1694 = x37 | n614 ;
  assign n1695 = n1110 & ~n1694 ;
  assign n1696 = n604 ^ x18 ^ 1'b0 ;
  assign n1697 = x110 & n1696 ;
  assign n1698 = n1697 ^ n224 ^ 1'b0 ;
  assign n1699 = ~n980 & n1698 ;
  assign n1700 = n134 | n1699 ;
  assign n1701 = n399 | n744 ;
  assign n1702 = n1700 | n1701 ;
  assign n1703 = ~n1695 & n1702 ;
  assign n1704 = ~n571 & n854 ;
  assign n1705 = n1033 ^ x23 ^ 1'b0 ;
  assign n1706 = n524 & ~n1705 ;
  assign n1707 = n1706 ^ n152 ^ 1'b0 ;
  assign n1708 = ~n510 & n937 ;
  assign n1709 = n1708 ^ n1352 ^ 1'b0 ;
  assign n1710 = n1059 & n1709 ;
  assign n1711 = ~n300 & n545 ;
  assign n1712 = n1711 ^ n1517 ^ 1'b0 ;
  assign n1713 = n266 & ~n1712 ;
  assign n1714 = n715 & n1106 ;
  assign n1715 = n1714 ^ n775 ^ 1'b0 ;
  assign n1716 = n1333 & ~n1715 ;
  assign n1717 = n1323 ^ n962 ^ 1'b0 ;
  assign n1718 = ~x106 & n1717 ;
  assign n1719 = n1188 & n1718 ;
  assign n1720 = n1719 ^ n355 ^ 1'b0 ;
  assign n1721 = n190 & n1652 ;
  assign n1722 = n1389 & n1721 ;
  assign n1723 = x14 & n276 ;
  assign n1724 = n1321 & ~n1723 ;
  assign n1725 = n1401 ^ n245 ^ 1'b0 ;
  assign n1726 = x123 & n1725 ;
  assign n1727 = n1726 ^ n1272 ^ 1'b0 ;
  assign n1728 = n721 | n1727 ;
  assign n1729 = n801 ^ n487 ^ 1'b0 ;
  assign n1730 = n731 | n1729 ;
  assign n1731 = n1730 ^ n1485 ^ 1'b0 ;
  assign n1732 = n213 & n956 ;
  assign n1734 = n1406 ^ n1002 ^ 1'b0 ;
  assign n1733 = n349 & ~n1247 ;
  assign n1735 = n1734 ^ n1733 ^ 1'b0 ;
  assign n1736 = n1732 & ~n1735 ;
  assign n1737 = n1011 & n1146 ;
  assign n1738 = n1737 ^ n866 ^ x106 ;
  assign n1746 = ~n689 & n729 ;
  assign n1740 = x4 & ~n568 ;
  assign n1741 = ~x39 & n1740 ;
  assign n1742 = n1741 ^ n394 ^ 1'b0 ;
  assign n1743 = n1646 | n1742 ;
  assign n1739 = n325 & ~n749 ;
  assign n1744 = n1743 ^ n1739 ^ 1'b0 ;
  assign n1745 = ~n1049 & n1744 ;
  assign n1747 = n1746 ^ n1745 ^ 1'b0 ;
  assign n1748 = n1268 ^ n1059 ^ n788 ;
  assign n1749 = x11 | n593 ;
  assign n1750 = n305 & n1749 ;
  assign n1751 = n1748 & n1750 ;
  assign n1752 = n535 & ~n1751 ;
  assign n1753 = n1752 ^ n832 ^ 1'b0 ;
  assign n1754 = ( n238 & ~n1325 ) | ( n238 & n1364 ) | ( ~n1325 & n1364 ) ;
  assign n1755 = n1754 ^ n131 ^ 1'b0 ;
  assign n1756 = ~n1185 & n1470 ;
  assign n1757 = n1517 ^ n1187 ^ 1'b0 ;
  assign n1758 = ~n406 & n1757 ;
  assign n1759 = n1758 ^ n1016 ^ n351 ;
  assign n1760 = n1759 ^ n1031 ^ n879 ;
  assign n1761 = n972 & ~n1760 ;
  assign n1762 = n1054 ^ n192 ^ 1'b0 ;
  assign n1763 = n360 | n445 ;
  assign n1764 = n1762 & ~n1763 ;
  assign n1765 = x109 & ~n146 ;
  assign n1766 = n1765 ^ n1264 ^ 1'b0 ;
  assign n1769 = x0 & n1131 ;
  assign n1767 = x24 & ~n574 ;
  assign n1768 = ~n283 & n1767 ;
  assign n1770 = n1769 ^ n1768 ^ 1'b0 ;
  assign n1771 = n1030 ^ n731 ^ 1'b0 ;
  assign n1772 = n705 & n1771 ;
  assign n1773 = n1772 ^ n1561 ^ 1'b0 ;
  assign n1774 = n717 ^ n297 ^ 1'b0 ;
  assign n1775 = n1342 ^ n1016 ^ 1'b0 ;
  assign n1776 = n1601 & ~n1775 ;
  assign n1777 = n459 | n1776 ;
  assign n1778 = x111 & n1087 ;
  assign n1779 = n302 & n1778 ;
  assign n1780 = ~n904 & n1180 ;
  assign n1781 = n1780 ^ n1240 ^ 1'b0 ;
  assign n1782 = n1221 ^ n1038 ^ 1'b0 ;
  assign n1783 = n1209 ^ n394 ^ 1'b0 ;
  assign n1784 = n616 & n1783 ;
  assign n1786 = n655 & ~n1508 ;
  assign n1787 = n701 & ~n1786 ;
  assign n1788 = n1787 ^ n885 ^ 1'b0 ;
  assign n1785 = x11 & ~n988 ;
  assign n1789 = n1788 ^ n1785 ^ 1'b0 ;
  assign n1790 = n1230 | n1287 ;
  assign n1791 = ~n1115 & n1422 ;
  assign n1792 = n1791 ^ n473 ^ 1'b0 ;
  assign n1793 = n1792 ^ x12 ^ 1'b0 ;
  assign n1794 = n983 | n1793 ;
  assign n1795 = n1794 ^ x61 ^ 1'b0 ;
  assign n1796 = x33 & n889 ;
  assign n1797 = n571 ^ n444 ^ 1'b0 ;
  assign n1798 = n562 & n1797 ;
  assign n1799 = ~n616 & n1798 ;
  assign n1800 = n1799 ^ n448 ^ 1'b0 ;
  assign n1801 = n1796 | n1800 ;
  assign n1802 = n1801 ^ n195 ^ 1'b0 ;
  assign n1803 = ~n450 & n1802 ;
  assign n1804 = n1795 & ~n1803 ;
  assign n1805 = n196 & n1804 ;
  assign n1806 = n533 | n1112 ;
  assign n1807 = n1265 & n1806 ;
  assign n1808 = n129 & ~n344 ;
  assign n1809 = n422 & ~n781 ;
  assign n1810 = ~n325 & n1809 ;
  assign n1811 = n1810 ^ n572 ^ 1'b0 ;
  assign n1812 = n1749 ^ n1634 ^ 1'b0 ;
  assign n1813 = n326 & ~n1812 ;
  assign n1814 = n1813 ^ n822 ^ 1'b0 ;
  assign n1815 = n270 & n531 ;
  assign n1816 = n1815 ^ n1235 ^ x99 ;
  assign n1817 = n1389 ^ n717 ^ 1'b0 ;
  assign n1818 = n1708 ^ n221 ^ 1'b0 ;
  assign n1819 = ~n924 & n1818 ;
  assign n1820 = x89 & ~n175 ;
  assign n1821 = n1820 ^ n248 ^ 1'b0 ;
  assign n1822 = n1821 ^ x98 ^ 1'b0 ;
  assign n1823 = n998 & ~n1822 ;
  assign n1827 = n1020 ^ n491 ^ n396 ;
  assign n1824 = x98 & n689 ;
  assign n1825 = ~n150 & n1824 ;
  assign n1826 = n770 | n1825 ;
  assign n1828 = n1827 ^ n1826 ^ 1'b0 ;
  assign n1829 = ( ~n252 & n671 ) | ( ~n252 & n1828 ) | ( n671 & n1828 ) ;
  assign n1830 = x44 | n636 ;
  assign n1831 = n1720 ^ n851 ^ 1'b0 ;
  assign n1832 = n660 | n778 ;
  assign n1833 = n538 & ~n1832 ;
  assign n1834 = ~n1055 & n1658 ;
  assign n1835 = n1437 & n1834 ;
  assign n1838 = n159 ^ x114 ^ 1'b0 ;
  assign n1836 = x94 & n1034 ;
  assign n1837 = n1836 ^ n1301 ^ 1'b0 ;
  assign n1839 = n1838 ^ n1837 ^ n1151 ;
  assign n1840 = n450 & n707 ;
  assign n1841 = n1840 ^ x69 ^ 1'b0 ;
  assign n1842 = n380 & ~n1841 ;
  assign n1843 = x12 | n354 ;
  assign n1844 = n153 & ~n1843 ;
  assign n1845 = ~n1842 & n1844 ;
  assign n1846 = ~n1272 & n1845 ;
  assign n1847 = n1076 & n1815 ;
  assign n1848 = n1847 ^ n1015 ^ 1'b0 ;
  assign n1849 = n1848 ^ n1270 ^ 1'b0 ;
  assign n1850 = n879 ^ x82 ^ 1'b0 ;
  assign n1851 = n1667 ^ n555 ^ 1'b0 ;
  assign n1852 = n1059 & ~n1519 ;
  assign n1853 = n1852 ^ n1048 ^ 1'b0 ;
  assign n1854 = n771 & n1051 ;
  assign n1855 = n1853 & n1854 ;
  assign n1856 = n638 | n1855 ;
  assign n1857 = n796 ^ n408 ^ 1'b0 ;
  assign n1858 = n800 ^ n522 ^ 1'b0 ;
  assign n1859 = n1033 | n1858 ;
  assign n1860 = n1857 & ~n1859 ;
  assign n1861 = n826 ^ n722 ^ 1'b0 ;
  assign n1862 = n1204 ^ x5 ^ 1'b0 ;
  assign n1863 = n1087 & ~n1862 ;
  assign n1864 = n1863 ^ n601 ^ 1'b0 ;
  assign n1865 = ~n711 & n1864 ;
  assign n1866 = n1002 ^ n800 ^ 1'b0 ;
  assign n1867 = n1120 ^ n169 ^ 1'b0 ;
  assign n1868 = ( ~n245 & n1071 ) | ( ~n245 & n1867 ) | ( n1071 & n1867 ) ;
  assign n1869 = x48 & n533 ;
  assign n1870 = n1869 ^ n163 ^ 1'b0 ;
  assign n1871 = n639 | n1468 ;
  assign n1872 = n413 ^ n296 ^ 1'b0 ;
  assign n1873 = n1872 ^ n516 ^ 1'b0 ;
  assign n1874 = n1839 & ~n1873 ;
  assign n1875 = n1177 ^ x127 ^ 1'b0 ;
  assign n1876 = n1875 ^ n801 ^ 1'b0 ;
  assign n1877 = n1876 ^ n931 ^ 1'b0 ;
  assign n1878 = n205 ^ x24 ^ 1'b0 ;
  assign n1879 = x41 & x112 ;
  assign n1880 = n700 & n1879 ;
  assign n1881 = n1185 | n1880 ;
  assign n1882 = n235 | n1881 ;
  assign n1883 = n455 | n1882 ;
  assign n1884 = ~n245 & n604 ;
  assign n1885 = ~n1179 & n1884 ;
  assign n1886 = n616 | n1885 ;
  assign n1887 = n1886 ^ n385 ^ 1'b0 ;
  assign n1888 = x30 & n1887 ;
  assign n1889 = n1422 ^ x53 ^ 1'b0 ;
  assign n1890 = n1888 & n1889 ;
  assign n1891 = n308 & ~n1890 ;
  assign n1892 = n1183 | n1680 ;
  assign n1893 = n529 ^ x34 ^ 1'b0 ;
  assign n1894 = x105 & ~n1893 ;
  assign n1895 = n487 ^ n158 ^ 1'b0 ;
  assign n1896 = n268 | n963 ;
  assign n1897 = n1895 & ~n1896 ;
  assign n1898 = n1467 | n1609 ;
  assign n1899 = n1534 ^ n1260 ^ 1'b0 ;
  assign n1900 = n954 ^ n768 ^ 1'b0 ;
  assign n1901 = n1040 ^ n614 ^ 1'b0 ;
  assign n1902 = n526 & n1901 ;
  assign n1903 = n1900 & n1902 ;
  assign n1904 = n1903 ^ n963 ^ 1'b0 ;
  assign n1905 = x119 & n524 ;
  assign n1906 = n1006 ^ n790 ^ 1'b0 ;
  assign n1907 = n1905 & ~n1906 ;
  assign n1908 = n320 | n579 ;
  assign n1909 = ( ~x43 & n179 ) | ( ~x43 & n610 ) | ( n179 & n610 ) ;
  assign n1910 = n1079 & ~n1909 ;
  assign n1911 = x57 & n1299 ;
  assign n1912 = n1910 & n1911 ;
  assign n1913 = ~n1664 & n1912 ;
  assign n1914 = n355 & n1128 ;
  assign n1915 = ( n1272 & ~n1487 ) | ( n1272 & n1914 ) | ( ~n1487 & n1914 ) ;
  assign n1916 = n634 & n1329 ;
  assign n1917 = n1103 ^ n287 ^ 1'b0 ;
  assign n1918 = n1025 ^ n273 ^ 1'b0 ;
  assign n1922 = n296 ^ x5 ^ 1'b0 ;
  assign n1923 = n583 & ~n1922 ;
  assign n1924 = n1923 ^ n967 ^ n418 ;
  assign n1919 = ( n200 & ~n272 ) | ( n200 & n376 ) | ( ~n272 & n376 ) ;
  assign n1920 = x126 ^ x104 ^ 1'b0 ;
  assign n1921 = ~n1919 & n1920 ;
  assign n1925 = n1924 ^ n1921 ^ 1'b0 ;
  assign n1926 = ~n1741 & n1827 ;
  assign n1927 = ~n450 & n1926 ;
  assign n1928 = n1163 | n1398 ;
  assign n1929 = n1927 | n1928 ;
  assign n1930 = n1929 ^ n1904 ^ 1'b0 ;
  assign n1931 = n375 | n510 ;
  assign n1932 = n1931 ^ n673 ^ 1'b0 ;
  assign n1933 = n574 | n1932 ;
  assign n1934 = n558 & ~n1933 ;
  assign n1935 = n1644 ^ x42 ^ 1'b0 ;
  assign n1936 = n1589 & n1632 ;
  assign n1937 = n1936 ^ n666 ^ 1'b0 ;
  assign n1943 = n1576 ^ x104 ^ 1'b0 ;
  assign n1944 = n904 | n1943 ;
  assign n1938 = n221 & ~n1006 ;
  assign n1939 = n571 & n1938 ;
  assign n1940 = n439 | n1885 ;
  assign n1941 = n1939 & ~n1940 ;
  assign n1942 = n893 | n1941 ;
  assign n1945 = n1944 ^ n1942 ^ 1'b0 ;
  assign n1946 = n1632 ^ n709 ^ 1'b0 ;
  assign n1947 = ~n806 & n1170 ;
  assign n1948 = n652 ^ n464 ^ 1'b0 ;
  assign n1949 = ~n613 & n981 ;
  assign n1950 = n1949 ^ x113 ^ 1'b0 ;
  assign n1951 = n1950 ^ n307 ^ 1'b0 ;
  assign n1952 = n825 & ~n1768 ;
  assign n1953 = n326 & ~n1005 ;
  assign n1954 = n1953 ^ n1374 ^ 1'b0 ;
  assign n1955 = n1680 ^ x15 ^ 1'b0 ;
  assign n1956 = x107 & ~n713 ;
  assign n1957 = n134 & n1956 ;
  assign n1958 = ~x53 & n870 ;
  assign n1959 = ~n898 & n1051 ;
  assign n1960 = n782 & n1022 ;
  assign n1961 = n1959 & n1960 ;
  assign n1962 = n1329 ^ n1054 ^ 1'b0 ;
  assign n1963 = n620 & ~n1962 ;
  assign n1967 = n1199 ^ n1192 ^ 1'b0 ;
  assign n1968 = n308 & ~n1967 ;
  assign n1969 = n558 & n1968 ;
  assign n1970 = n1969 ^ n747 ^ 1'b0 ;
  assign n1964 = n1080 & n1389 ;
  assign n1965 = ~n1423 & n1964 ;
  assign n1966 = n1965 ^ n579 ^ 1'b0 ;
  assign n1971 = n1970 ^ n1966 ^ 1'b0 ;
  assign n1972 = n1963 & n1971 ;
  assign n1973 = ( ~x119 & n200 ) | ( ~x119 & n623 ) | ( n200 & n623 ) ;
  assign n1974 = n1973 ^ n1655 ^ x77 ;
  assign n1975 = n1542 & ~n1974 ;
  assign n1976 = n433 ^ n339 ^ 1'b0 ;
  assign n1977 = n581 | n1845 ;
  assign n1978 = x112 & ~n261 ;
  assign n1979 = n1588 & n1978 ;
  assign n1980 = n1133 & ~n1185 ;
  assign n1981 = n242 & n1191 ;
  assign n1982 = n444 & ~n1012 ;
  assign n1983 = ~n194 & n220 ;
  assign n1984 = x14 & ~n1983 ;
  assign n1985 = x64 & ~n1984 ;
  assign n1986 = n1399 | n1537 ;
  assign n1987 = x54 & n1244 ;
  assign n1990 = ~n545 & n1191 ;
  assign n1991 = n493 | n1990 ;
  assign n1988 = n1547 ^ x71 ^ 1'b0 ;
  assign n1989 = ~n990 & n1988 ;
  assign n1992 = n1991 ^ n1989 ^ 1'b0 ;
  assign n1993 = n851 | n1444 ;
  assign n1994 = n424 | n1472 ;
  assign n1995 = ~n934 & n1994 ;
  assign n1996 = n259 & n1995 ;
  assign n1997 = ~n996 & n1726 ;
  assign n1998 = n998 & n1997 ;
  assign n1999 = ~n1527 & n1874 ;
  assign n2000 = n594 & n1284 ;
  assign n2001 = n1072 | n1107 ;
  assign n2002 = n2000 & ~n2001 ;
  assign n2003 = n163 & n1348 ;
  assign n2004 = n424 & ~n1277 ;
  assign n2005 = ~n1888 & n2004 ;
  assign n2006 = n1186 & ~n1385 ;
  assign n2007 = n1468 ^ n1467 ^ 1'b0 ;
  assign n2008 = n231 & n2007 ;
  assign n2009 = ~n1063 & n2008 ;
  assign n2010 = n468 | n2009 ;
  assign n2011 = n512 & ~n806 ;
  assign n2012 = n2011 ^ n879 ^ 1'b0 ;
  assign n2013 = ~n400 & n849 ;
  assign n2014 = n2013 ^ n632 ^ 1'b0 ;
  assign n2020 = n530 | n1144 ;
  assign n2017 = n1901 ^ n1209 ^ 1'b0 ;
  assign n2015 = ( n483 & ~n1204 ) | ( n483 & n1718 ) | ( ~n1204 & n1718 ) ;
  assign n2016 = n2015 ^ n1369 ^ 1'b0 ;
  assign n2018 = n2017 ^ n2016 ^ 1'b0 ;
  assign n2019 = n1378 & n2018 ;
  assign n2021 = n2020 ^ n2019 ^ 1'b0 ;
  assign n2022 = n1089 ^ n638 ^ 1'b0 ;
  assign n2023 = ~n892 & n2022 ;
  assign n2024 = n671 ^ n444 ^ 1'b0 ;
  assign n2025 = n261 | n2024 ;
  assign n2026 = n2025 ^ n1584 ^ 1'b0 ;
  assign n2027 = n1400 ^ n134 ^ 1'b0 ;
  assign n2028 = n567 | n2027 ;
  assign n2029 = ~n899 & n1453 ;
  assign n2030 = n2029 ^ n1708 ^ 1'b0 ;
  assign n2031 = n1637 & ~n2030 ;
  assign n2032 = n506 & n2031 ;
  assign n2033 = n2028 | n2032 ;
  assign n2034 = n2026 & ~n2033 ;
  assign n2035 = n391 & n1321 ;
  assign n2036 = n1748 | n2035 ;
  assign n2037 = n432 & ~n2036 ;
  assign n2038 = ~n1167 & n1973 ;
  assign n2039 = n665 ^ n134 ^ 1'b0 ;
  assign n2040 = ~n520 & n2039 ;
  assign n2041 = x14 & n2040 ;
  assign n2042 = n995 ^ n381 ^ 1'b0 ;
  assign n2043 = n1034 | n2042 ;
  assign n2044 = n1467 & ~n2043 ;
  assign n2052 = n496 ^ n390 ^ 1'b0 ;
  assign n2053 = ~n391 & n2052 ;
  assign n2046 = n240 & ~n300 ;
  assign n2047 = ~x6 & n2046 ;
  assign n2045 = ~n251 & n768 ;
  assign n2048 = n2047 ^ n2045 ^ 1'b0 ;
  assign n2049 = n2048 ^ x112 ^ 1'b0 ;
  assign n2050 = n1167 & ~n2049 ;
  assign n2051 = n893 & n2050 ;
  assign n2054 = n2053 ^ n2051 ^ 1'b0 ;
  assign n2055 = n1038 | n1760 ;
  assign n2056 = n446 ^ x96 ^ 1'b0 ;
  assign n2057 = x84 ^ x52 ^ 1'b0 ;
  assign n2058 = n2056 & n2057 ;
  assign n2059 = n1171 ^ n643 ^ 1'b0 ;
  assign n2060 = n2058 & ~n2059 ;
  assign n2061 = n911 & n2060 ;
  assign n2062 = n2061 ^ n1800 ^ 1'b0 ;
  assign n2063 = n537 | n648 ;
  assign n2064 = n2063 ^ n603 ^ 1'b0 ;
  assign n2065 = x67 & n2064 ;
  assign n2066 = n2065 ^ x3 ^ 1'b0 ;
  assign n2067 = n1177 & n2066 ;
  assign n2068 = x45 & n2067 ;
  assign n2069 = n846 & n2068 ;
  assign n2070 = n2069 ^ n1398 ^ 1'b0 ;
  assign n2071 = ~n392 & n932 ;
  assign n2072 = n2071 ^ n763 ^ 1'b0 ;
  assign n2073 = n2072 ^ n847 ^ 1'b0 ;
  assign n2074 = n1061 & ~n2073 ;
  assign n2075 = n277 & n640 ;
  assign n2076 = n2075 ^ n200 ^ 1'b0 ;
  assign n2079 = ( ~x17 & x70 ) | ( ~x17 & n1827 ) | ( x70 & n1827 ) ;
  assign n2077 = n1291 & ~n1932 ;
  assign n2078 = n2077 ^ x100 ^ 1'b0 ;
  assign n2080 = n2079 ^ n2078 ^ 1'b0 ;
  assign n2081 = n540 & ~n2080 ;
  assign n2082 = n2081 ^ x67 ^ 1'b0 ;
  assign n2083 = n600 ^ n567 ^ 1'b0 ;
  assign n2084 = n2083 ^ n960 ^ 1'b0 ;
  assign n2085 = n1792 & n2084 ;
  assign n2086 = n2082 & n2085 ;
  assign n2087 = n594 & n717 ;
  assign n2088 = n177 | n441 ;
  assign n2089 = n2088 ^ n1115 ^ 1'b0 ;
  assign n2090 = n2087 | n2089 ;
  assign n2091 = n891 & n1734 ;
  assign n2092 = ~n1091 & n2091 ;
  assign n2093 = n2092 ^ n1427 ^ 1'b0 ;
  assign n2094 = n1308 & ~n2093 ;
  assign n2095 = n399 | n1880 ;
  assign n2096 = n2095 ^ n512 ^ 1'b0 ;
  assign n2097 = n859 ^ n473 ^ 1'b0 ;
  assign n2098 = n1304 & ~n2097 ;
  assign n2099 = n2098 ^ n359 ^ 1'b0 ;
  assign n2100 = n489 ^ n216 ^ 1'b0 ;
  assign n2101 = x23 & n2100 ;
  assign n2102 = n1523 ^ n1194 ^ 1'b0 ;
  assign n2103 = n2101 & n2102 ;
  assign n2104 = n2103 ^ n1811 ^ 1'b0 ;
  assign n2105 = n1162 & ~n2104 ;
  assign n2106 = ~n1289 & n1828 ;
  assign n2107 = n2106 ^ n831 ^ 1'b0 ;
  assign n2108 = n937 ^ n891 ^ 1'b0 ;
  assign n2109 = n2107 | n2108 ;
  assign n2111 = x64 & ~n836 ;
  assign n2112 = n711 & n2111 ;
  assign n2110 = ~x127 & n952 ;
  assign n2113 = n2112 ^ n2110 ^ 1'b0 ;
  assign n2114 = n886 | n934 ;
  assign n2115 = n2114 ^ n237 ^ 1'b0 ;
  assign n2116 = n2113 & n2115 ;
  assign n2117 = n2116 ^ n858 ^ 1'b0 ;
  assign n2118 = n698 ^ n326 ^ 1'b0 ;
  assign n2119 = n564 & n2118 ;
  assign n2120 = ~n992 & n2119 ;
  assign n2121 = ~n955 & n2120 ;
  assign n2122 = x18 & ~n2121 ;
  assign n2123 = ~n153 & n266 ;
  assign n2124 = ~n885 & n1788 ;
  assign n2125 = n276 & n2124 ;
  assign n2126 = n2125 ^ n1653 ^ 1'b0 ;
  assign n2127 = ~n383 & n2126 ;
  assign n2128 = n435 | n1768 ;
  assign n2129 = n2127 | n2128 ;
  assign n2131 = n444 | n1006 ;
  assign n2132 = n1147 & ~n2131 ;
  assign n2130 = n834 | n1317 ;
  assign n2133 = n2132 ^ n2130 ^ 1'b0 ;
  assign n2134 = n1512 | n2133 ;
  assign n2135 = n2134 ^ x12 ^ 1'b0 ;
  assign n2136 = ~n1368 & n2135 ;
  assign n2137 = ~n1946 & n2136 ;
  assign n2138 = x35 & ~n995 ;
  assign n2139 = n2138 ^ n571 ^ 1'b0 ;
  assign n2140 = n1054 ^ n503 ^ 1'b0 ;
  assign n2141 = n207 & ~n2140 ;
  assign n2142 = n2141 ^ n1542 ^ 1'b0 ;
  assign n2143 = ( ~x105 & n266 ) | ( ~x105 & n604 ) | ( n266 & n604 ) ;
  assign n2144 = x80 & ~x88 ;
  assign n2145 = n739 & n2144 ;
  assign n2146 = n496 | n1854 ;
  assign n2147 = n790 ^ n324 ^ 1'b0 ;
  assign n2148 = n1397 & ~n2147 ;
  assign n2149 = n647 & n1306 ;
  assign n2150 = n962 ^ n273 ^ 1'b0 ;
  assign n2151 = n954 & ~n2150 ;
  assign n2152 = ~n973 & n2151 ;
  assign n2153 = n272 & n2152 ;
  assign n2154 = ~x48 & n1620 ;
  assign n2155 = n2154 ^ x109 ^ 1'b0 ;
  assign n2158 = x17 & n729 ;
  assign n2159 = n1289 & n2158 ;
  assign n2157 = n938 & n1663 ;
  assign n2160 = n2159 ^ n2157 ^ 1'b0 ;
  assign n2156 = n739 & ~n1267 ;
  assign n2161 = n2160 ^ n2156 ^ 1'b0 ;
  assign n2162 = n834 | n2161 ;
  assign n2163 = n231 | n2162 ;
  assign n2164 = n618 & n1493 ;
  assign n2165 = n1796 & n2164 ;
  assign n2166 = ~n243 & n262 ;
  assign n2167 = n1984 & ~n2108 ;
  assign n2168 = n1062 & n2167 ;
  assign n2169 = n1821 ^ n439 ^ 1'b0 ;
  assign n2170 = ~n427 & n2169 ;
  assign n2171 = n1064 & ~n2170 ;
  assign n2172 = ~n501 & n1400 ;
  assign n2173 = n1016 & n2172 ;
  assign n2174 = x39 & n300 ;
  assign n2175 = n336 & ~n2174 ;
  assign n2176 = n2173 & n2175 ;
  assign n2177 = n1928 | n2176 ;
  assign n2178 = n1352 ^ n1135 ^ 1'b0 ;
  assign n2179 = ( n2171 & ~n2177 ) | ( n2171 & n2178 ) | ( ~n2177 & n2178 ) ;
  assign n2180 = n356 | n482 ;
  assign n2181 = n1694 & ~n2180 ;
  assign n2182 = n1737 ^ n594 ^ 1'b0 ;
  assign n2183 = n385 & n1228 ;
  assign n2184 = n252 & ~n1914 ;
  assign n2185 = n2184 ^ n1547 ^ 1'b0 ;
  assign n2186 = ( x36 & n983 ) | ( x36 & n2185 ) | ( n983 & n2185 ) ;
  assign n2187 = n1057 ^ n516 ^ 1'b0 ;
  assign n2188 = ~n1167 & n2187 ;
  assign n2189 = ~n557 & n2188 ;
  assign n2190 = n2189 ^ x27 ^ 1'b0 ;
  assign n2191 = n1972 ^ n928 ^ 1'b0 ;
  assign n2192 = n873 | n958 ;
  assign n2193 = n2192 ^ n2075 ^ 1'b0 ;
  assign n2194 = n1667 ^ n1052 ^ n492 ;
  assign n2195 = n810 ^ n507 ^ 1'b0 ;
  assign n2196 = n2194 | n2195 ;
  assign n2197 = n562 & ~n1030 ;
  assign n2198 = ~n1697 & n2197 ;
  assign n2199 = n1214 ^ n613 ^ 1'b0 ;
  assign n2200 = n2198 & n2199 ;
  assign n2201 = ~n1207 & n1606 ;
  assign n2202 = n687 & n844 ;
  assign n2203 = n2202 ^ x47 ^ 1'b0 ;
  assign n2204 = n1034 | n2203 ;
  assign n2205 = n597 & n2166 ;
  assign n2206 = n2204 & n2205 ;
  assign n2207 = n1550 ^ n790 ^ 1'b0 ;
  assign n2208 = n1030 | n2207 ;
  assign n2209 = n293 & ~n2208 ;
  assign n2210 = n2209 ^ x44 ^ 1'b0 ;
  assign n2211 = n2210 ^ n1650 ^ 1'b0 ;
  assign n2212 = x87 & ~n2211 ;
  assign n2213 = n494 & n1264 ;
  assign n2214 = ~n574 & n604 ;
  assign n2215 = n2214 ^ n1986 ^ 1'b0 ;
  assign n2216 = n1769 ^ n988 ^ 1'b0 ;
  assign n2217 = x83 & ~n2216 ;
  assign n2218 = n2217 ^ n1067 ^ 1'b0 ;
  assign n2219 = ~n590 & n862 ;
  assign n2220 = n806 | n1845 ;
  assign n2221 = n2219 & ~n2220 ;
  assign n2222 = x12 | n2177 ;
  assign n2223 = n2020 & n2103 ;
  assign n2224 = ~n308 & n2223 ;
  assign n2225 = n960 | n2224 ;
  assign n2226 = n2225 ^ n1699 ^ 1'b0 ;
  assign n2227 = ~n575 & n1067 ;
  assign n2228 = x96 & n2156 ;
  assign n2229 = n2227 & n2228 ;
  assign n2230 = n254 & ~n1714 ;
  assign n2231 = n1293 ^ n1082 ^ 1'b0 ;
  assign n2232 = n161 | n344 ;
  assign n2233 = n2231 & ~n2232 ;
  assign n2234 = ~x12 & x75 ;
  assign n2235 = n946 | n1498 ;
  assign n2236 = n2234 | n2235 ;
  assign n2237 = ~x61 & n1331 ;
  assign n2238 = ( n262 & n786 ) | ( n262 & ~n2237 ) | ( n786 & ~n2237 ) ;
  assign n2239 = n1966 & ~n2238 ;
  assign n2240 = n1631 & n2239 ;
  assign n2241 = n1482 & ~n1753 ;
  assign n2242 = n482 ^ n250 ^ 1'b0 ;
  assign n2243 = n1321 ^ n246 ^ 1'b0 ;
  assign n2244 = n430 | n2243 ;
  assign n2245 = n1398 & ~n2244 ;
  assign n2246 = n749 & n2215 ;
  assign n2247 = n427 | n1897 ;
  assign n2248 = n2247 ^ n2163 ^ 1'b0 ;
  assign n2249 = n1341 ^ n420 ^ 1'b0 ;
  assign n2250 = n2248 & ~n2249 ;
  assign n2251 = ~x12 & n932 ;
  assign n2255 = n1665 ^ n1270 ^ 1'b0 ;
  assign n2252 = n542 & n1399 ;
  assign n2253 = n2252 ^ n713 ^ 1'b0 ;
  assign n2254 = n652 & n2253 ;
  assign n2256 = n2255 ^ n2254 ^ 1'b0 ;
  assign n2258 = x4 & ~n360 ;
  assign n2259 = ~x14 & n2258 ;
  assign n2257 = n1430 ^ n1017 ^ n445 ;
  assign n2260 = n2259 ^ n2257 ^ 1'b0 ;
  assign n2262 = n207 | n519 ;
  assign n2263 = n2262 ^ x0 ^ 1'b0 ;
  assign n2264 = ~n873 & n2263 ;
  assign n2261 = n412 & n728 ;
  assign n2265 = n2264 ^ n2261 ^ 1'b0 ;
  assign n2266 = n2260 & ~n2265 ;
  assign n2267 = n1589 ^ n1385 ^ 1'b0 ;
  assign n2268 = n2267 ^ n992 ^ 1'b0 ;
  assign n2269 = n1207 ^ n1176 ^ 1'b0 ;
  assign n2270 = n833 & n1697 ;
  assign n2271 = n1517 & n2270 ;
  assign n2272 = n888 ^ n837 ^ 1'b0 ;
  assign n2273 = n461 & ~n2272 ;
  assign n2274 = x6 & n2273 ;
  assign n2275 = n2274 ^ n134 ^ 1'b0 ;
  assign n2276 = n1012 ^ n485 ^ 1'b0 ;
  assign n2277 = n175 | n323 ;
  assign n2278 = n2277 ^ n2073 ^ 1'b0 ;
  assign n2279 = n424 ^ x82 ^ 1'b0 ;
  assign n2280 = n221 & n1697 ;
  assign n2281 = n788 & n2280 ;
  assign n2282 = n2281 ^ n2176 ^ 1'b0 ;
  assign n2283 = ~n177 & n2282 ;
  assign n2284 = n324 & n926 ;
  assign n2285 = n2284 ^ n890 ^ 1'b0 ;
  assign n2287 = ~n245 & n1026 ;
  assign n2288 = n1841 & n2287 ;
  assign n2289 = n627 & ~n2288 ;
  assign n2290 = n2289 ^ n1432 ^ x42 ;
  assign n2286 = x13 & ~n1588 ;
  assign n2291 = n2290 ^ n2286 ^ 1'b0 ;
  assign n2292 = n1317 ^ n607 ^ 1'b0 ;
  assign n2293 = ~x127 & n1057 ;
  assign n2294 = n2293 ^ n1604 ^ 1'b0 ;
  assign n2295 = n2198 | n2294 ;
  assign n2296 = ~n695 & n1365 ;
  assign n2297 = n2296 ^ n847 ^ 1'b0 ;
  assign n2298 = n998 & ~n1172 ;
  assign n2299 = n2298 ^ n533 ^ 1'b0 ;
  assign n2300 = x62 & n852 ;
  assign n2301 = n2299 & n2300 ;
  assign n2302 = n2259 | n2301 ;
  assign n2303 = n2302 ^ n2201 ^ 1'b0 ;
  assign n2304 = n1979 ^ n428 ^ 1'b0 ;
  assign n2305 = n355 & n2304 ;
  assign n2306 = ~n892 & n1194 ;
  assign n2307 = n2306 ^ n627 ^ 1'b0 ;
  assign n2308 = n221 & n2307 ;
  assign n2309 = x45 | n1418 ;
  assign n2310 = n905 | n1031 ;
  assign n2311 = n1963 & n2310 ;
  assign n2312 = n2311 ^ n1830 ^ 1'b0 ;
  assign n2313 = n1759 ^ n1188 ^ 1'b0 ;
  assign n2314 = n1393 & n2020 ;
  assign n2315 = n2068 ^ n1463 ^ 1'b0 ;
  assign n2316 = n433 ^ n240 ^ 1'b0 ;
  assign n2317 = n2315 & ~n2316 ;
  assign n2318 = n2030 & n2317 ;
  assign n2319 = n981 & n1880 ;
  assign n2320 = n342 & n381 ;
  assign n2321 = n2320 ^ x86 ^ 1'b0 ;
  assign n2322 = x55 & n1961 ;
  assign n2323 = n711 | n2257 ;
  assign n2324 = n2305 ^ n1132 ^ 1'b0 ;
  assign n2325 = n899 | n1447 ;
  assign n2326 = n2325 ^ n788 ^ 1'b0 ;
  assign n2327 = ~n577 & n2326 ;
  assign n2328 = ~n998 & n2327 ;
  assign n2329 = n1201 | n2328 ;
  assign n2330 = n1632 ^ n642 ^ 1'b0 ;
  assign n2331 = n1247 ^ x54 ^ 1'b0 ;
  assign n2332 = n169 | n2331 ;
  assign n2333 = n2330 | n2332 ;
  assign n2334 = n492 & n1329 ;
  assign n2335 = n2334 ^ x67 ^ 1'b0 ;
  assign n2336 = n134 | n2335 ;
  assign n2337 = n2336 ^ n1632 ^ 1'b0 ;
  assign n2339 = n858 ^ n346 ^ 1'b0 ;
  assign n2338 = n192 | n2284 ;
  assign n2340 = n2339 ^ n2338 ^ 1'b0 ;
  assign n2341 = ~n930 & n1913 ;
  assign n2342 = n2341 ^ x80 ^ 1'b0 ;
  assign n2343 = n766 | n898 ;
  assign n2344 = n2056 ^ n432 ^ x52 ;
  assign n2345 = n1484 & ~n2344 ;
  assign n2346 = n655 ^ n161 ^ 1'b0 ;
  assign n2347 = n1989 & ~n2346 ;
  assign n2348 = n547 & n2347 ;
  assign n2349 = n287 & n2348 ;
  assign n2350 = n1666 | n2299 ;
  assign n2351 = n1249 | n2350 ;
  assign n2352 = x112 | n1335 ;
  assign n2353 = n497 | n1053 ;
  assign n2354 = n2353 ^ n194 ^ 1'b0 ;
  assign n2355 = ~n671 & n2354 ;
  assign n2356 = n1273 & n2355 ;
  assign n2357 = ~n483 & n2356 ;
  assign n2358 = n2349 | n2357 ;
  assign n2359 = n586 & ~n593 ;
  assign n2360 = ~x40 & n2359 ;
  assign n2361 = n491 & n1170 ;
  assign n2362 = n1537 | n2361 ;
  assign n2363 = n2360 & ~n2362 ;
  assign n2364 = n2363 ^ n2232 ^ 1'b0 ;
  assign n2365 = n1861 ^ x81 ^ 1'b0 ;
  assign n2366 = n1700 & n2365 ;
  assign n2367 = n1542 ^ n1180 ^ 1'b0 ;
  assign n2368 = x6 & n822 ;
  assign n2369 = n506 & n2368 ;
  assign n2370 = ~n254 & n1422 ;
  assign n2371 = n2370 ^ n2293 ^ 1'b0 ;
  assign n2374 = n289 & n701 ;
  assign n2375 = n2374 ^ n830 ^ 1'b0 ;
  assign n2376 = n453 | n2375 ;
  assign n2377 = n1437 & ~n2376 ;
  assign n2372 = n2290 ^ n721 ^ 1'b0 ;
  assign n2373 = n725 & n2372 ;
  assign n2378 = n2377 ^ n2373 ^ n1235 ;
  assign n2380 = n984 & ~n1483 ;
  assign n2381 = n2380 ^ n383 ^ 1'b0 ;
  assign n2382 = n636 ^ n576 ^ 1'b0 ;
  assign n2383 = n2381 & ~n2382 ;
  assign n2379 = n823 & ~n1290 ;
  assign n2384 = n2383 ^ n2379 ^ 1'b0 ;
  assign n2385 = n510 & n739 ;
  assign n2386 = n1183 & n2385 ;
  assign n2391 = n1588 ^ n623 ^ 1'b0 ;
  assign n2388 = ( n320 & n342 ) | ( n320 & n992 ) | ( n342 & n992 ) ;
  assign n2387 = n851 | n1030 ;
  assign n2389 = n2388 ^ n2387 ^ 1'b0 ;
  assign n2390 = ( n433 & n2374 ) | ( n433 & ~n2389 ) | ( n2374 & ~n2389 ) ;
  assign n2392 = n2391 ^ n2390 ^ 1'b0 ;
  assign n2393 = ~n971 & n1624 ;
  assign n2394 = n2393 ^ n1469 ^ n870 ;
  assign n2395 = n2392 | n2394 ;
  assign n2396 = n1534 ^ n1151 ^ 1'b0 ;
  assign n2397 = n266 ^ n201 ^ 1'b0 ;
  assign n2398 = ~n2177 & n2397 ;
  assign n2399 = n1552 ^ x2 ^ 1'b0 ;
  assign n2400 = n949 ^ n524 ^ 1'b0 ;
  assign n2403 = n996 ^ x28 ^ 1'b0 ;
  assign n2404 = x83 & n2403 ;
  assign n2401 = x38 & n863 ;
  assign n2402 = n2401 ^ n1732 ^ 1'b0 ;
  assign n2405 = n2404 ^ n2402 ^ 1'b0 ;
  assign n2406 = n531 & ~n2161 ;
  assign n2407 = n2406 ^ n1365 ^ 1'b0 ;
  assign n2408 = n2407 ^ n305 ^ 1'b0 ;
  assign n2409 = n2257 ^ n1510 ^ 1'b0 ;
  assign n2410 = ~n983 & n1966 ;
  assign n2411 = n2409 & n2410 ;
  assign n2412 = n879 ^ n363 ^ 1'b0 ;
  assign n2413 = n2411 | n2412 ;
  assign n2414 = n369 | n1950 ;
  assign n2415 = n2414 ^ n1803 ^ 1'b0 ;
  assign n2416 = x22 & n288 ;
  assign n2417 = n240 | n1193 ;
  assign n2418 = n2416 & ~n2417 ;
  assign n2419 = n1625 ^ n1616 ^ 1'b0 ;
  assign n2420 = n1623 & n2419 ;
  assign n2421 = n2420 ^ n1323 ^ 1'b0 ;
  assign n2422 = ~n1295 & n2421 ;
  assign n2423 = n905 ^ n250 ^ 1'b0 ;
  assign n2424 = n581 | n614 ;
  assign n2425 = n724 & ~n2424 ;
  assign n2426 = ~n2423 & n2425 ;
  assign n2427 = n1061 ^ n922 ^ 1'b0 ;
  assign n2428 = n2427 ^ n1412 ^ 1'b0 ;
  assign n2429 = n453 | n1810 ;
  assign n2430 = n1010 & ~n2429 ;
  assign n2431 = n394 & ~n2430 ;
  assign n2432 = ~n246 & n2431 ;
  assign n2433 = n250 | n2432 ;
  assign n2434 = n526 & ~n1344 ;
  assign n2435 = x35 & n763 ;
  assign n2436 = n2435 ^ n1020 ^ 1'b0 ;
  assign n2437 = n1864 | n2436 ;
  assign n2438 = n2437 ^ n1049 ^ 1'b0 ;
  assign n2439 = x86 & n1135 ;
  assign n2440 = n2439 ^ n354 ^ 1'b0 ;
  assign n2441 = ~n245 & n1071 ;
  assign n2442 = n1345 ^ n579 ^ 1'b0 ;
  assign n2443 = ( n355 & n969 ) | ( n355 & ~n2229 ) | ( n969 & ~n2229 ) ;
  assign n2444 = x27 & n2178 ;
  assign n2445 = n2250 & n2444 ;
  assign n2446 = n153 ^ x106 ^ 1'b0 ;
  assign n2447 = n316 & n594 ;
  assign n2448 = n2447 ^ x109 ^ 1'b0 ;
  assign n2449 = n2448 ^ n1046 ^ 1'b0 ;
  assign n2450 = n832 & ~n2449 ;
  assign n2451 = n1335 & ~n1958 ;
  assign n2452 = n424 & ~n931 ;
  assign n2453 = x87 & ~x103 ;
  assign n2454 = n2453 ^ n1837 ^ n724 ;
  assign n2455 = n731 & n1157 ;
  assign n2456 = n2112 & n2455 ;
  assign n2457 = n2456 ^ n2065 ^ 1'b0 ;
  assign n2458 = n1226 | n2457 ;
  assign n2464 = n2030 ^ n320 ^ 1'b0 ;
  assign n2465 = n358 | n2464 ;
  assign n2459 = ~x105 & n1167 ;
  assign n2460 = n2459 ^ n862 ^ 1'b0 ;
  assign n2461 = n277 & n2460 ;
  assign n2462 = x48 & n2461 ;
  assign n2463 = ~n195 & n2462 ;
  assign n2466 = n2465 ^ n2463 ^ 1'b0 ;
  assign n2467 = ~n591 & n2466 ;
  assign n2468 = ~n885 & n1161 ;
  assign n2469 = n662 | n1958 ;
  assign n2470 = n1876 ^ n788 ^ 1'b0 ;
  assign n2474 = x83 & ~n380 ;
  assign n2475 = n2474 ^ n911 ^ 1'b0 ;
  assign n2471 = ~x9 & n725 ;
  assign n2472 = n1830 & ~n2471 ;
  assign n2473 = n2472 ^ n922 ^ 1'b0 ;
  assign n2476 = n2475 ^ n2473 ^ 1'b0 ;
  assign n2477 = ~n390 & n1901 ;
  assign n2478 = n391 & n2477 ;
  assign n2479 = ~n885 & n2478 ;
  assign n2480 = n2479 ^ n320 ^ 1'b0 ;
  assign n2481 = x17 & n1608 ;
  assign n2482 = n2105 & n2481 ;
  assign n2483 = ~n788 & n2156 ;
  assign n2484 = n2483 ^ n1941 ^ 1'b0 ;
  assign n2485 = x112 & n2484 ;
  assign n2486 = ~n1452 & n2485 ;
  assign n2487 = n880 | n1089 ;
  assign n2488 = n2487 ^ n696 ^ 1'b0 ;
  assign n2489 = n2488 ^ n1756 ^ 1'b0 ;
  assign n2490 = n1265 | n2489 ;
  assign n2491 = n1788 & ~n2113 ;
  assign n2492 = ~n770 & n2491 ;
  assign n2493 = ~n1022 & n2492 ;
  assign n2494 = n763 ^ n158 ^ 1'b0 ;
  assign n2495 = ~n961 & n2494 ;
  assign n2496 = ( n715 & ~n2373 ) | ( n715 & n2495 ) | ( ~n2373 & n2495 ) ;
  assign n2497 = n865 & ~n2328 ;
  assign n2498 = n528 & n1441 ;
  assign n2499 = ~n763 & n2498 ;
  assign n2500 = n934 ^ x91 ^ 1'b0 ;
  assign n2501 = x65 & ~n2500 ;
  assign n2502 = n729 & n937 ;
  assign n2503 = ~n1444 & n2502 ;
  assign n2504 = n1945 | n2503 ;
  assign n2505 = n2501 | n2504 ;
  assign n2506 = n696 ^ n266 ^ 1'b0 ;
  assign n2510 = ~n574 & n1470 ;
  assign n2507 = n194 & n632 ;
  assign n2508 = n2507 ^ n896 ^ 1'b0 ;
  assign n2509 = n1437 & n2508 ;
  assign n2511 = n2510 ^ n2509 ^ 1'b0 ;
  assign n2512 = ( n786 & n983 ) | ( n786 & ~n1741 ) | ( n983 & ~n1741 ) ;
  assign n2513 = n754 ^ n358 ^ n240 ;
  assign n2514 = ~n2512 & n2513 ;
  assign n2515 = n272 & n2514 ;
  assign n2516 = n404 | n2515 ;
  assign n2517 = ~n1030 & n1181 ;
  assign n2518 = n2517 ^ n1829 ^ 1'b0 ;
  assign n2519 = n1723 ^ n1508 ^ 1'b0 ;
  assign n2520 = n1235 | n2519 ;
  assign n2521 = n2520 ^ n707 ^ 1'b0 ;
  assign n2522 = n518 | n930 ;
  assign n2523 = n2522 ^ n918 ^ 1'b0 ;
  assign n2524 = n442 & n1842 ;
  assign n2525 = n2524 ^ n1329 ^ 1'b0 ;
  assign n2526 = n266 & ~n812 ;
  assign n2527 = n1405 ^ n571 ^ 1'b0 ;
  assign n2528 = n2527 ^ n1012 ^ 1'b0 ;
  assign n2529 = ~n2526 & n2528 ;
  assign n2530 = ~n1177 & n1589 ;
  assign n2531 = n1005 & n2530 ;
  assign n2532 = n2529 & n2531 ;
  assign n2533 = n135 | n273 ;
  assign n2534 = n627 & ~n2533 ;
  assign n2535 = ~n1147 & n2534 ;
  assign n2536 = n311 & n882 ;
  assign n2537 = n2536 ^ n1093 ^ 1'b0 ;
  assign n2538 = n583 & ~n2537 ;
  assign n2539 = n1586 & n2538 ;
  assign n2540 = n2539 ^ n1472 ^ 1'b0 ;
  assign n2541 = ~n2535 & n2540 ;
  assign n2542 = n806 ^ n739 ^ 1'b0 ;
  assign n2543 = n792 ^ x100 ^ 1'b0 ;
  assign n2544 = ~n2542 & n2543 ;
  assign n2545 = n2544 ^ n237 ^ 1'b0 ;
  assign n2546 = n1783 ^ n1692 ^ x53 ;
  assign n2548 = n340 | n1558 ;
  assign n2549 = n2548 ^ n1209 ^ 1'b0 ;
  assign n2550 = ~x35 & n2549 ;
  assign n2547 = n696 & n1432 ;
  assign n2551 = n2550 ^ n2547 ^ 1'b0 ;
  assign n2552 = n373 | n1191 ;
  assign n2553 = n1898 ^ n630 ^ 1'b0 ;
  assign n2554 = n2553 ^ n1162 ^ 1'b0 ;
  assign n2555 = ~n175 & n2051 ;
  assign n2557 = n558 & ~n1270 ;
  assign n2558 = n1909 & ~n2557 ;
  assign n2559 = n640 & n2558 ;
  assign n2560 = n1848 | n2559 ;
  assign n2556 = n1126 | n2384 ;
  assign n2561 = n2560 ^ n2556 ^ 1'b0 ;
  assign n2562 = n2549 ^ n1247 ^ 1'b0 ;
  assign n2563 = n1059 & n2562 ;
  assign n2564 = n2563 ^ n601 ^ x93 ;
  assign n2565 = n2564 ^ n2411 ^ n1327 ;
  assign n2566 = n717 & ~n1830 ;
  assign n2567 = n2176 | n2255 ;
  assign n2568 = n2566 & ~n2567 ;
  assign n2569 = n548 & n823 ;
  assign n2570 = n1568 ^ n1055 ^ 1'b0 ;
  assign n2571 = n2570 ^ n2003 ^ 1'b0 ;
  assign n2573 = n2049 ^ n497 ^ 1'b0 ;
  assign n2574 = n2573 ^ n1975 ^ 1'b0 ;
  assign n2572 = x2 & ~n2086 ;
  assign n2575 = n2574 ^ n2572 ^ 1'b0 ;
  assign n2576 = n1073 & ~n2259 ;
  assign n2577 = n1904 ^ n1137 ^ 1'b0 ;
  assign n2578 = ~x46 & n2577 ;
  assign n2579 = n2510 & ~n2578 ;
  assign n2580 = n1534 | n1993 ;
  assign n2581 = n2580 ^ n1135 ^ 1'b0 ;
  assign n2582 = ~n713 & n873 ;
  assign n2583 = ( x44 & n195 ) | ( x44 & n2582 ) | ( n195 & n2582 ) ;
  assign n2584 = n216 & ~n514 ;
  assign n2585 = n1941 | n2584 ;
  assign n2586 = n2585 ^ n724 ^ 1'b0 ;
  assign n2587 = n356 | n2586 ;
  assign n2588 = n1185 ^ n363 ^ 1'b0 ;
  assign n2589 = x41 & n2588 ;
  assign n2590 = ~n1483 & n2589 ;
  assign n2591 = n2587 & n2590 ;
  assign n2592 = n2583 | n2591 ;
  assign n2593 = n216 | n1028 ;
  assign n2594 = n427 & ~n2593 ;
  assign n2595 = n177 | n2594 ;
  assign n2596 = n2595 ^ n1748 ^ 1'b0 ;
  assign n2597 = n2596 ^ n703 ^ 1'b0 ;
  assign n2598 = n164 | n2597 ;
  assign n2599 = n972 ^ n412 ^ 1'b0 ;
  assign n2600 = n2399 & ~n2599 ;
  assign n2601 = n542 & n1656 ;
  assign n2602 = ~n2261 & n2601 ;
  assign n2603 = x37 | n1793 ;
  assign n2604 = n245 & ~n907 ;
  assign n2605 = n1393 ^ n233 ^ 1'b0 ;
  assign n2606 = n2604 & ~n2605 ;
  assign n2607 = ~n1707 & n2552 ;
  assign n2608 = ~n2606 & n2607 ;
  assign n2609 = n939 ^ n144 ^ 1'b0 ;
  assign n2610 = n771 & ~n2609 ;
  assign n2611 = n616 & n2267 ;
  assign n2612 = n1071 & n2611 ;
  assign n2613 = n1955 ^ x88 ^ 1'b0 ;
  assign n2614 = x40 & n2613 ;
  assign n2615 = ( n1188 & n1827 ) | ( n1188 & ~n2313 ) | ( n1827 & ~n2313 ) ;
  assign n2616 = n1391 ^ n480 ^ 1'b0 ;
  assign n2617 = n539 | n2616 ;
  assign n2618 = n1020 | n2617 ;
  assign n2619 = ~n839 & n2618 ;
  assign n2620 = n2619 ^ n806 ^ 1'b0 ;
  assign n2621 = n2440 ^ x22 ^ 1'b0 ;
  assign n2622 = n1316 & ~n1351 ;
  assign n2623 = ~n1853 & n2622 ;
  assign n2624 = x84 | n2623 ;
  assign n2625 = n163 | n428 ;
  assign n2626 = n571 & ~n2625 ;
  assign n2628 = n634 & n701 ;
  assign n2629 = n2628 ^ n1087 ^ 1'b0 ;
  assign n2630 = n2123 & ~n2629 ;
  assign n2627 = n1395 & ~n1554 ;
  assign n2631 = n2630 ^ n2627 ^ 1'b0 ;
  assign n2632 = n175 | n2631 ;
  assign n2633 = ~n208 & n1076 ;
  assign n2634 = n2633 ^ n473 ^ 1'b0 ;
  assign n2635 = ~n1133 & n2488 ;
  assign n2636 = n268 | n1240 ;
  assign n2637 = n2635 & ~n2636 ;
  assign n2638 = n1070 ^ x89 ^ 1'b0 ;
  assign n2639 = n2638 ^ n1133 ^ 1'b0 ;
  assign n2640 = n1067 | n1584 ;
  assign n2641 = n2640 ^ n270 ^ 1'b0 ;
  assign n2642 = n1832 ^ n890 ^ 1'b0 ;
  assign n2643 = n2584 ^ n2143 ^ 1'b0 ;
  assign n2644 = n1216 & n1221 ;
  assign n2645 = x41 & ~n1376 ;
  assign n2646 = n2645 ^ n1101 ^ 1'b0 ;
  assign n2647 = n141 & ~n2646 ;
  assign n2648 = n975 | n1880 ;
  assign n2649 = n365 | n2648 ;
  assign n2654 = x23 & ~n1186 ;
  assign n2655 = n2654 ^ n1291 ^ 1'b0 ;
  assign n2650 = n579 ^ x119 ^ 1'b0 ;
  assign n2651 = n1583 ^ n221 ^ 1'b0 ;
  assign n2652 = ~n2650 & n2651 ;
  assign n2653 = n1208 & n2652 ;
  assign n2656 = n2655 ^ n2653 ^ n1991 ;
  assign n2657 = n2649 & ~n2656 ;
  assign n2658 = n2089 & n2657 ;
  assign n2659 = n1923 & n2240 ;
  assign n2660 = ~n1927 & n2079 ;
  assign n2661 = n2660 ^ n1758 ^ 1'b0 ;
  assign n2662 = n1478 ^ n273 ^ 1'b0 ;
  assign n2663 = n1041 ^ x52 ^ 1'b0 ;
  assign n2664 = n2662 & ~n2663 ;
  assign n2665 = n409 & n2105 ;
  assign n2666 = ~n2664 & n2665 ;
  assign n2667 = ~x79 & n812 ;
  assign n2671 = n1180 ^ x77 ^ 1'b0 ;
  assign n2672 = x114 & n2671 ;
  assign n2673 = n1749 ^ n245 ^ 1'b0 ;
  assign n2674 = n618 & n2673 ;
  assign n2675 = n766 & n2674 ;
  assign n2676 = n2672 & ~n2675 ;
  assign n2677 = n960 & n2676 ;
  assign n2668 = x112 & ~n338 ;
  assign n2669 = ~n526 & n2668 ;
  assign n2670 = ~n1195 & n2669 ;
  assign n2678 = n2677 ^ n2670 ^ 1'b0 ;
  assign n2679 = n1663 & n2678 ;
  assign n2680 = n2679 ^ n782 ^ 1'b0 ;
  assign n2681 = n2667 & n2680 ;
  assign n2682 = ~x119 & n1385 ;
  assign n2685 = n492 ^ n207 ^ 1'b0 ;
  assign n2686 = n645 & ~n2685 ;
  assign n2687 = n1540 & ~n2686 ;
  assign n2683 = n2035 ^ n261 ^ n181 ;
  assign n2684 = n2683 ^ n965 ^ 1'b0 ;
  assign n2688 = n2687 ^ n2684 ^ 1'b0 ;
  assign n2689 = n2682 & n2688 ;
  assign n2690 = n2078 ^ n1919 ^ n784 ;
  assign n2691 = x108 & n1204 ;
  assign n2692 = ~n2219 & n2307 ;
  assign n2693 = n2256 & n2269 ;
  assign n2694 = x127 & n177 ;
  assign n2695 = n629 & ~n1351 ;
  assign n2696 = ~n1082 & n2695 ;
  assign n2697 = n2696 ^ n1558 ^ 1'b0 ;
  assign n2698 = n2697 ^ n243 ^ 1'b0 ;
  assign n2699 = n2694 & ~n2698 ;
  assign n2700 = n389 | n428 ;
  assign n2701 = n607 | n2700 ;
  assign n2702 = n1901 & n2701 ;
  assign n2703 = n242 & ~n737 ;
  assign n2704 = n2703 ^ n387 ^ 1'b0 ;
  assign n2705 = n1671 | n2704 ;
  assign n2714 = n467 & ~n1680 ;
  assign n2715 = ~n349 & n2714 ;
  assign n2708 = x23 & ~n1141 ;
  assign n2709 = n1180 ^ x22 ^ 1'b0 ;
  assign n2710 = n450 | n2709 ;
  assign n2711 = n2708 & n2710 ;
  assign n2706 = n221 & n475 ;
  assign n2707 = n2706 ^ n464 ^ 1'b0 ;
  assign n2712 = n2711 ^ n2707 ^ 1'b0 ;
  assign n2713 = ~n1950 & n2712 ;
  assign n2716 = n2715 ^ n2713 ^ n2309 ;
  assign n2717 = n213 & n531 ;
  assign n2718 = n2717 ^ n761 ^ 1'b0 ;
  assign n2719 = n2718 ^ n507 ^ 1'b0 ;
  assign n2720 = n2719 ^ n2016 ^ 1'b0 ;
  assign n2721 = n2295 | n2720 ;
  assign n2722 = n720 ^ n477 ^ 1'b0 ;
  assign n2723 = ~n572 & n1997 ;
  assign n2724 = ~n2722 & n2723 ;
  assign n2725 = n754 | n1048 ;
  assign n2726 = x53 | n2725 ;
  assign n2728 = n292 | n1049 ;
  assign n2729 = n2728 ^ n727 ^ 1'b0 ;
  assign n2727 = ~n1482 & n2188 ;
  assign n2730 = n2729 ^ n2727 ^ 1'b0 ;
  assign n2731 = n2726 & ~n2730 ;
  assign n2732 = n1932 & n2731 ;
  assign n2733 = n2724 & ~n2732 ;
  assign n2734 = n2381 ^ n1461 ^ 1'b0 ;
  assign n2735 = n2734 ^ n415 ^ 1'b0 ;
  assign n2736 = n1697 ^ n945 ^ 1'b0 ;
  assign n2737 = n2736 ^ n618 ^ 1'b0 ;
  assign n2738 = n607 & n2737 ;
  assign n2739 = n2358 ^ n139 ^ 1'b0 ;
  assign n2740 = x59 & n1167 ;
  assign n2741 = ~n618 & n2740 ;
  assign n2742 = n198 & ~n2741 ;
  assign n2743 = n1054 & n2742 ;
  assign n2744 = n2070 & ~n2743 ;
  assign n2745 = ( n407 & n1229 ) | ( n407 & ~n2744 ) | ( n1229 & ~n2744 ) ;
  assign n2746 = n1508 ^ n889 ^ 1'b0 ;
  assign n2747 = n2264 & n2707 ;
  assign n2748 = n427 & n2747 ;
  assign n2749 = n2746 & ~n2748 ;
  assign n2750 = x112 | n1550 ;
  assign n2754 = n741 ^ n633 ^ 1'b0 ;
  assign n2755 = n131 | n2754 ;
  assign n2751 = n1073 & ~n1267 ;
  assign n2752 = n2751 ^ n553 ^ 1'b0 ;
  assign n2753 = n1624 & ~n2752 ;
  assign n2756 = n2755 ^ n2753 ^ 1'b0 ;
  assign n2757 = n2467 & n2525 ;
  assign n2758 = n607 & ~n2021 ;
  assign n2759 = ~n2614 & n2758 ;
  assign n2760 = n866 ^ n412 ^ 1'b0 ;
  assign n2761 = n2760 ^ n2117 ^ 1'b0 ;
  assign n2762 = n522 | n1862 ;
  assign n2763 = n2762 ^ n1919 ^ 1'b0 ;
  assign n2764 = n2584 ^ x69 ^ 1'b0 ;
  assign n2765 = ~n2763 & n2764 ;
  assign n2766 = ~n1167 & n2765 ;
  assign n2767 = n1762 & n2766 ;
  assign n2768 = n292 | n1517 ;
  assign n2769 = n2416 & ~n2768 ;
  assign n2770 = ~n2767 & n2769 ;
  assign n2771 = n1023 | n1194 ;
  assign n2772 = n2771 ^ n1866 ^ 1'b0 ;
  assign n2773 = n399 | n2772 ;
  assign n2774 = n2773 ^ n1878 ^ 1'b0 ;
  assign n2775 = n1161 & ~n2156 ;
  assign n2776 = n972 & n1636 ;
  assign n2777 = n1861 ^ n346 ^ 1'b0 ;
  assign n2778 = n666 & n822 ;
  assign n2779 = n2778 ^ x108 ^ 1'b0 ;
  assign n2780 = n2667 | n2779 ;
  assign n2781 = n217 & ~n1011 ;
  assign n2782 = ~n994 & n2781 ;
  assign n2783 = n2782 ^ n1178 ^ 1'b0 ;
  assign n2784 = n2153 ^ n1372 ^ 1'b0 ;
  assign n2785 = n1588 | n2784 ;
  assign n2786 = n2367 | n2785 ;
  assign n2787 = n1980 ^ n571 ^ 1'b0 ;
  assign n2788 = ~x31 & n2787 ;
  assign n2789 = n776 & n2788 ;
  assign n2790 = n632 & n796 ;
  assign n2791 = n2790 ^ n1653 ^ 1'b0 ;
  assign n2792 = ~n2709 & n2791 ;
  assign n2799 = n1232 ^ n1137 ^ 1'b0 ;
  assign n2800 = n387 & ~n1162 ;
  assign n2801 = n2213 & n2800 ;
  assign n2802 = n2799 & n2801 ;
  assign n2793 = ~n305 & n613 ;
  assign n2794 = n2793 ^ n1195 ^ 1'b0 ;
  assign n2795 = ~n629 & n2794 ;
  assign n2796 = n2337 ^ n1827 ^ 1'b0 ;
  assign n2797 = n2795 & ~n2796 ;
  assign n2798 = ~n2321 & n2797 ;
  assign n2803 = n2802 ^ n2798 ^ 1'b0 ;
  assign n2804 = n1139 & n1741 ;
  assign n2805 = n408 & n642 ;
  assign n2806 = n1476 & n2805 ;
  assign n2807 = n1228 | n2806 ;
  assign n2808 = n1760 & ~n2807 ;
  assign n2809 = n834 | n972 ;
  assign n2810 = ~n2350 & n2809 ;
  assign n2811 = n2810 ^ n1317 ^ 1'b0 ;
  assign n2812 = n983 | n2811 ;
  assign n2813 = n806 & ~n2812 ;
  assign n2814 = n2808 | n2813 ;
  assign n2815 = n1563 & ~n2814 ;
  assign n2816 = n2444 & ~n2815 ;
  assign n2817 = n2816 ^ x24 ^ 1'b0 ;
  assign n2818 = n2817 ^ n2569 ^ 1'b0 ;
  assign n2819 = n707 & ~n1814 ;
  assign n2820 = n983 | n2173 ;
  assign n2821 = n2820 ^ n481 ^ 1'b0 ;
  assign n2822 = n2821 ^ n737 ^ x105 ;
  assign n2823 = n1449 ^ n1425 ^ 1'b0 ;
  assign n2824 = n1583 & n2823 ;
  assign n2825 = n1251 & ~n2559 ;
  assign n2826 = n2825 ^ x16 ^ 1'b0 ;
  assign n2827 = n2432 ^ n1374 ^ 1'b0 ;
  assign n2828 = n1366 | n1476 ;
  assign n2829 = n2389 | n2828 ;
  assign n2830 = n2829 ^ n1459 ^ 1'b0 ;
  assign n2831 = n1613 & ~n2830 ;
  assign n2832 = n203 & ~n2221 ;
  assign n2833 = n574 & n2832 ;
  assign n2834 = n974 ^ n510 ^ 1'b0 ;
  assign n2835 = ~n650 & n2834 ;
  assign n2836 = n1854 ^ n1393 ^ 1'b0 ;
  assign n2837 = n1333 & n2684 ;
  assign n2838 = n2836 & n2837 ;
  assign n2839 = n1609 & ~n2592 ;
  assign n2840 = n496 ^ n330 ^ 1'b0 ;
  assign n2841 = n410 & ~n2840 ;
  assign n2842 = n258 & n2841 ;
  assign n2843 = n1504 ^ n576 ^ 1'b0 ;
  assign n2845 = ~n788 & n1209 ;
  assign n2846 = n1049 & n2845 ;
  assign n2847 = n2846 ^ n152 ^ 1'b0 ;
  assign n2848 = n1849 | n2847 ;
  assign n2844 = ~n1369 & n1867 ;
  assign n2849 = n2848 ^ n2844 ^ 1'b0 ;
  assign n2850 = n1871 ^ n205 ^ 1'b0 ;
  assign n2852 = n2584 ^ n485 ^ n314 ;
  assign n2851 = n1103 & n2488 ;
  assign n2853 = n2852 ^ n2851 ^ 1'b0 ;
  assign n2854 = n1010 | n2853 ;
  assign n2855 = ~n1632 & n2854 ;
  assign n2856 = ~n2331 & n2722 ;
  assign n2857 = ~x63 & n2856 ;
  assign n2858 = n1994 ^ n1948 ^ 1'b0 ;
  assign n2859 = n2443 ^ n1149 ^ 1'b0 ;
  assign n2860 = n717 & ~n1558 ;
  assign n2861 = n1597 & n2860 ;
  assign n2862 = n2861 ^ n1648 ^ n375 ;
  assign n2863 = n914 | n1769 ;
  assign n2864 = n2863 ^ n2299 ^ 1'b0 ;
  assign n2865 = n2864 ^ n773 ^ 1'b0 ;
  assign n2866 = ~n2862 & n2865 ;
  assign n2867 = n2323 ^ n217 ^ 1'b0 ;
  assign n2870 = n1626 & ~n2032 ;
  assign n2871 = ~n2732 & n2870 ;
  assign n2868 = n747 | n899 ;
  assign n2869 = n537 | n2868 ;
  assign n2872 = n2871 ^ n2869 ^ 1'b0 ;
  assign n2873 = n2557 ^ n1167 ^ 1'b0 ;
  assign n2874 = n2873 ^ n2465 ^ n1932 ;
  assign n2875 = ( n492 & ~n1833 ) | ( n492 & n2874 ) | ( ~n1833 & n2874 ) ;
  assign n2876 = n445 & n2690 ;
  assign n2877 = ~n185 & n1057 ;
  assign n2878 = n2877 ^ n1374 ^ 1'b0 ;
  assign n2879 = ~n2408 & n2878 ;
  assign n2880 = n1550 & ~n2325 ;
  assign n2881 = n1474 ^ n952 ^ x98 ;
  assign n2882 = n210 & ~n2469 ;
  assign n2883 = n612 ^ n529 ^ 1'b0 ;
  assign n2884 = n358 & ~n2883 ;
  assign n2885 = n1331 ^ n378 ^ 1'b0 ;
  assign n2886 = n702 & n1623 ;
  assign n2887 = n2886 ^ n195 ^ 1'b0 ;
  assign n2888 = n2885 & ~n2887 ;
  assign n2889 = ~n633 & n2888 ;
  assign n2890 = n996 ^ n482 ^ 1'b0 ;
  assign n2891 = n894 | n2890 ;
  assign n2892 = n1984 & n2891 ;
  assign n2893 = n1173 & n2892 ;
  assign n2894 = n2893 ^ n2866 ^ 1'b0 ;
  assign n2895 = ~n2889 & n2894 ;
  assign n2896 = ~n2535 & n2702 ;
  assign n2897 = n693 ^ x106 ^ 1'b0 ;
  assign n2898 = n132 | n2897 ;
  assign n2899 = n759 | n2526 ;
  assign n2900 = n2079 ^ n190 ^ 1'b0 ;
  assign n2901 = x42 & ~n1324 ;
  assign n2902 = n2383 & ~n2458 ;
  assign n2903 = ~n2901 & n2902 ;
  assign n2904 = n604 & n715 ;
  assign n2905 = n560 & n2904 ;
  assign n2906 = ( n737 & n1673 ) | ( n737 & ~n2905 ) | ( n1673 & ~n2905 ) ;
  assign n2907 = n1470 & n1974 ;
  assign n2908 = ~n1661 & n2388 ;
  assign n2909 = n1268 ^ n153 ^ 1'b0 ;
  assign n2910 = n1515 & n2909 ;
  assign n2911 = n2910 ^ n724 ^ 1'b0 ;
  assign n2912 = n1272 | n2911 ;
  assign n2913 = n1457 & ~n2912 ;
  assign n2914 = n1941 ^ n321 ^ 1'b0 ;
  assign n2915 = n707 | n2914 ;
  assign n2916 = ~n724 & n2079 ;
  assign n2917 = n2916 ^ n1681 ^ 1'b0 ;
  assign n2918 = ~n662 & n741 ;
  assign n2919 = n2918 ^ n482 ^ 1'b0 ;
  assign n2920 = n2266 ^ n321 ^ 1'b0 ;
  assign n2921 = n716 & n2920 ;
  assign n2922 = ~n373 & n745 ;
  assign n2923 = n2922 ^ n343 ^ 1'b0 ;
  assign n2924 = n2923 ^ n1107 ^ 1'b0 ;
  assign n2925 = n634 ^ n339 ^ 1'b0 ;
  assign n2926 = n2925 ^ n2887 ^ n880 ;
  assign n2927 = n2926 ^ n2292 ^ 1'b0 ;
  assign n2928 = n1910 | n2927 ;
  assign n2930 = n2650 & ~n2887 ;
  assign n2929 = n727 & ~n1352 ;
  assign n2931 = n2930 ^ n2929 ^ 1'b0 ;
  assign n2932 = n1951 ^ x74 ^ 1'b0 ;
  assign n2933 = n2932 ^ n612 ^ 1'b0 ;
  assign n2934 = n1584 ^ n1452 ^ 1'b0 ;
  assign n2935 = ( n509 & ~n707 ) | ( n509 & n2934 ) | ( ~n707 & n2934 ) ;
  assign n2936 = x70 & n2935 ;
  assign n2937 = n1176 & n2461 ;
  assign n2938 = n354 & ~n2882 ;
  assign n2939 = n1389 | n2642 ;
  assign n2940 = n1703 & ~n2939 ;
  assign n2941 = n1786 ^ x17 ^ 1'b0 ;
  assign n2942 = n1615 & n2649 ;
  assign n2943 = ( x116 & ~n1026 ) | ( x116 & n1950 ) | ( ~n1026 & n1950 ) ;
  assign n2944 = n1212 | n2516 ;
  assign n2945 = n1692 | n2944 ;
  assign n2946 = n853 | n2113 ;
  assign n2947 = n1997 & ~n2946 ;
  assign n2948 = n2947 ^ n277 ^ 1'b0 ;
  assign n2949 = x47 & n956 ;
  assign n2950 = n163 & ~n1030 ;
  assign n2951 = n2950 ^ n1680 ^ 1'b0 ;
  assign n2952 = ~n571 & n2951 ;
  assign n2953 = n2952 ^ n1537 ^ 1'b0 ;
  assign n2954 = x28 & n2953 ;
  assign n2955 = n998 ^ n603 ^ 1'b0 ;
  assign n2956 = n1651 ^ n1502 ^ 1'b0 ;
  assign n2957 = ~n1402 & n2956 ;
  assign n2958 = n1399 & ~n2957 ;
  assign n2959 = ~n356 & n1815 ;
  assign n2960 = ~n911 & n1572 ;
  assign n2961 = n1260 & n2794 ;
  assign n2962 = x88 & ~n2081 ;
  assign n2963 = n2962 ^ x117 ^ 1'b0 ;
  assign n2964 = n2961 & ~n2963 ;
  assign n2965 = n2331 | n2955 ;
  assign n2966 = n2964 | n2965 ;
  assign n2967 = n1746 ^ n1040 ^ 1'b0 ;
  assign n2968 = n2868 ^ n2293 ^ 1'b0 ;
  assign n2969 = n2967 | n2968 ;
  assign n2970 = n1626 ^ n487 ^ 1'b0 ;
  assign n2971 = n2641 & ~n2970 ;
  assign n2972 = n1635 ^ n826 ^ 1'b0 ;
  assign n2973 = n905 & n2972 ;
  assign n2974 = n2973 ^ n1095 ^ 1'b0 ;
  assign n2975 = n2028 ^ n1671 ^ 1'b0 ;
  assign n2976 = n2975 ^ n658 ^ 1'b0 ;
  assign n2977 = ~n2974 & n2976 ;
  assign n2978 = n435 | n784 ;
  assign n2979 = n1452 & ~n2649 ;
  assign n2980 = n2979 ^ n1344 ^ 1'b0 ;
  assign n2981 = n2980 ^ n2130 ^ n975 ;
  assign n2982 = n2068 | n2981 ;
  assign n2983 = n2978 | n2982 ;
  assign n2984 = n1156 & n2461 ;
  assign n2985 = ~n2373 & n2984 ;
  assign n2986 = ~n294 & n1919 ;
  assign n2987 = n2986 ^ n995 ^ 1'b0 ;
  assign n2988 = n2987 ^ n233 ^ 1'b0 ;
  assign n2989 = n1948 ^ x55 ^ 1'b0 ;
  assign n2990 = ~n1493 & n2672 ;
  assign n2991 = ~n2174 & n2275 ;
  assign n2992 = ~n2990 & n2991 ;
  assign n2993 = n2992 ^ n153 ^ 1'b0 ;
  assign n2994 = ~n451 & n608 ;
  assign n2995 = ~n2349 & n2994 ;
  assign n2996 = n1832 ^ n647 ^ 1'b0 ;
  assign n2997 = ( n1793 & n2122 ) | ( n1793 & ~n2996 ) | ( n2122 & ~n2996 ) ;
  assign n2998 = n866 ^ x79 ^ 1'b0 ;
  assign n2999 = n1738 & n1855 ;
  assign n3001 = n1974 ^ n806 ^ 1'b0 ;
  assign n3002 = n1853 & n3001 ;
  assign n3000 = x59 & ~n2981 ;
  assign n3003 = n3002 ^ n3000 ^ 1'b0 ;
  assign n3004 = n3003 ^ n1013 ^ 1'b0 ;
  assign n3005 = n137 & n3004 ;
  assign n3006 = n2999 & n3005 ;
  assign n3007 = ~n884 & n3006 ;
  assign n3008 = n1540 ^ x29 ^ 1'b0 ;
  assign n3009 = ~n1543 & n3008 ;
  assign n3010 = n351 & n438 ;
  assign n3011 = n825 ^ n439 ^ 1'b0 ;
  assign n3012 = n3010 & ~n3011 ;
  assign n3013 = n3012 ^ n2079 ^ 1'b0 ;
  assign n3014 = ~n2555 & n3013 ;
  assign n3015 = n3009 & ~n3014 ;
  assign n3016 = n2669 ^ n494 ^ 1'b0 ;
  assign n3017 = n289 & ~n3016 ;
  assign n3018 = n2186 ^ n571 ^ 1'b0 ;
  assign n3019 = n1327 ^ x125 ^ 1'b0 ;
  assign n3020 = n1214 & ~n3019 ;
  assign n3021 = ~n3018 & n3020 ;
  assign n3022 = n2748 | n3021 ;
  assign n3023 = n404 & ~n3022 ;
  assign n3024 = n3017 & ~n3023 ;
  assign n3025 = n3024 ^ n2196 ^ 1'b0 ;
  assign n3026 = n1046 & n2647 ;
  assign n3027 = n1537 & n3026 ;
  assign n3028 = n604 & n1695 ;
  assign n3029 = n948 & ~n2650 ;
  assign n3030 = n373 | n3029 ;
  assign n3031 = n3030 ^ n3003 ^ 1'b0 ;
  assign n3032 = x99 ^ x93 ^ 1'b0 ;
  assign n3033 = n702 & n954 ;
  assign n3034 = ~n3032 & n3033 ;
  assign n3035 = n2679 | n3034 ;
  assign n3036 = n2383 ^ n1287 ^ 1'b0 ;
  assign n3037 = n747 | n3036 ;
  assign n3038 = n1650 | n3019 ;
  assign n3039 = ~n358 & n1038 ;
  assign n3040 = n3039 ^ n672 ^ 1'b0 ;
  assign n3041 = n1069 | n3040 ;
  assign n3042 = n3041 ^ n2875 ^ 1'b0 ;
  assign n3043 = n971 & n3042 ;
  assign n3044 = n1079 ^ n548 ^ 1'b0 ;
  assign n3045 = n1018 | n3044 ;
  assign n3046 = n1355 | n3045 ;
  assign n3047 = n1464 ^ x65 ^ 1'b0 ;
  assign n3048 = x15 & n1166 ;
  assign n3049 = n3048 ^ n318 ^ 1'b0 ;
  assign n3050 = ~n3047 & n3049 ;
  assign n3051 = ~n417 & n722 ;
  assign n3052 = n1287 & n3051 ;
  assign n3053 = n3052 ^ n2527 ^ 1'b0 ;
  assign n3055 = n473 | n707 ;
  assign n3056 = n3055 ^ n2196 ^ 1'b0 ;
  assign n3054 = n1293 | n1527 ;
  assign n3057 = n3056 ^ n3054 ^ 1'b0 ;
  assign n3058 = n567 | n2704 ;
  assign n3059 = n1963 | n3058 ;
  assign n3060 = ~n1472 & n3059 ;
  assign n3061 = ~n356 & n1236 ;
  assign n3062 = n3061 ^ n595 ^ 1'b0 ;
  assign n3063 = n3062 ^ n1728 ^ 1'b0 ;
  assign n3064 = n2390 ^ x22 ^ 1'b0 ;
  assign n3065 = n3064 ^ x4 ^ 1'b0 ;
  assign n3066 = n2603 & ~n3065 ;
  assign n3067 = n1102 & ~n2227 ;
  assign n3068 = n451 & ~n2337 ;
  assign n3069 = n1996 ^ n747 ^ 1'b0 ;
  assign n3070 = x103 ^ x47 ^ 1'b0 ;
  assign n3071 = n3070 ^ n1321 ^ 1'b0 ;
  assign n3072 = n1463 | n2097 ;
  assign n3073 = n1880 ^ n518 ^ n491 ;
  assign n3074 = n2303 & ~n3073 ;
  assign n3075 = n3074 ^ n1548 ^ 1'b0 ;
  assign n3076 = n504 ^ n250 ^ 1'b0 ;
  assign n3077 = n254 & n2484 ;
  assign n3078 = n847 | n1631 ;
  assign n3079 = n2253 ^ n2038 ^ 1'b0 ;
  assign n3080 = n1945 | n2065 ;
  assign n3081 = n3080 ^ n2373 ^ 1'b0 ;
  assign n3082 = n1010 | n3081 ;
  assign n3083 = n369 | n3082 ;
  assign n3084 = x29 & ~n711 ;
  assign n3085 = ~x35 & n3084 ;
  assign n3086 = n3085 ^ n2170 ^ n1599 ;
  assign n3087 = n3086 ^ n2509 ^ 1'b0 ;
  assign n3088 = n2884 & n3010 ;
  assign n3089 = ~n1508 & n3088 ;
  assign n3091 = ~n194 & n851 ;
  assign n3090 = n1597 ^ x126 ^ 1'b0 ;
  assign n3092 = n3091 ^ n3090 ^ 1'b0 ;
  assign n3093 = ~n1729 & n3092 ;
  assign n3094 = n2774 & n3093 ;
  assign n3095 = n2137 & ~n2186 ;
  assign n3096 = n3095 ^ n538 ^ 1'b0 ;
  assign n3097 = n855 & ~n3093 ;
  assign n3098 = n797 & n2250 ;
  assign n3099 = n1364 ^ n216 ^ 1'b0 ;
  assign n3100 = n1115 | n3099 ;
  assign n3101 = n841 & n1173 ;
  assign n3102 = n3101 ^ x114 ^ 1'b0 ;
  assign n3103 = ~n3100 & n3102 ;
  assign n3104 = n2326 ^ n575 ^ 1'b0 ;
  assign n3105 = n3047 ^ n1226 ^ 1'b0 ;
  assign n3106 = n2253 | n3105 ;
  assign n3107 = n252 & ~n1772 ;
  assign n3108 = n141 | n3107 ;
  assign n3109 = n652 ^ n221 ^ 1'b0 ;
  assign n3110 = x16 & n3109 ;
  assign n3111 = n2516 ^ n177 ^ 1'b0 ;
  assign n3112 = n261 & n3111 ;
  assign n3113 = n1907 ^ n1046 ^ 1'b0 ;
  assign n3114 = ~n1371 & n3113 ;
  assign n3115 = ~n3080 & n3114 ;
  assign n3116 = n512 & n3115 ;
  assign n3117 = ~n806 & n2119 ;
  assign n3118 = ~n311 & n3117 ;
  assign n3119 = n1079 & ~n1131 ;
  assign n3120 = n3119 ^ n711 ^ 1'b0 ;
  assign n3121 = n494 | n2943 ;
  assign n3122 = n353 | n879 ;
  assign n3123 = n3122 ^ x33 ^ 1'b0 ;
  assign n3124 = n1023 ^ x69 ^ 1'b0 ;
  assign n3125 = ~x46 & n550 ;
  assign n3126 = n3125 ^ n2337 ^ 1'b0 ;
  assign n3127 = n1162 ^ n390 ^ 1'b0 ;
  assign n3128 = n457 | n3127 ;
  assign n3129 = n601 & n703 ;
  assign n3130 = ~n237 & n3129 ;
  assign n3131 = n2782 | n3130 ;
  assign n3132 = n614 & ~n3131 ;
  assign n3133 = n1564 & ~n3132 ;
  assign n3134 = ~n414 & n3133 ;
  assign n3135 = n3134 ^ n1974 ^ n879 ;
  assign n3136 = ~n1151 & n2291 ;
  assign n3144 = n270 | n839 ;
  assign n3137 = n316 & ~n1206 ;
  assign n3138 = n3137 ^ n1817 ^ n238 ;
  assign n3139 = n1599 & n2067 ;
  assign n3140 = n1688 & n3139 ;
  assign n3141 = n425 & ~n3140 ;
  assign n3142 = ~n2621 & n3141 ;
  assign n3143 = n3138 | n3142 ;
  assign n3145 = n3144 ^ n3143 ^ 1'b0 ;
  assign n3146 = n1026 & n2395 ;
  assign n3147 = n3146 ^ n1981 ^ 1'b0 ;
  assign n3148 = x56 & ~n785 ;
  assign n3149 = n3148 ^ n773 ^ 1'b0 ;
  assign n3150 = n2388 | n3149 ;
  assign n3151 = n2404 ^ n1255 ^ 1'b0 ;
  assign n3152 = n3151 ^ n220 ^ 1'b0 ;
  assign n3153 = n3152 ^ n1391 ^ 1'b0 ;
  assign n3154 = x61 & n542 ;
  assign n3155 = n3154 ^ n1312 ^ 1'b0 ;
  assign n3156 = n373 & ~n3155 ;
  assign n3157 = n1203 ^ n978 ^ 1'b0 ;
  assign n3158 = ( x4 & n192 ) | ( x4 & ~n3157 ) | ( n192 & ~n3157 ) ;
  assign n3159 = n2056 ^ n1759 ^ 1'b0 ;
  assign n3160 = n360 | n3159 ;
  assign n3161 = x112 & ~n1807 ;
  assign n3162 = n2201 & n3161 ;
  assign n3163 = n3160 & n3162 ;
  assign n3164 = x110 & n583 ;
  assign n3165 = ~n483 & n3164 ;
  assign n3166 = n1629 | n3165 ;
  assign n3167 = n3166 ^ n1188 ^ x73 ;
  assign n3168 = n533 & ~n672 ;
  assign n3169 = n886 & n3168 ;
  assign n3170 = n3169 ^ n2194 ^ 1'b0 ;
  assign n3171 = n2601 & ~n2860 ;
  assign n3172 = n2409 | n3171 ;
  assign n3173 = n1703 | n3172 ;
  assign n3174 = n3173 ^ n2808 ^ 1'b0 ;
  assign n3175 = ~n1571 & n1888 ;
  assign n3176 = n2862 & n3175 ;
  assign n3177 = n1556 ^ n422 ^ 1'b0 ;
  assign n3178 = n3177 ^ n731 ^ 1'b0 ;
  assign n3179 = n1030 | n3178 ;
  assign n3180 = n1892 & ~n3179 ;
  assign n3181 = n1764 ^ n1636 ^ 1'b0 ;
  assign n3182 = ~n2934 & n3181 ;
  assign n3183 = n243 | n1887 ;
  assign n3184 = n3182 | n3183 ;
  assign n3185 = ~n1172 & n1173 ;
  assign n3186 = n3185 ^ n1149 ^ 1'b0 ;
  assign n3187 = ~n1244 & n3186 ;
  assign n3188 = ~n3184 & n3187 ;
  assign n3189 = n1069 ^ x57 ^ 1'b0 ;
  assign n3190 = n2198 | n3189 ;
  assign n3191 = n3190 ^ n1187 ^ 1'b0 ;
  assign n3192 = ~n809 & n2271 ;
  assign n3193 = n2049 ^ n1604 ^ 1'b0 ;
  assign n3194 = n3193 ^ x45 ^ 1'b0 ;
  assign n3195 = n577 | n1378 ;
  assign n3196 = ~n773 & n3195 ;
  assign n3197 = n292 ^ n189 ^ 1'b0 ;
  assign n3198 = x115 & n3197 ;
  assign n3199 = n1887 | n2149 ;
  assign n3200 = n2250 & ~n3199 ;
  assign n3201 = n3200 ^ n1630 ^ 1'b0 ;
  assign n3202 = ~n261 & n998 ;
  assign n3203 = n433 & n3202 ;
  assign n3204 = n445 & n1275 ;
  assign n3205 = x5 & ~n3204 ;
  assign n3206 = n3205 ^ n1044 ^ 1'b0 ;
  assign n3207 = n669 | n3206 ;
  assign n3208 = n2523 | n3207 ;
  assign n3209 = n2738 ^ n694 ^ 1'b0 ;
  assign n3210 = n3208 & ~n3209 ;
  assign n3211 = ~x24 & n1001 ;
  assign n3212 = n1601 ^ n456 ^ 1'b0 ;
  assign n3213 = ~n3211 & n3212 ;
  assign n3214 = n1589 ^ n790 ^ 1'b0 ;
  assign n3215 = x127 & n3214 ;
  assign n3216 = n2746 ^ n1924 ^ 1'b0 ;
  assign n3217 = x55 & ~n3216 ;
  assign n3218 = n1622 & n3217 ;
  assign n3219 = n3215 & n3218 ;
  assign n3220 = n243 & n3219 ;
  assign n3221 = n3220 ^ n2234 ^ 1'b0 ;
  assign n3222 = n1724 & ~n3068 ;
  assign n3223 = n2828 & n3222 ;
  assign n3224 = n1548 & n1837 ;
  assign n3225 = ~n1212 & n3224 ;
  assign n3226 = n3225 ^ n916 ^ 1'b0 ;
  assign n3227 = n1669 & ~n1671 ;
  assign n3228 = ~n504 & n3227 ;
  assign n3229 = n567 | n939 ;
  assign n3230 = n2515 ^ n747 ^ n251 ;
  assign n3231 = n2198 ^ n2015 ^ 1'b0 ;
  assign n3232 = n786 ^ n713 ^ 1'b0 ;
  assign n3233 = n2549 ^ n2103 ^ 1'b0 ;
  assign n3234 = n970 & n3233 ;
  assign n3235 = n2907 ^ n934 ^ 1'b0 ;
  assign n3236 = n3234 & ~n3235 ;
  assign n3237 = n2653 ^ n1185 ^ 1'b0 ;
  assign n3238 = n1167 & ~n1895 ;
  assign n3239 = n361 & n3238 ;
  assign n3240 = ~n1655 & n3239 ;
  assign n3241 = n3240 ^ n1631 ^ 1'b0 ;
  assign n3242 = n1515 & n3241 ;
  assign n3243 = ~n1666 & n2878 ;
  assign n3244 = n3243 ^ n192 ^ 1'b0 ;
  assign n3245 = n235 & n1491 ;
  assign n3246 = n3245 ^ n2099 ^ 1'b0 ;
  assign n3247 = ~n994 & n3246 ;
  assign n3248 = ~n169 & n256 ;
  assign n3249 = ~x58 & n3248 ;
  assign n3250 = n342 & ~n391 ;
  assign n3251 = n2430 & n3250 ;
  assign n3252 = n3019 | n3251 ;
  assign n3253 = n3249 & ~n3252 ;
  assign n3254 = n928 ^ x41 ^ 1'b0 ;
  assign n3255 = ~n3253 & n3254 ;
  assign n3256 = n909 & n1120 ;
  assign n3257 = n2213 & ~n3256 ;
  assign n3258 = n1979 & n3257 ;
  assign n3259 = x19 & n507 ;
  assign n3260 = ~n163 & n3259 ;
  assign n3261 = n3260 ^ n530 ^ 1'b0 ;
  assign n3262 = n2276 & ~n3261 ;
  assign n3263 = n3262 ^ n497 ^ 1'b0 ;
  assign n3264 = ~n3258 & n3263 ;
  assign n3265 = n1753 ^ x52 ^ 1'b0 ;
  assign n3266 = n2292 & ~n3265 ;
  assign n3267 = n1599 ^ n1314 ^ 1'b0 ;
  assign n3268 = n3266 & n3267 ;
  assign n3269 = n1952 & ~n3268 ;
  assign n3270 = n1769 ^ n1645 ^ n1147 ;
  assign n3273 = n1329 ^ n450 ^ 1'b0 ;
  assign n3274 = ~n1410 & n3273 ;
  assign n3272 = n976 ^ n867 ^ 1'b0 ;
  assign n3275 = n3274 ^ n3272 ^ 1'b0 ;
  assign n3271 = x35 & n358 ;
  assign n3276 = n3275 ^ n3271 ^ 1'b0 ;
  assign n3277 = n1830 ^ n514 ^ 1'b0 ;
  assign n3278 = ~n1793 & n3277 ;
  assign n3279 = n614 | n877 ;
  assign n3280 = x120 & n2074 ;
  assign n3281 = n3280 ^ n2227 ^ 1'b0 ;
  assign n3282 = n1803 ^ n439 ^ 1'b0 ;
  assign n3283 = ~n356 & n2690 ;
  assign n3284 = ~n1106 & n3283 ;
  assign n3285 = n3282 & n3284 ;
  assign n3287 = n1689 ^ x61 ^ 1'b0 ;
  assign n3288 = n2035 | n3287 ;
  assign n3289 = n2430 | n3288 ;
  assign n3286 = n1380 ^ n376 ^ 1'b0 ;
  assign n3290 = n3289 ^ n3286 ^ n2451 ;
  assign n3291 = x28 & n333 ;
  assign n3292 = n2818 & n3291 ;
  assign n3293 = n1073 & ~n1206 ;
  assign n3294 = ~n2745 & n2859 ;
  assign n3295 = ~n1602 & n3294 ;
  assign n3296 = n1163 ^ n1157 ^ 1'b0 ;
  assign n3297 = n771 & ~n3296 ;
  assign n3298 = ~n2815 & n3297 ;
  assign n3299 = n1245 | n1457 ;
  assign n3300 = ( n1310 & ~n2206 ) | ( n1310 & n3299 ) | ( ~n2206 & n3299 ) ;
  assign n3301 = n928 & n2587 ;
  assign n3302 = n1758 | n3301 ;
  assign n3303 = n165 & ~n1904 ;
  assign n3304 = n430 & n3303 ;
  assign n3305 = n219 | n266 ;
  assign n3306 = n3305 ^ x41 ^ 1'b0 ;
  assign n3307 = n177 & ~n3306 ;
  assign n3310 = n876 | n1336 ;
  assign n3308 = n2144 ^ n1425 ^ 1'b0 ;
  assign n3309 = n775 & ~n3308 ;
  assign n3311 = n3310 ^ n3309 ^ 1'b0 ;
  assign n3312 = ~n2704 & n3311 ;
  assign n3313 = n448 & ~n497 ;
  assign n3314 = n958 & n3313 ;
  assign n3315 = ~n2854 & n3314 ;
  assign n3316 = n1034 | n3315 ;
  assign n3317 = n2079 & ~n3316 ;
  assign n3318 = n1344 & n3317 ;
  assign n3320 = n972 ^ n316 ^ 1'b0 ;
  assign n3321 = n3320 ^ n1685 ^ 1'b0 ;
  assign n3322 = n1662 & ~n3321 ;
  assign n3323 = ~n1808 & n3322 ;
  assign n3324 = n1631 & n3323 ;
  assign n3319 = ~n1397 & n3010 ;
  assign n3325 = n3324 ^ n3319 ^ 1'b0 ;
  assign n3326 = n3325 ^ n1574 ^ 1'b0 ;
  assign n3327 = n2019 & n3326 ;
  assign n3328 = n1823 | n2767 ;
  assign n3329 = n595 & ~n720 ;
  assign n3330 = n2741 & n3329 ;
  assign n3332 = n579 | n1181 ;
  assign n3333 = n463 | n3332 ;
  assign n3331 = n684 & n2794 ;
  assign n3334 = n3333 ^ n3331 ^ 1'b0 ;
  assign n3335 = n552 & ~n607 ;
  assign n3336 = ~n3334 & n3335 ;
  assign n3337 = n355 & ~n783 ;
  assign n3338 = n3336 & n3337 ;
  assign n3339 = n2193 ^ n1677 ^ 1'b0 ;
  assign n3340 = n3339 ^ n3262 ^ 1'b0 ;
  assign n3341 = x80 & n1927 ;
  assign n3342 = n1769 | n3341 ;
  assign n3343 = n507 & ~n3342 ;
  assign n3344 = n766 & ~n3343 ;
  assign n3346 = n1485 | n2409 ;
  assign n3347 = n2990 | n3346 ;
  assign n3345 = x29 & ~n497 ;
  assign n3348 = n3347 ^ n3345 ^ 1'b0 ;
  assign n3352 = n756 & ~n2058 ;
  assign n3353 = n2179 & n3352 ;
  assign n3349 = x32 & n1333 ;
  assign n3350 = ~n2060 & n3349 ;
  assign n3351 = n1991 | n3350 ;
  assign n3354 = n3353 ^ n3351 ^ 1'b0 ;
  assign n3355 = n315 | n3354 ;
  assign n3356 = n215 & ~n3355 ;
  assign n3357 = n1187 ^ n330 ^ 1'b0 ;
  assign n3358 = n2501 & ~n3357 ;
  assign n3359 = n1444 & n3358 ;
  assign n3360 = n1037 & ~n2264 ;
  assign n3361 = n1049 | n1825 ;
  assign n3362 = n3361 ^ n1964 ^ 1'b0 ;
  assign n3363 = ~n3360 & n3362 ;
  assign n3364 = ~x6 & x108 ;
  assign n3365 = n448 & ~n1927 ;
  assign n3366 = ~n976 & n3365 ;
  assign n3367 = ~x92 & n229 ;
  assign n3368 = n3367 ^ n474 ^ 1'b0 ;
  assign n3369 = n439 | n3368 ;
  assign n3370 = n1541 | n3369 ;
  assign n3371 = n1741 & ~n3370 ;
  assign n3372 = n3366 | n3371 ;
  assign n3373 = n1958 & ~n3372 ;
  assign n3374 = n1882 ^ n304 ^ 1'b0 ;
  assign n3375 = n695 | n3374 ;
  assign n3376 = n3375 ^ n2726 ^ 1'b0 ;
  assign n3377 = n1371 & n1953 ;
  assign n3378 = x22 & n459 ;
  assign n3379 = ~n1939 & n2755 ;
  assign n3380 = n2732 | n2759 ;
  assign n3381 = n3380 ^ n3275 ^ 1'b0 ;
  assign n3382 = n1482 | n2936 ;
  assign n3386 = ~n2194 & n2525 ;
  assign n3383 = n1487 ^ n1073 ^ 1'b0 ;
  assign n3384 = n3383 ^ n2721 ^ 1'b0 ;
  assign n3385 = n2047 | n3384 ;
  assign n3387 = n3386 ^ n3385 ^ 1'b0 ;
  assign n3388 = ~n2413 & n3387 ;
  assign n3390 = n519 | n1915 ;
  assign n3391 = n3152 & ~n3390 ;
  assign n3389 = n1040 & n1405 ;
  assign n3392 = n3391 ^ n3389 ^ 1'b0 ;
  assign n3393 = n1366 & n3074 ;
  assign n3394 = ~n279 & n846 ;
  assign n3395 = ~n3393 & n3394 ;
  assign n3396 = n1107 | n3395 ;
  assign n3397 = n2347 ^ n2115 ^ 1'b0 ;
  assign n3398 = n428 & ~n606 ;
  assign n3399 = n250 & ~n3398 ;
  assign n3400 = ~x25 & n3399 ;
  assign n3401 = n2629 ^ n1179 ^ 1'b0 ;
  assign n3402 = n355 & ~n662 ;
  assign n3403 = ~n3401 & n3402 ;
  assign n3404 = n1267 | n2693 ;
  assign n3405 = n3404 ^ n2520 ^ 1'b0 ;
  assign n3406 = n3403 | n3405 ;
  assign n3407 = n2915 ^ n2550 ^ 1'b0 ;
  assign n3413 = ~x125 & n230 ;
  assign n3408 = n666 & ~n3352 ;
  assign n3409 = n3408 ^ n893 ^ 1'b0 ;
  assign n3410 = n190 & n3409 ;
  assign n3411 = n1849 & n3410 ;
  assign n3412 = n2473 & ~n3411 ;
  assign n3414 = n3413 ^ n3412 ^ 1'b0 ;
  assign n3415 = n3272 & ~n3414 ;
  assign n3416 = n1324 ^ n245 ^ n233 ;
  assign n3417 = ~n1471 & n3416 ;
  assign n3418 = ~n2852 & n3417 ;
  assign n3419 = n3418 ^ n1749 ^ 1'b0 ;
  assign n3420 = n604 & n3350 ;
  assign n3421 = ~n512 & n3420 ;
  assign n3422 = ~n939 & n3421 ;
  assign n3424 = n1838 | n3398 ;
  assign n3425 = n259 & ~n3424 ;
  assign n3423 = ~x106 & n3182 ;
  assign n3426 = n3425 ^ n3423 ^ 1'b0 ;
  assign n3427 = ~n3422 & n3426 ;
  assign n3428 = n3419 & n3427 ;
  assign n3429 = n634 | n3407 ;
  assign n3430 = n2551 ^ n293 ^ 1'b0 ;
  assign n3431 = n3341 ^ n1756 ^ 1'b0 ;
  assign n3432 = ~n1671 & n3124 ;
  assign n3433 = x38 | n741 ;
  assign n3434 = ~n1452 & n3433 ;
  assign n3435 = n340 | n2198 ;
  assign n3436 = x24 & ~n3435 ;
  assign n3437 = ~n164 & n365 ;
  assign n3438 = n360 & n3437 ;
  assign n3439 = n3438 ^ n1532 ^ 1'b0 ;
  assign n3440 = ~n960 & n3439 ;
  assign n3441 = n1107 & n3440 ;
  assign n3442 = n2672 ^ n969 ^ 1'b0 ;
  assign n3443 = n806 | n3442 ;
  assign n3446 = n2430 ^ n562 ^ 1'b0 ;
  assign n3444 = n2229 ^ n262 ^ 1'b0 ;
  assign n3445 = n2263 & ~n3444 ;
  assign n3447 = n3446 ^ n3445 ^ n2601 ;
  assign n3448 = n2206 ^ n2093 ^ 1'b0 ;
  assign n3449 = ~n1784 & n3448 ;
  assign n3450 = ~n2347 & n3449 ;
  assign n3451 = ~x100 & n3012 ;
  assign n3452 = n3451 ^ n3299 ^ 1'b0 ;
  assign n3453 = n2967 ^ n1207 ^ 1'b0 ;
  assign n3454 = n3453 ^ n1610 ^ 1'b0 ;
  assign n3455 = n813 & ~n3454 ;
  assign n3456 = n3455 ^ n2911 ^ 1'b0 ;
  assign n3459 = n2660 ^ x127 ^ 1'b0 ;
  assign n3457 = n392 | n446 ;
  assign n3458 = n3457 ^ x42 ^ 1'b0 ;
  assign n3460 = n3459 ^ n3458 ^ 1'b0 ;
  assign n3461 = ~n2525 & n3460 ;
  assign n3462 = x127 & ~n2121 ;
  assign n3463 = n221 & n547 ;
  assign n3464 = ~n248 & n3463 ;
  assign n3465 = n3464 ^ n1255 ^ 1'b0 ;
  assign n3466 = n2376 & n3465 ;
  assign n3467 = n2578 & ~n3466 ;
  assign n3468 = ~x60 & n3467 ;
  assign n3469 = n483 ^ n396 ^ 1'b0 ;
  assign n3470 = n3469 ^ n1693 ^ 1'b0 ;
  assign n3471 = n1366 & ~n2891 ;
  assign n3472 = n3471 ^ n3413 ^ 1'b0 ;
  assign n3473 = n3470 & ~n3472 ;
  assign n3474 = x1 & n163 ;
  assign n3475 = ( n1059 & ~n1781 ) | ( n1059 & n3474 ) | ( ~n1781 & n3474 ) ;
  assign n3476 = n590 ^ n290 ^ 1'b0 ;
  assign n3477 = n2458 | n3476 ;
  assign n3478 = x1 & ~n1133 ;
  assign n3479 = n3478 ^ n1245 ^ 1'b0 ;
  assign n3480 = n456 & n672 ;
  assign n3481 = n173 & ~n3480 ;
  assign n3482 = n1671 & ~n2582 ;
  assign n3483 = n1222 ^ n857 ^ 1'b0 ;
  assign n3484 = n240 & n1968 ;
  assign n3485 = ~n3483 & n3484 ;
  assign n3486 = ~n2461 & n3485 ;
  assign n3487 = ( n3481 & n3482 ) | ( n3481 & ~n3486 ) | ( n3482 & ~n3486 ) ;
  assign n3488 = n3199 | n3230 ;
  assign n3489 = ~n1613 & n1959 ;
  assign n3490 = x22 & ~n1805 ;
  assign n3491 = n3490 ^ n2925 ^ 1'b0 ;
  assign n3492 = ( ~x73 & n1576 ) | ( ~x73 & n2391 ) | ( n1576 & n2391 ) ;
  assign n3493 = n3439 ^ n764 ^ 1'b0 ;
  assign n3494 = ~n3492 & n3493 ;
  assign n3495 = n684 ^ n216 ^ 1'b0 ;
  assign n3496 = ~n344 & n3495 ;
  assign n3497 = n876 & n1534 ;
  assign n3498 = ~n2056 & n3497 ;
  assign n3499 = n3496 & ~n3498 ;
  assign n3500 = n1144 & n2090 ;
  assign n3501 = ~n1993 & n3500 ;
  assign n3502 = n3501 ^ n2573 ^ 1'b0 ;
  assign n3503 = ~n1543 & n3335 ;
  assign n3504 = n349 & ~n3503 ;
  assign n3505 = n1178 & ~n2792 ;
  assign n3506 = n794 & ~n2000 ;
  assign n3507 = n3506 ^ n828 ^ 1'b0 ;
  assign n3508 = n1766 ^ x73 ^ 1'b0 ;
  assign n3509 = n1228 | n3508 ;
  assign n3510 = n3507 | n3509 ;
  assign n3513 = n267 & ~n2453 ;
  assign n3514 = n3513 ^ n152 ^ 1'b0 ;
  assign n3511 = x69 ^ x55 ^ 1'b0 ;
  assign n3512 = n756 & n3511 ;
  assign n3515 = n3514 ^ n3512 ^ 1'b0 ;
  assign n3516 = n1366 & ~n3515 ;
  assign n3517 = n408 & n3516 ;
  assign n3518 = n3517 ^ n2478 ^ 1'b0 ;
  assign n3519 = n1344 & ~n1427 ;
  assign n3520 = n2125 ^ n1714 ^ 1'b0 ;
  assign n3521 = n1280 & n3520 ;
  assign n3522 = n3521 ^ n2827 ^ 1'b0 ;
  assign n3523 = n270 & ~n3522 ;
  assign n3524 = ~n970 & n2149 ;
  assign n3525 = n1919 & n3524 ;
  assign n3526 = n3290 ^ n750 ^ 1'b0 ;
  assign n3527 = x39 & ~n537 ;
  assign n3528 = ~n694 & n2513 ;
  assign n3529 = n1895 & n3528 ;
  assign n3530 = n3529 ^ n946 ^ 1'b0 ;
  assign n3531 = ~n614 & n3530 ;
  assign n3532 = n3334 & n3531 ;
  assign n3533 = n1406 | n2838 ;
  assign n3534 = n3533 ^ n1984 ^ 1'b0 ;
  assign n3535 = n1234 ^ n1057 ^ 1'b0 ;
  assign n3536 = n2003 | n3535 ;
  assign n3537 = n1918 | n3536 ;
  assign n3538 = n1651 & ~n1789 ;
  assign n3539 = ~n3537 & n3538 ;
  assign n3540 = ~n2083 & n3539 ;
  assign n3541 = n3540 ^ n594 ^ 1'b0 ;
  assign n3542 = n1697 ^ n526 ^ 1'b0 ;
  assign n3543 = n1718 & n2589 ;
  assign n3544 = n3543 ^ n1439 ^ 1'b0 ;
  assign n3545 = ( n577 & n3542 ) | ( n577 & ~n3544 ) | ( n3542 & ~n3544 ) ;
  assign n3546 = n3545 ^ n1704 ^ 1'b0 ;
  assign n3547 = n3079 & ~n3546 ;
  assign n3548 = ~n2159 & n3172 ;
  assign n3549 = n164 & n1073 ;
  assign n3550 = n3549 ^ n861 ^ 1'b0 ;
  assign n3551 = n3191 | n3550 ;
  assign n3552 = n3551 ^ n3211 ^ n537 ;
  assign n3553 = n965 & n2398 ;
  assign n3554 = ~x96 & n1240 ;
  assign n3555 = ~n3411 & n3554 ;
  assign n3556 = n3555 ^ n2446 ^ 1'b0 ;
  assign n3557 = n3545 & ~n3556 ;
  assign n3558 = n3121 ^ n2520 ^ 1'b0 ;
  assign n3559 = n2329 ^ n330 ^ n320 ;
  assign n3560 = ~n409 & n3559 ;
  assign n3561 = ~n795 & n3560 ;
  assign n3562 = ~n132 & n2583 ;
  assign n3563 = n3562 ^ x2 ^ 1'b0 ;
  assign n3564 = x41 | n3563 ;
  assign n3565 = n3564 ^ n1747 ^ 1'b0 ;
  assign n3566 = n744 ^ n305 ^ 1'b0 ;
  assign n3567 = n528 & ~n3566 ;
  assign n3568 = ~n2291 & n3567 ;
  assign n3569 = ~n3014 & n3568 ;
  assign n3570 = ~n842 & n1287 ;
  assign n3571 = n3570 ^ n859 ^ 1'b0 ;
  assign n3572 = n2108 | n3571 ;
  assign n3573 = n3572 ^ n753 ^ 1'b0 ;
  assign n3574 = n2735 ^ n604 ^ 1'b0 ;
  assign n3575 = n3573 & ~n3574 ;
  assign n3576 = n391 ^ x52 ^ 1'b0 ;
  assign n3577 = n2392 & ~n3576 ;
  assign n3578 = n972 & ~n1149 ;
  assign n3579 = n3578 ^ n3031 ^ 1'b0 ;
  assign n3580 = n3213 & n3527 ;
  assign n3581 = ~n564 & n1180 ;
  assign n3582 = ~n1843 & n3581 ;
  assign n3583 = n3582 ^ n2075 ^ 1'b0 ;
  assign n3584 = n3583 ^ n2265 ^ 1'b0 ;
  assign n3585 = n1865 | n1957 ;
  assign n3586 = n687 & ~n3446 ;
  assign n3587 = n1185 & n3586 ;
  assign n3588 = n1894 & ~n3587 ;
  assign n3589 = n3588 ^ n277 ^ 1'b0 ;
  assign n3590 = x36 & ~n1436 ;
  assign n3591 = n3590 ^ n1345 ^ 1'b0 ;
  assign n3592 = ~n1499 & n3591 ;
  assign n3593 = n613 & n1427 ;
  assign n3594 = ~n3592 & n3593 ;
  assign n3595 = n3594 ^ n904 ^ n167 ;
  assign n3596 = n2427 | n2491 ;
  assign n3597 = n3596 ^ n1267 ^ 1'b0 ;
  assign n3598 = n3249 ^ n1030 ^ 1'b0 ;
  assign n3599 = ~n2363 & n3598 ;
  assign n3600 = ~x104 & n634 ;
  assign n3601 = ~n1457 & n3600 ;
  assign n3602 = n3601 ^ n1156 ^ 1'b0 ;
  assign n3603 = x108 & n2563 ;
  assign n3604 = ~n1658 & n3603 ;
  assign n3605 = ~x55 & n2425 ;
  assign n3606 = n3019 ^ n473 ^ 1'b0 ;
  assign n3607 = n616 & n3606 ;
  assign n3608 = n3607 ^ n3177 ^ 1'b0 ;
  assign n3609 = n1015 | n3526 ;
  assign n3610 = x0 | n3609 ;
  assign n3612 = n296 | n2488 ;
  assign n3613 = n874 & ~n3612 ;
  assign n3611 = n1651 & n2860 ;
  assign n3614 = n3613 ^ n3611 ^ 1'b0 ;
  assign n3615 = n219 | n3614 ;
  assign n3617 = n612 & ~n1631 ;
  assign n3618 = n1537 & n3617 ;
  assign n3616 = ~n2842 & n3271 ;
  assign n3619 = n3618 ^ n3616 ^ 1'b0 ;
  assign n3620 = n262 & n1170 ;
  assign n3621 = ~n868 & n3620 ;
  assign n3622 = ~n177 & n3621 ;
  assign n3623 = n618 & ~n1897 ;
  assign n3624 = n3623 ^ n1279 ^ 1'b0 ;
  assign n3625 = n2606 ^ n2224 ^ 1'b0 ;
  assign n3626 = n1070 & ~n3625 ;
  assign n3627 = ~n3624 & n3626 ;
  assign n3628 = ( ~n1048 & n3622 ) | ( ~n1048 & n3627 ) | ( n3622 & n3627 ) ;
  assign n3629 = ~n1496 & n2402 ;
  assign n3630 = n3135 ^ n717 ^ 1'b0 ;
  assign n3631 = n1574 & n1828 ;
  assign n3632 = n3631 ^ n2349 ^ 1'b0 ;
  assign n3633 = ~n2144 & n3632 ;
  assign n3634 = ~n886 & n2079 ;
  assign n3636 = n735 ^ n466 ^ 1'b0 ;
  assign n3635 = n360 & n3420 ;
  assign n3637 = n3636 ^ n3635 ^ 1'b0 ;
  assign n3638 = n645 & ~n2065 ;
  assign n3647 = n213 & ~n2555 ;
  assign n3648 = ~n152 & n3647 ;
  assign n3639 = n1597 | n3177 ;
  assign n3640 = n3639 ^ n3029 ^ 1'b0 ;
  assign n3641 = n3341 ^ n2996 ^ 1'b0 ;
  assign n3642 = n378 | n3641 ;
  assign n3643 = n3642 ^ n1835 ^ 1'b0 ;
  assign n3644 = ~n3640 & n3643 ;
  assign n3645 = n3644 ^ n289 ^ 1'b0 ;
  assign n3646 = ( n1187 & n2923 ) | ( n1187 & ~n3645 ) | ( n2923 & ~n3645 ) ;
  assign n3649 = n3648 ^ n3646 ^ 1'b0 ;
  assign n3650 = n3638 | n3649 ;
  assign n3651 = n595 & ~n656 ;
  assign n3652 = ~n630 & n861 ;
  assign n3653 = ~n471 & n3652 ;
  assign n3654 = n3653 ^ n1837 ^ 1'b0 ;
  assign n3655 = n198 | n3654 ;
  assign n3656 = n315 | n2089 ;
  assign n3657 = n3656 ^ n3104 ^ 1'b0 ;
  assign n3658 = ~n2478 & n3657 ;
  assign n3659 = n1952 | n2284 ;
  assign n3660 = ~n3170 & n3659 ;
  assign n3661 = n3660 ^ n1026 ^ 1'b0 ;
  assign n3662 = n1821 ^ x68 ^ 1'b0 ;
  assign n3663 = ~n571 & n3662 ;
  assign n3664 = n315 & n3663 ;
  assign n3665 = n3664 ^ n642 ^ 1'b0 ;
  assign n3666 = n1131 ^ n662 ^ 1'b0 ;
  assign n3667 = n3666 ^ n1013 ^ n812 ;
  assign n3668 = n1556 & ~n2067 ;
  assign n3669 = n3667 & n3668 ;
  assign n3670 = n998 & ~n1329 ;
  assign n3671 = ~n891 & n3670 ;
  assign n3672 = ~n439 & n1663 ;
  assign n3673 = ~n877 & n2569 ;
  assign n3674 = n1663 | n1695 ;
  assign n3675 = n1325 & n1984 ;
  assign n3676 = n2729 ^ n1328 ^ 1'b0 ;
  assign n3677 = n2650 | n3676 ;
  assign n3678 = n506 & n2527 ;
  assign n3679 = n354 & n727 ;
  assign n3680 = n3679 ^ n1913 ^ 1'b0 ;
  assign n3691 = n194 & n912 ;
  assign n3686 = n972 ^ n753 ^ 1'b0 ;
  assign n3687 = x21 & n3686 ;
  assign n3685 = n851 | n1051 ;
  assign n3688 = n3687 ^ n3685 ^ 1'b0 ;
  assign n3681 = n2746 ^ n634 ^ 1'b0 ;
  assign n3682 = n2946 | n3681 ;
  assign n3683 = n3682 ^ n2755 ^ n594 ;
  assign n3684 = n1666 | n3683 ;
  assign n3689 = n3688 ^ n3684 ^ 1'b0 ;
  assign n3690 = ~n1841 & n3689 ;
  assign n3692 = n3691 ^ n3690 ^ 1'b0 ;
  assign n3693 = x87 & n3692 ;
  assign n3694 = n1841 & n3693 ;
  assign n3695 = n3694 ^ x8 ^ 1'b0 ;
  assign n3696 = ~n2972 & n3452 ;
  assign n3697 = n1268 ^ n1254 ^ 1'b0 ;
  assign n3698 = n3697 ^ n2484 ^ 1'b0 ;
  assign n3699 = n3698 ^ n250 ^ 1'b0 ;
  assign n3700 = n2847 | n3327 ;
  assign n3701 = n2229 ^ n1871 ^ 1'b0 ;
  assign n3702 = ~n1033 & n3701 ;
  assign n3703 = n3615 ^ n3027 ^ 1'b0 ;
  assign n3704 = n3702 & ~n3703 ;
  assign n3705 = n831 & n939 ;
  assign n3706 = ~n2201 & n3705 ;
  assign n3707 = n3706 ^ n1779 ^ 1'b0 ;
  assign n3708 = n880 ^ n501 ^ 1'b0 ;
  assign n3709 = n2357 ^ n1542 ^ 1'b0 ;
  assign n3710 = n3708 | n3709 ;
  assign n3711 = n1815 | n3710 ;
  assign n3712 = n2136 ^ n985 ^ 1'b0 ;
  assign n3713 = n1908 ^ x73 ^ 1'b0 ;
  assign n3714 = x75 | n3713 ;
  assign n3715 = ~n1107 & n3714 ;
  assign n3716 = n1800 & ~n2986 ;
  assign n3717 = n3400 | n3716 ;
  assign n3718 = ~n1226 & n3717 ;
  assign n3719 = n3343 ^ n922 ^ 1'b0 ;
  assign n3720 = n3719 ^ x106 ^ 1'b0 ;
  assign n3721 = ~n433 & n3720 ;
  assign n3722 = n148 & n1827 ;
  assign n3723 = n3722 ^ n2151 ^ 1'b0 ;
  assign n3724 = n2722 & n3094 ;
  assign n3725 = n3724 ^ x58 ^ 1'b0 ;
  assign n3726 = x12 | n240 ;
  assign n3727 = n277 & ~n638 ;
  assign n3728 = n3727 ^ n740 ^ 1'b0 ;
  assign n3729 = n1521 & ~n2345 ;
  assign n3730 = n481 & ~n1016 ;
  assign n3731 = x15 & ~n1154 ;
  assign n3732 = n2051 & n3731 ;
  assign n3733 = n1376 & n1414 ;
  assign n3734 = n2942 | n3733 ;
  assign n3735 = n165 & ~n669 ;
  assign n3736 = n2596 & n3735 ;
  assign n3737 = n830 & ~n1016 ;
  assign n3738 = n3737 ^ x109 ^ 1'b0 ;
  assign n3739 = n3736 | n3738 ;
  assign n3740 = n1627 & ~n1917 ;
  assign n3741 = n1020 & ~n1234 ;
  assign n3742 = n3741 ^ n1316 ^ 1'b0 ;
  assign n3743 = n1861 & ~n3742 ;
  assign n3744 = n1746 & n3743 ;
  assign n3745 = n2909 ^ n360 ^ 1'b0 ;
  assign n3746 = n1640 | n3745 ;
  assign n3747 = n3491 ^ n1080 ^ 1'b0 ;
  assign n3748 = ~n3746 & n3747 ;
  assign n3749 = n2859 ^ x110 ^ 1'b0 ;
  assign n3750 = x63 & n496 ;
  assign n3751 = ~n1854 & n3152 ;
  assign n3752 = n3751 ^ n3208 ^ 1'b0 ;
  assign n3753 = n3726 & ~n3752 ;
  assign n3754 = n3203 ^ n2839 ^ 1'b0 ;
  assign n3755 = n2107 | n3754 ;
  assign n3756 = n912 & ~n2859 ;
  assign n3757 = n3756 ^ n1905 ^ 1'b0 ;
  assign n3758 = x94 & n3757 ;
  assign n3759 = ~n1227 & n2948 ;
  assign n3760 = n245 | n390 ;
  assign n3761 = n2127 & ~n2480 ;
  assign n3762 = n3760 & n3761 ;
  assign n3763 = n2086 ^ n259 ^ 1'b0 ;
  assign n3764 = ~n1240 & n2409 ;
  assign n3765 = x72 & ~n3764 ;
  assign n3766 = ~n1451 & n3765 ;
  assign n3767 = ~n3765 & n3766 ;
  assign n3768 = n3172 | n3767 ;
  assign n3769 = n3172 & ~n3768 ;
  assign n3770 = n1597 & n2006 ;
  assign n3771 = n1716 & ~n3770 ;
  assign n3772 = n1959 & n3771 ;
  assign n3773 = n1010 & n3120 ;
  assign n3774 = x125 | n3199 ;
  assign n3775 = n975 | n2166 ;
  assign n3776 = x36 | n3775 ;
  assign n3777 = x6 & n1317 ;
  assign n3778 = ~n1193 & n3777 ;
  assign n3779 = n1105 | n2568 ;
  assign n3780 = n1864 & ~n3779 ;
  assign n3781 = n729 & n1209 ;
  assign n3782 = n1932 & n3781 ;
  assign n3783 = n2360 | n3782 ;
  assign n3784 = n3783 ^ n1358 ^ 1'b0 ;
  assign n3785 = n242 | n3784 ;
  assign n3786 = n2557 & n3785 ;
  assign n3787 = n2537 | n3786 ;
  assign n3788 = n1662 | n3787 ;
  assign n3789 = x110 ^ x17 ^ 1'b0 ;
  assign n3790 = n1380 & ~n1457 ;
  assign n3791 = n2944 | n3790 ;
  assign n3792 = ~n3789 & n3791 ;
  assign n3793 = n1262 ^ x66 ^ 1'b0 ;
  assign n3794 = n3060 ^ n1202 ^ 1'b0 ;
  assign n3795 = n2087 & ~n2101 ;
  assign n3796 = n258 | n3507 ;
  assign n3797 = n3728 | n3796 ;
  assign n3798 = n1240 ^ n205 ^ 1'b0 ;
  assign n3799 = n1374 | n3632 ;
  assign n3800 = n3798 | n3799 ;
  assign n3801 = n1681 & ~n2394 ;
  assign n3802 = n3801 ^ n616 ^ 1'b0 ;
  assign n3803 = n3401 ^ n1369 ^ 1'b0 ;
  assign n3804 = n1352 & ~n2981 ;
  assign n3809 = n1623 ^ n1086 ^ 1'b0 ;
  assign n3806 = n912 ^ n391 ^ 1'b0 ;
  assign n3807 = n988 | n3806 ;
  assign n3808 = n2238 | n3807 ;
  assign n3810 = n3809 ^ n3808 ^ 1'b0 ;
  assign n3811 = n2043 | n3810 ;
  assign n3812 = n3811 ^ n3023 ^ 1'b0 ;
  assign n3805 = n574 | n2962 ;
  assign n3813 = n3812 ^ n3805 ^ 1'b0 ;
  assign n3814 = n820 ^ n593 ^ 1'b0 ;
  assign n3815 = ~n753 & n3814 ;
  assign n3816 = n285 | n3815 ;
  assign n3817 = n1303 & ~n3816 ;
  assign n3818 = n3817 ^ n859 ^ 1'b0 ;
  assign n3819 = n1397 & ~n3417 ;
  assign n3820 = n1700 ^ x83 ^ 1'b0 ;
  assign n3821 = n3819 & n3820 ;
  assign n3822 = n507 | n2515 ;
  assign n3823 = n3822 ^ n1905 ^ 1'b0 ;
  assign n3824 = n1372 & ~n2763 ;
  assign n3825 = ~n3203 & n3824 ;
  assign n3826 = n1258 & n3825 ;
  assign n3827 = n3826 ^ n3350 ^ 1'b0 ;
  assign n3828 = n1564 & ~n3827 ;
  assign n3829 = n1613 & ~n3366 ;
  assign n3830 = x6 & n1530 ;
  assign n3831 = n315 & n3830 ;
  assign n3832 = n574 | n3199 ;
  assign n3833 = n3832 ^ n1208 ^ 1'b0 ;
  assign n3834 = n3833 ^ n1308 ^ 1'b0 ;
  assign n3835 = n1521 ^ x37 ^ 1'b0 ;
  assign n3836 = ~n1904 & n3835 ;
  assign n3837 = n2198 ^ n1321 ^ 1'b0 ;
  assign n3838 = ~n3267 & n3837 ;
  assign n3839 = n3453 | n3838 ;
  assign n3840 = n3839 ^ n169 ^ 1'b0 ;
  assign n3841 = n2980 ^ n667 ^ 1'b0 ;
  assign n3842 = ~n427 & n3841 ;
  assign n3843 = n2517 ^ n1903 ^ 1'b0 ;
  assign n3844 = ~n3842 & n3843 ;
  assign n3845 = n2643 ^ n2569 ^ 1'b0 ;
  assign n3846 = n1581 & n3845 ;
  assign n3847 = n3613 | n3846 ;
  assign n3851 = n673 | n2028 ;
  assign n3852 = n1810 & ~n3851 ;
  assign n3848 = ~n1059 & n2203 ;
  assign n3849 = n3848 ^ n2589 ^ 1'b0 ;
  assign n3850 = n2467 & ~n3849 ;
  assign n3853 = n3852 ^ n3850 ^ 1'b0 ;
  assign n3855 = n1329 & n1880 ;
  assign n3854 = ~n360 & n3754 ;
  assign n3856 = n3855 ^ n3854 ^ 1'b0 ;
  assign n3857 = n1892 ^ n845 ^ 1'b0 ;
  assign n3858 = n504 & ~n3857 ;
  assign n3859 = n3856 & ~n3858 ;
  assign n3860 = ( ~n837 & n2349 ) | ( ~n837 & n3859 ) | ( n2349 & n3859 ) ;
  assign n3861 = n3106 ^ n2090 ^ 1'b0 ;
  assign n3864 = n1829 & n3581 ;
  assign n3865 = n3864 ^ n2779 ^ 1'b0 ;
  assign n3862 = n1336 & n1980 ;
  assign n3863 = n3169 | n3862 ;
  assign n3866 = n3865 ^ n3863 ^ 1'b0 ;
  assign n3867 = n2915 ^ n2769 ^ 1'b0 ;
  assign n3868 = n1994 & ~n3867 ;
  assign n3871 = n828 | n3707 ;
  assign n3872 = n3871 ^ n1020 ^ 1'b0 ;
  assign n3869 = n173 | n2240 ;
  assign n3870 = n3869 ^ n287 ^ 1'b0 ;
  assign n3873 = n3872 ^ n3870 ^ 1'b0 ;
  assign n3874 = ( n177 & n407 ) | ( n177 & n1316 ) | ( n407 & n1316 ) ;
  assign n3875 = n3874 ^ n1420 ^ 1'b0 ;
  assign n3876 = n1434 ^ x119 ^ 1'b0 ;
  assign n3877 = n3876 ^ n478 ^ 1'b0 ;
  assign n3878 = n3292 ^ n2503 ^ n1939 ;
  assign n3879 = n1601 | n1832 ;
  assign n3880 = n3879 ^ n2930 ^ 1'b0 ;
  assign n3881 = ~n2782 & n3880 ;
  assign n3882 = ~n2482 & n3881 ;
  assign n3887 = n1477 & n3770 ;
  assign n3883 = ~n724 & n984 ;
  assign n3884 = n3883 ^ n1098 ^ 1'b0 ;
  assign n3885 = n3884 ^ n689 ^ 1'b0 ;
  assign n3886 = n1747 & ~n3885 ;
  assign n3888 = n3887 ^ n3886 ^ 1'b0 ;
  assign n3890 = n1829 & n2683 ;
  assign n3889 = n2971 ^ n2889 ^ n1833 ;
  assign n3891 = n3890 ^ n3889 ^ n430 ;
  assign n3892 = n1356 & n2271 ;
  assign n3893 = n3892 ^ n1918 ^ 1'b0 ;
  assign n3894 = ~n594 & n877 ;
  assign n3895 = n221 & ~n3894 ;
  assign n3896 = n3895 ^ n709 ^ 1'b0 ;
  assign n3897 = n1321 & n3896 ;
  assign n3898 = n450 | n489 ;
  assign n3899 = n1323 & n3898 ;
  assign n3900 = n3899 ^ x48 ^ 1'b0 ;
  assign n3901 = n3858 ^ n1829 ^ 1'b0 ;
  assign n3902 = n1147 & n3901 ;
  assign n3903 = n2623 ^ n1075 ^ 1'b0 ;
  assign n3904 = x66 | n3903 ;
  assign n3905 = n3544 & ~n3904 ;
  assign n3906 = n702 & n2021 ;
  assign n3907 = n3785 ^ n1243 ^ 1'b0 ;
  assign n3908 = ( n2330 & n2587 ) | ( n2330 & ~n3110 ) | ( n2587 & ~n3110 ) ;
  assign n3909 = x85 & n378 ;
  assign n3910 = ~n566 & n1955 ;
  assign n3911 = n3380 ^ n494 ^ 1'b0 ;
  assign n3912 = n324 | n600 ;
  assign n3913 = n324 & ~n3912 ;
  assign n3914 = n3756 & ~n3913 ;
  assign n3915 = n3911 & n3914 ;
  assign n3916 = n733 | n788 ;
  assign n3917 = n2263 ^ n1900 ^ n978 ;
  assign n3918 = n1728 ^ n1541 ^ 1'b0 ;
  assign n3919 = n1169 & n3918 ;
  assign n3920 = n837 ^ n809 ^ 1'b0 ;
  assign n3921 = n3919 & n3920 ;
  assign n3922 = n1713 & ~n3682 ;
  assign n3923 = n2306 & n2557 ;
  assign n3924 = n2582 | n3923 ;
  assign n3925 = n3924 ^ n1620 ^ 1'b0 ;
  assign n3926 = n2415 & n2923 ;
  assign n3927 = n3926 ^ n2739 ^ n2183 ;
  assign n3928 = n2892 ^ n2399 ^ 1'b0 ;
  assign n3929 = n1420 | n3928 ;
  assign n3930 = ~n484 & n3929 ;
  assign n3931 = n1635 & ~n3930 ;
  assign n3932 = n1394 ^ x59 ^ 1'b0 ;
  assign n3933 = n571 | n3932 ;
  assign n3934 = n3933 ^ n3689 ^ 1'b0 ;
  assign n3935 = n1693 ^ n1306 ^ 1'b0 ;
  assign n3936 = n2928 ^ n2091 ^ 1'b0 ;
  assign n3937 = ~n3935 & n3936 ;
  assign n3940 = n2024 ^ n439 ^ 1'b0 ;
  assign n3941 = n1883 & n3940 ;
  assign n3942 = n425 & n3941 ;
  assign n3943 = n3942 ^ n1695 ^ 1'b0 ;
  assign n3938 = n3548 ^ n3063 ^ 1'b0 ;
  assign n3939 = ~n1129 & n3938 ;
  assign n3944 = n3943 ^ n3939 ^ 1'b0 ;
  assign n3945 = n3818 ^ n1493 ^ 1'b0 ;
  assign n3946 = n3052 | n3945 ;
  assign n3947 = ( n200 & n557 ) | ( n200 & ~n2707 ) | ( n557 & ~n2707 ) ;
  assign n3948 = n3947 ^ n1329 ^ 1'b0 ;
  assign n3949 = ~n616 & n3784 ;
  assign n3951 = x20 & n2009 ;
  assign n3952 = n2840 & n3951 ;
  assign n3950 = n1935 | n2360 ;
  assign n3953 = n3952 ^ n3950 ^ 1'b0 ;
  assign n3954 = n1331 & ~n1348 ;
  assign n3955 = n3954 ^ n501 ^ 1'b0 ;
  assign n3957 = n1623 ^ n1517 ^ 1'b0 ;
  assign n3958 = n1005 & ~n3957 ;
  assign n3956 = n3544 ^ n1749 ^ 1'b0 ;
  assign n3959 = n3958 ^ n3956 ^ 1'b0 ;
  assign n3960 = n741 & ~n3959 ;
  assign n3961 = n3955 & n3960 ;
  assign n3962 = n3961 ^ n2314 ^ 1'b0 ;
  assign n3963 = n1129 ^ n464 ^ 1'b0 ;
  assign n3964 = n1035 & n3963 ;
  assign n3965 = n1226 ^ n830 ^ 1'b0 ;
  assign n3966 = ( ~n3583 & n3964 ) | ( ~n3583 & n3965 ) | ( n3964 & n3965 ) ;
  assign n3968 = n1412 ^ n811 ^ n516 ;
  assign n3967 = n880 & n1057 ;
  assign n3969 = n3968 ^ n3967 ^ n1443 ;
  assign n3970 = n2315 & n3969 ;
  assign n3971 = n920 ^ n387 ^ 1'b0 ;
  assign n3972 = ~n3929 & n3971 ;
  assign n3973 = ~n3070 & n3972 ;
  assign n3974 = n1654 & ~n3204 ;
  assign n3975 = n1222 & n3114 ;
  assign n3976 = n952 & n967 ;
  assign n3977 = n572 | n1561 ;
  assign n3978 = n1629 & n3179 ;
  assign n3980 = ~n776 & n788 ;
  assign n3981 = ~x84 & n3980 ;
  assign n3982 = n1129 ^ x104 ^ 1'b0 ;
  assign n3983 = n3981 | n3982 ;
  assign n3979 = n604 & ~n2107 ;
  assign n3984 = n3983 ^ n3979 ^ 1'b0 ;
  assign n3985 = ~n579 & n3984 ;
  assign n3986 = ~x105 & n418 ;
  assign n3987 = n3986 ^ x67 ^ 1'b0 ;
  assign n3988 = n1316 ^ x120 ^ 1'b0 ;
  assign n3989 = x36 & n3988 ;
  assign n3990 = ~n1941 & n3989 ;
  assign n3991 = n3990 ^ n1016 ^ 1'b0 ;
  assign n3992 = n1590 ^ n1414 ^ n642 ;
  assign n3993 = n3991 | n3992 ;
  assign n3994 = n3993 ^ n2591 ^ 1'b0 ;
  assign n3995 = n1842 ^ n689 ^ 1'b0 ;
  assign n3996 = n509 & n3995 ;
  assign n3997 = n1221 ^ n250 ^ 1'b0 ;
  assign n3998 = n3996 & n3997 ;
  assign n3999 = n3998 ^ n1023 ^ 1'b0 ;
  assign n4000 = n2309 | n3999 ;
  assign n4001 = n4000 ^ n2909 ^ 1'b0 ;
  assign n4002 = n2926 ^ n2440 ^ 1'b0 ;
  assign n4003 = n4002 ^ n2937 ^ 1'b0 ;
  assign n4004 = n3101 & ~n4003 ;
  assign n4005 = n4004 ^ x58 ^ 1'b0 ;
  assign n4006 = n2394 ^ x57 ^ 1'b0 ;
  assign n4007 = n2430 ^ n939 ^ x104 ;
  assign n4008 = n200 | n3177 ;
  assign n4009 = n4007 | n4008 ;
  assign n4010 = n4006 & n4009 ;
  assign n4011 = n4010 ^ n3484 ^ 1'b0 ;
  assign n4014 = n161 ^ x8 ^ 1'b0 ;
  assign n4012 = ~n696 & n1819 ;
  assign n4013 = ~n2289 & n4012 ;
  assign n4015 = n4014 ^ n4013 ^ 1'b0 ;
  assign n4016 = ~n3037 & n4015 ;
  assign n4024 = n693 ^ n672 ^ 1'b0 ;
  assign n4025 = n1983 & n4024 ;
  assign n4017 = n1947 & ~n2357 ;
  assign n4018 = ~n956 & n4017 ;
  assign n4019 = x114 & ~n1344 ;
  assign n4020 = ( n1525 & n3446 ) | ( n1525 & n4019 ) | ( n3446 & n4019 ) ;
  assign n4021 = n4020 ^ n3388 ^ 1'b0 ;
  assign n4022 = n4018 | n4021 ;
  assign n4023 = n2030 & ~n4022 ;
  assign n4026 = n4025 ^ n4023 ^ 1'b0 ;
  assign n4027 = n2678 & ~n4026 ;
  assign n4028 = n1635 & ~n3494 ;
  assign n4029 = ~n3419 & n3570 ;
  assign n4030 = n792 ^ x46 ^ 1'b0 ;
  assign n4031 = n1105 | n4030 ;
  assign n4032 = n4031 ^ x99 ^ 1'b0 ;
  assign n4033 = n939 & ~n1422 ;
  assign n4034 = ~n245 & n4033 ;
  assign n4035 = n3459 ^ n3401 ^ 1'b0 ;
  assign n4036 = ~n741 & n3196 ;
  assign n4037 = n4036 ^ n926 ^ 1'b0 ;
  assign n4038 = n824 & ~n4037 ;
  assign n4039 = n3101 ^ x53 ^ 1'b0 ;
  assign n4040 = n813 & n4039 ;
  assign n4041 = n1383 | n1989 ;
  assign n4042 = n4041 ^ n1228 ^ 1'b0 ;
  assign n4043 = n912 & n1351 ;
  assign n4044 = n2878 ^ n1270 ^ 1'b0 ;
  assign n4045 = n972 & n4044 ;
  assign n4046 = ~n2994 & n3012 ;
  assign n4047 = ~n4045 & n4046 ;
  assign n4048 = n131 & ~n811 ;
  assign n4049 = n1051 & n1756 ;
  assign n4050 = n3305 & n4049 ;
  assign n4051 = ~n189 & n608 ;
  assign n4052 = n3262 ^ n2125 ^ n893 ;
  assign n4053 = n4052 ^ n471 ^ 1'b0 ;
  assign n4054 = n4051 & n4053 ;
  assign n4058 = n1037 ^ x16 ^ 1'b0 ;
  assign n4059 = x10 & n4058 ;
  assign n4060 = ~n1723 & n4059 ;
  assign n4055 = n1204 & ~n1803 ;
  assign n4056 = n4055 ^ x22 ^ 1'b0 ;
  assign n4057 = n4056 ^ n2154 ^ 1'b0 ;
  assign n4061 = n4060 ^ n4057 ^ 1'b0 ;
  assign n4062 = n3450 ^ n741 ^ 1'b0 ;
  assign n4063 = n4062 ^ n3934 ^ 1'b0 ;
  assign n4064 = n2601 & n4063 ;
  assign n4065 = n481 & n1365 ;
  assign n4066 = n512 & ~n4065 ;
  assign n4067 = ~n3874 & n4066 ;
  assign n4068 = n2392 ^ n990 ^ 1'b0 ;
  assign n4069 = n4067 | n4068 ;
  assign n4070 = n2238 & n2573 ;
  assign n4071 = n2024 | n2947 ;
  assign n4072 = n1385 | n3819 ;
  assign n4073 = ~n3128 & n3785 ;
  assign n4074 = n4073 ^ n1737 ^ 1'b0 ;
  assign n4075 = ~n889 & n1658 ;
  assign n4076 = ~n595 & n4075 ;
  assign n4077 = n4076 ^ x14 ^ 1'b0 ;
  assign n4078 = n4077 ^ n3659 ^ n571 ;
  assign n4079 = n2456 ^ n339 ^ 1'b0 ;
  assign n4080 = n920 & ~n2151 ;
  assign n4081 = ~n2608 & n4080 ;
  assign n4082 = n518 | n2678 ;
  assign n4083 = n4082 ^ n2776 ^ 1'b0 ;
  assign n4084 = ~n806 & n3654 ;
  assign n4085 = n1552 ^ n1363 ^ 1'b0 ;
  assign n4086 = n1508 & ~n4085 ;
  assign n4087 = n4086 ^ n3651 ^ 1'b0 ;
  assign n4090 = n507 & ~n544 ;
  assign n4091 = n2946 & n4090 ;
  assign n4088 = n2115 & ~n2176 ;
  assign n4089 = n4088 ^ x39 ^ 1'b0 ;
  assign n4092 = n4091 ^ n4089 ^ 1'b0 ;
  assign n4093 = ~n3887 & n4092 ;
  assign n4094 = ~n2191 & n4032 ;
  assign n4095 = n380 & n4094 ;
  assign n4096 = n1474 ^ n294 ^ 1'b0 ;
  assign n4097 = n623 & ~n4096 ;
  assign n4098 = n4095 & n4097 ;
  assign n4099 = n4098 ^ n501 ^ 1'b0 ;
  assign n4100 = n4093 & n4099 ;
  assign n4105 = n474 | n1129 ;
  assign n4106 = n4105 ^ x82 ^ 1'b0 ;
  assign n4101 = n489 | n1586 ;
  assign n4102 = n4101 ^ n1823 ^ 1'b0 ;
  assign n4103 = n2966 ^ n1082 ^ 1'b0 ;
  assign n4104 = n4102 & ~n4103 ;
  assign n4107 = n4106 ^ n4104 ^ 1'b0 ;
  assign n4108 = n4096 ^ n3742 ^ 1'b0 ;
  assign n4109 = n632 & n4108 ;
  assign n4110 = n1046 & n2389 ;
  assign n4111 = n4110 ^ n2221 ^ n740 ;
  assign n4112 = n4111 ^ n3635 ^ 1'b0 ;
  assign n4113 = n266 & n2389 ;
  assign n4114 = n2705 | n4113 ;
  assign n4115 = n1319 | n3498 ;
  assign n4116 = n2208 | n2666 ;
  assign n4117 = n4116 ^ n1412 ^ 1'b0 ;
  assign n4118 = n2212 | n4117 ;
  assign n4119 = n1744 & ~n3290 ;
  assign n4120 = ~n3687 & n4119 ;
  assign n4121 = n632 ^ n427 ^ 1'b0 ;
  assign n4122 = n2003 | n4121 ;
  assign n4128 = n667 | n3031 ;
  assign n4123 = n2091 ^ n1470 ^ 1'b0 ;
  assign n4124 = ~n2868 & n4123 ;
  assign n4125 = n1994 & n2289 ;
  assign n4126 = ~n4124 & n4125 ;
  assign n4127 = n2079 & ~n4126 ;
  assign n4129 = n4128 ^ n4127 ^ 1'b0 ;
  assign n4130 = n1786 & n2109 ;
  assign n4131 = n4130 ^ n2722 ^ 1'b0 ;
  assign n4132 = n3818 & n4131 ;
  assign n4133 = n4132 ^ n1998 ^ 1'b0 ;
  assign n4134 = n629 ^ n571 ^ 1'b0 ;
  assign n4135 = n1335 | n4134 ;
  assign n4136 = n1800 ^ n1644 ^ 1'b0 ;
  assign n4137 = n806 | n2735 ;
  assign n4138 = n4136 & ~n4137 ;
  assign n4139 = n4138 ^ n1115 ^ 1'b0 ;
  assign n4140 = n2208 | n2962 ;
  assign n4141 = n4140 ^ n857 ^ 1'b0 ;
  assign n4142 = x25 & ~n2448 ;
  assign n4143 = n4142 ^ n1147 ^ 1'b0 ;
  assign n4144 = n2942 & n4143 ;
  assign n4145 = n813 & ~n2112 ;
  assign n4146 = n3862 & n4145 ;
  assign n4147 = n1537 & n2021 ;
  assign n4148 = n4146 | n4147 ;
  assign n4149 = n177 & n788 ;
  assign n4150 = n1329 & n4149 ;
  assign n4151 = n2355 ^ n1652 ^ 1'b0 ;
  assign n4152 = ~n1661 & n1747 ;
  assign n4153 = n3419 & n4152 ;
  assign n4154 = n3124 | n4153 ;
  assign n4155 = n4153 & ~n4154 ;
  assign n4156 = n1329 ^ n478 ^ 1'b0 ;
  assign n4157 = n1229 | n4156 ;
  assign n4158 = n4157 ^ n3046 ^ 1'b0 ;
  assign n4159 = n299 | n560 ;
  assign n4160 = x127 | n4159 ;
  assign n4161 = n427 | n1107 ;
  assign n4162 = n4160 | n4161 ;
  assign n4163 = n1982 | n4162 ;
  assign n4164 = n394 & n3049 ;
  assign n4165 = ~n4163 & n4164 ;
  assign n4166 = n2444 & ~n4165 ;
  assign n4167 = n4166 ^ n1349 ^ 1'b0 ;
  assign n4168 = n1498 ^ n1170 ^ 1'b0 ;
  assign n4169 = x123 & ~n4168 ;
  assign n4170 = n4169 ^ n2363 ^ 1'b0 ;
  assign n4171 = n852 ^ n571 ^ 1'b0 ;
  assign n4172 = n1808 & ~n4171 ;
  assign n4173 = n4172 ^ n2216 ^ 1'b0 ;
  assign n4174 = ~n1310 & n1415 ;
  assign n4175 = n1640 ^ n1147 ^ 1'b0 ;
  assign n4176 = n507 & ~n3091 ;
  assign n4177 = ~n4175 & n4176 ;
  assign n4178 = n207 | n4177 ;
  assign n4179 = n4174 | n4178 ;
  assign n4180 = n1247 & n4179 ;
  assign n4181 = ~n1281 & n4180 ;
  assign n4182 = n2488 ^ n2136 ^ 1'b0 ;
  assign n4183 = n4182 ^ n1606 ^ 1'b0 ;
  assign n4184 = n455 ^ n380 ^ 1'b0 ;
  assign n4185 = ~n830 & n4184 ;
  assign n4186 = n4185 ^ n2702 ^ 1'b0 ;
  assign n4187 = n2649 & ~n3812 ;
  assign n4188 = n4187 ^ n267 ^ 1'b0 ;
  assign n4189 = n1642 ^ n564 ^ x52 ;
  assign n4190 = ( ~n2230 & n3655 ) | ( ~n2230 & n3964 ) | ( n3655 & n3964 ) ;
  assign n4191 = ~n519 & n4190 ;
  assign n4192 = n2000 ^ n806 ^ 1'b0 ;
  assign n4193 = ~n3353 & n4192 ;
  assign n4195 = ~n200 & n965 ;
  assign n4196 = n1356 & ~n4195 ;
  assign n4197 = ( n1018 & n1193 ) | ( n1018 & n4196 ) | ( n1193 & n4196 ) ;
  assign n4194 = n1747 & n1948 ;
  assign n4198 = n4197 ^ n4194 ^ n2408 ;
  assign n4199 = n702 & n4198 ;
  assign n4200 = n406 & n4199 ;
  assign n4201 = ~n315 & n3763 ;
  assign n4202 = n4201 ^ n3175 ^ 1'b0 ;
  assign n4203 = ~n1084 & n1692 ;
  assign n4204 = n4203 ^ n1756 ^ 1'b0 ;
  assign n4205 = n3848 & n4204 ;
  assign n4206 = n853 ^ x112 ^ 1'b0 ;
  assign n4207 = n3531 & n4206 ;
  assign n4208 = ~n4205 & n4207 ;
  assign n4209 = n4020 | n4208 ;
  assign n4210 = n1887 & ~n4209 ;
  assign n4211 = n1199 & ~n1664 ;
  assign n4212 = ~n4196 & n4211 ;
  assign n4213 = n2677 ^ n1659 ^ 1'b0 ;
  assign n4214 = n3772 ^ n205 ^ 1'b0 ;
  assign n4215 = n3281 & n3795 ;
  assign n4216 = n1883 ^ x82 ^ 1'b0 ;
  assign n4217 = n463 & ~n876 ;
  assign n4218 = n3066 ^ n304 ^ 1'b0 ;
  assign n4219 = n2423 ^ n859 ^ 1'b0 ;
  assign n4220 = n3837 ^ n764 ^ 1'b0 ;
  assign n4221 = ~n1279 & n4220 ;
  assign n4222 = n3354 & n4221 ;
  assign n4223 = n414 ^ n216 ^ 1'b0 ;
  assign n4224 = n163 & ~n4223 ;
  assign n4225 = n2776 ^ n1579 ^ 1'b0 ;
  assign n4226 = n4224 & ~n4225 ;
  assign n4227 = n4226 ^ n1554 ^ 1'b0 ;
  assign n4236 = n1247 ^ n908 ^ 1'b0 ;
  assign n4237 = n262 | n459 ;
  assign n4238 = n1112 & ~n4237 ;
  assign n4239 = x58 | n4238 ;
  assign n4240 = n4236 & ~n4239 ;
  assign n4241 = ~n1345 & n4240 ;
  assign n4228 = n3937 ^ n3477 ^ 1'b0 ;
  assign n4232 = n289 ^ x121 ^ 1'b0 ;
  assign n4229 = n918 ^ n914 ^ 1'b0 ;
  assign n4230 = n415 & ~n4229 ;
  assign n4231 = ~n571 & n4230 ;
  assign n4233 = n4232 ^ n4231 ^ 1'b0 ;
  assign n4234 = n4233 ^ n2715 ^ 1'b0 ;
  assign n4235 = ~n4228 & n4234 ;
  assign n4242 = n4241 ^ n4235 ^ 1'b0 ;
  assign n4243 = n246 & ~n2789 ;
  assign n4244 = n4243 ^ n3986 ^ 1'b0 ;
  assign n4245 = ~n1187 & n2642 ;
  assign n4246 = n2847 ^ n2306 ^ 1'b0 ;
  assign n4247 = n2140 | n4246 ;
  assign n4248 = n1833 ^ n784 ^ x4 ;
  assign n4249 = x95 & ~n2426 ;
  assign n4250 = n725 & n2198 ;
  assign n4251 = n4250 ^ n3880 ^ 1'b0 ;
  assign n4252 = n3764 ^ n3279 ^ 1'b0 ;
  assign n4253 = ~n1443 & n1788 ;
  assign n4254 = n2198 ^ x94 ^ 1'b0 ;
  assign n4255 = n4254 ^ n620 ^ 1'b0 ;
  assign n4256 = n2075 & n4255 ;
  assign n4257 = x92 & ~n2181 ;
  assign n4258 = n3537 & n4257 ;
  assign n4259 = n4258 ^ n801 ^ 1'b0 ;
  assign n4260 = ~n292 & n3400 ;
  assign n4261 = n2669 & n4260 ;
  assign n4262 = n1065 | n1171 ;
  assign n4263 = n4262 ^ n1835 ^ 1'b0 ;
  assign n4264 = n4263 ^ n847 ^ 1'b0 ;
  assign n4265 = ~n1729 & n4264 ;
  assign n4266 = n805 | n1479 ;
  assign n4267 = n4266 ^ n3469 ^ 1'b0 ;
  assign n4268 = n3778 | n4267 ;
  assign n4269 = n722 & n2023 ;
  assign n4270 = ~n1864 & n2355 ;
  assign n4271 = n4270 ^ n1758 ^ 1'b0 ;
  assign n4272 = n3925 & ~n4271 ;
  assign n4273 = x69 & ~n1741 ;
  assign n4274 = ~n1157 & n4273 ;
  assign n4275 = n290 & ~n4274 ;
  assign n4276 = n4275 ^ n2440 ^ 1'b0 ;
  assign n4277 = n4276 ^ x82 ^ 1'b0 ;
  assign n4278 = n1327 & n4277 ;
  assign n4279 = n4278 ^ n4072 ^ 1'b0 ;
  assign n4280 = n200 | n1895 ;
  assign n4281 = n4031 | n4280 ;
  assign n4282 = n4281 ^ n571 ^ 1'b0 ;
  assign n4283 = n3007 ^ n2503 ^ 1'b0 ;
  assign n4284 = ~n1393 & n4283 ;
  assign n4286 = n203 ^ n137 ^ 1'b0 ;
  assign n4287 = ~n3107 & n4286 ;
  assign n4285 = n373 & n2062 ;
  assign n4288 = n4287 ^ n4285 ^ 1'b0 ;
  assign n4289 = x103 & ~n2283 ;
  assign n4290 = n698 & n1270 ;
  assign n4291 = ~n3503 & n4290 ;
  assign n4292 = n2818 | n4291 ;
  assign n4293 = n4289 & ~n4292 ;
  assign n4294 = ~n1167 & n2154 ;
  assign n4295 = n771 ^ n254 ^ 1'b0 ;
  assign n4296 = n444 | n4295 ;
  assign n4297 = x13 & ~n4296 ;
  assign n4298 = n539 & n4297 ;
  assign n4299 = n4298 ^ n3279 ^ 1'b0 ;
  assign n4300 = n1996 | n4299 ;
  assign n4301 = n1779 | n2469 ;
  assign n4302 = n1399 & n2257 ;
  assign n4303 = ~n1552 & n4302 ;
  assign n4304 = n4303 ^ n4148 ^ 1'b0 ;
  assign n4305 = n3391 ^ n2255 ^ 1'b0 ;
  assign n4306 = n1260 | n4305 ;
  assign n4307 = n2627 ^ n972 ^ 1'b0 ;
  assign n4308 = n485 | n3579 ;
  assign n4309 = n4308 ^ n3453 ^ 1'b0 ;
  assign n4310 = n4307 & ~n4309 ;
  assign n4311 = n1578 & ~n3124 ;
  assign n4312 = n4311 ^ n2383 ^ 1'b0 ;
  assign n4313 = x40 & n788 ;
  assign n4314 = n1436 ^ n1315 ^ 1'b0 ;
  assign n4315 = n4314 ^ n207 ^ 1'b0 ;
  assign n4316 = n1118 ^ x126 ^ 1'b0 ;
  assign n4317 = n2186 | n4316 ;
  assign n4318 = n3746 & ~n4317 ;
  assign n4319 = n2779 ^ n683 ^ 1'b0 ;
  assign n4320 = n742 | n4319 ;
  assign n4321 = n4320 ^ n709 ^ 1'b0 ;
  assign n4322 = n3567 ^ n1062 ^ 1'b0 ;
  assign n4323 = n1833 & ~n2743 ;
  assign n4326 = n2190 ^ n702 ^ 1'b0 ;
  assign n4324 = n1552 ^ n811 ^ 1'b0 ;
  assign n4325 = n2944 & ~n4324 ;
  assign n4327 = n4326 ^ n4325 ^ 1'b0 ;
  assign n4328 = ~n980 & n4327 ;
  assign n4329 = x7 & x122 ;
  assign n4330 = n4329 ^ n983 ^ 1'b0 ;
  assign n4331 = n1498 ^ n1253 ^ 1'b0 ;
  assign n4332 = ~n1513 & n4331 ;
  assign n4333 = ~x46 & n4332 ;
  assign n4334 = n2716 | n4333 ;
  assign n4335 = n300 | n2967 ;
  assign n4336 = n4335 ^ n3155 ^ 1'b0 ;
  assign n4337 = n2273 | n2734 ;
  assign n4338 = n2770 ^ n812 ^ 1'b0 ;
  assign n4339 = n512 & ~n3888 ;
  assign n4340 = n2439 ^ n1848 ^ 1'b0 ;
  assign n4341 = n1502 & n2155 ;
  assign n4342 = n877 ^ n134 ^ 1'b0 ;
  assign n4343 = n962 & ~n4342 ;
  assign n4344 = ~n4341 & n4343 ;
  assign n4345 = n3494 & n3874 ;
  assign n4346 = ( ~n775 & n955 ) | ( ~n775 & n2053 ) | ( n955 & n2053 ) ;
  assign n4347 = n1498 & n4346 ;
  assign n4348 = n3502 | n4347 ;
  assign n4349 = n3072 | n4348 ;
  assign n4350 = n2733 ^ n2426 ^ 1'b0 ;
  assign n4351 = n3134 ^ n896 ^ n731 ;
  assign n4352 = n1048 | n4351 ;
  assign n4353 = n4352 ^ x90 ^ 1'b0 ;
  assign n4354 = ~n414 & n2404 ;
  assign n4355 = n616 & ~n3032 ;
  assign n4356 = n579 & ~n1086 ;
  assign n4357 = n3805 ^ n1891 ^ 1'b0 ;
  assign n4358 = n336 & n620 ;
  assign n4359 = ~n1595 & n4358 ;
  assign n4360 = n4359 ^ n825 ^ 1'b0 ;
  assign n4361 = n4357 | n4360 ;
  assign n4363 = x111 & ~n504 ;
  assign n4362 = n330 & n2423 ;
  assign n4364 = n4363 ^ n4362 ^ 1'b0 ;
  assign n4365 = n1909 & n3721 ;
  assign n4366 = n391 & n4365 ;
  assign n4367 = n741 | n3247 ;
  assign n4368 = n4367 ^ n2086 ^ 1'b0 ;
  assign n4370 = n703 & ~n1477 ;
  assign n4369 = n2643 | n3169 ;
  assign n4371 = n4370 ^ n4369 ^ 1'b0 ;
  assign n4372 = n4371 ^ n3719 ^ 1'b0 ;
  assign n4373 = x72 & ~n2838 ;
  assign n4374 = n2718 ^ n830 ^ 1'b0 ;
  assign n4375 = ~n4371 & n4374 ;
  assign n4376 = n4343 ^ n359 ^ 1'b0 ;
  assign n4377 = x91 & ~n336 ;
  assign n4378 = n192 & n381 ;
  assign n4379 = ~n1868 & n4378 ;
  assign n4380 = n3762 & n4379 ;
  assign n4381 = n2618 & ~n4380 ;
  assign n4382 = ~n876 & n4381 ;
  assign n4383 = n4382 ^ n2915 ^ 1'b0 ;
  assign n4384 = x45 & n4383 ;
  assign n4385 = n2925 ^ n880 ^ 1'b0 ;
  assign n4386 = n156 & n4385 ;
  assign n4387 = ~n245 & n4386 ;
  assign n4388 = n2523 & ~n4387 ;
  assign n4389 = n2673 ^ n516 ^ 1'b0 ;
  assign n4390 = ~n3917 & n4389 ;
  assign n4391 = n3212 ^ x97 ^ 1'b0 ;
  assign n4392 = n425 ^ n230 ^ 1'b0 ;
  assign n4393 = x4 & n4392 ;
  assign n4394 = n4180 ^ n3153 ^ 1'b0 ;
  assign n4395 = n4393 & n4394 ;
  assign n4396 = n1636 ^ n707 ^ 1'b0 ;
  assign n4397 = n4395 & ~n4396 ;
  assign n4398 = n1728 | n2079 ;
  assign n4399 = n1341 ^ n508 ^ 1'b0 ;
  assign n4400 = n491 & n4399 ;
  assign n4401 = n2925 & n4400 ;
  assign n4402 = n4401 ^ n2134 ^ 1'b0 ;
  assign n4403 = ~n1265 & n4402 ;
  assign n4404 = n4403 ^ n3070 ^ 1'b0 ;
  assign n4405 = n2376 | n3642 ;
  assign n4406 = n4274 & ~n4405 ;
  assign n4407 = n3120 & ~n4406 ;
  assign n4408 = n4404 & n4407 ;
  assign n4409 = n4408 ^ n2578 ^ 1'b0 ;
  assign n4410 = n2385 & ~n4409 ;
  assign n4411 = n980 & ~n2776 ;
  assign n4412 = n1162 ^ n590 ^ 1'b0 ;
  assign n4413 = n4411 & ~n4412 ;
  assign n4414 = n3784 ^ n2201 ^ 1'b0 ;
  assign n4415 = ~n2635 & n4414 ;
  assign n4416 = n1880 & ~n4319 ;
  assign n4417 = n338 & n1599 ;
  assign n4418 = ~n3398 & n4417 ;
  assign n4419 = n4096 & n4418 ;
  assign n4420 = n1587 & n3790 ;
  assign n4421 = n4420 ^ n770 ^ 1'b0 ;
  assign n4422 = n1316 & n2345 ;
  assign n4423 = ~n4421 & n4422 ;
  assign n4424 = n4423 ^ n1329 ^ 1'b0 ;
  assign n4425 = n2982 | n4424 ;
  assign n4426 = n1710 & ~n2200 ;
  assign n4427 = n4426 ^ n1985 ^ 1'b0 ;
  assign n4428 = n836 | n4045 ;
  assign n4429 = n4427 & n4428 ;
  assign n4430 = n2279 ^ n1270 ^ 1'b0 ;
  assign n4431 = n4175 ^ n1467 ^ 1'b0 ;
  assign n4432 = n4430 & ~n4431 ;
  assign n4433 = n3189 & n4432 ;
  assign n4434 = n2967 ^ n2367 ^ n509 ;
  assign n4435 = n3893 ^ n3585 ^ 1'b0 ;
  assign n4436 = n652 & ~n4435 ;
  assign n4437 = n1808 ^ n371 ^ 1'b0 ;
  assign n4438 = n3503 & ~n4437 ;
  assign n4442 = n2028 ^ n365 ^ 1'b0 ;
  assign n4443 = n2278 | n4442 ;
  assign n4439 = n237 & ~n830 ;
  assign n4440 = n4439 ^ n1049 ^ 1'b0 ;
  assign n4441 = n1601 & n4440 ;
  assign n4444 = n4443 ^ n4441 ^ 1'b0 ;
  assign n4445 = n2442 ^ n2085 ^ 1'b0 ;
  assign n4446 = n155 | n1680 ;
  assign n4447 = n1968 | n4446 ;
  assign n4448 = n2602 & n4447 ;
  assign n4461 = n756 & n3027 ;
  assign n4449 = n4135 ^ n1400 ^ 1'b0 ;
  assign n4450 = n324 | n1161 ;
  assign n4452 = n335 & n537 ;
  assign n4453 = n277 & n739 ;
  assign n4454 = n4452 & n4453 ;
  assign n4451 = n788 & ~n1201 ;
  assign n4455 = n4454 ^ n4451 ^ 1'b0 ;
  assign n4456 = n4455 ^ n281 ^ 1'b0 ;
  assign n4457 = ~n4450 & n4456 ;
  assign n4458 = n4449 & n4457 ;
  assign n4459 = n1335 | n3589 ;
  assign n4460 = n4458 | n4459 ;
  assign n4462 = n4461 ^ n4460 ^ 1'b0 ;
  assign n4463 = x85 & n3558 ;
  assign n4464 = n4463 ^ n1875 ^ 1'b0 ;
  assign n4465 = n1856 ^ n1816 ^ 1'b0 ;
  assign n4466 = n503 ^ n290 ^ 1'b0 ;
  assign n4467 = ~n2325 & n4466 ;
  assign n4468 = ~n2653 & n4467 ;
  assign n4469 = n4468 ^ n2039 ^ 1'b0 ;
  assign n4470 = n3707 | n4469 ;
  assign n4471 = n4470 ^ n435 ^ 1'b0 ;
  assign n4472 = n2694 ^ x120 ^ 1'b0 ;
  assign n4473 = n1035 & ~n1201 ;
  assign n4474 = n4473 ^ x74 ^ 1'b0 ;
  assign n4475 = n1228 | n4474 ;
  assign n4476 = n4475 ^ n3935 ^ 1'b0 ;
  assign n4477 = n4472 & ~n4476 ;
  assign n4478 = n4477 ^ n666 ^ 1'b0 ;
  assign n4479 = n2019 & ~n4478 ;
  assign n4480 = ~n2399 & n4479 ;
  assign n4481 = n1868 | n3267 ;
  assign n4482 = n3715 & ~n4481 ;
  assign n4483 = x105 & ~n2486 ;
  assign n4484 = ~n3919 & n4483 ;
  assign n4485 = n3110 | n4484 ;
  assign n4486 = x1 & ~n1846 ;
  assign n4487 = n1510 & ~n2013 ;
  assign n4488 = n4487 ^ n3965 ^ n753 ;
  assign n4489 = n1025 ^ n307 ^ 1'b0 ;
  assign n4490 = n4489 ^ x54 ^ 1'b0 ;
  assign n4491 = n1832 | n4490 ;
  assign n4492 = n4488 | n4491 ;
  assign n4493 = n4492 ^ n4077 ^ n806 ;
  assign n4495 = n1800 | n2852 ;
  assign n4496 = n1035 | n4495 ;
  assign n4497 = n4496 ^ x96 ^ 1'b0 ;
  assign n4494 = n380 ^ x89 ^ 1'b0 ;
  assign n4498 = n4497 ^ n4494 ^ 1'b0 ;
  assign n4499 = n233 & n4498 ;
  assign n4500 = n3784 ^ n231 ^ 1'b0 ;
  assign n4501 = ~n3636 & n4500 ;
  assign n4502 = n3341 ^ n1107 ^ n477 ;
  assign n4503 = n4502 ^ n851 ^ 1'b0 ;
  assign n4504 = x16 & ~n2871 ;
  assign n4505 = n4504 ^ n1918 ^ 1'b0 ;
  assign n4506 = n2924 | n4505 ;
  assign n4507 = n614 | n2257 ;
  assign n4508 = n560 | n1028 ;
  assign n4509 = n4508 ^ n1948 ^ 1'b0 ;
  assign n4510 = n229 & n387 ;
  assign n4511 = n4510 ^ x11 ^ 1'b0 ;
  assign n4512 = ~n296 & n1154 ;
  assign n4513 = n4511 & n4512 ;
  assign n4514 = n1055 | n4513 ;
  assign n4515 = x26 | n4514 ;
  assign n4516 = n4515 ^ n3322 ^ 1'b0 ;
  assign n4517 = n4509 & n4516 ;
  assign n4518 = n2179 ^ n1008 ^ x78 ;
  assign n4519 = x41 & ~n4518 ;
  assign n4520 = n2148 & n4519 ;
  assign n4521 = n1636 ^ x91 ^ 1'b0 ;
  assign n4522 = n3158 | n4521 ;
  assign n4523 = n4522 ^ n533 ^ 1'b0 ;
  assign n4524 = n3396 ^ n1178 ^ 1'b0 ;
  assign n4525 = ( n2062 & ~n4016 ) | ( n2062 & n4524 ) | ( ~n4016 & n4524 ) ;
  assign n4526 = ~n2868 & n4525 ;
  assign n4527 = n4526 ^ n491 ^ 1'b0 ;
  assign n4528 = n507 & n2355 ;
  assign n4529 = n283 ^ x60 ^ 1'b0 ;
  assign n4530 = ~n960 & n4529 ;
  assign n4531 = n4530 ^ n439 ^ 1'b0 ;
  assign n4532 = n4528 & n4531 ;
  assign n4533 = x108 & n863 ;
  assign n4534 = ~x108 & n4533 ;
  assign n4535 = x87 & n1316 ;
  assign n4536 = ~x87 & n4535 ;
  assign n4537 = ~x106 & x114 ;
  assign n4538 = ~x114 & n4537 ;
  assign n4539 = ~n529 & n4538 ;
  assign n4540 = n195 & ~n4539 ;
  assign n4541 = n4539 & n4540 ;
  assign n4542 = n4536 | n4541 ;
  assign n4543 = n4536 & ~n4542 ;
  assign n4544 = ~n2363 & n4543 ;
  assign n4545 = n4534 & n4544 ;
  assign n4546 = n4314 ^ n634 ^ 1'b0 ;
  assign n4547 = n4545 & n4546 ;
  assign n4548 = n1758 & n4547 ;
  assign n4549 = n4548 ^ n3887 ^ 1'b0 ;
  assign n4550 = n272 | n1842 ;
  assign n4551 = n608 & n1361 ;
  assign n4552 = ~n747 & n1177 ;
  assign n4553 = ~n4551 & n4552 ;
  assign n4557 = n822 ^ n340 ^ 1'b0 ;
  assign n4556 = x125 | n1532 ;
  assign n4554 = ~x100 & n1655 ;
  assign n4555 = n1574 & n4554 ;
  assign n4558 = n4557 ^ n4556 ^ n4555 ;
  assign n4559 = n1395 ^ n507 ^ 1'b0 ;
  assign n4560 = n4559 ^ n451 ^ 1'b0 ;
  assign n4561 = n2049 & n3166 ;
  assign n4562 = n262 & ~n3196 ;
  assign n4563 = n1147 & n4562 ;
  assign n4564 = n4563 ^ n3654 ^ 1'b0 ;
  assign n4565 = n2667 & ~n4194 ;
  assign n4566 = n788 & ~n4565 ;
  assign n4567 = ~n1056 & n1341 ;
  assign n4568 = ~n381 & n2188 ;
  assign n4569 = n233 & n4205 ;
  assign n4570 = n3707 ^ n669 ^ 1'b0 ;
  assign n4571 = n259 | n1749 ;
  assign n4572 = n4418 & ~n4571 ;
  assign n4573 = n1183 | n2604 ;
  assign n4574 = n3425 & n4573 ;
  assign n4578 = ~n1189 & n2923 ;
  assign n4575 = n4195 ^ n1267 ^ 1'b0 ;
  assign n4576 = n1230 & ~n4575 ;
  assign n4577 = n3436 & n4576 ;
  assign n4579 = n4578 ^ n4577 ^ 1'b0 ;
  assign n4580 = x83 | n2836 ;
  assign n4583 = n740 ^ n728 ^ 1'b0 ;
  assign n4584 = x97 & ~n4583 ;
  assign n4581 = n647 & ~n1781 ;
  assign n4582 = n4581 ^ n1851 ^ 1'b0 ;
  assign n4585 = n4584 ^ n4582 ^ 1'b0 ;
  assign n4586 = n1075 ^ x40 ^ 1'b0 ;
  assign n4587 = ~x86 & n2843 ;
  assign n4588 = n1477 & ~n4587 ;
  assign n4589 = n4588 ^ n2146 ^ 1'b0 ;
  assign n4590 = n432 ^ n220 ^ 1'b0 ;
  assign n4591 = n998 & ~n2709 ;
  assign n4592 = ~n4590 & n4591 ;
  assign n4594 = n1534 & ~n2840 ;
  assign n4595 = n922 & n4594 ;
  assign n4596 = n4595 ^ x115 ^ 1'b0 ;
  assign n4597 = n4240 | n4596 ;
  assign n4593 = ~n854 & n2906 ;
  assign n4598 = n4597 ^ n4593 ^ 1'b0 ;
  assign n4599 = n1808 & n1819 ;
  assign n4600 = n4599 ^ n1480 ^ 1'b0 ;
  assign n4601 = n4600 ^ n3392 ^ 1'b0 ;
  assign n4602 = n2882 & ~n4601 ;
  assign n4603 = n400 & n3025 ;
  assign n4604 = n1455 | n1552 ;
  assign n4605 = n4487 | n4604 ;
  assign n4606 = n1279 | n3989 ;
  assign n4607 = x46 & ~n764 ;
  assign n4608 = n4607 ^ n1188 ^ 1'b0 ;
  assign n4609 = n1973 & ~n4608 ;
  assign n4610 = ~n4606 & n4609 ;
  assign n4611 = n2345 & ~n2385 ;
  assign n4612 = n1937 ^ n1508 ^ 1'b0 ;
  assign n4613 = n1342 ^ n1228 ^ 1'b0 ;
  assign n4614 = n375 & n3931 ;
  assign n4615 = n4614 ^ n1365 ^ 1'b0 ;
  assign n4616 = n1355 & n3425 ;
  assign n4617 = n4025 ^ n880 ^ 1'b0 ;
  assign n4618 = n4617 ^ n3112 ^ 1'b0 ;
  assign n4619 = n1240 & n2649 ;
  assign n4620 = n1017 ^ n446 ^ 1'b0 ;
  assign n4621 = n1002 | n4620 ;
  assign n4622 = n492 & ~n4621 ;
  assign n4623 = n484 & n4622 ;
  assign n4624 = n246 & ~n4623 ;
  assign n4625 = n4624 ^ n1030 ^ 1'b0 ;
  assign n4626 = n4625 ^ n775 ^ 1'b0 ;
  assign n4627 = n1456 & n4626 ;
  assign n4628 = n4627 ^ n1109 ^ 1'b0 ;
  assign n4629 = n1457 ^ x47 ^ 1'b0 ;
  assign n4630 = n1381 & n4629 ;
  assign n4631 = n4630 ^ n3450 ^ n1046 ;
  assign n4632 = n2227 | n4457 ;
  assign n4634 = n542 & ~n2416 ;
  assign n4635 = n4634 ^ n1457 ^ 1'b0 ;
  assign n4633 = x116 & ~n753 ;
  assign n4636 = n4635 ^ n4633 ^ 1'b0 ;
  assign n4638 = n1961 ^ n581 ^ 1'b0 ;
  assign n4637 = n1784 | n2833 ;
  assign n4639 = n4638 ^ n4637 ^ 1'b0 ;
  assign n4640 = n468 & n1428 ;
  assign n4641 = n161 & ~n1126 ;
  assign n4642 = n2035 ^ n1651 ^ 1'b0 ;
  assign n4643 = n4034 & ~n4642 ;
  assign n4644 = ~n4641 & n4643 ;
  assign n4645 = ~n4640 & n4644 ;
  assign n4646 = n624 | n4645 ;
  assign n4647 = n161 | n4646 ;
  assign n4648 = n1177 | n1395 ;
  assign n4649 = x12 & n1947 ;
  assign n4650 = ~n1508 & n4649 ;
  assign n4651 = n1126 | n1527 ;
  assign n4652 = n4650 & ~n4651 ;
  assign n4653 = n4652 ^ n1646 ^ 1'b0 ;
  assign n4654 = ~n909 & n4653 ;
  assign n4655 = n1170 & ~n1578 ;
  assign n4656 = n3179 | n4655 ;
  assign n4657 = n2948 ^ n2745 ^ 1'b0 ;
  assign n4658 = n385 | n564 ;
  assign n4659 = n4658 ^ n1868 ^ 1'b0 ;
  assign n4660 = ~n3267 & n4659 ;
  assign n4661 = ~n2710 & n3123 ;
  assign n4662 = n992 & ~n1561 ;
  assign n4663 = n143 ^ x22 ^ 1'b0 ;
  assign n4664 = ~n1406 & n4663 ;
  assign n4665 = ~n1234 & n2738 ;
  assign n4666 = ~n4664 & n4665 ;
  assign n4667 = n630 | n4666 ;
  assign n4668 = n4667 ^ n2526 ^ 1'b0 ;
  assign n4669 = n2859 ^ x26 ^ 1'b0 ;
  assign n4670 = n904 ^ n153 ^ 1'b0 ;
  assign n4671 = ~n1186 & n4670 ;
  assign n4672 = n797 ^ n279 ^ 1'b0 ;
  assign n4673 = n4671 & ~n4672 ;
  assign n4674 = n981 & n2399 ;
  assign n4675 = n2866 ^ n1702 ^ 1'b0 ;
  assign n4676 = n4674 & n4675 ;
  assign n4677 = ( ~n1776 & n1812 ) | ( ~n1776 & n4676 ) | ( n1812 & n4676 ) ;
  assign n4678 = n896 | n1061 ;
  assign n4679 = n1950 & ~n4678 ;
  assign n4680 = n700 | n4679 ;
  assign n4681 = n3880 | n4680 ;
  assign n4682 = x99 & n4681 ;
  assign n4683 = n1102 & n4682 ;
  assign n4684 = n3217 ^ x72 ^ 1'b0 ;
  assign n4685 = ~n3563 & n4684 ;
  assign n4686 = n2037 | n2632 ;
  assign n4687 = n4214 | n4686 ;
  assign n4688 = n1623 ^ x114 ^ 1'b0 ;
  assign n4689 = n1461 | n4688 ;
  assign n4690 = n3407 ^ n1354 ^ 1'b0 ;
  assign n4691 = n3651 ^ n867 ^ 1'b0 ;
  assign n4692 = n1732 & ~n2023 ;
  assign n4693 = n863 & ~n1080 ;
  assign n4697 = n825 ^ n131 ^ 1'b0 ;
  assign n4694 = n4454 ^ n2448 ^ 1'b0 ;
  assign n4695 = n1601 & n2710 ;
  assign n4696 = n4694 & n4695 ;
  assign n4698 = n4697 ^ n4696 ^ 1'b0 ;
  assign n4699 = n3644 & n4698 ;
  assign n4700 = ~n2709 & n3245 ;
  assign n4701 = n2014 & n4700 ;
  assign n4702 = n2732 | n4701 ;
  assign n4703 = n542 | n4702 ;
  assign n4704 = n4346 & n4448 ;
  assign n4705 = n2855 & n4704 ;
  assign n4706 = n245 | n4430 ;
  assign n4707 = n1262 ^ n895 ^ 1'b0 ;
  assign n4708 = ~n1483 & n2212 ;
  assign n4709 = n1737 & ~n3195 ;
  assign n4710 = n4709 ^ n4289 ^ 1'b0 ;
  assign n4711 = n4332 & ~n4710 ;
  assign n4712 = n181 & ~n770 ;
  assign n4713 = n4712 ^ n2230 ^ 1'b0 ;
  assign n4714 = n1456 ^ n1325 ^ 1'b0 ;
  assign n4715 = n3086 & n4714 ;
  assign n4716 = n339 & n4715 ;
  assign n4717 = ~n4713 & n4716 ;
  assign n4718 = n4717 ^ n4146 ^ 1'b0 ;
  assign n4719 = n1759 ^ n163 ^ 1'b0 ;
  assign n4720 = ~n3587 & n4719 ;
  assign n4722 = n584 | n2301 ;
  assign n4723 = n4722 ^ x9 ^ 1'b0 ;
  assign n4721 = n2171 ^ n492 ^ 1'b0 ;
  assign n4724 = n4723 ^ n4721 ^ 1'b0 ;
  assign n4725 = n954 & ~n4282 ;
  assign n4726 = ~n4724 & n4725 ;
  assign n4727 = n227 | n558 ;
  assign n4728 = n131 | n4727 ;
  assign n4729 = n4623 ^ n3584 ^ 1'b0 ;
  assign n4730 = n4729 ^ n3027 ^ 1'b0 ;
  assign n4732 = n950 | n3107 ;
  assign n4733 = n3107 & ~n4732 ;
  assign n4731 = ~n1749 & n3108 ;
  assign n4734 = n4733 ^ n4731 ^ n408 ;
  assign n4735 = n3589 & n4523 ;
  assign n4736 = x57 | n2344 ;
  assign n4737 = n1693 & n2293 ;
  assign n4738 = n4737 ^ n131 ^ 1'b0 ;
  assign n4739 = n2831 ^ n1216 ^ 1'b0 ;
  assign n4740 = n3654 | n4739 ;
  assign n4741 = n4740 ^ n1186 ^ 1'b0 ;
  assign n4742 = ~n4738 & n4741 ;
  assign n4743 = n3276 & n4009 ;
  assign n4744 = n1153 ^ n590 ^ 1'b0 ;
  assign n4745 = n1201 & n4744 ;
  assign n4746 = n776 ^ n227 ^ 1'b0 ;
  assign n4747 = n665 | n4746 ;
  assign n4748 = n733 & ~n4513 ;
  assign n4749 = ( x87 & ~n463 ) | ( x87 & n1620 ) | ( ~n463 & n1620 ) ;
  assign n4750 = n4748 & ~n4749 ;
  assign n4751 = n4750 ^ n3579 ^ 1'b0 ;
  assign n4752 = n4751 ^ x35 ^ 1'b0 ;
  assign n4753 = n2394 ^ n1523 ^ 1'b0 ;
  assign n4754 = n4087 & n4753 ;
  assign n4755 = n4754 ^ n865 ^ 1'b0 ;
  assign n4756 = n1634 & n2860 ;
  assign n4757 = n4756 ^ n336 ^ 1'b0 ;
  assign n4758 = n867 | n4757 ;
  assign n4759 = n2736 ^ n606 ^ 1'b0 ;
  assign n4760 = n3998 ^ n2357 ^ 1'b0 ;
  assign n4761 = n4182 | n4760 ;
  assign n4762 = n639 ^ n571 ^ 1'b0 ;
  assign n4763 = n718 | n4762 ;
  assign n4764 = n1356 & ~n4763 ;
  assign n4765 = n4764 ^ x15 ^ 1'b0 ;
  assign n4766 = n1162 & ~n4474 ;
  assign n4767 = n4766 ^ n1737 ^ 1'b0 ;
  assign n4768 = n1333 | n4767 ;
  assign n4769 = x119 & ~n836 ;
  assign n4770 = ~n567 & n4769 ;
  assign n4771 = n4770 ^ n194 ^ 1'b0 ;
  assign n4772 = n3731 & n4771 ;
  assign n4773 = n4772 ^ n851 ^ 1'b0 ;
  assign n4774 = n530 & ~n3579 ;
  assign n4775 = n3422 & n4774 ;
  assign n4776 = n3230 ^ n2101 ^ 1'b0 ;
  assign n4777 = n201 & n4776 ;
  assign n4779 = n3281 ^ n544 ^ 1'b0 ;
  assign n4778 = n1093 & n4310 ;
  assign n4780 = n4779 ^ n4778 ^ 1'b0 ;
  assign n4781 = n2566 | n4780 ;
  assign n4782 = n2942 & n4338 ;
  assign n4783 = n1937 & n4782 ;
  assign n4784 = n1443 | n4783 ;
  assign n4785 = n428 | n872 ;
  assign n4786 = n2986 | n4785 ;
  assign n4787 = n4786 ^ n2166 ^ n2130 ;
  assign n4788 = n1381 ^ n533 ^ 1'b0 ;
  assign n4789 = n4788 ^ n4375 ^ 1'b0 ;
  assign n4790 = ~n4787 & n4789 ;
  assign n4791 = n2563 ^ n2561 ^ 1'b0 ;
  assign n4792 = n1199 & n2245 ;
  assign n4793 = n3981 & n4792 ;
  assign n4795 = ~n1351 & n2851 ;
  assign n4796 = n1116 & n4795 ;
  assign n4794 = ~n3435 & n4618 ;
  assign n4797 = n4796 ^ n4794 ^ 1'b0 ;
  assign n4798 = x64 & n3998 ;
  assign n4799 = n574 | n2743 ;
  assign n4800 = n4799 ^ n4421 ^ 1'b0 ;
  assign n4801 = n4800 ^ n3213 ^ 1'b0 ;
  assign n4802 = n233 & ~n4801 ;
  assign n4803 = n2064 & n2618 ;
  assign n4804 = n4803 ^ n2851 ^ 1'b0 ;
  assign n4805 = ~n567 & n3987 ;
  assign n4806 = ~n508 & n4805 ;
  assign n4807 = n4748 ^ n3262 ^ n3147 ;
  assign n4808 = n1966 ^ n1786 ^ 1'b0 ;
  assign n4809 = ~n4807 & n4808 ;
  assign n4810 = n3328 ^ n2035 ^ 1'b0 ;
  assign n4811 = n1985 | n4810 ;
  assign n4812 = n828 | n1612 ;
  assign n4813 = n1217 ^ n385 ^ 1'b0 ;
  assign n4814 = n4812 | n4813 ;
  assign n4815 = n1312 & n2923 ;
  assign n4816 = n4815 ^ n3855 ^ 1'b0 ;
  assign n4817 = n812 & ~n4816 ;
  assign n4818 = n173 & n430 ;
  assign n4819 = n4818 ^ n1793 ^ 1'b0 ;
  assign n4820 = ~x56 & n2632 ;
  assign n4821 = ~n1054 & n1839 ;
  assign n4822 = ~n4091 & n4821 ;
  assign n4823 = n4822 ^ n3807 ^ 1'b0 ;
  assign n4824 = n2736 ^ n344 ^ 1'b0 ;
  assign n4825 = n129 | n2733 ;
  assign n4826 = n1993 & ~n3289 ;
  assign n4827 = n277 & ~n4826 ;
  assign n4828 = n4827 ^ n141 ^ 1'b0 ;
  assign n4829 = n1833 & ~n4218 ;
  assign n4830 = ~n2664 & n4829 ;
  assign n4831 = n996 & n1819 ;
  assign n4832 = n4831 ^ n163 ^ 1'b0 ;
  assign n4833 = x47 & n3890 ;
  assign n4834 = n4833 ^ n1993 ^ 1'b0 ;
  assign n4835 = n4832 & n4834 ;
  assign n4837 = ~n510 & n1412 ;
  assign n4836 = n3098 & n3989 ;
  assign n4838 = n4837 ^ n4836 ^ 1'b0 ;
  assign n4839 = n2196 ^ n886 ^ 1'b0 ;
  assign n4840 = n2797 & n4839 ;
  assign n4841 = n4234 & n4840 ;
  assign n4842 = ~x80 & n4841 ;
  assign n4843 = n3987 ^ n2644 ^ 1'b0 ;
  assign n4844 = n2967 & n3015 ;
  assign n4845 = ~n3677 & n4844 ;
  assign n4846 = n1005 & n3708 ;
  assign n4847 = n4846 ^ n3891 ^ 1'b0 ;
  assign n4848 = n4847 ^ n3445 ^ n686 ;
  assign n4849 = n4848 ^ n2198 ^ 1'b0 ;
  assign n4850 = ~n945 & n4849 ;
  assign n4851 = n3391 ^ n3338 ^ 1'b0 ;
  assign n4852 = n493 & ~n3091 ;
  assign n4853 = ~n1669 & n4852 ;
  assign n4854 = n1080 | n4853 ;
  assign n4855 = ~n2178 & n2395 ;
  assign n4856 = n1578 & n4855 ;
  assign n4857 = n3662 ^ n901 ^ 1'b0 ;
  assign n4858 = n1784 & n2678 ;
  assign n4859 = n1867 & ~n4858 ;
  assign n4860 = n2243 & ~n2470 ;
  assign n4861 = n2339 | n3458 ;
  assign n4862 = n3648 ^ x60 ^ 1'b0 ;
  assign n4863 = n169 & ~n1340 ;
  assign n4864 = n766 | n4863 ;
  assign n4865 = n4862 & ~n4864 ;
  assign n4870 = n2087 ^ n1512 ^ x8 ;
  assign n4866 = ~n904 & n1444 ;
  assign n4867 = n4866 ^ n663 ^ 1'b0 ;
  assign n4868 = n2210 | n2309 ;
  assign n4869 = n4867 | n4868 ;
  assign n4871 = n4870 ^ n4869 ^ 1'b0 ;
  assign n4872 = n4871 ^ n2743 ^ 1'b0 ;
  assign n4873 = ~n3474 & n4872 ;
  assign n4875 = n1380 | n1383 ;
  assign n4876 = n4875 ^ n1364 ^ 1'b0 ;
  assign n4874 = ~n1476 & n3182 ;
  assign n4877 = n4876 ^ n4874 ^ 1'b0 ;
  assign n4878 = n1807 ^ x124 ^ 1'b0 ;
  assign n4879 = ~n299 & n3955 ;
  assign n4880 = n4879 ^ n1158 ^ 1'b0 ;
  assign n4881 = ~n1314 & n4880 ;
  assign n4882 = n4881 ^ n1153 ^ 1'b0 ;
  assign n4890 = n1351 & ~n4076 ;
  assign n4891 = n4890 ^ n3503 ^ 1'b0 ;
  assign n4883 = n213 & ~n724 ;
  assign n4884 = x96 & ~n146 ;
  assign n4885 = n1781 & n4884 ;
  assign n4886 = n849 & n4885 ;
  assign n4887 = n844 & ~n4886 ;
  assign n4888 = ~n4883 & n4887 ;
  assign n4889 = n4669 | n4888 ;
  assign n4892 = n4891 ^ n4889 ^ n1201 ;
  assign n4893 = n2994 & n3383 ;
  assign n4894 = x124 & n951 ;
  assign n4895 = n4894 ^ n1703 ^ 1'b0 ;
  assign n4896 = n3961 ^ n1683 ^ 1'b0 ;
  assign n4897 = n3498 | n4896 ;
  assign n4898 = n4897 ^ n3110 ^ 1'b0 ;
  assign n4899 = n1993 & ~n3710 ;
  assign n4900 = n4240 ^ n4206 ^ n478 ;
  assign n4901 = n2694 | n2917 ;
  assign n4902 = n642 & ~n961 ;
  assign n4903 = n4901 & ~n4902 ;
  assign n4904 = n4900 & n4903 ;
  assign n4905 = n4904 ^ n361 ^ 1'b0 ;
  assign n4906 = n2864 | n4905 ;
  assign n4907 = n4771 ^ n3666 ^ 1'b0 ;
  assign n4908 = n436 & ~n2156 ;
  assign n4909 = ~n632 & n3573 ;
  assign n4910 = n4908 & n4909 ;
  assign n4911 = n2198 ^ n2097 ^ 1'b0 ;
  assign n4912 = n406 & ~n1699 ;
  assign n4913 = ~n4911 & n4912 ;
  assign n4914 = n2516 & n4913 ;
  assign n4915 = n376 | n2151 ;
  assign n4916 = ~n288 & n1973 ;
  assign n4917 = n3581 ^ n2040 ^ 1'b0 ;
  assign n4918 = n634 & n4917 ;
  assign n4919 = n2265 & n4918 ;
  assign n4920 = x62 & ~n4919 ;
  assign n4921 = n1031 & ~n1675 ;
  assign n4923 = n2553 ^ x60 ^ 1'b0 ;
  assign n4922 = n3902 & n3964 ;
  assign n4924 = n4923 ^ n4922 ^ 1'b0 ;
  assign n4925 = ~n4921 & n4924 ;
  assign n4926 = n155 & n4925 ;
  assign n4927 = n1866 ^ n143 ^ 1'b0 ;
  assign n4928 = ~n839 & n4927 ;
  assign n4929 = n2686 & ~n3066 ;
  assign n4930 = n339 | n2394 ;
  assign n4931 = n4930 ^ n3563 ^ 1'b0 ;
  assign n4932 = n3731 ^ n1395 ^ 1'b0 ;
  assign n4933 = n4931 | n4932 ;
  assign n4934 = n1270 & ~n1880 ;
  assign n4935 = ~n1329 & n4934 ;
  assign n4936 = n2743 | n4935 ;
  assign n4937 = n4936 ^ n2285 ^ 1'b0 ;
  assign n4938 = n4937 ^ n950 ^ 1'b0 ;
  assign n4939 = n221 & ~n4938 ;
  assign n4940 = ~n1468 & n4939 ;
  assign n4941 = ~n594 & n4940 ;
  assign n4942 = n1211 ^ n687 ^ 1'b0 ;
  assign n4945 = n1015 ^ n721 ^ 1'b0 ;
  assign n4946 = n632 & n4945 ;
  assign n4943 = n4747 ^ n1588 ^ 1'b0 ;
  assign n4944 = x37 & ~n4943 ;
  assign n4947 = n4946 ^ n4944 ^ 1'b0 ;
  assign n4948 = n3840 & n4009 ;
  assign n4950 = n512 ^ n394 ^ 1'b0 ;
  assign n4951 = ~n428 & n4950 ;
  assign n4952 = n729 & n3865 ;
  assign n4953 = ~n4951 & n4952 ;
  assign n4949 = ~n3135 & n4019 ;
  assign n4954 = n4953 ^ n4949 ^ 1'b0 ;
  assign n4955 = x126 & n305 ;
  assign n4956 = n4018 & n4955 ;
  assign n4957 = n3414 & ~n4098 ;
  assign n4958 = n4957 ^ n3544 ^ 1'b0 ;
  assign n4959 = n137 & ~n2392 ;
  assign n4960 = n4959 ^ n1461 ^ x44 ;
  assign n4961 = ( n4636 & n4958 ) | ( n4636 & ~n4960 ) | ( n4958 & ~n4960 ) ;
  assign n4962 = n3542 | n3714 ;
  assign n4963 = ~n1436 & n2367 ;
  assign n4964 = n4962 & n4963 ;
  assign n4965 = n528 ^ x52 ^ 1'b0 ;
  assign n4966 = n1327 ^ n1224 ^ 1'b0 ;
  assign n4967 = x114 & ~n1463 ;
  assign n4968 = ~x118 & n3094 ;
  assign n4969 = n1004 | n4964 ;
  assign n4970 = n788 | n4969 ;
  assign n4971 = n2101 ^ n857 ^ 1'b0 ;
  assign n4972 = n2592 & n4971 ;
  assign n4973 = n2679 ^ n642 ^ 1'b0 ;
  assign n4974 = n4972 & ~n4973 ;
  assign n4975 = n333 & ~n632 ;
  assign n4976 = n677 & n4975 ;
  assign n4977 = n4976 ^ n2694 ^ 1'b0 ;
  assign n4978 = n985 | n4977 ;
  assign n4980 = n926 ^ n707 ^ 1'b0 ;
  assign n4979 = n163 & n1064 ;
  assign n4981 = n4980 ^ n4979 ^ 1'b0 ;
  assign n4982 = n2697 ^ n1609 ^ 1'b0 ;
  assign n4983 = n763 & ~n4982 ;
  assign n4984 = n4059 & n4983 ;
  assign n4985 = n4757 & n4984 ;
  assign n4986 = n4985 ^ n1428 ^ 1'b0 ;
  assign n4987 = n139 | n4986 ;
  assign n4988 = n3007 ^ n132 ^ 1'b0 ;
  assign n4989 = ~n4987 & n4988 ;
  assign n4990 = n4989 ^ n2981 ^ 1'b0 ;
  assign n4991 = n2168 ^ n1160 ^ 1'b0 ;
  assign n4992 = n3327 & ~n4991 ;
  assign n4993 = n793 & n3291 ;
  assign n4994 = ~n1694 & n4993 ;
  assign n4995 = ~n3613 & n4994 ;
  assign n4996 = n978 & ~n3272 ;
  assign n4997 = n3210 ^ n1756 ^ 1'b0 ;
  assign n4998 = n806 & ~n4997 ;
  assign n5000 = n566 | n877 ;
  assign n4999 = n4296 ^ n453 ^ 1'b0 ;
  assign n5001 = n5000 ^ n4999 ^ 1'b0 ;
  assign n5002 = ~n936 & n5001 ;
  assign n5003 = n1823 ^ n358 ^ 1'b0 ;
  assign n5004 = n2148 | n2981 ;
  assign n5005 = n2598 ^ n2264 ^ n1673 ;
  assign n5006 = ~n4908 & n5005 ;
  assign n5007 = n360 & n5006 ;
  assign n5008 = n542 ^ x65 ^ 1'b0 ;
  assign n5009 = x17 & ~n5008 ;
  assign n5010 = ~n1079 & n5009 ;
  assign n5011 = n3271 ^ n2194 ^ n890 ;
  assign n5012 = n2989 ^ n2041 ^ 1'b0 ;
  assign n5013 = n2441 & ~n5012 ;
  assign n5014 = ~n1932 & n5013 ;
  assign n5015 = ~n1613 & n5014 ;
  assign n5016 = n5015 ^ n2186 ^ 1'b0 ;
  assign n5017 = n2176 ^ n528 ^ 1'b0 ;
  assign n5018 = x37 & ~n5017 ;
  assign n5019 = n3514 ^ n967 ^ 1'b0 ;
  assign n5020 = n1542 & ~n5019 ;
  assign n5021 = n613 | n2361 ;
  assign n5022 = n3708 & ~n5021 ;
  assign n5023 = n1428 ^ n508 ^ 1'b0 ;
  assign n5024 = n992 | n5023 ;
  assign n5025 = n2079 | n5024 ;
  assign n5026 = ~n5022 & n5025 ;
  assign n5027 = n5026 ^ n2344 ^ 1'b0 ;
  assign n5028 = n793 & n5027 ;
  assign n5029 = ( ~n684 & n5020 ) | ( ~n684 & n5028 ) | ( n5020 & n5028 ) ;
  assign n5030 = n5029 ^ n2516 ^ 1'b0 ;
  assign n5031 = n2366 & ~n5030 ;
  assign n5032 = ~n2822 & n3960 ;
  assign n5033 = ~n1637 & n5032 ;
  assign n5034 = n4796 | n5033 ;
  assign n5035 = n5034 ^ n2210 ^ 1'b0 ;
  assign n5036 = n5035 ^ n4107 ^ 1'b0 ;
  assign n5037 = n2694 ^ n285 ^ 1'b0 ;
  assign n5038 = n2020 ^ n639 ^ 1'b0 ;
  assign n5039 = ~n2741 & n5038 ;
  assign n5040 = n535 | n1811 ;
  assign n5041 = n2263 & ~n2789 ;
  assign n5042 = n5041 ^ n1491 ^ 1'b0 ;
  assign n5044 = n4341 ^ n2765 ^ 1'b0 ;
  assign n5045 = ~n427 & n5044 ;
  assign n5043 = n2734 ^ n487 ^ 1'b0 ;
  assign n5046 = n5045 ^ n5043 ^ 1'b0 ;
  assign n5047 = n3414 & ~n4713 ;
  assign n5048 = n5046 & n5047 ;
  assign n5049 = n572 ^ n432 ^ 1'b0 ;
  assign n5050 = n387 & ~n5049 ;
  assign n5051 = n2144 | n2872 ;
  assign n5052 = n5050 | n5051 ;
  assign n5053 = n311 & n1817 ;
  assign n5054 = ~n5052 & n5053 ;
  assign n5055 = n409 & ~n1349 ;
  assign n5056 = n1606 & n5055 ;
  assign n5057 = n5056 ^ n1631 ^ 1'b0 ;
  assign n5058 = n593 | n2037 ;
  assign n5059 = n5058 ^ n478 ^ 1'b0 ;
  assign n5060 = n5059 ^ n159 ^ 1'b0 ;
  assign n5061 = n1262 & n2264 ;
  assign n5062 = ~n251 & n5061 ;
  assign n5063 = n5062 ^ n499 ^ 1'b0 ;
  assign n5064 = n1452 & n5063 ;
  assign n5065 = n5064 ^ n3874 ^ 1'b0 ;
  assign n5066 = n2893 & ~n3165 ;
  assign n5067 = n811 & n5066 ;
  assign n5068 = n2994 ^ n717 ^ 1'b0 ;
  assign n5069 = n177 | n1340 ;
  assign n5070 = n5069 ^ n4282 ^ 1'b0 ;
  assign n5071 = n2833 | n5070 ;
  assign n5072 = n5068 & ~n5071 ;
  assign n5073 = n4019 & n4937 ;
  assign n5074 = ~n1042 & n5073 ;
  assign n5075 = n2692 ^ n2517 ^ 1'b0 ;
  assign n5076 = n359 & ~n5075 ;
  assign n5077 = n2160 | n2601 ;
  assign n5078 = n2532 | n4113 ;
  assign n5079 = n4113 & ~n5078 ;
  assign n5080 = n4253 & ~n5079 ;
  assign n5081 = n5079 & n5080 ;
  assign n5082 = n5077 & ~n5081 ;
  assign n5083 = ~n5077 & n5082 ;
  assign n5084 = n1580 & ~n5083 ;
  assign n5085 = n4323 & n5084 ;
  assign n5086 = ~n1071 & n4521 ;
  assign n5087 = n1372 & n1843 ;
  assign n5088 = n2201 ^ n1914 ^ 1'b0 ;
  assign n5089 = n1985 | n5088 ;
  assign n5090 = ~n5011 & n5089 ;
  assign n5091 = ~n3132 & n3182 ;
  assign n5092 = n1856 ^ n667 ^ 1'b0 ;
  assign n5093 = n2374 & n5092 ;
  assign n5094 = ~n698 & n1968 ;
  assign n5095 = n5094 ^ x114 ^ 1'b0 ;
  assign n5096 = n237 & ~n5095 ;
  assign n5097 = n5096 ^ n4346 ^ 1'b0 ;
  assign n5098 = ~n1158 & n2285 ;
  assign n5099 = n4289 ^ n3431 ^ 1'b0 ;
  assign n5100 = n1710 ^ n510 ^ 1'b0 ;
  assign n5101 = n1502 | n5100 ;
  assign n5102 = n4816 ^ n3174 ^ 1'b0 ;
  assign n5103 = n4325 ^ n2237 ^ 1'b0 ;
  assign n5104 = ~n1878 & n2155 ;
  assign n5105 = n2735 | n5104 ;
  assign n5106 = n4671 ^ n310 ^ 1'b0 ;
  assign n5107 = ~n1513 & n4557 ;
  assign n5108 = n5107 ^ n2163 ^ 1'b0 ;
  assign n5109 = n5108 ^ n2321 ^ 1'b0 ;
  assign n5110 = ~n1975 & n5109 ;
  assign n5111 = n469 | n1932 ;
  assign n5112 = n1456 | n5111 ;
  assign n5113 = n2582 | n3900 ;
  assign n5114 = n5112 & ~n5113 ;
  assign n5115 = ~n3400 & n5114 ;
  assign n5116 = x87 & ~n238 ;
  assign n5117 = n5116 ^ n625 ^ 1'b0 ;
  assign n5118 = n5117 ^ n996 ^ 1'b0 ;
  assign n5119 = n5118 ^ n4106 ^ n728 ;
  assign n5120 = n931 | n5119 ;
  assign n5121 = ~n2130 & n4457 ;
  assign n5122 = n4749 ^ x23 ^ 1'b0 ;
  assign n5123 = x19 & ~n2017 ;
  assign n5124 = n2099 & n2543 ;
  assign n5125 = n5124 ^ n2323 ^ 1'b0 ;
  assign n5126 = n5125 ^ n3698 ^ 1'b0 ;
  assign n5127 = n4990 & n5126 ;
  assign n5128 = n1361 | n3853 ;
  assign n5129 = n4048 ^ n1832 ^ 1'b0 ;
  assign n5130 = n623 & ~n5129 ;
  assign n5131 = n1950 ^ n939 ^ 1'b0 ;
  assign n5132 = n781 | n5131 ;
  assign n5139 = ~n235 & n2729 ;
  assign n5134 = ~n974 & n1170 ;
  assign n5135 = ~n1986 & n5134 ;
  assign n5136 = n5135 ^ n2855 ^ 1'b0 ;
  assign n5133 = n1212 | n1532 ;
  assign n5137 = n5136 ^ n5133 ^ 1'b0 ;
  assign n5138 = x57 & n5137 ;
  assign n5140 = n5139 ^ n5138 ^ 1'b0 ;
  assign n5141 = ~n300 & n1663 ;
  assign n5142 = n5141 ^ n2394 ^ 1'b0 ;
  assign n5143 = n5142 ^ n901 ^ 1'b0 ;
  assign n5151 = n1733 & n3220 ;
  assign n5144 = n414 ^ n262 ^ 1'b0 ;
  assign n5145 = n5061 ^ n3170 ^ 1'b0 ;
  assign n5146 = n2108 | n5145 ;
  assign n5147 = n5146 ^ n3251 ^ 1'b0 ;
  assign n5148 = ~x39 & n5147 ;
  assign n5149 = n5148 ^ n245 ^ 1'b0 ;
  assign n5150 = ~n5144 & n5149 ;
  assign n5152 = n5151 ^ n5150 ^ 1'b0 ;
  assign n5154 = x61 & ~n2906 ;
  assign n5153 = n358 | n2281 ;
  assign n5155 = n5154 ^ n5153 ^ 1'b0 ;
  assign n5156 = ~x17 & n5155 ;
  assign n5157 = n161 & n1308 ;
  assign n5158 = n3614 & n5157 ;
  assign n5159 = n296 & ~n4592 ;
  assign n5160 = n1588 | n3746 ;
  assign n5161 = n1758 & ~n5160 ;
  assign n5162 = n1827 & n4194 ;
  assign n5163 = ~n2308 & n5162 ;
  assign n5164 = n507 & ~n3969 ;
  assign n5165 = n4450 & n5164 ;
  assign n5166 = n5165 ^ n3722 ^ 1'b0 ;
  assign n5167 = n5166 ^ n2009 ^ 1'b0 ;
  assign n5168 = ~n5163 & n5167 ;
  assign n5169 = x5 & ~n2852 ;
  assign n5170 = ~n835 & n5169 ;
  assign n5171 = n2975 ^ n1493 ^ 1'b0 ;
  assign n5172 = n5170 | n5171 ;
  assign n5174 = n2763 ^ n2309 ^ 1'b0 ;
  assign n5175 = n1146 & n5174 ;
  assign n5173 = n582 | n2161 ;
  assign n5176 = n5175 ^ n5173 ^ 1'b0 ;
  assign n5177 = n439 | n2533 ;
  assign n5178 = n233 | n5177 ;
  assign n5179 = n3157 & n3403 ;
  assign n5180 = n1001 & n3892 ;
  assign n5181 = n1420 & n5180 ;
  assign n5182 = n4746 & ~n5181 ;
  assign n5183 = n2982 ^ n650 ^ 1'b0 ;
  assign n5184 = n5183 ^ n4415 ^ 1'b0 ;
  assign n5187 = n570 ^ n321 ^ 1'b0 ;
  assign n5188 = n1724 | n3587 ;
  assign n5189 = n5187 & ~n5188 ;
  assign n5185 = n607 & n1280 ;
  assign n5186 = n5185 ^ n2086 ^ 1'b0 ;
  assign n5190 = n5189 ^ n5186 ^ 1'b0 ;
  assign n5191 = n3810 | n5190 ;
  assign n5192 = n5191 ^ n2900 ^ 1'b0 ;
  assign n5193 = n937 & ~n5192 ;
  assign n5194 = n2343 & n3077 ;
  assign n5195 = n5194 ^ n4708 ^ 1'b0 ;
  assign n5196 = n2091 ^ n1883 ^ 1'b0 ;
  assign n5197 = n4765 ^ n2692 ^ n775 ;
  assign n5198 = n2427 ^ n2269 ^ 1'b0 ;
  assign n5199 = n4455 ^ n3047 ^ 1'b0 ;
  assign n5200 = ~n5119 & n5199 ;
  assign n5201 = x3 & n2919 ;
  assign n5202 = ~n1790 & n5201 ;
  assign n5203 = n1882 & n5202 ;
  assign n5204 = n5203 ^ n4472 ^ n601 ;
  assign n5205 = n5204 ^ x92 ^ 1'b0 ;
  assign n5206 = n1142 & n1848 ;
  assign n5207 = n5206 ^ n245 ^ 1'b0 ;
  assign n5208 = n150 & n5207 ;
  assign n5209 = n797 & n5208 ;
  assign n5210 = ~n1590 & n5209 ;
  assign n5211 = n2094 | n5210 ;
  assign n5212 = n1052 ^ x42 ^ 1'b0 ;
  assign n5213 = x117 & ~n5212 ;
  assign n5214 = n1072 & ~n4204 ;
  assign n5215 = n5213 & n5214 ;
  assign n5216 = n1156 ^ n980 ^ 1'b0 ;
  assign n5217 = n1854 | n5216 ;
  assign n5218 = n1376 | n3655 ;
  assign n5219 = n3213 & ~n5218 ;
  assign n5220 = n909 & ~n2335 ;
  assign n5222 = ( n1782 & n2385 ) | ( n1782 & n3425 ) | ( n2385 & n3425 ) ;
  assign n5221 = n1264 | n2847 ;
  assign n5223 = n5222 ^ n5221 ^ 1'b0 ;
  assign n5224 = n1749 ^ x40 ^ 1'b0 ;
  assign n5225 = ~n4638 & n5224 ;
  assign n5226 = ~n5223 & n5225 ;
  assign n5227 = n1788 ^ n640 ^ 1'b0 ;
  assign n5228 = n1315 ^ x23 ^ 1'b0 ;
  assign n5229 = ( n2307 & n5227 ) | ( n2307 & ~n5228 ) | ( n5227 & ~n5228 ) ;
  assign n5230 = n4716 & n5229 ;
  assign n5231 = n3091 ^ x52 ^ 1'b0 ;
  assign n5232 = n3608 & n3794 ;
  assign n5233 = n540 & n2402 ;
  assign n5234 = n2505 ^ n1661 ^ 1'b0 ;
  assign n5235 = n189 | n3333 ;
  assign n5236 = n404 | n5235 ;
  assign n5237 = n5236 ^ n150 ^ 1'b0 ;
  assign n5238 = n865 | n2526 ;
  assign n5239 = ( n3662 & n4846 ) | ( n3662 & n5238 ) | ( n4846 & n5238 ) ;
  assign n5240 = n4318 & ~n5239 ;
  assign n5241 = n1786 ^ n455 ^ 1'b0 ;
  assign n5242 = ~n1841 & n5186 ;
  assign n5243 = n373 & ~n686 ;
  assign n5244 = n1277 ^ n542 ^ 1'b0 ;
  assign n5245 = n1635 & ~n5244 ;
  assign n5246 = n3764 ^ n912 ^ 1'b0 ;
  assign n5247 = n1209 & ~n5243 ;
  assign n5248 = n1636 | n3320 ;
  assign n5249 = n2935 ^ n2864 ^ 1'b0 ;
  assign n5250 = n442 & ~n448 ;
  assign n5251 = ~n4489 & n5250 ;
  assign n5252 = n304 | n707 ;
  assign n5253 = n4787 ^ n4343 ^ n1545 ;
  assign n5254 = n3403 ^ n1795 ^ 1'b0 ;
  assign n5255 = n1470 & ~n2139 ;
  assign n5256 = n3742 | n5255 ;
  assign n5257 = n4853 & ~n5256 ;
  assign n5258 = x116 & ~n3782 ;
  assign n5259 = n1959 ^ n134 ^ 1'b0 ;
  assign n5260 = n1290 & ~n2655 ;
  assign n5261 = n2404 & n2623 ;
  assign n5262 = n5261 ^ n1905 ^ 1'b0 ;
  assign n5263 = n5260 & n5262 ;
  assign n5264 = n754 ^ n425 ^ 1'b0 ;
  assign n5265 = ( n1854 & n3220 ) | ( n1854 & ~n4513 ) | ( n3220 & ~n4513 ) ;
  assign n5266 = n4650 | n5265 ;
  assign n5267 = n1697 | n5266 ;
  assign n5268 = n5264 & ~n5267 ;
  assign n5269 = n3966 ^ n1694 ^ 1'b0 ;
  assign n5270 = n4309 | n5269 ;
  assign n5271 = n1983 & ~n5270 ;
  assign n5272 = x94 & n2681 ;
  assign n5273 = n5272 ^ n1930 ^ 1'b0 ;
  assign n5274 = n4608 ^ n1418 ^ 1'b0 ;
  assign n5275 = n808 & n1478 ;
  assign n5276 = ~n5274 & n5275 ;
  assign n5277 = n5276 ^ n4941 ^ 1'b0 ;
  assign n5278 = n998 & n5277 ;
  assign n5279 = n1788 & ~n4370 ;
  assign n5280 = n4775 & n5279 ;
  assign n5281 = n3124 | n4933 ;
  assign n5282 = n1654 & ~n5281 ;
  assign n5283 = n1807 ^ n1749 ^ 1'b0 ;
  assign n5289 = x113 & ~n4490 ;
  assign n5285 = n645 & ~n1601 ;
  assign n5286 = n5285 ^ n262 ^ 1'b0 ;
  assign n5284 = n1914 ^ n310 ^ 1'b0 ;
  assign n5287 = n5286 ^ n5284 ^ 1'b0 ;
  assign n5288 = n4016 & n5287 ;
  assign n5290 = n5289 ^ n5288 ^ 1'b0 ;
  assign n5291 = n1788 ^ n1146 ^ n932 ;
  assign n5292 = ( n1251 & n2989 ) | ( n1251 & n5291 ) | ( n2989 & n5291 ) ;
  assign n5293 = x73 & n2337 ;
  assign n5294 = ~n222 & n1310 ;
  assign n5295 = n3823 & ~n5294 ;
  assign n5296 = n5293 & n5295 ;
  assign n5297 = ~n1281 & n5296 ;
  assign n5298 = n1707 ^ n361 ^ 1'b0 ;
  assign n5299 = n5298 ^ n4423 ^ 1'b0 ;
  assign n5300 = n575 | n5299 ;
  assign n5301 = n4041 & n4744 ;
  assign n5302 = n5301 ^ n3242 ^ 1'b0 ;
  assign n5303 = ~n640 & n1012 ;
  assign n5304 = ~n3470 & n5303 ;
  assign n5305 = n717 | n5304 ;
  assign n5306 = n5305 ^ n3439 ^ 1'b0 ;
  assign n5307 = n5306 ^ n4457 ^ 1'b0 ;
  assign n5308 = n3700 & ~n5307 ;
  assign n5309 = n1336 & ~n4559 ;
  assign n5310 = n3917 ^ n739 ^ 1'b0 ;
  assign n5311 = n279 | n2026 ;
  assign n5312 = n5311 ^ n267 ^ 1'b0 ;
  assign n5313 = n5312 ^ n2635 ^ n2143 ;
  assign n5314 = n1485 | n2584 ;
  assign n5315 = n4282 & ~n5314 ;
  assign n5316 = n2034 ^ n636 ^ 1'b0 ;
  assign n5317 = n3275 & n5316 ;
  assign n5318 = n5317 ^ n4282 ^ 1'b0 ;
  assign n5319 = n1041 ^ n782 ^ 1'b0 ;
  assign n5320 = n4895 & ~n5319 ;
  assign n5321 = n1342 ^ n169 ^ 1'b0 ;
  assign n5322 = n1366 | n1703 ;
  assign n5323 = n159 & n277 ;
  assign n5324 = n5322 & n5323 ;
  assign n5326 = n620 & ~n1812 ;
  assign n5327 = ~n2707 & n5326 ;
  assign n5325 = n970 & n1980 ;
  assign n5328 = n5327 ^ n5325 ^ 1'b0 ;
  assign n5329 = n2560 ^ n1228 ^ 1'b0 ;
  assign n5330 = n2815 ^ n2145 ^ n231 ;
  assign n5331 = n5330 ^ n1832 ^ 1'b0 ;
  assign n5332 = n908 & n5331 ;
  assign n5333 = ~n358 & n1087 ;
  assign n5334 = n1659 ^ n558 ^ 1'b0 ;
  assign n5335 = ~n675 & n5334 ;
  assign n5336 = n5335 ^ n1796 ^ 1'b0 ;
  assign n5337 = n2428 & n5336 ;
  assign n5339 = n3492 ^ n1979 ^ 1'b0 ;
  assign n5340 = ~n2705 & n5339 ;
  assign n5338 = n4062 ^ n1114 ^ 1'b0 ;
  assign n5341 = n5340 ^ n5338 ^ 1'b0 ;
  assign n5344 = n837 | n3124 ;
  assign n5345 = n814 | n5344 ;
  assign n5342 = n5165 ^ n786 ^ 1'b0 ;
  assign n5343 = ~n990 & n5342 ;
  assign n5346 = n5345 ^ n5343 ^ 1'b0 ;
  assign n5347 = n2602 & ~n3395 ;
  assign n5348 = n3592 ^ n753 ^ 1'b0 ;
  assign n5349 = n4444 & n5348 ;
  assign n5350 = n4489 ^ n338 ^ 1'b0 ;
  assign n5351 = n4263 ^ n2987 ^ 1'b0 ;
  assign n5352 = ~n5350 & n5351 ;
  assign n5353 = n2897 & ~n5352 ;
  assign n5354 = n557 | n1590 ;
  assign n5355 = n5354 ^ n2475 ^ 1'b0 ;
  assign n5356 = ~n5353 & n5355 ;
  assign n5357 = n1161 & ~n1928 ;
  assign n5358 = n5357 ^ n4298 ^ 1'b0 ;
  assign n5359 = n1480 ^ n722 ^ 1'b0 ;
  assign n5360 = ~n1993 & n5359 ;
  assign n5361 = n2852 ^ n1504 ^ 1'b0 ;
  assign n5362 = n5142 ^ n1747 ^ 1'b0 ;
  assign n5363 = n603 & ~n5362 ;
  assign n5364 = n3091 ^ n1312 ^ 1'b0 ;
  assign n5365 = n920 & ~n1082 ;
  assign n5366 = ~n1656 & n1720 ;
  assign n5367 = n1389 & ~n5366 ;
  assign n5368 = n3275 ^ n524 ^ 1'b0 ;
  assign n5369 = ~n5367 & n5368 ;
  assign n5370 = ~n5365 & n5369 ;
  assign n5371 = n5370 ^ n361 ^ 1'b0 ;
  assign n5372 = ~n5364 & n5371 ;
  assign n5373 = n972 ^ x97 ^ 1'b0 ;
  assign n5374 = n1232 ^ n165 ^ 1'b0 ;
  assign n5375 = n4397 ^ x55 ^ 1'b0 ;
  assign n5376 = n5374 & n5375 ;
  assign n5377 = n375 | n5376 ;
  assign n5378 = n853 ^ x97 ^ 1'b0 ;
  assign n5379 = ~n865 & n1920 ;
  assign n5380 = n5379 ^ n3687 ^ 1'b0 ;
  assign n5381 = n2733 & ~n5380 ;
  assign n5382 = x111 & n5381 ;
  assign n5383 = n781 & n5382 ;
  assign n5384 = n1865 & ~n5383 ;
  assign n5385 = n5384 ^ n3064 ^ 1'b0 ;
  assign n5386 = n307 & n5385 ;
  assign n5387 = n5386 ^ n5330 ^ 1'b0 ;
  assign n5388 = ~n2053 & n2391 ;
  assign n5389 = n2669 & ~n5139 ;
  assign n5390 = n3407 & n5389 ;
  assign n5391 = n5091 ^ n830 ^ 1'b0 ;
  assign n5392 = n4233 | n5391 ;
  assign n5393 = n4697 ^ n342 ^ 1'b0 ;
  assign n5394 = n1166 ^ n279 ^ 1'b0 ;
  assign n5395 = n5393 & ~n5394 ;
  assign n5396 = n3629 ^ n2707 ^ 1'b0 ;
  assign n5397 = n5395 & ~n5396 ;
  assign n5398 = n5377 ^ n2775 ^ 1'b0 ;
  assign n5399 = n4775 | n5398 ;
  assign n5400 = n412 | n2339 ;
  assign n5402 = n277 & ~n346 ;
  assign n5403 = ~n806 & n5402 ;
  assign n5401 = n2073 & ~n2985 ;
  assign n5404 = n5403 ^ n5401 ^ 1'b0 ;
  assign n5405 = n2643 ^ n2094 ^ n198 ;
  assign n5406 = n2828 ^ n1589 ^ n1463 ;
  assign n5407 = n5406 ^ n2630 ^ 1'b0 ;
  assign n5408 = n1563 | n5407 ;
  assign n5409 = n5408 ^ n1185 ^ 1'b0 ;
  assign n5410 = n5405 & n5409 ;
  assign n5411 = ~n1738 & n1964 ;
  assign n5412 = n2155 ^ n1393 ^ x61 ;
  assign n5413 = n5412 ^ n2056 ^ 1'b0 ;
  assign n5414 = n5413 ^ n451 ^ 1'b0 ;
  assign n5415 = ~n1623 & n2800 ;
  assign n5416 = n955 ^ n593 ^ 1'b0 ;
  assign n5417 = ~n2969 & n5416 ;
  assign n5418 = ~n656 & n3790 ;
  assign n5419 = ~n1240 & n5418 ;
  assign n5420 = ~n4751 & n5419 ;
  assign n5421 = n307 & n1157 ;
  assign n5422 = n5421 ^ n408 ^ 1'b0 ;
  assign n5423 = ~n2475 & n5422 ;
  assign n5424 = n5423 ^ n3717 ^ 1'b0 ;
  assign n5425 = n2381 ^ n1944 ^ 1'b0 ;
  assign n5426 = n2954 & ~n5425 ;
  assign n5427 = x73 & n3279 ;
  assign n5428 = n5427 ^ n1086 ^ 1'b0 ;
  assign n5429 = n5426 & ~n5428 ;
  assign n5430 = n2716 ^ n671 ^ 1'b0 ;
  assign n5431 = ~n1406 & n3260 ;
  assign n5432 = n5150 & ~n5431 ;
  assign n5435 = ~n2661 & n3500 ;
  assign n5433 = n131 & n1589 ;
  assign n5434 = n5433 ^ n2243 ^ 1'b0 ;
  assign n5436 = n5435 ^ n5434 ^ 1'b0 ;
  assign n5437 = n3218 & ~n3465 ;
  assign n5438 = n1779 & ~n2557 ;
  assign n5439 = n784 ^ x15 ^ 1'b0 ;
  assign n5440 = n3196 ^ n788 ^ 1'b0 ;
  assign n5441 = n2459 ^ n238 ^ 1'b0 ;
  assign n5442 = ~n444 & n5441 ;
  assign n5443 = ( x33 & n1052 ) | ( x33 & n5442 ) | ( n1052 & n5442 ) ;
  assign n5444 = ~x84 & n5443 ;
  assign n5445 = n4458 & n5444 ;
  assign n5446 = x70 & ~n2887 ;
  assign n5447 = n5446 ^ n849 ^ 1'b0 ;
  assign n5448 = x52 | n1020 ;
  assign n5449 = n842 | n5448 ;
  assign n5450 = n5447 & ~n5449 ;
  assign n5451 = n1177 & n1470 ;
  assign n5452 = n410 & n2303 ;
  assign n5453 = ~n1747 & n5452 ;
  assign n5454 = n135 & n3989 ;
  assign n5455 = ~n262 & n5454 ;
  assign n5456 = n4198 ^ n2692 ^ n1013 ;
  assign n5457 = ~n5455 & n5456 ;
  assign n5458 = ~n1381 & n5457 ;
  assign n5459 = n5453 | n5458 ;
  assign n5460 = n5459 ^ n2847 ^ 1'b0 ;
  assign n5461 = n165 & ~n656 ;
  assign n5462 = ~n874 & n5461 ;
  assign n5463 = n5462 ^ n4954 ^ 1'b0 ;
  assign n5464 = n2226 ^ n1552 ^ 1'b0 ;
  assign n5465 = ~n2926 & n3730 ;
  assign n5466 = n5465 ^ n1808 ^ 1'b0 ;
  assign n5467 = ~n2569 & n3570 ;
  assign n5468 = n2156 & ~n2669 ;
  assign n5469 = n5468 ^ n583 ^ 1'b0 ;
  assign n5470 = n3393 | n5469 ;
  assign n5472 = n496 | n1499 ;
  assign n5473 = n2323 & ~n5472 ;
  assign n5474 = n5181 & n5473 ;
  assign n5471 = n558 & n4816 ;
  assign n5475 = n5474 ^ n5471 ^ 1'b0 ;
  assign n5476 = n1400 | n1671 ;
  assign n5477 = n158 | n799 ;
  assign n5478 = n4631 ^ n4153 ^ 1'b0 ;
  assign n5479 = n5477 & n5478 ;
  assign n5480 = n2136 ^ n739 ^ 1'b0 ;
  assign n5481 = ~n868 & n5480 ;
  assign n5482 = ~n266 & n5481 ;
  assign n5483 = n144 | n2364 ;
  assign n5484 = n3195 ^ n2704 ^ 1'b0 ;
  assign n5485 = n4671 & n5484 ;
  assign n5486 = n5485 ^ n1537 ^ 1'b0 ;
  assign n5487 = n1580 ^ n776 ^ 1'b0 ;
  assign n5488 = n5487 ^ n5364 ^ 1'b0 ;
  assign n5489 = n4564 | n5488 ;
  assign n5490 = n5486 & ~n5489 ;
  assign n5491 = n5490 ^ n4992 ^ 1'b0 ;
  assign n5492 = n1858 | n3128 ;
  assign n5493 = x8 & n316 ;
  assign n5494 = ~n316 & n5493 ;
  assign n5495 = x94 & n5494 ;
  assign n5496 = n639 & n5495 ;
  assign n5497 = ~n3514 & n5496 ;
  assign n5498 = n1950 & ~n5497 ;
  assign n5505 = x56 & ~n1832 ;
  assign n5506 = ~x56 & n5505 ;
  assign n5507 = ~n485 & n1833 ;
  assign n5508 = n5506 & n5507 ;
  assign n5503 = n363 | n4652 ;
  assign n5499 = n2257 & n4346 ;
  assign n5500 = n2677 & n5499 ;
  assign n5501 = n5500 ^ n2112 ^ 1'b0 ;
  assign n5502 = ~n3807 & n5501 ;
  assign n5504 = n5503 ^ n5502 ^ 1'b0 ;
  assign n5509 = n5508 ^ n5504 ^ 1'b0 ;
  assign n5510 = n5498 | n5509 ;
  assign n5511 = n2923 & ~n4303 ;
  assign n5512 = n5511 ^ n1913 ^ 1'b0 ;
  assign n5513 = ( n811 & ~n1258 ) | ( n811 & n5512 ) | ( ~n1258 & n5512 ) ;
  assign n5514 = n171 & n1961 ;
  assign n5515 = n5514 ^ n3680 ^ 1'b0 ;
  assign n5516 = n5513 | n5515 ;
  assign n5517 = n3557 | n4304 ;
  assign n5518 = n487 | n5327 ;
  assign n5519 = n5518 ^ n2664 ^ 1'b0 ;
  assign n5520 = n1387 | n1394 ;
  assign n5521 = n800 & ~n5520 ;
  assign n5522 = ~n5519 & n5521 ;
  assign n5523 = n5492 | n5522 ;
  assign n5524 = n3433 & ~n5523 ;
  assign n5525 = n356 & n1788 ;
  assign n5526 = n5525 ^ n1340 ^ 1'b0 ;
  assign n5527 = n1786 & n2347 ;
  assign n5528 = ~n4210 & n5527 ;
  assign n5529 = ~n3525 & n5395 ;
  assign n5530 = n5529 ^ n1205 ^ 1'b0 ;
  assign n5531 = n2010 & ~n4600 ;
  assign n5532 = n5531 ^ n1443 ^ 1'b0 ;
  assign n5533 = n1487 | n5532 ;
  assign n5534 = n5530 & ~n5533 ;
  assign n5535 = n830 & ~n2882 ;
  assign n5536 = n5535 ^ n1642 ^ 1'b0 ;
  assign n5537 = n616 | n3218 ;
  assign n5538 = n2325 ^ n999 ^ 1'b0 ;
  assign n5539 = n5538 ^ n1290 ^ 1'b0 ;
  assign n5540 = n3525 | n5539 ;
  assign n5541 = n5103 ^ n2692 ^ n2009 ;
  assign n5547 = n1499 ^ n489 ^ 1'b0 ;
  assign n5548 = n2137 & n5547 ;
  assign n5543 = n3151 ^ n2381 ^ 1'b0 ;
  assign n5544 = n1367 ^ n1080 ^ 1'b0 ;
  assign n5545 = n5543 & ~n5544 ;
  assign n5542 = n251 | n1990 ;
  assign n5546 = n5545 ^ n5542 ^ 1'b0 ;
  assign n5549 = n5548 ^ n5546 ^ 1'b0 ;
  assign n5550 = n4529 ^ n3138 ^ n2749 ;
  assign n5551 = n2953 | n3602 ;
  assign n5552 = n3664 & n5551 ;
  assign n5553 = n1724 ^ n570 ^ 1'b0 ;
  assign n5554 = n694 | n3764 ;
  assign n5555 = n5553 | n5554 ;
  assign n5556 = n4179 ^ n2208 ^ 1'b0 ;
  assign n5557 = n1331 ^ n623 ^ 1'b0 ;
  assign n5558 = n5557 ^ n235 ^ 1'b0 ;
  assign n5559 = n1456 | n1537 ;
  assign n5560 = n601 ^ n478 ^ 1'b0 ;
  assign n5561 = n1437 | n3416 ;
  assign n5562 = n5561 ^ x91 ^ 1'b0 ;
  assign n5563 = n293 ^ n213 ^ 1'b0 ;
  assign n5564 = n992 & n3398 ;
  assign n5565 = n5563 & n5564 ;
  assign n5566 = n5565 ^ n3238 ^ 1'b0 ;
  assign n5567 = n960 ^ x35 ^ 1'b0 ;
  assign n5568 = n1489 & ~n5567 ;
  assign n5569 = n790 & n5568 ;
  assign n5570 = n1055 & n5569 ;
  assign n5571 = n4177 & ~n5570 ;
  assign n5572 = ( n4298 & n4878 ) | ( n4298 & n5571 ) | ( n4878 & n5571 ) ;
  assign n5573 = n1738 ^ n616 ^ 1'b0 ;
  assign n5574 = n5341 ^ n4505 ^ 1'b0 ;
  assign n5575 = n2149 & n4179 ;
  assign n5577 = n194 & n2109 ;
  assign n5578 = n5577 ^ x59 ^ 1'b0 ;
  assign n5576 = ~n741 & n3837 ;
  assign n5579 = n5578 ^ n5576 ^ 1'b0 ;
  assign n5580 = n3654 ^ n2885 ^ 1'b0 ;
  assign n5581 = n3195 ^ n938 ^ 1'b0 ;
  assign n5582 = ~n4341 & n5581 ;
  assign n5583 = ~n786 & n5582 ;
  assign n5584 = n1909 ^ n353 ^ 1'b0 ;
  assign n5585 = n3009 & n3041 ;
  assign n5586 = n5585 ^ n3071 ^ 1'b0 ;
  assign n5587 = n3147 & n5586 ;
  assign n5588 = x57 & n5587 ;
  assign n5589 = n1728 | n5412 ;
  assign n5590 = n2946 & n3186 ;
  assign n5591 = n728 & n1315 ;
  assign n5592 = n5591 ^ n2317 ^ 1'b0 ;
  assign n5593 = ~n5532 & n5592 ;
  assign n5594 = n3866 ^ n1240 ^ 1'b0 ;
  assign n5595 = n2702 & n4190 ;
  assign n5596 = ~n880 & n1041 ;
  assign n5597 = n5596 ^ n1402 ^ 1'b0 ;
  assign n5598 = ~n272 & n5597 ;
  assign n5599 = ~n2789 & n5598 ;
  assign n5600 = ~n5595 & n5599 ;
  assign n5601 = n889 ^ n213 ^ 1'b0 ;
  assign n5602 = n1052 | n5601 ;
  assign n5603 = n5602 ^ n5235 ^ 1'b0 ;
  assign n5604 = ~n5132 & n5603 ;
  assign n5605 = ~n1042 & n5604 ;
  assign n5606 = n320 | n1554 ;
  assign n5607 = n3559 ^ n131 ^ 1'b0 ;
  assign n5608 = n3894 & n5607 ;
  assign n5609 = n3967 ^ n175 ^ 1'b0 ;
  assign n5610 = n4573 & n4820 ;
  assign n5611 = n5609 & n5610 ;
  assign n5612 = n5070 | n5611 ;
  assign n5613 = n5612 ^ n1510 ^ 1'b0 ;
  assign n5614 = n2393 ^ n895 ^ 1'b0 ;
  assign n5615 = n2173 | n5614 ;
  assign n5618 = x104 & x125 ;
  assign n5619 = n3290 | n5618 ;
  assign n5620 = n2942 | n5619 ;
  assign n5616 = n2521 ^ n1628 ^ 1'b0 ;
  assign n5617 = ~n2933 & n5616 ;
  assign n5621 = n5620 ^ n5617 ^ 1'b0 ;
  assign n5622 = n5621 ^ n4087 ^ n3900 ;
  assign n5623 = n1808 & n2374 ;
  assign n5624 = ~n238 & n1656 ;
  assign n5625 = ~x104 & n5624 ;
  assign n5626 = n5625 ^ n1578 ^ 1'b0 ;
  assign n5627 = n5626 ^ n5249 ^ 1'b0 ;
  assign n5628 = ~n1051 & n5627 ;
  assign n5629 = n5628 ^ n1659 ^ 1'b0 ;
  assign n5633 = ~n1428 & n1478 ;
  assign n5630 = n2383 & n5239 ;
  assign n5631 = ~n1133 & n1534 ;
  assign n5632 = n5630 & n5631 ;
  assign n5634 = n5633 ^ n5632 ^ n1183 ;
  assign n5635 = n869 & ~n3340 ;
  assign n5636 = n3116 | n5635 ;
  assign n5637 = n5636 ^ n200 ^ 1'b0 ;
  assign n5638 = ~n824 & n5637 ;
  assign n5639 = n177 | n2371 ;
  assign n5640 = n3502 ^ n2384 ^ 1'b0 ;
  assign n5641 = n1046 & n5640 ;
  assign n5642 = n5639 | n5641 ;
  assign n5643 = ( x94 & n1691 ) | ( x94 & ~n3754 ) | ( n1691 & ~n3754 ) ;
  assign n5644 = n189 | n1301 ;
  assign n5645 = n3169 & ~n5644 ;
  assign n5646 = n606 | n5645 ;
  assign n5647 = n2171 & ~n5646 ;
  assign n5648 = n304 & n5647 ;
  assign n5649 = n5621 ^ n2708 ^ 1'b0 ;
  assign n5650 = n1827 ^ n1694 ^ 1'b0 ;
  assign n5651 = n4188 & ~n5650 ;
  assign n5652 = x73 | n571 ;
  assign n5653 = n1427 & ~n5652 ;
  assign n5654 = n1627 & ~n3548 ;
  assign n5656 = ~n2480 & n3374 ;
  assign n5655 = x83 & ~n512 ;
  assign n5657 = n5656 ^ n5655 ^ 1'b0 ;
  assign n5658 = n5657 ^ n1695 ^ n326 ;
  assign n5659 = ~n1340 & n3268 ;
  assign n5660 = n383 | n1385 ;
  assign n5661 = n5660 ^ n5485 ^ 1'b0 ;
  assign n5662 = n2972 & ~n5461 ;
  assign n5663 = ~n4857 & n5662 ;
  assign n5664 = n1329 | n3195 ;
  assign n5665 = n5664 ^ n3431 ^ 1'b0 ;
  assign n5666 = n3157 & ~n5665 ;
  assign n5667 = n5666 ^ n4730 ^ 1'b0 ;
  assign n5668 = x94 & n3322 ;
  assign n5669 = n5668 ^ n2629 ^ 1'b0 ;
  assign n5670 = n5669 ^ n4086 ^ n2292 ;
  assign n5671 = n3100 | n5670 ;
  assign n5672 = n720 & ~n5671 ;
  assign n5673 = n888 & ~n1013 ;
  assign n5674 = ~n1783 & n5673 ;
  assign n5675 = n2351 | n3029 ;
  assign n5676 = n5674 & ~n5675 ;
  assign n5677 = ~x52 & n1713 ;
  assign n5678 = n1214 & n5677 ;
  assign n5679 = n5678 ^ n1620 ^ 1'b0 ;
  assign n5680 = ~n4013 & n5679 ;
  assign n5681 = n5680 ^ n766 ^ 1'b0 ;
  assign n5682 = n2573 & ~n5681 ;
  assign n5683 = n4202 | n5682 ;
  assign n5684 = x52 & n1837 ;
  assign n5685 = n992 & n5684 ;
  assign n5686 = x3 & n683 ;
  assign n5687 = n2573 & ~n5686 ;
  assign n5688 = n880 & n1328 ;
  assign n5689 = n5688 ^ n2678 ^ 1'b0 ;
  assign n5690 = n949 & ~n5689 ;
  assign n5691 = n5690 ^ n4037 ^ 1'b0 ;
  assign n5692 = x41 & ~n3544 ;
  assign n5693 = n2833 ^ n1321 ^ 1'b0 ;
  assign n5694 = n256 & n533 ;
  assign n5695 = n5022 & n5694 ;
  assign n5696 = n4282 & ~n5695 ;
  assign n5697 = n5387 & ~n5696 ;
  assign n5698 = ~n882 & n5697 ;
  assign n5699 = n3614 ^ n516 ^ 1'b0 ;
  assign n5700 = n3362 & ~n5699 ;
  assign n5701 = n1180 & ~n1563 ;
  assign n5702 = n1959 & n5701 ;
  assign n5703 = n1161 & n4019 ;
  assign n5704 = n5702 & n5703 ;
  assign n5705 = n438 | n5704 ;
  assign n5707 = n2980 & ~n4513 ;
  assign n5708 = n5707 ^ n4487 ^ 1'b0 ;
  assign n5706 = n1979 | n3678 ;
  assign n5709 = n5708 ^ n5706 ^ 1'b0 ;
  assign n5711 = n3675 ^ n3334 ^ 1'b0 ;
  assign n5710 = ~n924 & n2260 ;
  assign n5712 = n5711 ^ n5710 ^ n1629 ;
  assign n5713 = n3620 & ~n5712 ;
  assign n5714 = n3486 | n4282 ;
  assign n5715 = n1724 | n5714 ;
  assign n5716 = n5715 ^ n1080 ^ 1'b0 ;
  assign n5717 = n3486 ^ n3224 ^ 1'b0 ;
  assign n5718 = n428 | n5717 ;
  assign n5719 = ~n867 & n3958 ;
  assign n5720 = x94 | n5719 ;
  assign n5721 = ~n2049 & n3275 ;
  assign n5722 = n5249 | n5721 ;
  assign n5723 = n481 ^ n349 ^ 1'b0 ;
  assign n5724 = ~x54 & n5723 ;
  assign n5725 = n5724 ^ n4937 ^ 1'b0 ;
  assign n5726 = ~n2146 & n5725 ;
  assign n5727 = n2424 ^ n1566 ^ 1'b0 ;
  assign n5728 = n3009 & ~n3179 ;
  assign n5729 = n2430 & n5728 ;
  assign n5731 = n1864 & ~n4303 ;
  assign n5730 = n2862 | n3927 ;
  assign n5732 = n5731 ^ n5730 ^ n5176 ;
  assign n5733 = n3251 ^ n1162 ^ 1'b0 ;
  assign n5734 = n351 ^ x46 ^ 1'b0 ;
  assign n5735 = ~n613 & n5734 ;
  assign n5736 = n880 | n1437 ;
  assign n5737 = n1062 & n1064 ;
  assign n5738 = n5736 & n5737 ;
  assign n5739 = ~n2667 & n5738 ;
  assign n5740 = n702 & n1686 ;
  assign n5741 = ~n4753 & n5740 ;
  assign n5742 = n5741 ^ n279 ^ 1'b0 ;
  assign n5743 = ~n5739 & n5742 ;
  assign n5744 = n5743 ^ n2324 ^ 1'b0 ;
  assign n5745 = n5735 & n5744 ;
  assign n5746 = n1865 & n5005 ;
  assign n5747 = n3791 | n3882 ;
  assign n5748 = ( n1169 & n1759 ) | ( n1169 & ~n5747 ) | ( n1759 & ~n5747 ) ;
  assign n5749 = n1498 ^ n361 ^ n143 ;
  assign n5750 = n5748 & ~n5749 ;
  assign n5751 = n3019 & n5750 ;
  assign n5752 = n4865 | n5751 ;
  assign n5753 = n5752 ^ n1952 ^ 1'b0 ;
  assign n5754 = ( n219 & ~n1723 ) | ( n219 & n5679 ) | ( ~n1723 & n5679 ) ;
  assign n5755 = n5754 ^ n4621 ^ 1'b0 ;
  assign n5756 = ~n1781 & n3388 ;
  assign n5757 = n5756 ^ x104 ^ 1'b0 ;
  assign n5758 = n5437 ^ n4569 ^ 1'b0 ;
  assign n5759 = n3380 ^ n2256 ^ 1'b0 ;
  assign n5760 = n5759 ^ n981 ^ 1'b0 ;
  assign n5761 = n1080 | n2075 ;
  assign n5762 = n2101 ^ n749 ^ 1'b0 ;
  assign n5763 = n2776 | n5762 ;
  assign n5764 = n4602 ^ n1825 ^ 1'b0 ;
  assign n5765 = ~n1957 & n2308 ;
  assign n5766 = n2948 & n5765 ;
  assign n5767 = n2604 & ~n3952 ;
  assign n5768 = n5766 & n5767 ;
  assign n5769 = n689 | n4147 ;
  assign n5770 = n1002 | n5769 ;
  assign n5771 = n5770 ^ n2942 ^ 1'b0 ;
  assign n5772 = x32 & x94 ;
  assign n5773 = ~x32 & n5772 ;
  assign n5774 = x127 & ~n250 ;
  assign n5775 = n250 & n5774 ;
  assign n5776 = n1080 | n5775 ;
  assign n5777 = n5773 | n5776 ;
  assign n5778 = n5777 ^ n4855 ^ 1'b0 ;
  assign n5779 = n4148 ^ n3112 ^ 1'b0 ;
  assign n5780 = n353 & ~n1645 ;
  assign n5781 = n4888 | n5780 ;
  assign n5782 = n5781 ^ n5291 ^ 1'b0 ;
  assign n5783 = ( x97 & n1552 ) | ( x97 & n4676 ) | ( n1552 & n4676 ) ;
  assign n5784 = ~n577 & n2879 ;
  assign n5785 = ~n2879 & n5784 ;
  assign n5786 = n5317 & ~n5785 ;
  assign n5787 = n5783 & n5786 ;
  assign n5788 = ~n1098 & n3482 ;
  assign n5789 = n5788 ^ x53 ^ 1'b0 ;
  assign n5790 = n3902 & n5789 ;
  assign n5791 = ~n3292 & n5790 ;
  assign n5792 = n433 & ~n2174 ;
  assign n5793 = n5792 ^ n1034 ^ 1'b0 ;
  assign n5794 = n4811 | n5793 ;
  assign n5795 = ~n299 & n4310 ;
  assign n5796 = n5795 ^ n4482 ^ 1'b0 ;
  assign n5800 = ( n1451 & n2295 ) | ( n1451 & n3728 ) | ( n2295 & n3728 ) ;
  assign n5797 = x81 & ~n2450 ;
  assign n5798 = n880 | n5797 ;
  assign n5799 = n4487 & n5798 ;
  assign n5801 = n5800 ^ n5799 ^ 1'b0 ;
  assign n5802 = ( ~n1365 & n4135 ) | ( ~n1365 & n4632 ) | ( n4135 & n4632 ) ;
  assign n5803 = n3482 & ~n5377 ;
  assign n5804 = ~n5802 & n5803 ;
  assign n5805 = x21 & ~n1132 ;
  assign n5806 = n5139 & n5805 ;
  assign n5807 = n5806 ^ n2732 ^ 1'b0 ;
  assign n5808 = n414 & ~n3282 ;
  assign n5809 = ~n365 & n5808 ;
  assign n5810 = n564 & ~n790 ;
  assign n5811 = n1321 & ~n5810 ;
  assign n5812 = n5811 ^ n2501 ^ 1'b0 ;
  assign n5813 = n1069 & ~n5812 ;
  assign n5814 = n4318 & n5813 ;
  assign n5815 = ~n251 & n4267 ;
  assign n5816 = n5815 ^ n638 ^ 1'b0 ;
  assign n5817 = n3876 & n5816 ;
  assign n5818 = n1668 ^ n1030 ^ n700 ;
  assign n5819 = n1474 ^ n444 ^ 1'b0 ;
  assign n5820 = ~n5818 & n5819 ;
  assign n5821 = n5820 ^ n1419 ^ 1'b0 ;
  assign n5822 = n731 ^ x68 ^ 1'b0 ;
  assign n5824 = ~n680 & n2385 ;
  assign n5825 = n5824 ^ n1900 ^ 1'b0 ;
  assign n5823 = x76 & ~n1958 ;
  assign n5826 = n5825 ^ n5823 ^ 1'b0 ;
  assign n5831 = x104 | n356 ;
  assign n5832 = n5831 ^ n2345 ^ 1'b0 ;
  assign n5830 = n336 & n3538 ;
  assign n5833 = n5832 ^ n5830 ^ 1'b0 ;
  assign n5827 = x118 & ~n753 ;
  assign n5828 = n5827 ^ x94 ^ 1'b0 ;
  assign n5829 = n5828 ^ n192 ^ 1'b0 ;
  assign n5834 = n5833 ^ n5829 ^ n3714 ;
  assign n5835 = ~n2759 & n2957 ;
  assign n5836 = n3683 & n5835 ;
  assign n5837 = n869 ^ n279 ^ 1'b0 ;
  assign n5838 = n2601 | n3706 ;
  assign n5839 = n1249 | n1366 ;
  assign n5840 = n5839 ^ n1861 ^ 1'b0 ;
  assign n5841 = n3320 ^ n394 ^ 1'b0 ;
  assign n5842 = n2738 & ~n5841 ;
  assign n5843 = n344 | n1663 ;
  assign n5844 = n5843 ^ n2491 ^ 1'b0 ;
  assign n5845 = n4296 | n5844 ;
  assign n5846 = ~n2299 & n5845 ;
  assign n5847 = n5846 ^ n3010 ^ 1'b0 ;
  assign n5848 = n5847 ^ n5453 ^ 1'b0 ;
  assign n5849 = ~n4597 & n5848 ;
  assign n5850 = n5849 ^ n3074 ^ 1'b0 ;
  assign n5851 = ~n568 & n1209 ;
  assign n5852 = n5851 ^ n1290 ^ 1'b0 ;
  assign n5853 = n5852 ^ n851 ^ 1'b0 ;
  assign n5854 = n5850 & n5853 ;
  assign n5855 = n3664 ^ n2360 ^ 1'b0 ;
  assign n5856 = n3348 ^ n531 ^ 1'b0 ;
  assign n5857 = n3702 & ~n5856 ;
  assign n5858 = n2196 ^ n1508 ^ 1'b0 ;
  assign n5859 = n792 & ~n5858 ;
  assign n5860 = ( ~n2049 & n2882 ) | ( ~n2049 & n2903 ) | ( n2882 & n2903 ) ;
  assign n5861 = n1707 & n5860 ;
  assign n5862 = ( ~n4314 & n5859 ) | ( ~n4314 & n5861 ) | ( n5859 & n5861 ) ;
  assign n5863 = n2432 ^ n2166 ^ 1'b0 ;
  assign n5864 = ( n924 & n5525 ) | ( n924 & n5863 ) | ( n5525 & n5863 ) ;
  assign n5865 = n5336 | n5864 ;
  assign n5866 = n4151 & n4503 ;
  assign n5867 = ~n1616 & n2696 ;
  assign n5868 = ~n2682 & n3192 ;
  assign n5869 = n2242 | n4350 ;
  assign n5870 = n5868 | n5869 ;
  assign n5871 = ~n3156 & n5870 ;
  assign n5872 = n1861 & ~n2889 ;
  assign n5873 = n2215 & n5872 ;
  assign n5874 = ~n5094 & n5873 ;
  assign n5875 = n950 ^ n811 ^ 1'b0 ;
  assign n5876 = n3732 ^ x62 ^ 1'b0 ;
  assign n5877 = n4503 ^ n1502 ^ 1'b0 ;
  assign n5878 = x1 & n5877 ;
  assign n5879 = n3232 ^ n2399 ^ 1'b0 ;
  assign n5880 = n5879 ^ n2911 ^ 1'b0 ;
  assign n5881 = n2156 & n2257 ;
  assign n5882 = ~n4304 & n5881 ;
  assign n5883 = n3446 ^ n897 ^ 1'b0 ;
  assign n5884 = n2675 ^ n707 ^ 1'b0 ;
  assign n5885 = n5883 | n5884 ;
  assign n5886 = n3916 & ~n5885 ;
  assign n5887 = n5886 ^ n1766 ^ n1295 ;
  assign n5888 = ( n481 & n810 ) | ( n481 & ~n2604 ) | ( n810 & ~n2604 ) ;
  assign n5889 = n2446 & ~n5888 ;
  assign n5890 = ~n820 & n5150 ;
  assign n5891 = n4729 & n5878 ;
  assign n5893 = n3754 ^ n1214 ^ n962 ;
  assign n5892 = n2967 & ~n3613 ;
  assign n5894 = n5893 ^ n5892 ^ 1'b0 ;
  assign n5895 = n2921 | n5365 ;
  assign n5896 = n314 & n5895 ;
  assign n5897 = n5896 ^ n1972 ^ 1'b0 ;
  assign n5898 = n510 & n1452 ;
  assign n5899 = n638 | n5503 ;
  assign n5900 = n5898 & n5899 ;
  assign n5901 = ~n2709 & n4356 ;
  assign n5902 = ~x79 & n5901 ;
  assign n5903 = n2026 | n5902 ;
  assign n5904 = n5438 ^ n1786 ^ 1'b0 ;
  assign n5905 = n717 | n3952 ;
  assign n5906 = n717 & ~n5905 ;
  assign n5907 = ( ~n3544 & n3846 ) | ( ~n3544 & n5906 ) | ( n3846 & n5906 ) ;
  assign n5908 = n5907 ^ n1472 ^ 1'b0 ;
  assign n5909 = n1909 & ~n5908 ;
  assign n5910 = n5708 ^ n3080 ^ 1'b0 ;
  assign n5911 = n5910 ^ n5797 ^ 1'b0 ;
  assign n5912 = n5055 & ~n5911 ;
  assign n5913 = n861 & ~n2312 ;
  assign n5914 = x48 & ~n614 ;
  assign n5915 = n614 & n5914 ;
  assign n5916 = n5915 ^ n3656 ^ 1'b0 ;
  assign n5917 = n1244 | n5916 ;
  assign n5918 = n5913 & ~n5917 ;
  assign n5919 = ~x75 & n5909 ;
  assign n5920 = ~n3721 & n5919 ;
  assign n5921 = n3514 ^ x125 ^ x88 ;
  assign n5922 = n2306 & n5921 ;
  assign n5923 = n4582 & n5922 ;
  assign n5924 = n1115 & n5413 ;
  assign n5925 = ~n1694 & n2354 ;
  assign n5926 = n5925 ^ n1588 ^ 1'b0 ;
  assign n5927 = n750 ^ n725 ^ 1'b0 ;
  assign n5928 = n608 & ~n5927 ;
  assign n5929 = ~n814 & n5928 ;
  assign n5930 = n5929 ^ n2091 ^ 1'b0 ;
  assign n5931 = n343 & ~n5930 ;
  assign n5932 = n4064 & ~n5719 ;
  assign n5933 = n5932 ^ n724 ^ 1'b0 ;
  assign n5934 = n4524 ^ n3733 ^ 1'b0 ;
  assign n5935 = n5154 & ~n5934 ;
  assign n5936 = n825 ^ n314 ^ 1'b0 ;
  assign n5937 = n308 & n5936 ;
  assign n5938 = ( n607 & n639 ) | ( n607 & ~n5937 ) | ( n639 & ~n5937 ) ;
  assign n5939 = n1622 ^ n1122 ^ 1'b0 ;
  assign n5940 = n2529 | n5939 ;
  assign n5941 = n3754 ^ n165 ^ 1'b0 ;
  assign n5942 = n1905 & ~n5941 ;
  assign n5943 = ~n5940 & n5942 ;
  assign n5944 = n3615 ^ n294 ^ 1'b0 ;
  assign n5945 = x127 ^ x83 ^ 1'b0 ;
  assign n5946 = n296 | n5945 ;
  assign n5947 = n830 | n1482 ;
  assign n5948 = n3468 ^ n487 ^ 1'b0 ;
  assign n5949 = n2201 & ~n5948 ;
  assign n5950 = n315 & n5949 ;
  assign n5951 = n3789 | n4177 ;
  assign n5952 = n2297 ^ n1957 ^ 1'b0 ;
  assign n5953 = n3575 & n5952 ;
  assign n5954 = n1065 | n5953 ;
  assign n5955 = n5954 ^ n3019 ^ 1'b0 ;
  assign n5956 = n237 & ~n5955 ;
  assign n5957 = n5159 & n5387 ;
  assign n5958 = n5957 ^ n5437 ^ 1'b0 ;
  assign n5961 = ~n2107 & n2517 ;
  assign n5962 = n1888 | n5961 ;
  assign n5959 = ~n355 & n4674 ;
  assign n5960 = n3615 | n5959 ;
  assign n5963 = n5962 ^ n5960 ^ 1'b0 ;
  assign n5964 = n2266 & ~n5963 ;
  assign n5965 = n5964 ^ n4215 ^ 1'b0 ;
  assign n5966 = n2598 ^ n820 ^ 1'b0 ;
  assign n5971 = ( n487 & ~n2811 ) | ( n487 & n3498 ) | ( ~n2811 & n3498 ) ;
  assign n5972 = n5971 ^ n3782 ^ 1'b0 ;
  assign n5967 = ~n882 & n965 ;
  assign n5968 = n3247 & ~n5967 ;
  assign n5969 = n5968 ^ n2608 ^ 1'b0 ;
  assign n5970 = n3218 & ~n5969 ;
  assign n5973 = n5972 ^ n5970 ^ 1'b0 ;
  assign n5974 = n2006 & ~n4412 ;
  assign n5975 = n1939 | n5242 ;
  assign n5976 = n2885 ^ n636 ^ 1'b0 ;
  assign n5977 = n851 | n5976 ;
  assign n5978 = n2213 ^ n1383 ^ 1'b0 ;
  assign n5979 = n1894 & ~n5978 ;
  assign n5980 = n2535 & ~n4443 ;
  assign n5981 = n1211 & ~n4074 ;
  assign n5982 = n4126 ^ n387 ^ 1'b0 ;
  assign n5983 = n846 & n5982 ;
  assign n5984 = n5983 ^ n2564 ^ 1'b0 ;
  assign n5985 = n5245 ^ n3257 ^ 1'b0 ;
  assign n5986 = ~n2979 & n5985 ;
  assign n5987 = n492 | n1640 ;
  assign n5988 = n207 | n1270 ;
  assign n5989 = n5988 ^ n2733 ^ 1'b0 ;
  assign n5990 = n531 | n5989 ;
  assign n5991 = n245 | n2635 ;
  assign n5992 = n5991 ^ n3264 ^ 1'b0 ;
  assign n5993 = n1312 & ~n5992 ;
  assign n5994 = n5990 & n5993 ;
  assign n5995 = n5994 ^ n896 ^ 1'b0 ;
  assign n5996 = ~n5987 & n5995 ;
  assign n5997 = ~n1292 & n3480 ;
  assign n5998 = n4146 & n5997 ;
  assign n5999 = n5998 ^ n378 ^ 1'b0 ;
  assign n6000 = n5418 & ~n5999 ;
  assign n6001 = ~n2109 & n6000 ;
  assign n6002 = n972 & ~n2321 ;
  assign n6003 = n2227 & ~n6002 ;
  assign n6004 = n6003 ^ n1897 ^ 1'b0 ;
  assign n6009 = n1838 ^ n1493 ^ 1'b0 ;
  assign n6010 = n4163 & ~n6009 ;
  assign n6011 = n6010 ^ n962 ^ 1'b0 ;
  assign n6005 = n2951 ^ x108 ^ 1'b0 ;
  assign n6006 = n1470 & n6005 ;
  assign n6007 = n6006 ^ n1733 ^ 1'b0 ;
  assign n6008 = n3846 & n6007 ;
  assign n6012 = n6011 ^ n6008 ^ 1'b0 ;
  assign n6013 = n203 & ~n5447 ;
  assign n6014 = n6013 ^ n1093 ^ 1'b0 ;
  assign n6015 = n1049 | n6014 ;
  assign n6016 = n6015 ^ n1861 ^ 1'b0 ;
  assign n6017 = n1534 | n3075 ;
  assign n6018 = ~n584 & n1758 ;
  assign n6019 = ~n3461 & n4106 ;
  assign n6020 = n5819 ^ n4638 ^ 1'b0 ;
  assign n6022 = n1737 ^ n970 ^ 1'b0 ;
  assign n6021 = ~n1561 & n4946 ;
  assign n6023 = n6022 ^ n6021 ^ 1'b0 ;
  assign n6024 = n430 | n2047 ;
  assign n6025 = n3764 ^ n707 ^ 1'b0 ;
  assign n6026 = ~n397 & n6025 ;
  assign n6027 = n6024 & n6026 ;
  assign n6028 = n2804 ^ n782 ^ 1'b0 ;
  assign n6029 = n6028 ^ n3611 ^ 1'b0 ;
  assign n6030 = n1380 & n6029 ;
  assign n6031 = n828 ^ n288 ^ 1'b0 ;
  assign n6032 = n3409 & ~n6031 ;
  assign n6033 = n6032 ^ n2854 ^ 1'b0 ;
  assign n6034 = n2070 & ~n6033 ;
  assign n6035 = n4608 ^ n1950 ^ 1'b0 ;
  assign n6036 = n6034 & n6035 ;
  assign n6037 = ~n390 & n494 ;
  assign n6038 = n6037 ^ n5527 ^ n4271 ;
  assign n6039 = n6038 ^ n2289 ^ n493 ;
  assign n6040 = n6039 ^ n2512 ^ 1'b0 ;
  assign n6041 = n2091 & n6040 ;
  assign n6044 = n3180 & n3758 ;
  assign n6042 = ~n3583 & n4051 ;
  assign n6043 = n1983 | n6042 ;
  assign n6045 = n6044 ^ n6043 ^ 1'b0 ;
  assign n6046 = n2486 & ~n3541 ;
  assign n6047 = n200 | n250 ;
  assign n6048 = n1317 | n2606 ;
  assign n6049 = n5689 ^ n510 ^ 1'b0 ;
  assign n6050 = n6048 & n6049 ;
  assign n6053 = n2123 ^ n531 ^ 1'b0 ;
  assign n6051 = n1630 | n5416 ;
  assign n6052 = n2065 & ~n6051 ;
  assign n6054 = n6053 ^ n6052 ^ 1'b0 ;
  assign n6056 = x99 & ~n1349 ;
  assign n6055 = n2633 & ~n3244 ;
  assign n6057 = n6056 ^ n6055 ^ n3580 ;
  assign n6061 = n4652 ^ n502 ^ 1'b0 ;
  assign n6058 = n3450 & ~n3551 ;
  assign n6059 = n930 & n6058 ;
  assign n6060 = n185 | n6059 ;
  assign n6062 = n6061 ^ n6060 ^ 1'b0 ;
  assign n6063 = n725 & n742 ;
  assign n6064 = n3257 | n6063 ;
  assign n6065 = ( n1556 & n3573 ) | ( n1556 & n4298 ) | ( n3573 & n4298 ) ;
  assign n6066 = n499 | n2591 ;
  assign n6067 = n6065 | n6066 ;
  assign n6068 = n562 & ~n5522 ;
  assign n6069 = n886 & n6068 ;
  assign n6070 = n4454 ^ n3462 ^ n928 ;
  assign n6071 = n3354 | n3966 ;
  assign n6073 = n724 ^ x27 ^ 1'b0 ;
  assign n6072 = x5 & ~n3981 ;
  assign n6074 = n6073 ^ n6072 ^ 1'b0 ;
  assign n6075 = n2371 | n6074 ;
  assign n6076 = n266 & ~n1293 ;
  assign n6077 = n741 & n6076 ;
  assign n6078 = n3585 & ~n6077 ;
  assign n6079 = ~n4267 & n6078 ;
  assign n6080 = n6079 ^ n3584 ^ 1'b0 ;
  assign n6081 = n4694 ^ n1631 ^ 1'b0 ;
  assign n6082 = n1228 ^ n873 ^ 1'b0 ;
  assign n6083 = n6081 | n6082 ;
  assign n6084 = n497 | n4574 ;
  assign n6085 = n4788 ^ n4464 ^ 1'b0 ;
  assign n6086 = n3335 & n6085 ;
  assign n6087 = n542 & n2687 ;
  assign n6088 = n6087 ^ n1146 ^ 1'b0 ;
  assign n6089 = n870 & n6088 ;
  assign n6090 = n4307 ^ n3439 ^ 1'b0 ;
  assign n6091 = n290 & ~n6090 ;
  assign n6092 = n3105 ^ n946 ^ 1'b0 ;
  assign n6093 = n1939 | n2653 ;
  assign n6094 = n4598 | n6093 ;
  assign n6095 = n156 & ~n1982 ;
  assign n6096 = n1808 | n6095 ;
  assign n6097 = ~n2281 & n3195 ;
  assign n6098 = n3343 & n6097 ;
  assign n6099 = n6098 ^ x58 ^ 1'b0 ;
  assign n6100 = n2385 & n6099 ;
  assign n6101 = n5028 & n6100 ;
  assign n6102 = n830 | n931 ;
  assign n6103 = n1170 & n4397 ;
  assign n6104 = ~n1179 & n6103 ;
  assign n6105 = n3559 & ~n6104 ;
  assign n6106 = n6105 ^ n299 ^ 1'b0 ;
  assign n6107 = n687 ^ x125 ^ 1'b0 ;
  assign n6108 = n1888 & n6107 ;
  assign n6109 = n4193 ^ n2932 ^ 1'b0 ;
  assign n6110 = n3452 & n6109 ;
  assign n6111 = n1407 & n6110 ;
  assign n6112 = n6111 ^ n1371 ^ 1'b0 ;
  assign n6113 = x62 & n1534 ;
  assign n6114 = ~n932 & n6113 ;
  assign n6115 = n1823 | n5442 ;
  assign n6116 = ~n2732 & n6115 ;
  assign n6117 = n1654 | n4892 ;
  assign n6118 = n1126 & ~n1857 ;
  assign n6119 = n6118 ^ n2266 ^ 1'b0 ;
  assign n6120 = n4592 | n6119 ;
  assign n6121 = n6120 ^ n1957 ^ 1'b0 ;
  assign n6122 = x52 & n346 ;
  assign n6123 = n4217 & ~n6122 ;
  assign n6124 = n6123 ^ n2828 ^ 1'b0 ;
  assign n6125 = x2 | n566 ;
  assign n6126 = x66 | n6125 ;
  assign n6127 = ~n1226 & n6126 ;
  assign n6128 = n6127 ^ n4559 ^ 1'b0 ;
  assign n6129 = ~n6124 & n6128 ;
  assign n6130 = n5825 ^ n3053 ^ 1'b0 ;
  assign n6131 = n4821 & ~n6130 ;
  assign n6132 = n2565 & ~n5115 ;
  assign n6133 = x43 & ~n1048 ;
  assign n6134 = ~x43 & n6133 ;
  assign n6135 = x39 & ~n6134 ;
  assign n6136 = ~x39 & n6135 ;
  assign n6137 = x92 & ~n6136 ;
  assign n6138 = n6136 & n6137 ;
  assign n6139 = ~n1423 & n2266 ;
  assign n6140 = ~n2266 & n6139 ;
  assign n6141 = n6138 | n6140 ;
  assign n6142 = n6138 & ~n6141 ;
  assign n6143 = n2849 ^ n754 ^ 1'b0 ;
  assign n6144 = n1472 | n6143 ;
  assign n6145 = n4311 ^ n444 ^ 1'b0 ;
  assign n6146 = n6145 ^ n1161 ^ 1'b0 ;
  assign n6147 = ~n4282 & n6146 ;
  assign n6148 = n420 & n3865 ;
  assign n6149 = n6148 ^ n2373 ^ 1'b0 ;
  assign n6150 = n1975 | n3195 ;
  assign n6151 = n6150 ^ n3544 ^ 1'b0 ;
  assign n6152 = n6151 ^ n4904 ^ 1'b0 ;
  assign n6153 = ~n268 & n6152 ;
  assign n6154 = ~n702 & n2012 ;
  assign n6155 = ~n375 & n6154 ;
  assign n6157 = n240 & n1833 ;
  assign n6158 = n1314 & n6157 ;
  assign n6156 = n4041 ^ n1788 ^ 1'b0 ;
  assign n6159 = n6158 ^ n6156 ^ 1'b0 ;
  assign n6160 = n1035 & n4271 ;
  assign n6161 = ~n2892 & n6160 ;
  assign n6162 = n6161 ^ n3812 ^ 1'b0 ;
  assign n6163 = n3188 ^ n3035 ^ 1'b0 ;
  assign n6164 = n6163 ^ n5638 ^ 1'b0 ;
  assign n6165 = n2476 ^ n1188 ^ 1'b0 ;
  assign n6166 = n2743 | n6165 ;
  assign n6169 = x36 & ~n945 ;
  assign n6170 = n6169 ^ n485 ^ 1'b0 ;
  assign n6167 = n502 | n884 ;
  assign n6168 = ~n2512 & n6167 ;
  assign n6171 = n6170 ^ n6168 ^ 1'b0 ;
  assign n6172 = n1297 | n3840 ;
  assign n6173 = n4661 & ~n6172 ;
  assign n6174 = n1920 & ~n6173 ;
  assign n6175 = n6174 ^ n4574 ^ 1'b0 ;
  assign n6176 = n604 | n3121 ;
  assign n6177 = n5844 & n6176 ;
  assign n6178 = n6177 ^ n5870 ^ 1'b0 ;
  assign n6179 = n3262 ^ n839 ^ 1'b0 ;
  assign n6180 = n978 & n6179 ;
  assign n6181 = n6180 ^ n2687 ^ n613 ;
  assign n6182 = n768 & n6009 ;
  assign n6183 = n6181 | n6182 ;
  assign n6184 = n1970 | n6183 ;
  assign n6185 = n3717 & n6184 ;
  assign n6186 = n6185 ^ x23 ^ 1'b0 ;
  assign n6187 = n2570 | n5351 ;
  assign n6188 = n6187 ^ n3549 ^ 1'b0 ;
  assign n6189 = n1857 ^ n1275 ^ 1'b0 ;
  assign n6190 = n1901 & ~n2121 ;
  assign n6191 = n5404 & n6190 ;
  assign n6192 = n6189 & n6191 ;
  assign n6193 = ~n1601 & n1815 ;
  assign n6194 = n3715 ^ n2718 ^ n652 ;
  assign n6195 = ~n2096 & n6194 ;
  assign n6196 = n6195 ^ n978 ^ 1'b0 ;
  assign n6197 = ~n3319 & n6196 ;
  assign n6199 = x104 ^ x75 ^ 1'b0 ;
  assign n6200 = n6199 ^ n4571 ^ 1'b0 ;
  assign n6201 = n1316 & ~n6200 ;
  assign n6202 = ~n2759 & n6201 ;
  assign n6203 = n6202 ^ n1726 ^ 1'b0 ;
  assign n6204 = n2634 | n6203 ;
  assign n6205 = n6204 ^ n970 ^ 1'b0 ;
  assign n6198 = n3865 & ~n5097 ;
  assign n6206 = n6205 ^ n6198 ^ 1'b0 ;
  assign n6207 = ~n4037 & n4659 ;
  assign n6208 = n3702 ^ n2161 ^ 1'b0 ;
  assign n6210 = n1630 | n2395 ;
  assign n6209 = n2315 & n3868 ;
  assign n6211 = n6210 ^ n6209 ^ 1'b0 ;
  assign n6212 = n4197 ^ n2852 ^ 1'b0 ;
  assign n6213 = n1328 | n3788 ;
  assign n6214 = ~n5000 & n5551 ;
  assign n6215 = n6214 ^ n4163 ^ 1'b0 ;
  assign n6216 = n3823 & n6215 ;
  assign n6217 = ~n6213 & n6216 ;
  assign n6218 = n3165 ^ n2478 ^ 1'b0 ;
  assign n6219 = n5731 | n6218 ;
  assign n6220 = n6219 ^ n5059 ^ n2241 ;
  assign n6221 = n4100 ^ n375 ^ 1'b0 ;
  assign n6222 = n6221 ^ n5613 ^ 1'b0 ;
  assign n6223 = x90 | n1945 ;
  assign n6224 = x31 | n4788 ;
  assign n6225 = n1478 & ~n3592 ;
  assign n6226 = n1163 | n6225 ;
  assign n6227 = n3198 ^ n211 ^ 1'b0 ;
  assign n6228 = n2815 | n3266 ;
  assign n6229 = n1642 | n6228 ;
  assign n6230 = n731 | n6229 ;
  assign n6231 = n6230 ^ n1329 ^ 1'b0 ;
  assign n6232 = n4998 & n6231 ;
  assign n6233 = ~n3721 & n6232 ;
  assign n6234 = n3059 | n3656 ;
  assign n6235 = n2246 & ~n4361 ;
  assign n6236 = n6234 & ~n6235 ;
  assign n6237 = n3253 ^ n2999 ^ 1'b0 ;
  assign n6238 = x75 & n800 ;
  assign n6239 = n6238 ^ n571 ^ 1'b0 ;
  assign n6240 = n4202 ^ n245 ^ 1'b0 ;
  assign n6241 = n1689 & ~n2216 ;
  assign n6242 = n2176 | n2574 ;
  assign n6243 = ~x66 & n3687 ;
  assign n6244 = ~n576 & n6243 ;
  assign n6245 = n526 | n6244 ;
  assign n6246 = n6245 ^ n1930 ^ 1'b0 ;
  assign n6247 = ~n6114 & n6246 ;
  assign n6248 = n1784 ^ n478 ^ 1'b0 ;
  assign n6249 = x73 & ~n6248 ;
  assign n6250 = n3320 | n6249 ;
  assign n6251 = n6250 ^ n1724 ^ 1'b0 ;
  assign n6252 = n2204 | n4911 ;
  assign n6253 = n198 & n3422 ;
  assign n6254 = n6252 | n6253 ;
  assign n6255 = n2996 | n6254 ;
  assign n6256 = n6255 ^ n2241 ^ 1'b0 ;
  assign n6257 = n2129 | n5596 ;
  assign n6258 = n6257 ^ n893 ^ 1'b0 ;
  assign n6259 = n6258 ^ n2087 ^ 1'b0 ;
  assign n6260 = n2821 ^ n1816 ^ 1'b0 ;
  assign n6261 = ~n2961 & n5410 ;
  assign n6262 = n2445 ^ n430 ^ 1'b0 ;
  assign n6263 = n5317 & ~n6262 ;
  assign n6264 = n4370 ^ n4183 ^ 1'b0 ;
  assign n6265 = n2649 & n6264 ;
  assign n6266 = n1632 & ~n6265 ;
  assign n6267 = n6266 ^ n2895 ^ 1'b0 ;
  assign n6268 = n694 & ~n6267 ;
  assign n6269 = n2395 & n3784 ;
  assign n6270 = n6269 ^ n216 ^ 1'b0 ;
  assign n6271 = n315 | n2148 ;
  assign n6272 = ( n672 & n4648 ) | ( n672 & n6271 ) | ( n4648 & n6271 ) ;
  assign n6273 = ~n2430 & n2851 ;
  assign n6274 = ~n538 & n6273 ;
  assign n6275 = n620 | n6274 ;
  assign n6276 = n2911 | n6275 ;
  assign n6277 = n6276 ^ n2942 ^ 1'b0 ;
  assign n6278 = n4217 & ~n6277 ;
  assign n6279 = ~n1868 & n3086 ;
  assign n6280 = ~n2068 & n6279 ;
  assign n6281 = n1636 & ~n6280 ;
  assign n6282 = n1064 & ~n1163 ;
  assign n6283 = n6282 ^ n1030 ^ 1'b0 ;
  assign n6285 = n992 & ~n4282 ;
  assign n6284 = n1415 | n1484 ;
  assign n6286 = n6285 ^ n6284 ^ 1'b0 ;
  assign n6287 = n3215 ^ n1861 ^ 1'b0 ;
  assign n6288 = n3097 | n6287 ;
  assign n6292 = n4636 | n5450 ;
  assign n6293 = n2012 | n6292 ;
  assign n6289 = n4671 ^ n1841 ^ n250 ;
  assign n6290 = n3353 ^ n1293 ^ 1'b0 ;
  assign n6291 = ~n6289 & n6290 ;
  assign n6294 = n6293 ^ n6291 ^ 1'b0 ;
  assign n6298 = n558 & n796 ;
  assign n6295 = n518 | n3838 ;
  assign n6296 = n2581 & ~n6295 ;
  assign n6297 = n3723 & ~n6296 ;
  assign n6299 = n6298 ^ n6297 ^ 1'b0 ;
  assign n6300 = n415 & n3803 ;
  assign n6301 = n6300 ^ n1427 ^ 1'b0 ;
  assign n6302 = n1714 & n1947 ;
  assign n6303 = n1631 & n6302 ;
  assign n6304 = ( n4048 & ~n6301 ) | ( n4048 & n6303 ) | ( ~n6301 & n6303 ) ;
  assign n6305 = n6304 ^ n261 ^ 1'b0 ;
  assign n6306 = ~n2436 & n6305 ;
  assign n6307 = n2224 ^ n1008 ^ 1'b0 ;
  assign n6308 = ~n4738 & n5360 ;
  assign n6309 = ~n1829 & n6308 ;
  assign n6310 = n1464 ^ n242 ^ 1'b0 ;
  assign n6311 = n6310 ^ n237 ^ 1'b0 ;
  assign n6312 = n6311 ^ n2013 ^ 1'b0 ;
  assign n6313 = ~n5101 & n6312 ;
  assign n6314 = n320 & ~n717 ;
  assign n6315 = n6002 & n6314 ;
  assign n6316 = n6182 | n6315 ;
  assign n6317 = n6316 ^ n5527 ^ 1'b0 ;
  assign n6318 = n3204 ^ n1842 ^ 1'b0 ;
  assign n6319 = ( n1480 & n2491 ) | ( n1480 & ~n2659 ) | ( n2491 & ~n2659 ) ;
  assign n6320 = n5050 & n6206 ;
  assign n6321 = n920 ^ n167 ^ 1'b0 ;
  assign n6322 = ( n2459 & ~n4579 ) | ( n2459 & n6214 ) | ( ~n4579 & n6214 ) ;
  assign n6323 = n2241 | n5408 ;
  assign n6324 = n6323 ^ n3195 ^ 1'b0 ;
  assign n6325 = ~n2661 & n3289 ;
  assign n6326 = x27 & n6325 ;
  assign n6327 = ~n799 & n2638 ;
  assign n6328 = ~n6326 & n6327 ;
  assign n6329 = ~n2307 & n2800 ;
  assign n6330 = ~n4494 & n6329 ;
  assign n6331 = n1680 & n1842 ;
  assign n6332 = n6331 ^ n4430 ^ 1'b0 ;
  assign n6333 = ~n4521 & n6332 ;
  assign n6334 = n3496 & n4769 ;
  assign n6335 = ~n6333 & n6334 ;
  assign n6336 = ~n328 & n2780 ;
  assign n6337 = n2047 ^ n1328 ^ 1'b0 ;
  assign n6338 = n2554 & ~n3195 ;
  assign n6339 = n6338 ^ n6304 ^ 1'b0 ;
  assign n6340 = n6337 & n6339 ;
  assign n6341 = n3893 ^ n1798 ^ 1'b0 ;
  assign n6347 = n731 & ~n1793 ;
  assign n6348 = ~n205 & n6347 ;
  assign n6343 = n612 & n1829 ;
  assign n6342 = n519 | n1537 ;
  assign n6344 = n6343 ^ n6342 ^ 1'b0 ;
  assign n6345 = ~n5151 & n6344 ;
  assign n6346 = n4364 & n6345 ;
  assign n6349 = n6348 ^ n6346 ^ 1'b0 ;
  assign n6350 = n2961 & n6349 ;
  assign n6351 = x75 | n3464 ;
  assign n6352 = n6351 ^ n1504 ^ 1'b0 ;
  assign n6353 = n2948 & ~n4796 ;
  assign n6354 = n932 & ~n6353 ;
  assign n6355 = ~n859 & n6354 ;
  assign n6356 = n6352 & ~n6355 ;
  assign n6357 = n129 & n6356 ;
  assign n6358 = n1321 & n3671 ;
  assign n6359 = ~n721 & n5289 ;
  assign n6360 = n6359 ^ n614 ^ 1'b0 ;
  assign n6361 = n1816 & ~n4296 ;
  assign n6362 = ~n745 & n3884 ;
  assign n6364 = n2710 ^ n1226 ^ 1'b0 ;
  assign n6365 = n2091 & ~n6364 ;
  assign n6363 = n2112 | n4631 ;
  assign n6366 = n6365 ^ n6363 ^ 1'b0 ;
  assign n6369 = n3932 ^ n402 ^ n132 ;
  assign n6367 = ( n224 & n230 ) | ( n224 & ~n2603 ) | ( n230 & ~n2603 ) ;
  assign n6368 = n2218 & n6367 ;
  assign n6370 = n6369 ^ n6368 ^ 1'b0 ;
  assign n6371 = n427 | n3581 ;
  assign n6372 = n2384 ^ n293 ^ 1'b0 ;
  assign n6373 = n6371 | n6372 ;
  assign n6375 = n866 | n1363 ;
  assign n6376 = n983 & ~n6375 ;
  assign n6374 = n358 & n1683 ;
  assign n6377 = n6376 ^ n6374 ^ 1'b0 ;
  assign n6383 = n1046 & n2933 ;
  assign n6384 = n6383 ^ n1181 ^ 1'b0 ;
  assign n6378 = n2357 ^ n1071 ^ 1'b0 ;
  assign n6379 = ~n4592 & n6378 ;
  assign n6380 = n859 & ~n1479 ;
  assign n6381 = n6380 ^ n6190 ^ 1'b0 ;
  assign n6382 = n6379 & ~n6381 ;
  assign n6385 = n6384 ^ n6382 ^ 1'b0 ;
  assign n6386 = ~n2363 & n5479 ;
  assign n6387 = n6386 ^ n4727 ^ 1'b0 ;
  assign n6388 = n5970 & ~n6387 ;
  assign n6389 = n2183 ^ n1811 ^ 1'b0 ;
  assign n6390 = n446 & ~n4122 ;
  assign n6391 = n6390 ^ n1699 ^ 1'b0 ;
  assign n6392 = n5395 & n6036 ;
  assign n6393 = n6392 ^ n1470 ^ 1'b0 ;
  assign n6394 = n5483 ^ n5474 ^ 1'b0 ;
  assign n6395 = n952 & ~n1680 ;
  assign n6396 = ~n1470 & n6395 ;
  assign n6397 = n5189 | n6396 ;
  assign n6398 = n2493 & ~n6397 ;
  assign n6399 = n6398 ^ n1959 ^ 1'b0 ;
  assign n6400 = n2136 | n6399 ;
  assign n6401 = ~n1487 & n6400 ;
  assign n6402 = n2887 & n4648 ;
  assign n6403 = ~n3228 & n5491 ;
  assign n6404 = n6403 ^ n824 ^ 1'b0 ;
  assign n6405 = n960 | n4095 ;
  assign n6406 = n6405 ^ n931 ^ n512 ;
  assign n6407 = n4515 ^ n1625 ^ 1'b0 ;
  assign n6408 = n1872 & ~n6407 ;
  assign n6409 = n978 | n1176 ;
  assign n6410 = n6409 ^ n2028 ^ 1'b0 ;
  assign n6411 = ~n1934 & n5345 ;
  assign n6412 = n6411 ^ n385 ^ 1'b0 ;
  assign n6413 = ~n1345 & n6412 ;
  assign n6414 = n6410 & n6413 ;
  assign n6416 = n911 ^ n428 ^ 1'b0 ;
  assign n6417 = n753 | n6416 ;
  assign n6415 = n259 | n5469 ;
  assign n6418 = n6417 ^ n6415 ^ 1'b0 ;
  assign n6419 = n2702 ^ n2377 ^ 1'b0 ;
  assign n6420 = n1589 & n2765 ;
  assign n6421 = ( n1401 & ~n2179 ) | ( n1401 & n6420 ) | ( ~n2179 & n6420 ) ;
  assign n6422 = n2191 | n6421 ;
  assign n6423 = n456 & ~n5617 ;
  assign n6424 = n6311 ^ n4858 ^ 1'b0 ;
  assign n6425 = n6423 | n6424 ;
  assign n6426 = n996 ^ n594 ^ 1'b0 ;
  assign n6427 = n5122 & n6426 ;
  assign n6428 = ( n2702 & n3981 ) | ( n2702 & ~n4354 ) | ( n3981 & ~n4354 ) ;
  assign n6429 = n3120 ^ n2603 ^ 1'b0 ;
  assign n6430 = n4077 ^ n2982 ^ 1'b0 ;
  assign n6431 = n6430 ^ n1908 ^ n930 ;
  assign n6432 = n1526 | n6431 ;
  assign n6433 = n5001 ^ n859 ^ 1'b0 ;
  assign n6434 = n2154 ^ n1170 ^ n1048 ;
  assign n6435 = ( ~n620 & n4003 ) | ( ~n620 & n6434 ) | ( n4003 & n6434 ) ;
  assign n6436 = n6435 ^ n1917 ^ n473 ;
  assign n6437 = ~n861 & n5186 ;
  assign n6438 = n6437 ^ n4193 ^ 1'b0 ;
  assign n6439 = n1702 ^ x30 ^ 1'b0 ;
  assign n6440 = ~n3977 & n6439 ;
  assign n6441 = n6438 & n6440 ;
  assign n6442 = n2323 & ~n3931 ;
  assign n6443 = n1782 ^ n1552 ^ 1'b0 ;
  assign n6444 = ~n2746 & n6443 ;
  assign n6445 = n3090 ^ x43 ^ 1'b0 ;
  assign n6446 = ~n4288 & n4823 ;
  assign n6447 = n739 & n6446 ;
  assign n6448 = n6447 ^ n5890 ^ n4052 ;
  assign n6449 = n1443 & ~n3262 ;
  assign n6453 = n2852 ^ n2771 ^ 1'b0 ;
  assign n6454 = n6453 ^ n3635 ^ 1'b0 ;
  assign n6450 = n4102 & n5425 ;
  assign n6451 = n6450 ^ n1732 ^ 1'b0 ;
  assign n6452 = ~n1222 & n6451 ;
  assign n6455 = n6454 ^ n6452 ^ 1'b0 ;
  assign n6456 = n4014 ^ n1537 ^ 1'b0 ;
  assign n6457 = ( n991 & n4746 ) | ( n991 & ~n6456 ) | ( n4746 & ~n6456 ) ;
  assign n6458 = n2107 ^ n1212 ^ 1'b0 ;
  assign n6459 = n735 | n945 ;
  assign n6460 = ( n2343 & ~n6458 ) | ( n2343 & n6459 ) | ( ~n6458 & n6459 ) ;
  assign n6461 = n3083 ^ n1361 ^ x54 ;
  assign n6462 = n6461 ^ n1321 ^ 1'b0 ;
  assign n6463 = n5376 & ~n6462 ;
  assign n6464 = n6463 ^ n1992 ^ 1'b0 ;
  assign n6465 = ~n6348 & n6464 ;
  assign n6466 = ~n4158 & n6465 ;
  assign n6467 = ~n6460 & n6466 ;
  assign n6468 = n1579 & n3244 ;
  assign n6469 = n6468 ^ n165 ^ 1'b0 ;
  assign n6470 = n2010 & n6217 ;
  assign n6471 = n690 & ~n6070 ;
  assign n6472 = n1167 ^ x32 ^ 1'b0 ;
  assign n6473 = n1342 & ~n6472 ;
  assign n6474 = n6473 ^ n1308 ^ 1'b0 ;
  assign n6475 = n6474 ^ n1905 ^ 1'b0 ;
  assign n6476 = n2704 | n6475 ;
  assign n6479 = ~n1102 & n1446 ;
  assign n6480 = n4994 & n6479 ;
  assign n6477 = n4996 ^ n359 ^ 1'b0 ;
  assign n6478 = n420 & n6477 ;
  assign n6481 = n6480 ^ n6478 ^ 1'b0 ;
  assign n6482 = n6476 | n6481 ;
  assign n6483 = n339 & ~n2827 ;
  assign n6484 = n6483 ^ n4647 ^ 1'b0 ;
  assign n6485 = n5475 & n6484 ;
  assign n6486 = n1974 ^ x84 ^ 1'b0 ;
  assign n6487 = n4222 ^ n131 ^ 1'b0 ;
  assign n6488 = ~n2624 & n6487 ;
  assign n6489 = n261 & ~n5876 ;
  assign n6490 = n4579 & n6489 ;
  assign n6491 = n6490 ^ n1179 ^ 1'b0 ;
  assign n6492 = n6488 & n6491 ;
  assign n6493 = n2808 ^ n1430 ^ 1'b0 ;
  assign n6494 = n3604 & ~n4141 ;
  assign n6495 = n614 | n3789 ;
  assign n6496 = n6212 ^ n5689 ^ 1'b0 ;
  assign n6497 = n5367 ^ x78 ^ 1'b0 ;
  assign n6504 = n2366 ^ n570 ^ 1'b0 ;
  assign n6501 = n2560 ^ n473 ^ 1'b0 ;
  assign n6498 = n763 & n1270 ;
  assign n6499 = n6498 ^ n782 ^ 1'b0 ;
  assign n6500 = n3228 | n6499 ;
  assign n6502 = n6501 ^ n6500 ^ 1'b0 ;
  assign n6503 = n3064 & ~n6502 ;
  assign n6505 = n6504 ^ n6503 ^ 1'b0 ;
  assign n6506 = n5632 ^ n277 ^ 1'b0 ;
  assign n6507 = n1664 | n6506 ;
  assign n6508 = n215 | n6095 ;
  assign n6509 = n1989 & ~n5857 ;
  assign n6510 = n3604 | n4143 ;
  assign n6511 = n6510 ^ n939 ^ 1'b0 ;
  assign n6512 = n5548 & n6511 ;
  assign n6513 = n237 & n2385 ;
  assign n6514 = ~n1623 & n6513 ;
  assign n6515 = n6514 ^ n1842 ^ 1'b0 ;
  assign n6516 = n2907 ^ n1107 ^ 1'b0 ;
  assign n6517 = n6515 & ~n6516 ;
  assign n6518 = n2787 & n4567 ;
  assign n6519 = ~n3480 & n6518 ;
  assign n6520 = n640 & ~n6519 ;
  assign n6521 = n2470 | n2488 ;
  assign n6522 = n2408 | n6521 ;
  assign n6523 = ~n4280 & n6522 ;
  assign n6524 = n4449 | n6523 ;
  assign n6525 = n6524 ^ n1240 ^ 1'b0 ;
  assign n6526 = ( n2564 & ~n2985 ) | ( n2564 & n4767 ) | ( ~n2985 & n4767 ) ;
  assign n6527 = n6526 ^ n6026 ^ 1'b0 ;
  assign n6528 = n2293 ^ n720 ^ 1'b0 ;
  assign n6529 = n2598 ^ x108 ^ 1'b0 ;
  assign n6530 = n6528 & ~n6529 ;
  assign n6531 = n5156 ^ n711 ^ 1'b0 ;
  assign n6532 = ~n4177 & n6531 ;
  assign n6533 = n6532 ^ n3477 ^ 1'b0 ;
  assign n6534 = x44 & x120 ;
  assign n6535 = n363 & ~n6534 ;
  assign n6536 = n6535 ^ n425 ^ 1'b0 ;
  assign n6537 = n5068 ^ n3145 ^ 1'b0 ;
  assign n6538 = n6536 | n6537 ;
  assign n6539 = n6538 ^ n884 ^ 1'b0 ;
  assign n6540 = n1135 ^ x107 ^ 1'b0 ;
  assign n6541 = n3772 | n6540 ;
  assign n6542 = n6541 ^ n6522 ^ 1'b0 ;
  assign n6547 = n1245 | n2210 ;
  assign n6543 = ~n330 & n1548 ;
  assign n6544 = n6543 ^ n4635 ^ 1'b0 ;
  assign n6545 = n1630 | n6544 ;
  assign n6546 = n6545 ^ n1918 ^ 1'b0 ;
  assign n6548 = n6547 ^ n6546 ^ 1'b0 ;
  assign n6549 = n6343 & n6548 ;
  assign n6550 = n4929 ^ n2957 ^ 1'b0 ;
  assign n6551 = n2360 | n4727 ;
  assign n6552 = n6551 ^ n1618 ^ 1'b0 ;
  assign n6553 = ~n6550 & n6552 ;
  assign n6554 = n6553 ^ n137 ^ 1'b0 ;
  assign n6555 = n3629 ^ n612 ^ 1'b0 ;
  assign n6556 = n311 & n2687 ;
  assign n6557 = ~n3234 & n6556 ;
  assign n6558 = n5163 ^ n3454 ^ 1'b0 ;
  assign n6559 = n6558 ^ n2198 ^ 1'b0 ;
  assign n6560 = ~n2828 & n4032 ;
  assign n6561 = ~n1077 & n6560 ;
  assign n6562 = n1475 & n6561 ;
  assign n6563 = n1208 ^ n210 ^ 1'b0 ;
  assign n6564 = ~n2839 & n3339 ;
  assign n6565 = n4871 ^ n4457 ^ n1221 ;
  assign n6566 = n6565 ^ n3177 ^ 1'b0 ;
  assign n6567 = n2585 & ~n2693 ;
  assign n6568 = n3312 & n6567 ;
  assign n6569 = n892 & n6568 ;
  assign n6570 = n417 & n4753 ;
  assign n6571 = n5487 ^ n3788 ^ 1'b0 ;
  assign n6572 = n5545 & ~n6571 ;
  assign n6573 = n1632 & ~n6572 ;
  assign n6574 = n6570 | n6573 ;
  assign n6575 = n1772 | n6574 ;
  assign n6576 = n432 & n2884 ;
  assign n6577 = n2306 & ~n6576 ;
  assign n6578 = n6577 ^ n358 ^ 1'b0 ;
  assign n6579 = n1283 ^ n1209 ^ 1'b0 ;
  assign n6580 = n4395 | n6579 ;
  assign n6581 = n2584 & ~n6580 ;
  assign n6582 = n4169 | n6313 ;
  assign n6583 = n2171 | n6257 ;
  assign n6584 = n1428 & ~n4452 ;
  assign n6585 = ~n3824 & n6584 ;
  assign n6586 = n5257 | n6585 ;
  assign n6587 = n6586 ^ n508 ^ 1'b0 ;
  assign n6588 = ~n3526 & n3821 ;
  assign n6589 = n6588 ^ n2123 ^ 1'b0 ;
  assign n6590 = n3906 | n6079 ;
  assign n6591 = n2324 ^ n504 ^ 1'b0 ;
  assign n6592 = n4163 & ~n6591 ;
  assign n6593 = n2604 & ~n3629 ;
  assign n6594 = n6593 ^ n243 ^ 1'b0 ;
  assign n6595 = n6594 ^ x116 ^ 1'b0 ;
  assign n6596 = n6592 & ~n6595 ;
  assign n6597 = n2499 ^ n2293 ^ 1'b0 ;
  assign n6598 = n2486 | n6597 ;
  assign n6599 = ~n961 & n2293 ;
  assign n6600 = ~x7 & n6599 ;
  assign n6601 = n6600 ^ n1401 ^ 1'b0 ;
  assign n6602 = n1070 & n1650 ;
  assign n6603 = n6602 ^ n3401 ^ 1'b0 ;
  assign n6604 = n351 | n6603 ;
  assign n6605 = n3429 & n6604 ;
  assign n6607 = n603 & n1292 ;
  assign n6606 = n1172 & ~n5431 ;
  assign n6608 = n6607 ^ n6606 ^ n6370 ;
  assign n6609 = x4 | n2962 ;
  assign n6610 = n3184 | n6609 ;
  assign n6611 = n6610 ^ n624 ^ 1'b0 ;
  assign n6612 = n4817 & n6611 ;
  assign n6613 = n5938 & ~n6244 ;
  assign n6614 = ~n1495 & n6613 ;
  assign n6615 = ~n373 & n528 ;
  assign n6616 = n6615 ^ n788 ^ 1'b0 ;
  assign n6617 = ~n1443 & n6616 ;
  assign n6618 = ( n1574 & ~n3302 ) | ( n1574 & n6617 ) | ( ~n3302 & n6617 ) ;
  assign n6619 = n4080 ^ n1234 ^ 1'b0 ;
  assign n6620 = x109 & ~n6619 ;
  assign n6621 = ~n4087 & n6620 ;
  assign n6622 = n2650 ^ n1166 ^ 1'b0 ;
  assign n6623 = ( x100 & n2473 ) | ( x100 & n6622 ) | ( n2473 & n6622 ) ;
  assign n6624 = n2974 ^ n2800 ^ 1'b0 ;
  assign n6625 = n3253 | n6624 ;
  assign n6626 = n2344 & ~n6625 ;
  assign n6627 = n5132 ^ n4924 ^ 1'b0 ;
  assign n6628 = n5615 ^ n1551 ^ 1'b0 ;
  assign n6629 = n6627 & ~n6628 ;
  assign n6630 = n1891 | n2166 ;
  assign n6631 = n6630 ^ n1329 ^ 1'b0 ;
  assign n6632 = n2992 & n6631 ;
  assign n6634 = n3184 ^ n2082 ^ 1'b0 ;
  assign n6635 = n5480 | n6634 ;
  assign n6633 = n2233 | n2255 ;
  assign n6636 = n6635 ^ n6633 ^ 1'b0 ;
  assign n6637 = n509 ^ n135 ^ 1'b0 ;
  assign n6638 = ~x106 & n6637 ;
  assign n6639 = n1178 & n6638 ;
  assign n6640 = n6639 ^ n507 ^ 1'b0 ;
  assign n6641 = n6640 ^ n4296 ^ 1'b0 ;
  assign n6642 = n1301 & n6641 ;
  assign n6643 = ( n1703 & n2850 ) | ( n1703 & ~n6642 ) | ( n2850 & ~n6642 ) ;
  assign n6644 = x67 & ~n831 ;
  assign n6645 = n4202 ^ n299 ^ 1'b0 ;
  assign n6646 = ~n5280 & n6645 ;
  assign n6647 = n4448 ^ n3976 ^ 1'b0 ;
  assign n6648 = x125 | n6647 ;
  assign n6649 = n5345 & n6648 ;
  assign n6651 = ( n499 & ~n1129 ) | ( n499 & n3302 ) | ( ~n1129 & n3302 ) ;
  assign n6650 = n996 & ~n4775 ;
  assign n6652 = n6651 ^ n6650 ^ 1'b0 ;
  assign n6653 = n4274 | n4387 ;
  assign n6654 = n211 & ~n6653 ;
  assign n6655 = ~n302 & n6085 ;
  assign n6659 = n2585 ^ n323 ^ 1'b0 ;
  assign n6660 = n847 | n6659 ;
  assign n6656 = n799 | n902 ;
  assign n6657 = n2227 & ~n6656 ;
  assign n6658 = n311 & n6657 ;
  assign n6661 = n6660 ^ n6658 ^ 1'b0 ;
  assign n6662 = ~n2773 & n3794 ;
  assign n6663 = n6661 & n6662 ;
  assign n6664 = n6655 & n6663 ;
  assign n6665 = n215 & ~n2705 ;
  assign n6666 = n2337 & n6665 ;
  assign n6667 = n6666 ^ n894 ^ 1'b0 ;
  assign n6669 = n6579 ^ n1552 ^ 1'b0 ;
  assign n6668 = x48 & ~n1080 ;
  assign n6670 = n6669 ^ n6668 ^ 1'b0 ;
  assign n6671 = n2096 ^ n1163 ^ 1'b0 ;
  assign n6672 = n3398 ^ n790 ^ 1'b0 ;
  assign n6673 = n6671 & ~n6672 ;
  assign n6674 = n3602 | n5991 ;
  assign n6675 = n6674 ^ n4985 ^ 1'b0 ;
  assign n6676 = n4459 & ~n4781 ;
  assign n6677 = n1631 & n6676 ;
  assign n6678 = n5195 ^ n3992 ^ 1'b0 ;
  assign n6679 = n6677 | n6678 ;
  assign n6682 = x3 | n3258 ;
  assign n6683 = n6682 ^ n1558 ^ 1'b0 ;
  assign n6684 = n5562 & ~n6683 ;
  assign n6680 = ~n1934 & n5755 ;
  assign n6681 = n3803 & n6680 ;
  assign n6685 = n6684 ^ n6681 ^ 1'b0 ;
  assign n6686 = n4696 ^ n3130 ^ 1'b0 ;
  assign n6687 = n5258 & n6686 ;
  assign n6688 = n2667 & n3642 ;
  assign n6689 = n6055 | n6369 ;
  assign n6690 = n6688 | n6689 ;
  assign n6691 = n5330 ^ n4122 ^ 1'b0 ;
  assign n6692 = ~n3725 & n6691 ;
  assign n6693 = n1606 & n3234 ;
  assign n6694 = n1060 & n6693 ;
  assign n6695 = n6694 ^ n5814 ^ 1'b0 ;
  assign n6696 = n4385 & n6695 ;
  assign n6697 = n1918 & ~n2037 ;
  assign n6698 = ~n6696 & n6697 ;
  assign n6699 = n1532 ^ n911 ^ 1'b0 ;
  assign n6700 = n6699 ^ n3538 ^ n593 ;
  assign n6701 = n1476 | n6700 ;
  assign n6702 = n5200 | n6701 ;
  assign n6703 = n6702 ^ n5046 ^ 1'b0 ;
  assign n6704 = n1340 ^ n770 ^ 1'b0 ;
  assign n6705 = n1770 & ~n6704 ;
  assign n6706 = n4584 ^ n3665 ^ n2612 ;
  assign n6707 = n623 & ~n6706 ;
  assign n6708 = n6705 & n6707 ;
  assign n6709 = n450 & n1001 ;
  assign n6710 = ~n1737 & n6709 ;
  assign n6711 = n4580 ^ n3186 ^ 1'b0 ;
  assign n6712 = n308 | n469 ;
  assign n6713 = x70 & ~n6712 ;
  assign n6714 = n6713 ^ n666 ^ 1'b0 ;
  assign n6715 = n6714 ^ n222 ^ 1'b0 ;
  assign n6716 = ~n2459 & n6715 ;
  assign n6717 = n459 & ~n6716 ;
  assign n6718 = n6717 ^ n3823 ^ 1'b0 ;
  assign n6719 = n6718 ^ n5302 ^ 1'b0 ;
  assign n6720 = n2711 ^ n519 ^ 1'b0 ;
  assign n6721 = n6181 | n6720 ;
  assign n6722 = n1839 | n5022 ;
  assign n6723 = n6722 ^ n6318 ^ 1'b0 ;
  assign n6724 = n4835 ^ n3764 ^ 1'b0 ;
  assign n6725 = n6723 & ~n6724 ;
  assign n6726 = n3577 ^ n1640 ^ 1'b0 ;
  assign n6727 = n1749 & n2630 ;
  assign n6728 = n6727 ^ n6180 ^ 1'b0 ;
  assign n6729 = ( n392 & ~n3611 ) | ( n392 & n3837 ) | ( ~n3611 & n3837 ) ;
  assign n6730 = n4845 | n6729 ;
  assign n6731 = n3393 & n6296 ;
  assign n6732 = n3419 ^ n1355 ^ n1207 ;
  assign n6733 = n5249 ^ n153 ^ 1'b0 ;
  assign n6734 = ~n3908 & n6733 ;
  assign n6735 = n3428 & n6562 ;
  assign n6736 = ~n965 & n4602 ;
  assign n6737 = n1073 & ~n1935 ;
  assign n6738 = ~n3021 & n6737 ;
  assign n6739 = n5827 ^ n3217 ^ 1'b0 ;
  assign n6740 = ~n252 & n2149 ;
  assign n6741 = n6739 & n6740 ;
  assign n6742 = ~n6739 & n6741 ;
  assign n6743 = n2062 & ~n6742 ;
  assign n6744 = n6743 ^ n5425 ^ 1'b0 ;
  assign n6745 = n5603 ^ n387 ^ 1'b0 ;
  assign n6746 = ~n5367 & n6745 ;
  assign n6747 = n6632 ^ n425 ^ 1'b0 ;
  assign n6748 = n867 | n2321 ;
  assign n6749 = n867 & ~n6748 ;
  assign n6750 = n2673 & n6749 ;
  assign n6751 = n6750 ^ n4393 ^ 1'b0 ;
  assign n6752 = ~n6705 & n6751 ;
  assign n6753 = n6752 ^ n2604 ^ 1'b0 ;
  assign n6754 = n1351 & ~n3950 ;
  assign n6755 = n749 | n761 ;
  assign n6756 = n1843 & ~n6755 ;
  assign n6757 = n6754 & n6756 ;
  assign n6758 = n1064 ^ n896 ^ 1'b0 ;
  assign n6759 = n678 & n6758 ;
  assign n6760 = n3875 & n6759 ;
  assign n6761 = n1315 | n6760 ;
  assign n6762 = n4771 | n6761 ;
  assign n6763 = ~n259 & n6762 ;
  assign n6764 = ~n2606 & n6763 ;
  assign n6765 = x23 & n1635 ;
  assign n6766 = n6765 ^ n2493 ^ 1'b0 ;
  assign n6767 = n6766 ^ n5381 ^ 1'b0 ;
  assign n6768 = n3539 & n6767 ;
  assign n6769 = n6768 ^ n5929 ^ 1'b0 ;
  assign n6771 = n5282 ^ n4338 ^ 1'b0 ;
  assign n6772 = n1904 | n6771 ;
  assign n6770 = n1854 ^ n1808 ^ 1'b0 ;
  assign n6773 = n6772 ^ n6770 ^ 1'b0 ;
  assign n6774 = n3093 ^ n1208 ^ 1'b0 ;
  assign n6775 = n1312 & n6774 ;
  assign n6776 = n6074 & n6775 ;
  assign n6779 = n346 | n461 ;
  assign n6777 = x44 | n2470 ;
  assign n6778 = ~n5527 & n6777 ;
  assign n6780 = n6779 ^ n6778 ^ 1'b0 ;
  assign n6781 = ~n790 & n6003 ;
  assign n6782 = n834 & n6781 ;
  assign n6783 = n4112 | n4616 ;
  assign n6784 = n5548 ^ n1703 ^ 1'b0 ;
  assign n6785 = n6784 ^ n5550 ^ 1'b0 ;
  assign n6786 = n5864 & ~n6785 ;
  assign n6787 = n3396 ^ n597 ^ 1'b0 ;
  assign n6788 = n1624 & ~n6343 ;
  assign n6789 = n1568 ^ n1005 ^ 1'b0 ;
  assign n6790 = ~n3700 & n6789 ;
  assign n6791 = n4330 & ~n4628 ;
  assign n6792 = n6791 ^ n6406 ^ 1'b0 ;
  assign n6793 = ~n2177 & n4560 ;
  assign n6794 = n2026 & ~n3063 ;
  assign n6795 = n501 | n2623 ;
  assign n6796 = n2543 | n6795 ;
  assign n6797 = x73 & ~n277 ;
  assign n6798 = n2761 | n3085 ;
  assign n6799 = n6797 & ~n6798 ;
  assign n6800 = x28 & n2390 ;
  assign n6801 = ~n4193 & n6800 ;
  assign n6802 = n3793 & n6801 ;
  assign n6803 = ( n3650 & n4172 ) | ( n3650 & ~n6802 ) | ( n4172 & ~n6802 ) ;
  assign n6804 = ~n3978 & n4230 ;
  assign n6805 = n6804 ^ n2221 ^ 1'b0 ;
  assign n6806 = ~n686 & n6805 ;
  assign n6807 = n310 & n6806 ;
  assign n6808 = n6807 ^ n2749 ^ 1'b0 ;
  assign n6809 = n396 | n6808 ;
  assign n6810 = n6809 ^ n1830 ^ 1'b0 ;
  assign n6811 = ~n1552 & n6810 ;
  assign n6812 = n2576 & n3894 ;
  assign n6813 = n6812 ^ n1683 ^ 1'b0 ;
  assign n6814 = n4701 ^ n4185 ^ 1'b0 ;
  assign n6815 = n5211 & ~n6814 ;
  assign n6816 = n6815 ^ n1161 ^ 1'b0 ;
  assign n6817 = n3072 | n3969 ;
  assign n6820 = ~n1219 & n4467 ;
  assign n6821 = n6820 ^ n671 ^ 1'b0 ;
  assign n6818 = n210 & n1876 ;
  assign n6819 = n6197 & n6818 ;
  assign n6822 = n6821 ^ n6819 ^ 1'b0 ;
  assign n6823 = n907 | n2543 ;
  assign n6824 = n3161 & ~n6430 ;
  assign n6825 = ( n3280 & n6823 ) | ( n3280 & n6824 ) | ( n6823 & n6824 ) ;
  assign n6826 = n2529 & ~n3680 ;
  assign n6827 = ~n2315 & n6826 ;
  assign n6828 = n137 & ~n2635 ;
  assign n6829 = n6828 ^ n2136 ^ 1'b0 ;
  assign n6830 = x27 & ~n6829 ;
  assign n6831 = n6830 ^ n336 ^ 1'b0 ;
  assign n6832 = n2404 ^ n1986 ^ 1'b0 ;
  assign n6833 = ( ~n307 & n741 ) | ( ~n307 & n5358 ) | ( n741 & n5358 ) ;
  assign n6834 = n5749 ^ n4042 ^ 1'b0 ;
  assign n6835 = n6801 & ~n6834 ;
  assign n6836 = n5736 ^ n3758 ^ 1'b0 ;
  assign n6837 = n1842 & n6836 ;
  assign n6838 = n1659 ^ n1469 ^ 1'b0 ;
  assign n6839 = n3790 & n6838 ;
  assign n6840 = n2251 & n6839 ;
  assign n6841 = n311 & ~n3299 ;
  assign n6842 = ( n600 & n2218 ) | ( n600 & ~n6841 ) | ( n2218 & ~n6841 ) ;
  assign n6843 = n4287 ^ n2858 ^ 1'b0 ;
  assign n6844 = n4310 & n6843 ;
  assign n6845 = n6844 ^ n139 ^ 1'b0 ;
  assign n6846 = n5226 | n6845 ;
  assign n6847 = n4301 ^ n971 ^ 1'b0 ;
  assign n6848 = n945 & ~n2072 ;
  assign n6849 = n6848 ^ n487 ^ 1'b0 ;
  assign n6850 = n1979 | n6849 ;
  assign n6851 = n2615 & n4113 ;
  assign n6852 = n496 | n3678 ;
  assign n6853 = n6851 & ~n6852 ;
  assign n6854 = n6850 | n6853 ;
  assign n6855 = n6847 & ~n6854 ;
  assign n6856 = ( n3507 & n4730 ) | ( n3507 & ~n6855 ) | ( n4730 & ~n6855 ) ;
  assign n6857 = x100 & n2238 ;
  assign n6858 = n369 | n6857 ;
  assign n6859 = n4128 & ~n6858 ;
  assign n6860 = ~n353 & n5365 ;
  assign n6861 = ~n938 & n2861 ;
  assign n6862 = ( n2245 & ~n2897 ) | ( n2245 & n6861 ) | ( ~n2897 & n6861 ) ;
  assign n6863 = x17 & ~n1062 ;
  assign n6864 = n3722 & n6863 ;
  assign n6865 = n6864 ^ n5072 ^ 1'b0 ;
  assign n6866 = n6862 & n6865 ;
  assign n6867 = n750 & ~n2174 ;
  assign n6868 = n484 & n6867 ;
  assign n6869 = ( n3218 & n5267 ) | ( n3218 & n6458 ) | ( n5267 & n6458 ) ;
  assign n6870 = ~n6868 & n6869 ;
  assign n6871 = n6870 ^ n3862 ^ 1'b0 ;
  assign n6872 = n6871 ^ n601 ^ 1'b0 ;
  assign n6873 = ~n3339 & n6872 ;
  assign n6874 = n363 | n4011 ;
  assign n6875 = ~n3855 & n4084 ;
  assign n6876 = ( ~n4444 & n4658 ) | ( ~n4444 & n6875 ) | ( n4658 & n6875 ) ;
  assign n6877 = n535 & ~n891 ;
  assign n6878 = n4641 ^ x21 ^ 1'b0 ;
  assign n6879 = n1563 | n1903 ;
  assign n6880 = n2704 & ~n6879 ;
  assign n6881 = n6880 ^ n604 ^ 1'b0 ;
  assign n6882 = n304 & ~n4769 ;
  assign n6883 = n6882 ^ n2215 ^ 1'b0 ;
  assign n6884 = n1129 | n4901 ;
  assign n6885 = n1209 ^ n318 ^ 1'b0 ;
  assign n6886 = n404 | n6885 ;
  assign n6887 = n1554 | n4169 ;
  assign n6888 = ~n2779 & n6887 ;
  assign n6889 = n6886 & n6888 ;
  assign n6890 = n6884 & ~n6889 ;
  assign n6891 = n5575 | n6890 ;
  assign n6892 = n994 & n2667 ;
  assign n6893 = ~n1046 & n6892 ;
  assign n6894 = n1802 ^ n229 ^ 1'b0 ;
  assign n6895 = n6894 ^ n1770 ^ 1'b0 ;
  assign n6896 = n6893 | n6895 ;
  assign n6897 = n6896 ^ n2549 ^ 1'b0 ;
  assign n6898 = n3665 ^ n980 ^ 1'b0 ;
  assign n6899 = x2 | n6898 ;
  assign n6900 = n6899 ^ n3231 ^ 1'b0 ;
  assign n6901 = n1872 & n6900 ;
  assign n6902 = ~n4233 & n4506 ;
  assign n6903 = n2760 ^ n1468 ^ 1'b0 ;
  assign n6904 = ~n5282 & n6903 ;
  assign n6905 = n1427 ^ n173 ^ 1'b0 ;
  assign n6906 = n185 & ~n3240 ;
  assign n6907 = n1386 & n6906 ;
  assign n6908 = n4939 | n6907 ;
  assign n6911 = ~n1122 & n5937 ;
  assign n6909 = n3120 ^ n3062 ^ 1'b0 ;
  assign n6910 = ~n828 & n6909 ;
  assign n6912 = n6911 ^ n6910 ^ 1'b0 ;
  assign n6913 = n481 ^ x93 ^ 1'b0 ;
  assign n6914 = ~n1574 & n1708 ;
  assign n6915 = n6914 ^ n704 ^ 1'b0 ;
  assign n6916 = ~n2998 & n6915 ;
  assign n6917 = n6913 | n6916 ;
  assign n6918 = n4958 | n6706 ;
  assign n6919 = n6918 ^ n6605 ^ 1'b0 ;
  assign n6920 = n5072 ^ n704 ^ 1'b0 ;
  assign n6921 = n2681 & n6920 ;
  assign n6922 = n6921 ^ n1051 ^ 1'b0 ;
  assign n6923 = n2056 ^ n1924 ^ 1'b0 ;
  assign n6924 = n6923 ^ n496 ^ 1'b0 ;
  assign n6925 = ~n2044 & n6924 ;
  assign n6926 = n6925 ^ n1545 ^ 1'b0 ;
  assign n6927 = ~n2322 & n2422 ;
  assign n6928 = n6927 ^ n2038 ^ 1'b0 ;
  assign n6929 = n1817 & ~n2941 ;
  assign n6930 = n6544 & n6929 ;
  assign n6932 = n2151 & n3350 ;
  assign n6931 = n4459 ^ n2505 ^ 1'b0 ;
  assign n6933 = n6932 ^ n6931 ^ 1'b0 ;
  assign n6934 = n3157 ^ n2000 ^ n1664 ;
  assign n6935 = n6934 ^ n6032 ^ 1'b0 ;
  assign n6936 = n1079 | n1192 ;
  assign n6937 = n6935 & ~n6936 ;
  assign n6938 = n2604 & ~n5763 ;
  assign n6939 = ~n609 & n6938 ;
  assign n6940 = ( n499 & n3697 ) | ( n499 & ~n4267 ) | ( n3697 & ~n4267 ) ;
  assign n6941 = n336 & ~n1277 ;
  assign n6942 = n6941 ^ n310 ^ 1'b0 ;
  assign n6943 = n998 & n6117 ;
  assign n6947 = n4947 & n5298 ;
  assign n6944 = n2836 ^ n1497 ^ 1'b0 ;
  assign n6945 = x108 & ~n6944 ;
  assign n6946 = ~n6062 & n6945 ;
  assign n6948 = n6947 ^ n6946 ^ 1'b0 ;
  assign n6952 = n2630 & n6277 ;
  assign n6953 = n3411 & n6952 ;
  assign n6949 = n1713 & ~n4806 ;
  assign n6950 = ~n869 & n6949 ;
  assign n6951 = n4659 & ~n6950 ;
  assign n6954 = n6953 ^ n6951 ^ 1'b0 ;
  assign n6955 = ~n1130 & n4867 ;
  assign n6956 = n6955 ^ n5163 ^ 1'b0 ;
  assign n6957 = ( n886 & ~n4083 ) | ( n886 & n6956 ) | ( ~n4083 & n6956 ) ;
  assign n6958 = ~n3472 & n4434 ;
  assign n6959 = ~n3648 & n4268 ;
  assign n6960 = n6959 ^ n555 ^ 1'b0 ;
  assign n6961 = n6958 & ~n6960 ;
  assign n6962 = ~n3452 & n3819 ;
  assign n6963 = n1908 | n3090 ;
  assign n6964 = n6963 ^ n4527 ^ 1'b0 ;
  assign n6965 = n6473 ^ n639 ^ 1'b0 ;
  assign n6966 = n4042 ^ n1894 ^ 1'b0 ;
  assign n6967 = n6965 | n6966 ;
  assign n6968 = n6967 ^ n3740 ^ 1'b0 ;
  assign n6969 = n839 | n6968 ;
  assign n6970 = n4693 & n6871 ;
  assign n6971 = n6970 ^ n2539 ^ 1'b0 ;
  assign n6972 = ( n529 & ~n757 ) | ( n529 & n1982 ) | ( ~n757 & n1982 ) ;
  assign n6973 = n5664 ^ n3047 ^ n2765 ;
  assign n6974 = ~n292 & n6973 ;
  assign n6975 = ~n4102 & n6974 ;
  assign n6976 = n711 | n1419 ;
  assign n6977 = n1422 | n6976 ;
  assign n6978 = ~n245 & n1674 ;
  assign n6979 = ~n1165 & n6978 ;
  assign n6980 = n6977 & n6979 ;
  assign n6981 = n1768 ^ n1037 ^ 1'b0 ;
  assign n6982 = n3272 & n6981 ;
  assign n6983 = n2560 | n6982 ;
  assign n6984 = n4502 ^ n928 ^ 1'b0 ;
  assign n6985 = n359 & ~n5438 ;
  assign n6986 = n2433 ^ n568 ^ 1'b0 ;
  assign n6987 = n1414 & n6986 ;
  assign n6988 = n2683 | n4597 ;
  assign n6989 = n2967 ^ n2585 ^ 1'b0 ;
  assign n6990 = ~n1287 & n6989 ;
  assign n6992 = n1367 & n1983 ;
  assign n6991 = ~n245 & n711 ;
  assign n6993 = n6992 ^ n6991 ^ 1'b0 ;
  assign n6994 = n4238 | n6993 ;
  assign n6995 = n5801 ^ n1904 ^ 1'b0 ;
  assign n6996 = n4885 ^ n2929 ^ 1'b0 ;
  assign n6997 = ~n1908 & n6996 ;
  assign n6998 = n1201 & n6997 ;
  assign n6999 = n1023 & n6737 ;
  assign n7000 = ~n5825 & n6999 ;
  assign n7001 = n961 & n4840 ;
  assign n7002 = n2392 & n2913 ;
  assign n7003 = n4723 & ~n6383 ;
  assign n7004 = ~n5264 & n7003 ;
  assign n7005 = n2041 ^ x2 ^ 1'b0 ;
  assign n7006 = n7004 | n7005 ;
  assign n7007 = n2974 ^ n262 ^ 1'b0 ;
  assign n7008 = n7007 ^ n3393 ^ 1'b0 ;
  assign n7009 = ~n2480 & n7008 ;
  assign n7010 = n1491 & ~n2874 ;
  assign n7011 = ~n7009 & n7010 ;
  assign n7012 = n4105 ^ n1240 ^ 1'b0 ;
  assign n7013 = n1618 & ~n7012 ;
  assign n7014 = n2989 | n7013 ;
  assign n7015 = n7014 ^ n1206 ^ 1'b0 ;
  assign n7017 = n1744 & n1860 ;
  assign n7018 = n866 | n7017 ;
  assign n7019 = n1228 | n7018 ;
  assign n7016 = n639 | n5818 ;
  assign n7020 = n7019 ^ n7016 ^ n4288 ;
  assign n7021 = n574 & n757 ;
  assign n7022 = x14 & n1329 ;
  assign n7023 = n1049 & n7022 ;
  assign n7024 = n1365 & ~n1651 ;
  assign n7025 = n7024 ^ n267 ^ 1'b0 ;
  assign n7026 = n7023 | n7025 ;
  assign n7027 = n7021 & ~n7026 ;
  assign n7029 = ~n1683 & n3875 ;
  assign n7028 = ~n773 & n4494 ;
  assign n7030 = n7029 ^ n7028 ^ 1'b0 ;
  assign n7031 = ~n7027 & n7030 ;
  assign n7032 = n1376 | n6737 ;
  assign n7033 = n3155 ^ n1671 ^ 1'b0 ;
  assign n7034 = n7033 ^ n5913 ^ 1'b0 ;
  assign n7035 = n7032 & n7034 ;
  assign n7036 = x78 & n7035 ;
  assign n7037 = n7036 ^ n6355 ^ 1'b0 ;
  assign n7038 = n775 ^ n717 ^ 1'b0 ;
  assign n7039 = n7038 ^ n2394 ^ 1'b0 ;
  assign n7040 = n7037 & n7039 ;
  assign n7041 = n404 & n2236 ;
  assign n7042 = n7041 ^ n4484 ^ 1'b0 ;
  assign n7043 = n1870 & n7042 ;
  assign n7044 = n7043 ^ n5237 ^ n4212 ;
  assign n7045 = n4804 ^ n675 ^ 1'b0 ;
  assign n7046 = n5350 | n7045 ;
  assign n7047 = n1212 | n6802 ;
  assign n7048 = n735 | n1042 ;
  assign n7049 = n5801 | n7048 ;
  assign n7050 = n7049 ^ n4332 ^ 1'b0 ;
  assign n7051 = n1295 | n3142 ;
  assign n7052 = n7051 ^ n1997 ^ 1'b0 ;
  assign n7053 = n1551 ^ n1527 ^ 1'b0 ;
  assign n7054 = n7052 & ~n7053 ;
  assign n7055 = n3482 ^ n1668 ^ 1'b0 ;
  assign n7056 = n5874 | n7055 ;
  assign n7057 = n2934 & ~n7056 ;
  assign n7058 = n2521 ^ n1361 ^ 1'b0 ;
  assign n7059 = n795 & ~n7058 ;
  assign n7060 = n7059 ^ n4169 ^ 1'b0 ;
  assign n7061 = n6694 ^ n5393 ^ n4723 ;
  assign n7062 = ~n3017 & n7061 ;
  assign n7065 = n3050 & ~n4636 ;
  assign n7066 = ~n2638 & n7065 ;
  assign n7067 = n5243 & ~n7066 ;
  assign n7068 = n7067 ^ x36 ^ 1'b0 ;
  assign n7063 = n6454 ^ n3145 ^ 1'b0 ;
  assign n7064 = n6815 & ~n7063 ;
  assign n7069 = n7068 ^ n7064 ^ 1'b0 ;
  assign n7070 = n163 & n2575 ;
  assign n7071 = n484 & n7070 ;
  assign n7072 = n7071 ^ n2512 ^ 1'b0 ;
  assign n7073 = n1427 & n7072 ;
  assign n7074 = n863 & n1170 ;
  assign n7075 = n7074 ^ n2471 ^ 1'b0 ;
  assign n7076 = n3298 & n7075 ;
  assign n7077 = ~n6281 & n7076 ;
  assign n7078 = ~n1414 & n7077 ;
  assign n7079 = ( ~n1668 & n2545 ) | ( ~n1668 & n6645 ) | ( n2545 & n6645 ) ;
  assign n7080 = n3348 | n4865 ;
  assign n7081 = n2409 & ~n7080 ;
  assign n7082 = x116 & n7081 ;
  assign n7087 = n2705 & ~n4992 ;
  assign n7088 = n2565 | n7087 ;
  assign n7083 = ( ~n847 & n962 ) | ( ~n847 & n972 ) | ( n962 & n972 ) ;
  assign n7084 = n304 & n7083 ;
  assign n7085 = n1260 & n7084 ;
  assign n7086 = n5184 & ~n7085 ;
  assign n7089 = n7088 ^ n7086 ^ 1'b0 ;
  assign n7090 = n2822 ^ n1105 ^ 1'b0 ;
  assign n7091 = n3842 ^ n2145 ^ 1'b0 ;
  assign n7092 = n4674 & ~n7091 ;
  assign n7093 = n4366 | n7092 ;
  assign n7094 = n3510 & n7093 ;
  assign n7095 = ~n2408 & n2803 ;
  assign n7096 = n1993 | n5027 ;
  assign n7097 = ~n3564 & n4455 ;
  assign n7098 = n6048 & ~n7097 ;
  assign n7099 = n134 | n7098 ;
  assign n7100 = x1 & ~n7099 ;
  assign n7101 = ( n972 & n2051 ) | ( n972 & ~n2068 ) | ( n2051 & ~n2068 ) ;
  assign n7102 = n7101 ^ n526 ^ 1'b0 ;
  assign n7103 = x37 | n931 ;
  assign n7104 = n7103 ^ n5794 ^ 1'b0 ;
  assign n7105 = n4007 | n4361 ;
  assign n7106 = n4179 ^ n2716 ^ 1'b0 ;
  assign n7107 = n3859 & ~n7106 ;
  assign n7108 = n6371 ^ n4397 ^ 1'b0 ;
  assign n7109 = n3362 & n7108 ;
  assign n7110 = n974 & ~n6180 ;
  assign n7111 = n3381 | n4238 ;
  assign n7123 = n1287 & ~n2093 ;
  assign n7112 = n261 ^ n201 ^ 1'b0 ;
  assign n7116 = n2818 & n6540 ;
  assign n7117 = n662 | n1260 ;
  assign n7118 = n7116 | n7117 ;
  assign n7113 = n1540 & ~n4608 ;
  assign n7114 = n7113 ^ n1394 ^ 1'b0 ;
  assign n7115 = n7114 ^ n507 ^ 1'b0 ;
  assign n7119 = n7118 ^ n7115 ^ 1'b0 ;
  assign n7120 = n877 & ~n7119 ;
  assign n7121 = ( n4937 & n7112 ) | ( n4937 & ~n7120 ) | ( n7112 & ~n7120 ) ;
  assign n7122 = n2794 & ~n7121 ;
  assign n7124 = n7123 ^ n7122 ^ 1'b0 ;
  assign n7125 = n5061 ^ n3073 ^ 1'b0 ;
  assign n7126 = n346 | n707 ;
  assign n7127 = ~n2868 & n7126 ;
  assign n7128 = n7127 ^ n6104 ^ n5713 ;
  assign n7129 = n4902 ^ n1444 ^ 1'b0 ;
  assign n7137 = n427 | n1733 ;
  assign n7130 = n6610 ^ n2989 ^ 1'b0 ;
  assign n7131 = n7130 ^ n3354 ^ n1908 ;
  assign n7132 = ~n6296 & n7131 ;
  assign n7133 = n2582 & n5538 ;
  assign n7134 = n7133 ^ n1153 ^ 1'b0 ;
  assign n7135 = n5099 & ~n7134 ;
  assign n7136 = n7132 & ~n7135 ;
  assign n7138 = n7137 ^ n7136 ^ 1'b0 ;
  assign n7139 = n1001 ^ n246 ^ 1'b0 ;
  assign n7140 = n134 | n2140 ;
  assign n7141 = n7140 ^ n7031 ^ 1'b0 ;
  assign n7142 = n5739 ^ n4135 ^ 1'b0 ;
  assign n7143 = n1179 & ~n4310 ;
  assign n7145 = n4454 ^ n3040 ^ 1'b0 ;
  assign n7146 = x120 & ~n7145 ;
  assign n7147 = n1189 & n7146 ;
  assign n7148 = n1002 & n7147 ;
  assign n7149 = n2642 ^ n1694 ^ 1'b0 ;
  assign n7150 = n7148 | n7149 ;
  assign n7151 = n4783 ^ n724 ^ 1'b0 ;
  assign n7152 = n7150 | n7151 ;
  assign n7144 = n1829 & ~n6648 ;
  assign n7153 = n7152 ^ n7144 ^ 1'b0 ;
  assign n7154 = n564 & ~n4319 ;
  assign n7155 = ~n7153 & n7154 ;
  assign n7156 = n4682 & n6289 ;
  assign n7157 = n3862 & ~n6158 ;
  assign n7162 = n2198 ^ n2155 ^ n1412 ;
  assign n7158 = n3005 ^ n2813 ^ 1'b0 ;
  assign n7159 = x36 & ~n1645 ;
  assign n7160 = n7159 ^ n2561 ^ 1'b0 ;
  assign n7161 = n7158 & n7160 ;
  assign n7163 = n7162 ^ n7161 ^ 1'b0 ;
  assign n7164 = n3325 ^ n3028 ^ 1'b0 ;
  assign n7165 = n1321 & ~n7164 ;
  assign n7166 = n4076 & n7165 ;
  assign n7167 = n2776 & ~n5639 ;
  assign n7168 = x7 | n4914 ;
  assign n7169 = n1839 ^ n427 ^ 1'b0 ;
  assign n7170 = n7169 ^ n2759 ^ 1'b0 ;
  assign n7171 = n1628 & ~n3262 ;
  assign n7172 = n7171 ^ n6180 ^ 1'b0 ;
  assign n7174 = n643 ^ n360 ^ 1'b0 ;
  assign n7175 = n7174 ^ n1303 ^ 1'b0 ;
  assign n7173 = ~n6328 & n6627 ;
  assign n7176 = n7175 ^ n7173 ^ 1'b0 ;
  assign n7177 = x109 & n5741 ;
  assign n7178 = n7177 ^ x22 ^ 1'b0 ;
  assign n7179 = n729 & ~n7178 ;
  assign n7180 = ( x7 & ~n1329 ) | ( x7 & n3689 ) | ( ~n1329 & n3689 ) ;
  assign n7181 = n3948 ^ n2559 ^ 1'b0 ;
  assign n7182 = n339 | n7181 ;
  assign n7183 = n671 & n3906 ;
  assign n7184 = n7182 & n7183 ;
  assign n7185 = ( n1517 & n2442 ) | ( n1517 & n6840 ) | ( n2442 & n6840 ) ;
  assign n7186 = n1883 | n6367 ;
  assign n7187 = n989 | n6537 ;
  assign n7188 = n1331 | n7187 ;
  assign n7189 = n1766 | n2653 ;
  assign n7190 = n3149 | n7189 ;
  assign n7191 = n1800 ^ n854 ^ 1'b0 ;
  assign n7192 = n2571 & n7191 ;
  assign n7193 = n5466 & n7192 ;
  assign n7194 = n2861 | n4713 ;
  assign n7195 = n4052 & ~n6173 ;
  assign n7196 = n7195 ^ n4558 ^ 1'b0 ;
  assign n7197 = n6263 ^ n5330 ^ 1'b0 ;
  assign n7198 = n1602 & ~n7197 ;
  assign n7199 = n1867 | n7198 ;
  assign n7200 = ~n2928 & n6148 ;
  assign n7201 = ~n1806 & n7200 ;
  assign n7202 = ~n3435 & n7201 ;
  assign n7203 = n630 & n1628 ;
  assign n7204 = n5146 & n7203 ;
  assign n7205 = n858 & n2684 ;
  assign n7206 = n2083 & n7205 ;
  assign n7207 = n7206 ^ n6337 ^ 1'b0 ;
  assign n7208 = n3661 | n7207 ;
  assign n7209 = n1623 & ~n6714 ;
  assign n7210 = n469 & n7209 ;
  assign n7211 = n741 & n7210 ;
  assign n7212 = n7177 ^ n3611 ^ 1'b0 ;
  assign n7213 = n5048 ^ n2887 ^ 1'b0 ;
  assign n7214 = ~n1754 & n6447 ;
  assign n7215 = n7214 ^ n6563 ^ n4573 ;
  assign n7216 = n2091 | n3147 ;
  assign n7217 = n2433 ^ n1178 ^ 1'b0 ;
  assign n7218 = ~n983 & n1542 ;
  assign n7219 = n7218 ^ n4480 ^ 1'b0 ;
  assign n7220 = n3739 | n5998 ;
  assign n7221 = n2409 & ~n7220 ;
  assign n7222 = n2257 & ~n6387 ;
  assign n7223 = n131 | n1013 ;
  assign n7224 = n1616 & ~n7223 ;
  assign n7225 = ~n2043 & n7224 ;
  assign n7226 = ~n6962 & n7225 ;
  assign n7227 = ( n1329 & n5376 ) | ( n1329 & ~n6170 ) | ( n5376 & ~n6170 ) ;
  assign n7228 = n1980 & ~n4697 ;
  assign n7229 = ~n6445 & n7228 ;
  assign n7230 = n6661 ^ n6104 ^ n922 ;
  assign n7231 = n1792 & ~n5023 ;
  assign n7232 = n711 | n7231 ;
  assign n7233 = n790 | n7232 ;
  assign n7234 = n4230 ^ n1838 ^ 1'b0 ;
  assign n7235 = n2964 & ~n7234 ;
  assign n7236 = n1472 | n7235 ;
  assign n7237 = n1878 | n5647 ;
  assign n7238 = n5132 ^ n1383 ^ 1'b0 ;
  assign n7239 = n7237 & ~n7238 ;
  assign n7240 = n4002 | n6710 ;
  assign n7241 = n2945 | n7240 ;
  assign n7242 = n2436 & n5434 ;
  assign n7243 = n7242 ^ n5367 ^ 1'b0 ;
  assign n7244 = n7241 & ~n7243 ;
  assign n7245 = n806 & ~n7201 ;
  assign n7246 = n294 & n2055 ;
  assign n7247 = ~n3353 & n5010 ;
  assign n7248 = n5829 & n7247 ;
  assign n7249 = ~n4805 & n7248 ;
  assign n7250 = n155 | n4282 ;
  assign n7251 = n4180 ^ n3784 ^ 1'b0 ;
  assign n7252 = ~n2857 & n7251 ;
  assign n7253 = ~n5260 & n7252 ;
  assign n7254 = n1031 | n5488 ;
  assign n7255 = n4001 & ~n7254 ;
  assign n7256 = n7255 ^ n7019 ^ 1'b0 ;
  assign n7257 = n2490 & ~n7256 ;
  assign n7258 = x52 & ~n995 ;
  assign n7259 = ~n6688 & n7258 ;
  assign n7260 = n4137 ^ n3548 ^ 1'b0 ;
  assign n7261 = ~n7259 & n7260 ;
  assign n7262 = n7261 ^ n824 ^ 1'b0 ;
  assign n7263 = ~n660 & n2055 ;
  assign n7264 = ~n854 & n6226 ;
  assign n7265 = ~n308 & n7264 ;
  assign n7266 = n1228 & ~n5792 ;
  assign n7268 = n469 ^ n307 ^ 1'b0 ;
  assign n7267 = n645 & ~n5139 ;
  assign n7269 = n7268 ^ n7267 ^ 1'b0 ;
  assign n7270 = n944 ^ n702 ^ 1'b0 ;
  assign n7271 = n7270 ^ n1416 ^ 1'b0 ;
  assign n7272 = n5741 ^ n2966 ^ 1'b0 ;
  assign n7273 = n4615 | n7272 ;
  assign n7274 = ~n2911 & n3030 ;
  assign n7275 = n7274 ^ n1615 ^ 1'b0 ;
  assign n7276 = n4584 & ~n4966 ;
  assign n7277 = n1685 ^ n1139 ^ 1'b0 ;
  assign n7278 = n776 & ~n1321 ;
  assign n7279 = ~n1821 & n6725 ;
  assign n7280 = n7279 ^ n1996 ^ 1'b0 ;
  assign n7281 = ~n292 & n1806 ;
  assign n7282 = n7281 ^ n3091 ^ 1'b0 ;
  assign n7283 = n7282 ^ n1630 ^ 1'b0 ;
  assign n7284 = n5019 | n5363 ;
  assign n7285 = n4761 ^ n1147 ^ 1'b0 ;
  assign n7286 = ~n1130 & n5243 ;
  assign n7287 = n7286 ^ n2969 ^ 1'b0 ;
  assign n7291 = n1828 ^ n1762 ^ 1'b0 ;
  assign n7292 = n3398 | n7291 ;
  assign n7288 = n4351 ^ n2322 ^ n996 ;
  assign n7289 = ( n1080 & n2739 ) | ( n1080 & n7288 ) | ( n2739 & n7288 ) ;
  assign n7290 = n3330 | n7289 ;
  assign n7293 = n7292 ^ n7290 ^ 1'b0 ;
  assign n7294 = n141 & n311 ;
  assign n7295 = ~n766 & n7294 ;
  assign n7296 = n7295 ^ n1628 ^ 1'b0 ;
  assign n7297 = n4740 ^ n2072 ^ n1395 ;
  assign n7298 = n7297 ^ n1618 ^ 1'b0 ;
  assign n7299 = n7298 ^ n175 ^ 1'b0 ;
  assign n7300 = n5170 & n5243 ;
  assign n7301 = n2200 | n6186 ;
  assign n7302 = n3923 & ~n7301 ;
  assign n7303 = n4850 & ~n4939 ;
  assign n7304 = n6039 ^ n3074 ^ 1'b0 ;
  assign n7305 = n7304 ^ n6077 ^ n5730 ;
  assign n7306 = n2641 ^ n273 ^ 1'b0 ;
  assign n7307 = n413 | n5315 ;
  assign n7308 = n5791 ^ n5210 ^ 1'b0 ;
  assign n7309 = n2545 | n2843 ;
  assign n7310 = n7309 ^ n4763 ^ 1'b0 ;
  assign n7330 = ~n356 & n1284 ;
  assign n7331 = n356 & n7330 ;
  assign n7332 = n1741 | n7331 ;
  assign n7333 = n1741 & ~n7332 ;
  assign n7311 = ~n1020 & n5773 ;
  assign n7312 = x23 & ~n351 ;
  assign n7313 = ~x23 & n7312 ;
  assign n7314 = n7311 & ~n7313 ;
  assign n7315 = ~x120 & n7314 ;
  assign n7316 = n1432 & n2064 ;
  assign n7317 = ~n2064 & n7316 ;
  assign n7318 = n7317 ^ x127 ^ 1'b0 ;
  assign n7319 = x26 & ~n5773 ;
  assign n7320 = ~x26 & n7319 ;
  assign n7321 = n994 & ~n7320 ;
  assign n7322 = n7320 & n7321 ;
  assign n7323 = n1909 & ~n7322 ;
  assign n7324 = n7322 & n7323 ;
  assign n7325 = n7318 | n7324 ;
  assign n7326 = n7318 & ~n7325 ;
  assign n7327 = n1875 | n3253 ;
  assign n7328 = n7326 & ~n7327 ;
  assign n7329 = n7315 | n7328 ;
  assign n7334 = n7333 ^ n7329 ^ 1'b0 ;
  assign n7335 = n508 | n3299 ;
  assign n7336 = n7335 ^ n518 ^ 1'b0 ;
  assign n7337 = ~n6876 & n7336 ;
  assign n7338 = n5144 & n7092 ;
  assign n7339 = n4817 & n7338 ;
  assign n7340 = n571 | n1147 ;
  assign n7341 = n7340 ^ n3339 ^ 1'b0 ;
  assign n7342 = n2592 & ~n7341 ;
  assign n7343 = n7342 ^ n586 ^ 1'b0 ;
  assign n7344 = ~n4414 & n4919 ;
  assign n7345 = ~n5103 & n7344 ;
  assign n7346 = n3604 | n6213 ;
  assign n7347 = n3739 & ~n7346 ;
  assign n7348 = ~n6848 & n7347 ;
  assign n7349 = ~n806 & n1185 ;
  assign n7350 = ( ~n2330 & n3943 ) | ( ~n2330 & n7349 ) | ( n3943 & n7349 ) ;
  assign n7352 = n571 ^ x42 ^ 1'b0 ;
  assign n7353 = n5160 | n7352 ;
  assign n7354 = n590 & ~n7353 ;
  assign n7351 = ~n1387 & n4440 ;
  assign n7355 = n7354 ^ n7351 ^ 1'b0 ;
  assign n7356 = ~n6352 & n7355 ;
  assign n7357 = n3288 | n7356 ;
  assign n7358 = x61 | n7357 ;
  assign n7359 = n1290 | n2236 ;
  assign n7360 = ( n3754 & ~n5814 ) | ( n3754 & n7359 ) | ( ~n5814 & n7359 ) ;
  assign n7361 = n375 & n1201 ;
  assign n7362 = n2858 & ~n3722 ;
  assign n7363 = ~n1892 & n3919 ;
  assign n7364 = n7363 ^ n2130 ^ 1'b0 ;
  assign n7365 = ( n1841 & ~n6801 ) | ( n1841 & n7364 ) | ( ~n6801 & n7364 ) ;
  assign n7366 = n2117 | n7365 ;
  assign n7367 = n5020 | n7366 ;
  assign n7368 = n6303 ^ n1489 ^ 1'b0 ;
  assign n7369 = n2090 ^ x94 ^ 1'b0 ;
  assign n7370 = n2919 & ~n6542 ;
  assign n7371 = n181 & ~n5006 ;
  assign n7372 = ~n3516 & n5195 ;
  assign n7373 = n3392 & ~n5923 ;
  assign n7374 = ~n3865 & n7373 ;
  assign n7375 = n7374 ^ n4279 ^ 1'b0 ;
  assign n7376 = n4953 ^ n3257 ^ 1'b0 ;
  assign n7377 = n1177 & n1221 ;
  assign n7378 = n7377 ^ n1169 ^ 1'b0 ;
  assign n7380 = n5736 ^ x89 ^ 1'b0 ;
  assign n7379 = n1361 | n2855 ;
  assign n7381 = n7380 ^ n7379 ^ 1'b0 ;
  assign n7382 = ~n2705 & n6326 ;
  assign n7383 = n7382 ^ n6285 ^ 1'b0 ;
  assign n7384 = n1482 | n1998 ;
  assign n7385 = n1998 & ~n7384 ;
  assign n7386 = n7385 ^ n1663 ^ 1'b0 ;
  assign n7387 = n3644 & n7386 ;
  assign n7388 = ~n1669 & n7387 ;
  assign n7389 = n7388 ^ n1183 ^ 1'b0 ;
  assign n7390 = n1806 & n2707 ;
  assign n7391 = n1141 & n7390 ;
  assign n7392 = n4204 ^ n711 ^ 1'b0 ;
  assign n7393 = n3278 & n7392 ;
  assign n7394 = n7393 ^ x100 ^ 1'b0 ;
  assign n7395 = n3874 & n7394 ;
  assign n7396 = n912 & n7395 ;
  assign n7397 = n7391 & n7396 ;
  assign n7398 = n1900 | n7292 ;
  assign n7399 = n1875 & ~n7398 ;
  assign n7400 = n7399 ^ n3880 ^ 1'b0 ;
  assign n7401 = n4492 & ~n7400 ;
  assign n7402 = n2525 & ~n4096 ;
  assign n7403 = n7402 ^ n5374 ^ 1'b0 ;
  assign n7404 = n7401 & n7403 ;
  assign n7405 = n6369 ^ n2297 ^ n2232 ;
  assign n7406 = n5059 | n7405 ;
  assign n7407 = x67 | n7406 ;
  assign n7408 = ~n5836 & n7407 ;
  assign n7409 = n3992 ^ x123 ^ 1'b0 ;
  assign n7410 = n3479 | n7409 ;
  assign n7411 = n4319 & ~n7410 ;
  assign n7412 = n3714 ^ n786 ^ 1'b0 ;
  assign n7413 = n1890 & n7412 ;
  assign n7414 = n7413 ^ n805 ^ 1'b0 ;
  assign n7415 = n7414 ^ n4212 ^ 1'b0 ;
  assign n7416 = n7411 | n7415 ;
  assign n7417 = n1355 & n3469 ;
  assign n7418 = n7417 ^ n4800 ^ 1'b0 ;
  assign n7419 = n1604 ^ n545 ^ 1'b0 ;
  assign n7420 = n1452 & ~n7419 ;
  assign n7421 = n7420 ^ n6197 ^ 1'b0 ;
  assign n7422 = n1930 & ~n4271 ;
  assign n7423 = n1344 | n7422 ;
  assign n7424 = n5821 & n7422 ;
  assign n7425 = n159 & n5343 ;
  assign n7426 = n1226 & n7425 ;
  assign n7429 = n1098 | n3484 ;
  assign n7427 = n3301 ^ n2994 ^ 1'b0 ;
  assign n7428 = n879 & ~n7427 ;
  assign n7430 = n7429 ^ n7428 ^ 1'b0 ;
  assign n7431 = n7423 | n7430 ;
  assign n7432 = n7426 & ~n7431 ;
  assign n7433 = ( ~n614 & n1529 ) | ( ~n614 & n1613 ) | ( n1529 & n1613 ) ;
  assign n7434 = n2687 & n4784 ;
  assign n7435 = ~n7433 & n7434 ;
  assign n7436 = n7155 | n7435 ;
  assign n7437 = n542 & n895 ;
  assign n7438 = ( n4054 & n4638 ) | ( n4054 & ~n7437 ) | ( n4638 & ~n7437 ) ;
  assign n7439 = n7044 ^ n1013 ^ 1'b0 ;
  assign n7440 = n7438 & ~n7439 ;
  assign n7441 = n3244 ^ n2630 ^ 1'b0 ;
  assign n7442 = ~n1383 & n1699 ;
  assign n7443 = n7442 ^ n391 ^ 1'b0 ;
  assign n7444 = ~n304 & n7443 ;
  assign n7445 = n7444 ^ n7007 ^ 1'b0 ;
  assign n7446 = ~n666 & n6056 ;
  assign n7448 = n1651 ^ n638 ^ 1'b0 ;
  assign n7449 = n1366 & ~n7448 ;
  assign n7450 = n849 & ~n872 ;
  assign n7451 = ~n7449 & n7450 ;
  assign n7452 = n7451 ^ n4310 ^ 1'b0 ;
  assign n7453 = ~n5350 & n7452 ;
  assign n7447 = n841 & ~n5847 ;
  assign n7454 = n7453 ^ n7447 ^ 1'b0 ;
  assign n7455 = n4496 ^ n3581 ^ 1'b0 ;
  assign n7456 = ~n1532 & n7455 ;
  assign n7457 = n448 ^ x22 ^ 1'b0 ;
  assign n7458 = n2809 ^ n2436 ^ 1'b0 ;
  assign n7459 = n972 & ~n7458 ;
  assign n7460 = n1293 ^ n601 ^ 1'b0 ;
  assign n7461 = n1216 & ~n1264 ;
  assign n7462 = n1004 & n7461 ;
  assign n7463 = ~n7460 & n7462 ;
  assign n7464 = n5736 ^ n4916 ^ 1'b0 ;
  assign n7465 = n7463 | n7464 ;
  assign n7466 = n7465 ^ n1554 ^ 1'b0 ;
  assign n7467 = n1437 | n7466 ;
  assign n7468 = ( n825 & ~n3428 ) | ( n825 & n4057 ) | ( ~n3428 & n4057 ) ;
  assign n7469 = n5144 ^ n4319 ^ 1'b0 ;
  assign n7470 = n2123 ^ n886 ^ 1'b0 ;
  assign n7471 = n852 & ~n7470 ;
  assign n7472 = n7471 ^ n3318 ^ 1'b0 ;
  assign n7473 = n2248 & ~n7472 ;
  assign n7474 = n6387 & ~n7473 ;
  assign n7475 = n3052 ^ n2930 ^ 1'b0 ;
  assign n7476 = ( n1994 & n4288 ) | ( n1994 & ~n5117 ) | ( n4288 & ~n5117 ) ;
  assign n7477 = n4735 ^ n4249 ^ 1'b0 ;
  assign n7478 = n2857 | n7477 ;
  assign n7479 = ~n1517 & n3975 ;
  assign n7482 = n3465 ^ n1827 ^ 1'b0 ;
  assign n7483 = x46 | n2016 ;
  assign n7484 = n7482 | n7483 ;
  assign n7485 = n1795 ^ n192 ^ 1'b0 ;
  assign n7486 = n7484 & n7485 ;
  assign n7480 = x107 & n1983 ;
  assign n7481 = n7480 ^ n3729 ^ 1'b0 ;
  assign n7487 = n7486 ^ n7481 ^ 1'b0 ;
  assign n7488 = n296 | n6118 ;
  assign n7489 = n4796 ^ n2896 ^ 1'b0 ;
  assign n7490 = ~n482 & n7489 ;
  assign n7491 = n3170 & ~n5513 ;
  assign n7492 = n7491 ^ n485 ^ 1'b0 ;
  assign n7493 = ~n963 & n1954 ;
  assign n7494 = n7493 ^ n1419 ^ 1'b0 ;
  assign n7495 = x46 & ~n7494 ;
  assign n7496 = n6308 ^ n3503 ^ 1'b0 ;
  assign n7497 = n6975 | n7496 ;
  assign n7498 = n1908 ^ n882 ^ 1'b0 ;
  assign n7499 = ~x40 & n3123 ;
  assign n7500 = ~n165 & n7499 ;
  assign n7501 = n7500 ^ n544 ^ 1'b0 ;
  assign n7502 = ~n7498 & n7501 ;
  assign n7503 = ( x109 & n633 ) | ( x109 & n1592 ) | ( n633 & n1592 ) ;
  assign n7504 = ~n2989 & n7503 ;
  assign n7505 = ~n7502 & n7504 ;
  assign n7506 = n1998 ^ n1173 ^ 1'b0 ;
  assign n7507 = n1668 & n4162 ;
  assign n7508 = n7507 ^ n5170 ^ 1'b0 ;
  assign n7509 = n5602 & n7508 ;
  assign n7510 = ~n363 & n6781 ;
  assign n7511 = n7509 & n7510 ;
  assign n7512 = n7511 ^ n4037 ^ 1'b0 ;
  assign n7515 = n5818 ^ x93 ^ 1'b0 ;
  assign n7516 = n261 & n7515 ;
  assign n7517 = n7516 ^ n4336 ^ 1'b0 ;
  assign n7513 = ~n1467 & n1663 ;
  assign n7514 = n150 & ~n7513 ;
  assign n7518 = n7517 ^ n7514 ^ 1'b0 ;
  assign n7519 = n7518 ^ n1095 ^ 1'b0 ;
  assign n7520 = n937 & n3948 ;
  assign n7521 = n3360 & n7520 ;
  assign n7522 = n7521 ^ n4146 ^ 1'b0 ;
  assign n7523 = n4497 ^ n2140 ^ 1'b0 ;
  assign n7524 = n4499 | n4911 ;
  assign n7525 = ~n1452 & n2079 ;
  assign n7526 = ~n360 & n5477 ;
  assign n7527 = n7526 ^ n5989 ^ 1'b0 ;
  assign n7528 = x54 & n1534 ;
  assign n7529 = n7528 ^ n608 ^ 1'b0 ;
  assign n7530 = n245 & n7027 ;
  assign n7531 = n7530 ^ n950 ^ 1'b0 ;
  assign n7532 = n1580 & n3874 ;
  assign n7533 = n7532 ^ n1345 ^ 1'b0 ;
  assign n7534 = ~n250 & n1397 ;
  assign n7535 = ~n7533 & n7534 ;
  assign n7536 = n4641 ^ n2818 ^ 1'b0 ;
  assign n7537 = n3425 ^ n1851 ^ 1'b0 ;
  assign n7538 = n1547 & n1948 ;
  assign n7539 = n7538 ^ n299 ^ 1'b0 ;
  assign n7540 = n6011 ^ n2616 ^ 1'b0 ;
  assign n7541 = n7539 & n7540 ;
  assign n7542 = ~n894 & n7541 ;
  assign n7543 = n7537 & n7542 ;
  assign n7544 = n2998 & n5629 ;
  assign n7545 = n2426 & n5295 ;
  assign n7546 = n2646 ^ n549 ^ 1'b0 ;
  assign n7547 = n3089 | n7546 ;
  assign n7548 = n5086 ^ n400 ^ 1'b0 ;
  assign n7549 = n2091 & ~n7548 ;
  assign n7550 = n2245 ^ n788 ^ 1'b0 ;
  assign n7551 = n888 & ~n7405 ;
  assign n7552 = n7551 ^ n6454 ^ 1'b0 ;
  assign n7553 = n4415 | n6166 ;
  assign n7554 = n7552 & ~n7553 ;
  assign n7555 = n5483 | n7554 ;
  assign n7556 = n361 | n7555 ;
  assign n7557 = ~n2478 & n5558 ;
  assign n7558 = ~n1400 & n7557 ;
  assign n7561 = x7 & ~n1875 ;
  assign n7562 = n7561 ^ n1830 ^ 1'b0 ;
  assign n7559 = n3194 | n5789 ;
  assign n7560 = n7559 ^ n2560 ^ 1'b0 ;
  assign n7563 = n7562 ^ n7560 ^ n1323 ;
  assign n7564 = n4666 & n7563 ;
  assign n7565 = n7564 ^ n7268 ^ 1'b0 ;
  assign n7566 = ~n7465 & n7565 ;
  assign n7567 = n3128 | n7566 ;
  assign n7568 = n3819 ^ n3675 ^ 1'b0 ;
  assign n7569 = ~n4234 & n7568 ;
  assign n7570 = n1315 ^ n988 ^ 1'b0 ;
  assign n7571 = n7570 ^ n3074 ^ 1'b0 ;
  assign n7572 = n7569 & n7571 ;
  assign n7573 = n2321 | n7572 ;
  assign n7574 = n1245 | n7573 ;
  assign n7575 = n1989 ^ n1079 ^ 1'b0 ;
  assign n7576 = n1221 | n7575 ;
  assign n7577 = ~n1833 & n2664 ;
  assign n7578 = ~n2664 & n7577 ;
  assign n7579 = ~n5469 & n6978 ;
  assign n7580 = n5469 & n7579 ;
  assign n7581 = n7580 ^ n4579 ^ 1'b0 ;
  assign n7582 = ~n7578 & n7581 ;
  assign n7583 = ~n1107 & n7582 ;
  assign n7584 = ~n7582 & n7583 ;
  assign n7585 = n1853 & n1905 ;
  assign n7586 = n6417 ^ n1052 ^ 1'b0 ;
  assign n7587 = n7585 & ~n7586 ;
  assign n7588 = n7587 ^ n2983 ^ 1'b0 ;
  assign n7589 = ~n4078 & n7588 ;
  assign n7590 = n7589 ^ n3553 ^ 1'b0 ;
  assign n7591 = n6546 ^ n248 ^ 1'b0 ;
  assign n7592 = ~n7590 & n7591 ;
  assign n7593 = x72 | n886 ;
  assign n7594 = n1453 & n2354 ;
  assign n7595 = ~n4696 & n7594 ;
  assign n7596 = n4765 & ~n7595 ;
  assign n7597 = n4590 & ~n7596 ;
  assign n7598 = n4304 ^ n1756 ^ n889 ;
  assign n7599 = ~n2035 & n3600 ;
  assign n7600 = n254 & n7599 ;
  assign n7601 = ~n6053 & n6504 ;
  assign n7602 = ~n3661 & n5954 ;
  assign n7603 = n425 & ~n3773 ;
  assign n7604 = n6064 ^ n3721 ^ 1'b0 ;
  assign n7605 = n909 | n7604 ;
  assign n7606 = n5483 & n7605 ;
  assign n7607 = n7603 & n7606 ;
  assign n7608 = ( ~n402 & n2020 ) | ( ~n402 & n7607 ) | ( n2020 & n7607 ) ;
  assign n7609 = n137 & ~n2503 ;
  assign n7610 = ~n1692 & n7609 ;
  assign n7611 = n1862 | n7610 ;
  assign n7612 = n3996 | n7611 ;
  assign n7613 = n333 & ~n1167 ;
  assign n7614 = n1010 ^ n400 ^ x102 ;
  assign n7615 = n266 | n1724 ;
  assign n7616 = ( n2000 & n7614 ) | ( n2000 & ~n7615 ) | ( n7614 & ~n7615 ) ;
  assign n7617 = n353 & n825 ;
  assign n7618 = n7617 ^ n1436 ^ 1'b0 ;
  assign n7619 = ~n371 & n1099 ;
  assign n7620 = ~n6675 & n7619 ;
  assign n7621 = n7620 ^ n1141 ^ 1'b0 ;
  assign n7622 = n7618 & n7621 ;
  assign n7625 = n2523 ^ n2486 ^ 1'b0 ;
  assign n7623 = n1519 | n1541 ;
  assign n7624 = n7623 ^ n4258 ^ 1'b0 ;
  assign n7626 = n7625 ^ n7624 ^ 1'b0 ;
  assign n7627 = n1572 | n3253 ;
  assign n7628 = n471 | n7627 ;
  assign n7629 = n7628 ^ n6449 ^ 1'b0 ;
  assign n7630 = n1423 | n6850 ;
  assign n7631 = n7630 ^ n207 ^ 1'b0 ;
  assign n7632 = n2495 ^ n939 ^ 1'b0 ;
  assign n7633 = ~n7631 & n7632 ;
  assign n7634 = n1185 ^ x50 ^ 1'b0 ;
  assign n7635 = n1183 & ~n1762 ;
  assign n7636 = n790 & ~n7635 ;
  assign n7637 = n7634 & n7636 ;
  assign n7638 = ~n4886 & n6311 ;
  assign n7639 = n3027 & n7638 ;
  assign n7640 = n1372 | n6636 ;
  assign n7641 = n1153 & ~n2808 ;
  assign n7642 = n2505 & ~n3615 ;
  assign n7643 = n1973 & n7642 ;
  assign n7644 = n739 & n7292 ;
  assign n7645 = n3498 | n4098 ;
  assign n7646 = n7645 ^ n6788 ^ 1'b0 ;
  assign n7647 = n652 & n2493 ;
  assign n7648 = n4005 & n7647 ;
  assign n7649 = n1829 | n5927 ;
  assign n7650 = n7649 ^ n1470 ^ 1'b0 ;
  assign n7651 = n7650 ^ n1139 ^ 1'b0 ;
  assign n7652 = ~n3545 & n7651 ;
  assign n7653 = n2932 ^ n788 ^ 1'b0 ;
  assign n7655 = n2371 ^ n934 ^ 1'b0 ;
  assign n7654 = n3377 ^ n2980 ^ n2440 ;
  assign n7656 = n7655 ^ n7654 ^ 1'b0 ;
  assign n7657 = n1579 & n7656 ;
  assign n7658 = n867 & n7188 ;
  assign n7659 = n3422 | n5292 ;
  assign n7660 = n1069 | n5535 ;
  assign n7661 = n1566 & n5570 ;
  assign n7662 = n5558 & ~n7661 ;
  assign n7663 = n3773 ^ n2395 ^ 1'b0 ;
  assign n7664 = n1310 | n7663 ;
  assign n7665 = n6023 ^ n1628 ^ 1'b0 ;
  assign n7666 = ~n7664 & n7665 ;
  assign n7667 = n707 & n4883 ;
  assign n7668 = ~n2010 & n7667 ;
  assign n7669 = ~n3432 & n4571 ;
  assign n7670 = n7669 ^ n2446 ^ 1'b0 ;
  assign n7671 = n1018 ^ n230 ^ 1'b0 ;
  assign n7672 = n3719 & n7671 ;
  assign n7673 = n6017 & ~n7672 ;
  assign n7674 = n7378 & n7673 ;
  assign n7675 = n7674 ^ n3585 ^ 1'b0 ;
  assign n7676 = n1814 ^ n1253 ^ 1'b0 ;
  assign n7677 = n7369 ^ n1532 ^ 1'b0 ;
  assign n7678 = ~n7676 & n7677 ;
  assign n7679 = n4147 ^ n3797 ^ 1'b0 ;
  assign n7680 = n708 | n5818 ;
  assign n7681 = n7680 ^ n181 ^ 1'b0 ;
  assign n7682 = n3005 & n7681 ;
  assign n7683 = n7682 ^ n2669 ^ 1'b0 ;
  assign n7684 = n1193 ^ n1158 ^ 1'b0 ;
  assign n7685 = n7683 & ~n7684 ;
  assign n7686 = n7685 ^ n4946 ^ 1'b0 ;
  assign n7687 = ~n650 & n1076 ;
  assign n7688 = ~n701 & n7687 ;
  assign n7689 = ~n468 & n2701 ;
  assign n7690 = n7689 ^ n6809 ^ 1'b0 ;
  assign n7691 = ~n7688 & n7690 ;
  assign n7692 = n7691 ^ n2878 ^ 1'b0 ;
  assign n7693 = ~n1348 & n1716 ;
  assign n7694 = n7693 ^ x44 ^ 1'b0 ;
  assign n7695 = n7694 ^ n2101 ^ 1'b0 ;
  assign n7696 = n1862 | n6534 ;
  assign n7697 = n6114 & ~n7696 ;
  assign n7701 = ~n711 & n1808 ;
  assign n7698 = n3682 ^ n3327 ^ 1'b0 ;
  assign n7699 = x39 & ~n7698 ;
  assign n7700 = ~n2345 & n7699 ;
  assign n7702 = n7701 ^ n7700 ^ 1'b0 ;
  assign n7703 = n2349 & n7702 ;
  assign n7704 = n6155 & n7618 ;
  assign n7705 = n3193 & ~n6391 ;
  assign n7706 = n1394 & ~n6716 ;
  assign n7707 = n5057 ^ n2755 ^ 1'b0 ;
  assign n7708 = n466 | n5766 ;
  assign n7709 = n4652 | n7471 ;
  assign n7710 = n1391 ^ n692 ^ 1'b0 ;
  assign n7711 = n2016 | n7710 ;
  assign n7712 = n7711 ^ n1153 ^ 1'b0 ;
  assign n7714 = n3077 | n3844 ;
  assign n7715 = n2618 | n7714 ;
  assign n7713 = ~x4 & n6131 ;
  assign n7716 = n7715 ^ n7713 ^ 1'b0 ;
  assign n7717 = ~n2889 & n4571 ;
  assign n7718 = ~n4102 & n7717 ;
  assign n7719 = n7718 ^ n4393 ^ 1'b0 ;
  assign n7720 = n6071 ^ n5593 ^ 1'b0 ;
  assign n7721 = ~n7033 & n7720 ;
  assign n7722 = n5609 & n5845 ;
  assign n7723 = n2404 & n7722 ;
  assign n7724 = n6449 ^ n1161 ^ 1'b0 ;
  assign n7725 = n5223 ^ n4760 ^ n1056 ;
  assign n7726 = n835 ^ n430 ^ 1'b0 ;
  assign n7727 = n2800 & n7726 ;
  assign n7728 = n6945 ^ n5411 ^ 1'b0 ;
  assign n7729 = n4948 & n7728 ;
  assign n7730 = n7637 ^ n3487 ^ 1'b0 ;
  assign n7731 = n1351 & n7730 ;
  assign n7732 = n5801 ^ n2899 ^ 1'b0 ;
  assign n7733 = n6225 ^ n4848 ^ 1'b0 ;
  assign n7738 = n908 & n1245 ;
  assign n7739 = n7738 ^ n1035 ^ 1'b0 ;
  assign n7734 = n568 | n806 ;
  assign n7735 = n3367 | n7734 ;
  assign n7736 = n7735 ^ x71 ^ 1'b0 ;
  assign n7737 = n6077 | n7736 ;
  assign n7740 = n7739 ^ n7737 ^ 1'b0 ;
  assign n7741 = n6048 ^ n5745 ^ 1'b0 ;
  assign n7742 = n2458 & ~n2475 ;
  assign n7743 = n5235 & ~n7742 ;
  assign n7744 = n7743 ^ n5937 ^ 1'b0 ;
  assign n7746 = n1315 | n5253 ;
  assign n7747 = n7746 ^ n2208 ^ 1'b0 ;
  assign n7745 = n3898 ^ n3041 ^ n1063 ;
  assign n7748 = n7747 ^ n7745 ^ 1'b0 ;
  assign n7749 = n5096 | n7748 ;
  assign n7750 = ~x46 & n262 ;
  assign n7751 = n984 & n3182 ;
  assign n7752 = n7751 ^ n3425 ^ 1'b0 ;
  assign n7753 = ~n2469 & n7752 ;
  assign n7754 = n1736 & n6541 ;
  assign n7755 = n7754 ^ n1126 ^ 1'b0 ;
  assign n7756 = n5679 ^ n5146 ^ 1'b0 ;
  assign n7757 = n2091 ^ n221 ^ 1'b0 ;
  assign n7758 = ~n7756 & n7757 ;
  assign n7759 = n4893 ^ x107 ^ 1'b0 ;
  assign n7760 = n4482 | n7759 ;
  assign n7761 = n1072 | n7760 ;
  assign n7762 = n608 | n7761 ;
  assign n7763 = ~n2574 & n4689 ;
  assign n7764 = ~n757 & n1714 ;
  assign n7765 = ~n360 & n6283 ;
  assign n7766 = n7765 ^ n980 ^ 1'b0 ;
  assign n7767 = ~n2325 & n4641 ;
  assign n7768 = ~n862 & n6824 ;
  assign n7769 = n7768 ^ n6716 ^ 1'b0 ;
  assign n7770 = n1154 & ~n1290 ;
  assign n7771 = n2256 & ~n5930 ;
  assign n7772 = n7771 ^ n4430 ^ 1'b0 ;
  assign n7773 = n2616 & ~n7772 ;
  assign n7774 = ~n2808 & n3255 ;
  assign n7775 = n859 & n6448 ;
  assign n7776 = ~n7774 & n7775 ;
  assign n7777 = n7776 ^ n7017 ^ 1'b0 ;
  assign n7778 = ( n430 & n2039 ) | ( n430 & n4557 ) | ( n2039 & n4557 ) ;
  assign n7779 = n7778 ^ n3052 ^ 1'b0 ;
  assign n7780 = n4833 & n7779 ;
  assign n7781 = n1180 | n1393 ;
  assign n7782 = n4135 ^ n4126 ^ n806 ;
  assign n7783 = n7781 & ~n7782 ;
  assign n7784 = n7783 ^ n1900 ^ 1'b0 ;
  assign n7785 = n2333 & n2452 ;
  assign n7786 = x70 | n5941 ;
  assign n7787 = n5769 | n7786 ;
  assign n7788 = n7785 | n7787 ;
  assign n7789 = n2190 & ~n3302 ;
  assign n7790 = n571 ^ n307 ^ 1'b0 ;
  assign n7791 = ~n7789 & n7790 ;
  assign n7792 = n2818 ^ n307 ^ 1'b0 ;
  assign n7793 = ~x75 & n1966 ;
  assign n7794 = n4109 & ~n6827 ;
  assign n7795 = n5623 ^ n4149 ^ 1'b0 ;
  assign n7796 = n227 & n3420 ;
  assign n7797 = n2119 & ~n7739 ;
  assign n7798 = n7797 ^ n2662 ^ 1'b0 ;
  assign n7799 = n2366 & n7798 ;
  assign n7800 = n7156 ^ n4861 ^ 1'b0 ;
  assign n7801 = n7799 & n7800 ;
  assign n7802 = x89 | n6271 ;
  assign n7803 = n5397 & n7802 ;
  assign n7804 = n3169 ^ n1122 ^ x47 ;
  assign n7805 = x91 & ~n3629 ;
  assign n7806 = ~n7804 & n7805 ;
  assign n7807 = n7806 ^ n6129 ^ 1'b0 ;
  assign n7808 = n3723 & ~n7807 ;
  assign n7809 = n1854 & n7808 ;
  assign n7810 = n1035 ^ n258 ^ 1'b0 ;
  assign n7811 = n3210 & n6241 ;
  assign n7812 = n7811 ^ n5859 ^ 1'b0 ;
  assign n7813 = n2535 | n3862 ;
  assign n7814 = n1714 & ~n7813 ;
  assign n7815 = n7158 | n7814 ;
  assign n7816 = n3049 ^ n2636 ^ 1'b0 ;
  assign n7817 = n5070 ^ n3330 ^ 1'b0 ;
  assign n7818 = ~n3978 & n7817 ;
  assign n7819 = n7818 ^ n2409 ^ 1'b0 ;
  assign n7820 = x53 & ~n963 ;
  assign n7821 = n7820 ^ n4576 ^ 1'b0 ;
  assign n7822 = n642 | n7821 ;
  assign n7823 = n7822 ^ x13 ^ 1'b0 ;
  assign n7824 = n2999 ^ n216 ^ 1'b0 ;
  assign n7828 = ~n983 & n1610 ;
  assign n7829 = n7828 ^ n7739 ^ 1'b0 ;
  assign n7830 = ~n5543 & n7829 ;
  assign n7825 = n914 ^ n877 ^ 1'b0 ;
  assign n7826 = n2396 & n7825 ;
  assign n7827 = ~n3376 & n7826 ;
  assign n7831 = n7830 ^ n7827 ^ 1'b0 ;
  assign n7832 = n7824 | n7831 ;
  assign n7833 = n858 & ~n7832 ;
  assign n7834 = ~n7823 & n7833 ;
  assign n7835 = n4037 ^ n510 ^ 1'b0 ;
  assign n7836 = n5048 | n6118 ;
  assign n7837 = n2134 ^ n877 ^ 1'b0 ;
  assign n7838 = n7837 ^ n970 ^ 1'b0 ;
  assign n7839 = n7798 | n7838 ;
  assign n7840 = n6296 | n7839 ;
  assign n7841 = n7840 ^ n1746 ^ 1'b0 ;
  assign n7842 = n1080 | n7841 ;
  assign n7843 = n3072 | n7842 ;
  assign n7844 = n7593 & n7843 ;
  assign n7845 = n7844 ^ n211 ^ 1'b0 ;
  assign n7846 = n4744 ^ n4454 ^ 1'b0 ;
  assign n7847 = n2303 & ~n7846 ;
  assign n7848 = ( ~n1031 & n1558 ) | ( ~n1031 & n7847 ) | ( n1558 & n7847 ) ;
  assign n7849 = ( x57 & n1107 ) | ( x57 & n2885 ) | ( n1107 & n2885 ) ;
  assign n7850 = n2958 & n7849 ;
  assign n7851 = ~n7848 & n7850 ;
  assign n7852 = n7498 & ~n7627 ;
  assign n7853 = n7852 ^ n7140 ^ 1'b0 ;
  assign n7854 = ( n267 & n1463 ) | ( n267 & ~n5864 ) | ( n1463 & ~n5864 ) ;
  assign n7855 = n7854 ^ n195 ^ 1'b0 ;
  assign n7856 = ~n1147 & n4324 ;
  assign n7857 = n7856 ^ n506 ^ 1'b0 ;
  assign n7859 = n2626 & ~n6716 ;
  assign n7860 = ~n3299 & n6739 ;
  assign n7861 = ~n6739 & n7860 ;
  assign n7862 = n1502 & ~n7861 ;
  assign n7863 = n7859 & n7862 ;
  assign n7858 = n831 & ~n3817 ;
  assign n7864 = n7863 ^ n7858 ^ 1'b0 ;
  assign n7865 = ~n1456 & n5159 ;
  assign n7866 = n5469 ^ n1560 ^ 1'b0 ;
  assign n7867 = n7865 | n7866 ;
  assign n7868 = n3536 & ~n3607 ;
  assign n7869 = ~n3481 & n4744 ;
  assign n7870 = n7869 ^ n144 ^ 1'b0 ;
  assign n7871 = n3052 ^ n2093 ^ 1'b0 ;
  assign n7872 = n7870 & ~n7871 ;
  assign n7873 = n4796 & n7872 ;
  assign n7874 = n4305 ^ n2392 ^ 1'b0 ;
  assign n7875 = n865 ^ n491 ^ 1'b0 ;
  assign n7876 = n446 & n2857 ;
  assign n7877 = n3228 ^ n2889 ^ 1'b0 ;
  assign n7878 = n7876 & n7877 ;
  assign n7879 = n7875 & n7878 ;
  assign n7880 = n574 | n805 ;
  assign n7881 = n805 & ~n7880 ;
  assign n7882 = ~n1957 & n7881 ;
  assign n7883 = n2423 & n6193 ;
  assign n7884 = n7883 ^ n2926 ^ 1'b0 ;
  assign n7885 = n7882 & n7884 ;
  assign n7886 = n7885 ^ n5013 ^ 1'b0 ;
  assign n7887 = ~n1253 & n4461 ;
  assign n7888 = ~n3837 & n7887 ;
  assign n7889 = n4157 | n5463 ;
  assign n7891 = n2215 & n2702 ;
  assign n7890 = n6239 & ~n6542 ;
  assign n7892 = n7891 ^ n7890 ^ 1'b0 ;
  assign n7893 = n2702 & ~n6271 ;
  assign n7894 = n1552 & n7893 ;
  assign n7895 = n4467 & ~n7894 ;
  assign n7896 = n1260 & n7895 ;
  assign n7897 = n4610 ^ n2710 ^ 1'b0 ;
  assign n7898 = n183 | n7897 ;
  assign n7899 = n1217 & n5248 ;
  assign n7900 = ~n1107 & n7899 ;
  assign n7901 = n3542 ^ n2732 ^ 1'b0 ;
  assign n7902 = ~n5972 & n7901 ;
  assign n7903 = n6414 ^ n1510 ^ 1'b0 ;
  assign n7904 = n7903 ^ n1913 ^ 1'b0 ;
  assign n7905 = n3777 & ~n4117 ;
  assign n7906 = x42 & ~n2198 ;
  assign n7907 = ~x42 & n7906 ;
  assign n7908 = ~n1349 & n7907 ;
  assign n7909 = n4664 & n7908 ;
  assign n7910 = n514 & ~n7909 ;
  assign n7911 = n3371 ^ n538 ^ 1'b0 ;
  assign n7912 = ~n7910 & n7911 ;
  assign n7913 = n830 & n7912 ;
  assign n7914 = n978 | n5568 ;
  assign n7915 = n7914 ^ n1728 ^ 1'b0 ;
  assign n7916 = n3038 & ~n3722 ;
  assign n7917 = ~n812 & n7916 ;
  assign n7918 = n2896 ^ n1748 ^ 1'b0 ;
  assign n7919 = n2157 | n7918 ;
  assign n7920 = n6669 & ~n7919 ;
  assign n7921 = n7920 ^ n2143 ^ 1'b0 ;
  assign n7922 = n7917 | n7921 ;
  assign n7923 = n1120 & ~n3895 ;
  assign n7924 = n7923 ^ n3060 ^ 1'b0 ;
  assign n7925 = n5322 ^ n2694 ^ 1'b0 ;
  assign n7926 = n2739 & n5977 ;
  assign n7927 = n1020 & n7232 ;
  assign n7928 = n1188 & ~n3172 ;
  assign n7929 = n7928 ^ n2513 ^ 1'b0 ;
  assign n7930 = n2555 & n3038 ;
  assign n7931 = ~n5115 & n5492 ;
  assign n7932 = ~n1951 & n7931 ;
  assign n7933 = n1910 & ~n7129 ;
  assign n7934 = n553 & n6128 ;
  assign n7935 = n7595 ^ n2584 ^ 1'b0 ;
  assign n7936 = n6190 ^ n1558 ^ 1'b0 ;
  assign n7937 = n1714 ^ n1513 ^ 1'b0 ;
  assign n7938 = n6461 | n7937 ;
  assign n7939 = ~n5436 & n6511 ;
  assign n7940 = ~n1534 & n7939 ;
  assign n7941 = n5522 ^ n2208 ^ 1'b0 ;
  assign n7942 = ~n177 & n905 ;
  assign n7943 = n7942 ^ n1992 ^ 1'b0 ;
  assign n7944 = n5578 ^ n2470 ^ 1'b0 ;
  assign n7945 = ~n3193 & n4205 ;
  assign n7946 = n173 & n7945 ;
  assign n7947 = n7946 ^ n778 ^ 1'b0 ;
  assign n7948 = n7172 & n7947 ;
  assign n7949 = ( n562 & n1601 ) | ( n562 & n7739 ) | ( n1601 & n7739 ) ;
  assign n7950 = n2087 ^ n1983 ^ 1'b0 ;
  assign n7951 = n7949 & ~n7950 ;
  assign n7952 = n1972 | n6857 ;
  assign n7953 = n1655 ^ n315 ^ 1'b0 ;
  assign n7954 = n6932 & n7953 ;
  assign n7955 = ~n6210 & n7954 ;
  assign n7956 = ~n5649 & n7955 ;
  assign n7957 = n1191 & ~n1923 ;
  assign n7958 = n884 & n4448 ;
  assign n7959 = n7958 ^ n2981 ^ 1'b0 ;
  assign n7960 = n5042 ^ n662 ^ 1'b0 ;
  assign n7961 = n7959 & n7960 ;
  assign n7962 = n5832 ^ n2026 ^ n514 ;
  assign n7963 = n1290 | n7962 ;
  assign n7964 = n3859 & ~n4482 ;
  assign n7965 = ~n1397 & n7964 ;
  assign n7966 = ~n1360 & n7198 ;
  assign n7967 = n7966 ^ n3076 ^ 1'b0 ;
  assign n7968 = ( n537 & n6416 ) | ( n537 & ~n7356 ) | ( n6416 & ~n7356 ) ;
  assign n7969 = n2115 & n4985 ;
  assign n7970 = n7969 ^ n3298 ^ n717 ;
  assign n7971 = n2951 | n3003 ;
  assign n7972 = n189 & ~n958 ;
  assign n7973 = n3494 ^ n464 ^ 1'b0 ;
  assign n7974 = n7972 & n7973 ;
  assign n7975 = n1308 ^ n632 ^ 1'b0 ;
  assign n7976 = n161 | n7975 ;
  assign n7977 = n4692 | n6091 ;
  assign n7978 = ~n5907 & n7977 ;
  assign n7981 = n725 & n1919 ;
  assign n7982 = n4343 & ~n7981 ;
  assign n7983 = n483 & n2615 ;
  assign n7984 = n7982 & n7983 ;
  assign n7979 = n954 & ~n969 ;
  assign n7980 = ~n5793 & n7979 ;
  assign n7985 = n7984 ^ n7980 ^ 1'b0 ;
  assign n7986 = n1669 & ~n7985 ;
  assign n7987 = n533 & n2101 ;
  assign n7988 = n707 ^ x51 ^ 1'b0 ;
  assign n7989 = n336 & ~n7988 ;
  assign n7990 = n7989 ^ n7653 ^ 1'b0 ;
  assign n7991 = n7075 & ~n7990 ;
  assign n7993 = n7169 | n7839 ;
  assign n7994 = n3296 & ~n7993 ;
  assign n7992 = n702 & n2919 ;
  assign n7995 = n7994 ^ n7992 ^ 1'b0 ;
  assign n7996 = n2989 ^ n2099 ^ 1'b0 ;
  assign n7997 = n2694 & n3238 ;
  assign n7998 = ~n7760 & n7997 ;
  assign n7999 = n7998 ^ n2791 ^ 1'b0 ;
  assign n8004 = x72 & ~n3585 ;
  assign n8000 = ~n3419 & n3826 ;
  assign n8001 = n4234 ^ n618 ^ 1'b0 ;
  assign n8002 = n8000 & n8001 ;
  assign n8003 = ~n1550 & n8002 ;
  assign n8005 = n8004 ^ n8003 ^ 1'b0 ;
  assign n8006 = n4666 | n8005 ;
  assign n8007 = n8006 ^ x55 ^ 1'b0 ;
  assign n8008 = x15 & n809 ;
  assign n8009 = x17 & n3289 ;
  assign n8010 = n3292 | n8009 ;
  assign n8011 = n8010 ^ n3300 ^ 1'b0 ;
  assign n8012 = x37 | n1451 ;
  assign n8013 = n7997 ^ x126 ^ 1'b0 ;
  assign n8014 = n8012 & n8013 ;
  assign n8016 = n262 & n3169 ;
  assign n8017 = n8016 ^ n3930 ^ 1'b0 ;
  assign n8018 = n4505 | n8017 ;
  assign n8015 = n851 | n3089 ;
  assign n8019 = n8018 ^ n8015 ^ 1'b0 ;
  assign n8020 = n4823 | n7081 ;
  assign n8021 = n2015 ^ n512 ^ 1'b0 ;
  assign n8022 = n2948 & n8021 ;
  assign n8023 = n8022 ^ n1558 ^ 1'b0 ;
  assign n8024 = ~n1964 & n8023 ;
  assign n8025 = n6837 ^ n1574 ^ 1'b0 ;
  assign n8026 = ~n2440 & n8025 ;
  assign n8027 = n333 & ~n2000 ;
  assign n8028 = ~n359 & n8027 ;
  assign n8029 = n8028 ^ n5411 ^ 1'b0 ;
  assign n8030 = n3196 ^ n2517 ^ 1'b0 ;
  assign n8031 = n5308 & n8030 ;
  assign n8032 = n8031 ^ n1992 ^ 1'b0 ;
  assign n8033 = n1427 & ~n1716 ;
  assign n8034 = n5965 ^ n2146 ^ 1'b0 ;
  assign n8035 = n1695 | n5735 ;
  assign n8036 = ~n307 & n5974 ;
  assign n8037 = ~n8035 & n8036 ;
  assign n8038 = n1249 ^ n776 ^ 1'b0 ;
  assign n8039 = x29 & n8038 ;
  assign n8040 = n8039 ^ n3210 ^ 1'b0 ;
  assign n8041 = n6631 & n7162 ;
  assign n8042 = n5626 & n8041 ;
  assign n8043 = n8042 ^ n414 ^ 1'b0 ;
  assign n8044 = n530 ^ x62 ^ 1'b0 ;
  assign n8045 = n8044 ^ n3189 ^ 1'b0 ;
  assign n8046 = n1697 & ~n8045 ;
  assign n8047 = n1380 & ~n3791 ;
  assign n8048 = ~n1551 & n8047 ;
  assign n8049 = n6159 ^ n5611 ^ 1'b0 ;
  assign n8050 = n158 & ~n8049 ;
  assign n8051 = n7162 ^ n1179 ^ 1'b0 ;
  assign n8052 = n4901 & n8051 ;
  assign n8053 = n8052 ^ n2405 ^ 1'b0 ;
  assign n8054 = ~x22 & n8053 ;
  assign n8055 = ~x125 & n5820 ;
  assign n8056 = n7152 ^ n7017 ^ 1'b0 ;
  assign n8057 = n4110 | n5898 ;
  assign n8058 = n854 | n5863 ;
  assign n8059 = n2943 & ~n8058 ;
  assign n8060 = n8057 & n8059 ;
  assign n8061 = ~n5594 & n8060 ;
  assign n8062 = n6931 & ~n8061 ;
  assign n8063 = n8062 ^ n4858 ^ 1'b0 ;
  assign n8064 = n2893 & ~n8063 ;
  assign n8065 = n173 & n438 ;
  assign n8066 = n3770 | n7610 ;
  assign n8067 = n8066 ^ x17 ^ 1'b0 ;
  assign n8068 = ~n1640 & n8067 ;
  assign n8069 = n6399 & n8068 ;
  assign n8070 = n3858 & ~n4553 ;
  assign n8071 = n4553 & n8070 ;
  assign n8072 = ~n4775 & n8071 ;
  assign n8073 = ~x47 & n932 ;
  assign n8074 = x47 & n8073 ;
  assign n8075 = ~n3338 & n8074 ;
  assign n8076 = ~n8072 & n8075 ;
  assign n8077 = n8072 & n8076 ;
  assign n8078 = n1484 & n7423 ;
  assign n8079 = ~n2478 & n6704 ;
  assign n8080 = ( n1361 & n2371 ) | ( n1361 & n8079 ) | ( n2371 & n8079 ) ;
  assign n8081 = n7829 ^ n6206 ^ n2481 ;
  assign n8082 = n2585 | n3474 ;
  assign n8083 = ~n8081 & n8082 ;
  assign n8084 = n4897 & ~n8083 ;
  assign n8085 = n806 & n2337 ;
  assign n8086 = n8085 ^ n2592 ^ 1'b0 ;
  assign n8087 = n3977 | n8086 ;
  assign n8088 = n3281 | n4204 ;
  assign n8089 = n359 & n2312 ;
  assign n8090 = n8089 ^ n7776 ^ 1'b0 ;
  assign n8091 = n1596 | n4718 ;
  assign n8092 = n8091 ^ x90 ^ 1'b0 ;
  assign n8093 = n1310 & n5435 ;
  assign n8094 = n5626 & n6823 ;
  assign n8095 = ~n8093 & n8094 ;
  assign n8096 = n8095 ^ n3171 ^ 1'b0 ;
  assign n8097 = n4280 ^ x70 ^ 1'b0 ;
  assign n8098 = n8097 ^ n809 ^ 1'b0 ;
  assign n8100 = n5724 ^ n2125 ^ 1'b0 ;
  assign n8101 = n3868 & ~n8100 ;
  assign n8099 = n4395 & ~n5532 ;
  assign n8102 = n8101 ^ n8099 ^ 1'b0 ;
  assign n8105 = n7590 ^ n7451 ^ 1'b0 ;
  assign n8106 = n8086 & n8105 ;
  assign n8103 = ~n3228 & n3838 ;
  assign n8104 = x98 & ~n8103 ;
  assign n8107 = n8106 ^ n8104 ^ 1'b0 ;
  assign n8108 = n1574 & n1776 ;
  assign n8109 = n2290 & n8108 ;
  assign n8110 = ~n7424 & n8109 ;
  assign n8111 = n4749 ^ n3417 ^ 1'b0 ;
  assign n8112 = n5148 & ~n8111 ;
  assign n8113 = n3833 ^ n3553 ^ 1'b0 ;
  assign n8114 = ~n3262 & n7471 ;
  assign n8115 = n8113 & n8114 ;
  assign n8116 = n985 & n4612 ;
  assign n8117 = ~n3897 & n7473 ;
  assign n8118 = n4031 ^ n1087 ^ 1'b0 ;
  assign n8119 = n6998 ^ n2729 ^ 1'b0 ;
  assign n8120 = n1484 & ~n8119 ;
  assign n8121 = n1238 & n1534 ;
  assign n8122 = n2925 ^ n2232 ^ 1'b0 ;
  assign n8123 = n8122 ^ n701 ^ 1'b0 ;
  assign n8124 = n3488 & ~n8123 ;
  assign n8125 = n1580 ^ n392 ^ 1'b0 ;
  assign n8126 = n5118 ^ n4632 ^ n574 ;
  assign n8127 = n1122 & n3880 ;
  assign n8128 = n3210 & n8127 ;
  assign n8129 = n8128 ^ n2516 ^ 1'b0 ;
  assign n8130 = n6435 ^ n3465 ^ 1'b0 ;
  assign n8131 = n8129 & ~n8130 ;
  assign n8132 = n5731 ^ n2471 ^ 1'b0 ;
  assign n8133 = ~n3674 & n8132 ;
  assign n8134 = n2176 ^ n2079 ^ 1'b0 ;
  assign n8135 = n613 & ~n8134 ;
  assign n8136 = n5886 & n8135 ;
  assign n8137 = n750 & ~n1781 ;
  assign n8138 = n7615 & n8137 ;
  assign n8139 = n5255 ^ n634 ^ 1'b0 ;
  assign n8140 = ~n3661 & n8139 ;
  assign n8141 = ~n304 & n5207 ;
  assign n8142 = n3661 & n8141 ;
  assign n8143 = n2456 | n8142 ;
  assign n8144 = n8140 | n8143 ;
  assign n8145 = n6275 ^ n3396 ^ 1'b0 ;
  assign n8146 = n2579 | n8145 ;
  assign n8147 = n2405 ^ n1482 ^ 1'b0 ;
  assign n8148 = n1189 & ~n8147 ;
  assign n8151 = n169 | n2885 ;
  assign n8149 = ( n1126 & n1951 ) | ( n1126 & n1986 ) | ( n1951 & n1986 ) ;
  assign n8150 = n5232 & ~n8149 ;
  assign n8152 = n8151 ^ n8150 ^ 1'b0 ;
  assign n8153 = n4035 & n8152 ;
  assign n8154 = n8148 & n8153 ;
  assign n8155 = n3699 ^ n1589 ^ 1'b0 ;
  assign n8156 = ~n259 & n6205 ;
  assign n8157 = n8156 ^ n485 ^ 1'b0 ;
  assign n8158 = n3204 ^ n1010 ^ 1'b0 ;
  assign n8159 = n5944 & n8158 ;
  assign n8160 = ~n8157 & n8159 ;
  assign n8161 = ( n1202 & n1741 ) | ( n1202 & n2549 ) | ( n1741 & n2549 ) ;
  assign n8162 = ~n8137 & n8161 ;
  assign n8163 = n8162 ^ n5827 ^ 1'b0 ;
  assign n8164 = n2013 | n2278 ;
  assign n8165 = n4095 | n5637 ;
  assign n8166 = n8165 ^ n2006 ^ 1'b0 ;
  assign n8167 = n8166 ^ n3454 ^ 1'b0 ;
  assign n8168 = n1281 & ~n8167 ;
  assign n8169 = ~n4415 & n8168 ;
  assign n8170 = n6517 ^ n1662 ^ 1'b0 ;
  assign n8171 = ~n766 & n7083 ;
  assign n8172 = n8171 ^ n1534 ^ 1'b0 ;
  assign n8173 = ~n1459 & n8172 ;
  assign n8174 = n1950 ^ n1301 ^ 1'b0 ;
  assign n8175 = n5606 & n8174 ;
  assign n8176 = n1786 & ~n5809 ;
  assign n8177 = n3950 ^ n2746 ^ 1'b0 ;
  assign n8178 = n8177 ^ n2724 ^ 1'b0 ;
  assign n8179 = n4378 ^ n1226 ^ 1'b0 ;
  assign n8180 = ~n522 & n3080 ;
  assign n8181 = n307 & n8180 ;
  assign n8182 = n8179 & n8181 ;
  assign n8183 = n2003 ^ n324 ^ 1'b0 ;
  assign n8184 = ~n2411 & n6067 ;
  assign n8185 = ~n7847 & n8184 ;
  assign n8186 = n8052 ^ n233 ^ 1'b0 ;
  assign n8187 = ~n2032 & n6572 ;
  assign n8188 = ~n2972 & n8187 ;
  assign n8189 = n8188 ^ n504 ^ 1'b0 ;
  assign n8190 = x7 & ~n8189 ;
  assign n8191 = n2159 & n3066 ;
  assign n8192 = ~n3620 & n8191 ;
  assign n8193 = n2601 ^ x77 ^ 1'b0 ;
  assign n8194 = n6175 & ~n8193 ;
  assign n8195 = x22 & n2815 ;
  assign n8196 = n3179 & n8195 ;
  assign n8197 = n8196 ^ n195 ^ 1'b0 ;
  assign n8198 = n6818 & ~n8197 ;
  assign n8199 = n221 & n5751 ;
  assign n8200 = n7776 ^ n7414 ^ 1'b0 ;
  assign n8201 = n5341 & ~n5986 ;
  assign n8202 = n6923 | n8201 ;
  assign n8203 = n8202 ^ n2584 ^ 1'b0 ;
  assign n8204 = n4387 ^ n2756 ^ 1'b0 ;
  assign n8205 = n4197 ^ n2505 ^ 1'b0 ;
  assign n8206 = n1816 ^ n542 ^ 1'b0 ;
  assign n8207 = n8206 ^ n2445 ^ 1'b0 ;
  assign n8208 = ~n8205 & n8207 ;
  assign n8209 = n8208 ^ n1389 ^ 1'b0 ;
  assign n8214 = n761 & n3450 ;
  assign n8213 = n673 | n4825 ;
  assign n8215 = n8214 ^ n8213 ^ 1'b0 ;
  assign n8210 = n701 | n1468 ;
  assign n8211 = n1588 & ~n8210 ;
  assign n8212 = ~n5566 & n8211 ;
  assign n8216 = n8215 ^ n8212 ^ 1'b0 ;
  assign n8217 = n4319 ^ n582 ^ 1'b0 ;
  assign n8218 = n8217 ^ n7643 ^ 1'b0 ;
  assign n8219 = n728 & n1874 ;
  assign n8223 = n1724 & ~n2587 ;
  assign n8220 = n5500 ^ n1203 ^ 1'b0 ;
  assign n8221 = n1170 & n8220 ;
  assign n8222 = ~n4485 & n8221 ;
  assign n8224 = n8223 ^ n8222 ^ 1'b0 ;
  assign n8225 = n6268 ^ n4914 ^ 1'b0 ;
  assign n8226 = n909 | n7700 ;
  assign n8227 = n8226 ^ n2603 ^ 1'b0 ;
  assign n8228 = n845 ^ x94 ^ 1'b0 ;
  assign n8229 = n8227 & n8228 ;
  assign n8230 = ~n3789 & n8229 ;
  assign n8231 = n3629 ^ n2373 ^ 1'b0 ;
  assign n8232 = ~n2683 & n8231 ;
  assign n8233 = n1751 | n3828 ;
  assign n8234 = n3269 ^ n2800 ^ 1'b0 ;
  assign n8235 = x108 & n8234 ;
  assign n8236 = ~n8061 & n8235 ;
  assign n8237 = n8233 & n8236 ;
  assign n8241 = n3078 & n3610 ;
  assign n8242 = n2591 | n6003 ;
  assign n8243 = n3840 | n8242 ;
  assign n8244 = n2090 | n8243 ;
  assign n8245 = n8241 & n8244 ;
  assign n8238 = ~n2411 & n7690 ;
  assign n8239 = n1499 & n8238 ;
  assign n8240 = x22 | n8239 ;
  assign n8246 = n8245 ^ n8240 ^ 1'b0 ;
  assign n8247 = n1419 & n3629 ;
  assign n8248 = n1093 & n5166 ;
  assign n8249 = n8248 ^ n4942 ^ 1'b0 ;
  assign n8250 = ~n1149 & n8249 ;
  assign n8251 = ( n6328 & n6698 ) | ( n6328 & ~n6756 ) | ( n6698 & ~n6756 ) ;
  assign n8252 = n2808 & ~n7812 ;
  assign n8253 = n4248 & n8252 ;
  assign n8254 = n859 | n1498 ;
  assign n8255 = n4230 ^ n1631 ^ 1'b0 ;
  assign n8256 = n2673 & ~n8255 ;
  assign n8257 = n3696 & n8256 ;
  assign n8258 = ~n5096 & n8257 ;
  assign n8259 = n3086 | n8258 ;
  assign n8260 = n590 | n4287 ;
  assign n8261 = n8260 ^ n5070 ^ n1899 ;
  assign n8262 = x31 | n1920 ;
  assign n8263 = n2176 & ~n2724 ;
  assign n8264 = n8263 ^ n6026 ^ 1'b0 ;
  assign n8265 = n6240 & ~n8264 ;
  assign n8266 = n6337 ^ x77 ^ 1'b0 ;
  assign n8267 = n7552 ^ n380 ^ 1'b0 ;
  assign n8268 = n8266 | n8267 ;
  assign n8269 = n4761 ^ n4217 ^ 1'b0 ;
  assign n8270 = n6731 & ~n8269 ;
  assign n8271 = n6727 ^ n2363 ^ 1'b0 ;
  assign n8272 = n1972 & n8021 ;
  assign n8273 = n8271 & n8272 ;
  assign n8274 = n365 | n8273 ;
  assign n8277 = n1861 & ~n7718 ;
  assign n8278 = n8277 ^ n4901 ^ 1'b0 ;
  assign n8275 = n6547 ^ n5687 ^ 1'b0 ;
  assign n8276 = ~n3986 & n8275 ;
  assign n8279 = n8278 ^ n8276 ^ 1'b0 ;
  assign n8280 = n2702 & n8279 ;
  assign n8281 = ~n4636 & n7116 ;
  assign n8282 = n8281 ^ n2486 ^ 1'b0 ;
  assign n8283 = n962 | n1854 ;
  assign n8284 = n4226 & n8283 ;
  assign n8285 = ~n5403 & n8182 ;
  assign n8286 = x9 & n1541 ;
  assign n8287 = n7903 & ~n8286 ;
  assign n8288 = n8287 ^ n5248 ^ 1'b0 ;
  assign n8289 = n2276 & n3858 ;
  assign n8290 = n158 | n4417 ;
  assign n8291 = n8290 ^ n2159 ^ 1'b0 ;
  assign n8292 = n7664 & n8291 ;
  assign n8293 = n1959 | n4077 ;
  assign n8294 = n8293 ^ n1827 ^ 1'b0 ;
  assign n8295 = n6259 & n8294 ;
  assign n8296 = n242 & n3150 ;
  assign n8297 = n8296 ^ n2624 ^ 1'b0 ;
  assign n8298 = n1011 ^ x103 ^ 1'b0 ;
  assign n8299 = ~n8177 & n8298 ;
  assign n8300 = ~n8297 & n8299 ;
  assign n8301 = n2241 ^ n728 ^ 1'b0 ;
  assign n8302 = n1675 | n8301 ;
  assign n8303 = n1240 | n8302 ;
  assign n8304 = n8303 ^ n5953 ^ 1'b0 ;
  assign n8305 = ( n392 & ~n817 ) | ( n392 & n975 ) | ( ~n817 & n975 ) ;
  assign n8306 = ( n1165 & n4513 ) | ( n1165 & n8305 ) | ( n4513 & n8305 ) ;
  assign n8307 = ~n4280 & n7536 ;
  assign n8308 = n6531 & ~n6893 ;
  assign n8309 = n1487 & n8308 ;
  assign n8310 = n3312 & ~n4459 ;
  assign n8312 = n2371 | n2828 ;
  assign n8313 = n8312 ^ n5745 ^ 1'b0 ;
  assign n8311 = n786 | n4423 ;
  assign n8314 = n8313 ^ n8311 ^ 1'b0 ;
  assign n8315 = n1920 ^ n1206 ^ 1'b0 ;
  assign n8316 = n5213 ^ n4523 ^ 1'b0 ;
  assign n8317 = ~n4037 & n6473 ;
  assign n8318 = ~n8316 & n8317 ;
  assign n8319 = n3544 ^ n153 ^ 1'b0 ;
  assign n8320 = n1692 & n8319 ;
  assign n8324 = n3855 ^ n2351 ^ 1'b0 ;
  assign n8325 = n954 | n1062 ;
  assign n8326 = n8324 | n8325 ;
  assign n8322 = n2073 ^ n1875 ^ 1'b0 ;
  assign n8321 = n4647 & ~n5482 ;
  assign n8323 = n8322 ^ n8321 ^ 1'b0 ;
  assign n8327 = n8326 ^ n8323 ^ n7904 ;
  assign n8328 = n1419 | n5488 ;
  assign n8329 = n2321 | n8328 ;
  assign n8330 = n2392 & ~n8329 ;
  assign n8331 = n7971 ^ n3062 ^ 1'b0 ;
  assign n8332 = n3882 | n8331 ;
  assign n8333 = ~n2501 & n5096 ;
  assign n8334 = n159 & n167 ;
  assign n8335 = ~n442 & n8334 ;
  assign n8336 = n457 | n8335 ;
  assign n8337 = n8336 ^ n2919 ^ 1'b0 ;
  assign n8338 = n8337 ^ n3192 ^ 1'b0 ;
  assign n8339 = n3246 ^ n1255 ^ 1'b0 ;
  assign n8340 = ~n4347 & n8339 ;
  assign n8341 = n8340 ^ n320 ^ 1'b0 ;
  assign n8342 = n446 & n8341 ;
  assign n8343 = n826 & ~n8148 ;
  assign n8344 = ~n510 & n1328 ;
  assign n8345 = n8344 ^ n5405 ^ 1'b0 ;
  assign n8346 = n5035 | n5704 ;
  assign n8347 = n7884 | n8346 ;
  assign n8348 = n1890 ^ n810 ^ 1'b0 ;
  assign n8349 = n5613 | n8348 ;
  assign n8350 = n8349 ^ n150 ^ 1'b0 ;
  assign n8351 = n2868 ^ n2733 ^ 1'b0 ;
  assign n8352 = ~n512 & n8351 ;
  assign n8353 = n5883 & n8352 ;
  assign n8354 = n8353 ^ n623 ^ 1'b0 ;
  assign n8355 = n3981 | n7335 ;
  assign n8356 = n1013 | n8355 ;
  assign n8357 = n8356 ^ n373 ^ 1'b0 ;
  assign n8358 = n8354 & ~n8357 ;
  assign n8359 = ~n4980 & n5937 ;
  assign n8360 = n3149 & ~n8359 ;
  assign n8361 = ~n2981 & n5369 ;
  assign n8362 = ~n3544 & n8361 ;
  assign n8363 = n3687 & n5434 ;
  assign n8364 = ~n1033 & n6528 ;
  assign n8365 = n2407 & n8364 ;
  assign n8366 = n1631 | n8365 ;
  assign n8367 = n5350 & ~n8366 ;
  assign n8368 = ~n254 & n8367 ;
  assign n8369 = n1002 ^ n148 ^ 1'b0 ;
  assign n8370 = n3309 & ~n3353 ;
  assign n8371 = n7500 ^ n4305 ^ 1'b0 ;
  assign n8372 = n5632 ^ n5251 ^ 1'b0 ;
  assign n8373 = n6815 & ~n8372 ;
  assign n8374 = ( ~n3992 & n6034 ) | ( ~n3992 & n8373 ) | ( n6034 & n8373 ) ;
  assign n8375 = n2851 & n7719 ;
  assign n8376 = ~n7719 & n8375 ;
  assign n8377 = n1741 ^ n992 ^ 1'b0 ;
  assign n8378 = n272 & n2119 ;
  assign n8379 = ~n5317 & n8378 ;
  assign n8381 = n8129 ^ n510 ^ 1'b0 ;
  assign n8382 = n6011 | n8381 ;
  assign n8383 = n8210 | n8382 ;
  assign n8384 = n8383 ^ n5337 ^ 1'b0 ;
  assign n8380 = n874 | n2291 ;
  assign n8385 = n8384 ^ n8380 ^ 1'b0 ;
  assign n8386 = n1927 ^ n1371 ^ 1'b0 ;
  assign n8387 = n1861 & n8386 ;
  assign n8388 = ~n4656 & n5232 ;
  assign n8389 = n510 & n8388 ;
  assign n8390 = n4870 ^ n2940 ^ 1'b0 ;
  assign n8391 = n6515 ^ n3071 ^ 1'b0 ;
  assign n8392 = n1089 | n8391 ;
  assign n8393 = n2276 ^ n1485 ^ 1'b0 ;
  assign n8394 = ~n198 & n5889 ;
  assign n8395 = ~n3697 & n8394 ;
  assign n8396 = n604 & n786 ;
  assign n8397 = n528 & n8396 ;
  assign n8398 = n7355 ^ n2582 ^ 1'b0 ;
  assign n8399 = x33 & ~n296 ;
  assign n8400 = ~n1262 & n8399 ;
  assign n8401 = n8400 ^ n161 ^ 1'b0 ;
  assign n8402 = ~n3140 & n3637 ;
  assign n8403 = n8401 & n8402 ;
  assign n8404 = ~n8401 & n8403 ;
  assign n8405 = n902 | n1830 ;
  assign n8406 = n508 & ~n8405 ;
  assign n8407 = n2953 & n8406 ;
  assign n8408 = n5645 ^ n5208 ^ 1'b0 ;
  assign n8409 = n8407 | n8408 ;
  assign n8410 = n1867 | n5036 ;
  assign n8411 = n2962 & ~n8410 ;
  assign n8412 = ~n6450 & n7887 ;
  assign n8413 = n8412 ^ n805 ^ 1'b0 ;
  assign n8414 = n4941 ^ n2591 ^ 1'b0 ;
  assign n8415 = n3587 | n4323 ;
  assign n8416 = n8415 ^ n2183 ^ 1'b0 ;
  assign n8417 = n5304 ^ n1340 ^ 1'b0 ;
  assign n8418 = ~n8416 & n8417 ;
  assign n8419 = n2603 | n4040 ;
  assign n8420 = n3567 ^ n1838 ^ x6 ;
  assign n8421 = n8420 ^ n2089 ^ 1'b0 ;
  assign n8422 = ~n3288 & n6034 ;
  assign n8423 = ~n8421 & n8422 ;
  assign n8424 = n5306 ^ n4489 ^ 1'b0 ;
  assign n8425 = x85 & n8424 ;
  assign n8426 = n177 | n302 ;
  assign n8427 = n192 | n8426 ;
  assign n8428 = n8427 ^ n1230 ^ 1'b0 ;
  assign n8429 = n8425 & ~n8428 ;
  assign n8430 = n8407 ^ n2324 ^ 1'b0 ;
  assign n8431 = ~n926 & n5666 ;
  assign n8432 = n4711 & n6759 ;
  assign n8433 = ~n4525 & n8432 ;
  assign n8434 = n3407 | n5067 ;
  assign n8435 = n8434 ^ n6319 ^ 1'b0 ;
  assign n8436 = ~n5395 & n8435 ;
  assign n8437 = n3834 ^ x66 ^ 1'b0 ;
  assign n8438 = n1601 & ~n3541 ;
  assign n8439 = ~n1846 & n8438 ;
  assign n8440 = n6110 | n7735 ;
  assign n8441 = n4038 & n4824 ;
  assign n8443 = ~n2591 & n3420 ;
  assign n8444 = ~n1976 & n8443 ;
  assign n8442 = n159 | n4376 ;
  assign n8445 = n8444 ^ n8442 ^ 1'b0 ;
  assign n8446 = n8129 ^ n6170 ^ 1'b0 ;
  assign n8447 = n4791 ^ n3232 ^ 1'b0 ;
  assign n8448 = n4126 ^ n658 ^ 1'b0 ;
  assign n8449 = n2039 & ~n8448 ;
  assign n8450 = n590 & n5442 ;
  assign n8451 = n3717 & n8450 ;
  assign n8452 = ~n8449 & n8451 ;
  assign n8453 = n6759 ^ n6201 ^ 1'b0 ;
  assign n8454 = n3047 & n8453 ;
  assign n8455 = ~n4775 & n7083 ;
  assign n8456 = n8455 ^ n7688 ^ 1'b0 ;
  assign n8457 = n7468 ^ x20 ^ 1'b0 ;
  assign n8458 = n2143 & n8457 ;
  assign n8460 = n3034 | n4188 ;
  assign n8459 = n1843 ^ x106 ^ 1'b0 ;
  assign n8461 = n8460 ^ n8459 ^ 1'b0 ;
  assign n8462 = n1161 & n4641 ;
  assign n8463 = x94 & ~n307 ;
  assign n8464 = n942 & n8400 ;
  assign n8465 = n1837 ^ x51 ^ 1'b0 ;
  assign n8466 = n5139 ^ n1630 ^ 1'b0 ;
  assign n8467 = ~n8465 & n8466 ;
  assign n8468 = n4318 & n8467 ;
  assign n8469 = n2259 | n6953 ;
  assign n8470 = n1888 | n8469 ;
  assign n8471 = ~n466 & n8470 ;
  assign n8472 = n8468 & n8471 ;
  assign n8473 = n7681 ^ n1107 ^ 1'b0 ;
  assign n8474 = n8473 ^ n7438 ^ 1'b0 ;
  assign n8475 = n3142 | n3706 ;
  assign n8476 = n3695 | n8475 ;
  assign n8477 = x25 & n1776 ;
  assign n8478 = ~n1776 & n8477 ;
  assign n8479 = n2301 | n8478 ;
  assign n8480 = n2301 & ~n8479 ;
  assign n8481 = n7217 & ~n8480 ;
  assign n8482 = ~n696 & n6045 ;
  assign n8483 = n696 & n8482 ;
  assign n8484 = n876 | n8483 ;
  assign n8485 = ~n5588 & n8484 ;
  assign n8486 = ~n8481 & n8485 ;
  assign n8487 = ~n4005 & n6241 ;
  assign n8488 = ~n1819 & n6837 ;
  assign n8489 = n8487 & n8488 ;
  assign n8490 = ~n5213 & n8489 ;
  assign n8491 = n6456 & ~n6547 ;
  assign n8492 = ( n1037 & n4306 ) | ( n1037 & ~n6313 ) | ( n4306 & ~n6313 ) ;
  assign n8493 = ~n3636 & n4571 ;
  assign n8494 = n8493 ^ n2333 ^ 1'b0 ;
  assign n8500 = n1973 & ~n3305 ;
  assign n8501 = ~n2797 & n8500 ;
  assign n8502 = n1832 | n8501 ;
  assign n8495 = n1177 & n6234 ;
  assign n8496 = n5072 & n8495 ;
  assign n8497 = n8496 ^ n7433 ^ 1'b0 ;
  assign n8498 = n4858 | n8497 ;
  assign n8499 = n4310 | n8498 ;
  assign n8503 = n8502 ^ n8499 ^ 1'b0 ;
  assign n8504 = n5548 & ~n8503 ;
  assign n8505 = n444 | n844 ;
  assign n8506 = ~n430 & n8505 ;
  assign n8508 = ~n567 & n574 ;
  assign n8507 = n2672 & ~n4506 ;
  assign n8509 = n8508 ^ n8507 ^ 1'b0 ;
  assign n8510 = n3777 | n8509 ;
  assign n8511 = n989 | n4465 ;
  assign n8512 = n1683 & n5122 ;
  assign n8513 = n8512 ^ n5735 ^ 1'b0 ;
  assign n8514 = n4284 | n5442 ;
  assign n8515 = n7383 ^ n3544 ^ 1'b0 ;
  assign n8516 = n8515 ^ n3223 ^ 1'b0 ;
  assign n8517 = n8514 & ~n8516 ;
  assign n8518 = ~n1249 & n3274 ;
  assign n8519 = n6581 ^ n3309 ^ 1'b0 ;
  assign n8520 = n2806 ^ n2434 ^ n1141 ;
  assign n8521 = n7610 ^ n1035 ^ 1'b0 ;
  assign n8522 = n1919 | n8521 ;
  assign n8523 = n8144 ^ n3035 ^ 1'b0 ;
  assign n8524 = n5651 & ~n8523 ;
  assign n8525 = n7829 ^ n1691 ^ 1'b0 ;
  assign n8526 = n5716 & ~n8525 ;
  assign n8527 = n3196 | n8109 ;
  assign n8528 = n3615 & ~n8527 ;
  assign n8529 = ~n2583 & n8528 ;
  assign n8530 = n8529 ^ n7139 ^ n134 ;
  assign n8531 = n1240 ^ n624 ^ 1'b0 ;
  assign n8532 = n8531 ^ n4942 ^ 1'b0 ;
  assign n8533 = ~n6651 & n8532 ;
  assign n8534 = n1900 | n2994 ;
  assign n8535 = n2030 & ~n8534 ;
  assign n8536 = n5028 | n6932 ;
  assign n8539 = x81 & x93 ;
  assign n8540 = ~x93 & n8539 ;
  assign n8541 = ~x46 & x58 ;
  assign n8542 = n8540 & n8541 ;
  assign n8543 = ~n2911 & n8542 ;
  assign n8537 = n970 ^ n934 ^ 1'b0 ;
  assign n8538 = n557 & ~n8537 ;
  assign n8544 = n8543 ^ n8538 ^ 1'b0 ;
  assign n8560 = x93 & ~n385 ;
  assign n8561 = n385 & n8560 ;
  assign n8562 = n2746 | n8561 ;
  assign n8545 = x125 & n266 ;
  assign n8546 = ~n266 & n8545 ;
  assign n8547 = x93 & n240 ;
  assign n8548 = ~x93 & n8547 ;
  assign n8549 = n8548 ^ n753 ^ 1'b0 ;
  assign n8550 = n8546 & n8549 ;
  assign n8551 = ~n894 & n1205 ;
  assign n8552 = ~n1205 & n8551 ;
  assign n8553 = n1781 | n8552 ;
  assign n8554 = n8550 | n8553 ;
  assign n8555 = n8550 & ~n8554 ;
  assign n8556 = n1020 | n8555 ;
  assign n8557 = n8555 & ~n8556 ;
  assign n8558 = n3484 & ~n8557 ;
  assign n8559 = n8557 & n8558 ;
  assign n8563 = n8562 ^ n8559 ^ 1'b0 ;
  assign n8564 = ~n8544 & n8563 ;
  assign n8565 = n526 | n3732 ;
  assign n8566 = x125 & n8565 ;
  assign n8567 = n8566 ^ n320 ^ 1'b0 ;
  assign n8568 = n2591 | n6257 ;
  assign n8569 = n5119 | n8568 ;
  assign n8570 = n8569 ^ n4784 ^ 1'b0 ;
  assign n8571 = x114 & ~n945 ;
  assign n8572 = n3418 & n6128 ;
  assign n8573 = n8572 ^ n1861 ^ 1'b0 ;
  assign n8574 = n7604 & ~n8573 ;
  assign n8575 = n8574 ^ n595 ^ 1'b0 ;
  assign n8576 = n1378 & ~n8575 ;
  assign n8577 = n8571 & ~n8576 ;
  assign n8578 = n1299 & n2323 ;
  assign n8579 = ~n353 & n5982 ;
  assign n8580 = n2806 & n8579 ;
  assign n8581 = n4296 | n8359 ;
  assign n8582 = n5754 ^ n2009 ^ 1'b0 ;
  assign n8583 = n1480 ^ n344 ^ 1'b0 ;
  assign n8584 = n8211 & ~n8583 ;
  assign n8585 = ~n3240 & n5304 ;
  assign n8586 = n3193 ^ n2666 ^ 1'b0 ;
  assign n8587 = ~n3285 & n8586 ;
  assign n8588 = n6631 ^ n2949 ^ 1'b0 ;
  assign n8589 = n851 ^ n340 ^ 1'b0 ;
  assign n8590 = n1979 ^ n1455 ^ 1'b0 ;
  assign n8591 = n8589 | n8590 ;
  assign n8592 = n8588 & ~n8591 ;
  assign n8593 = ~n1808 & n3108 ;
  assign n8594 = ~n2378 & n8593 ;
  assign n8595 = ~n5826 & n7517 ;
  assign n8596 = ~n7002 & n7529 ;
  assign n8597 = n7272 ^ n1419 ^ 1'b0 ;
  assign n8598 = n1194 ^ n724 ^ 1'b0 ;
  assign n8599 = n6525 & n8598 ;
  assign n8602 = n1563 ^ n1395 ^ n718 ;
  assign n8600 = n4298 ^ n2062 ^ 1'b0 ;
  assign n8601 = n4040 & ~n8600 ;
  assign n8603 = n8602 ^ n8601 ^ 1'b0 ;
  assign n8604 = n8603 ^ n2385 ^ 1'b0 ;
  assign n8605 = n7918 ^ n2204 ^ 1'b0 ;
  assign n8608 = n4576 ^ n2851 ^ n1996 ;
  assign n8609 = n660 & n8608 ;
  assign n8606 = n3354 ^ n185 ^ 1'b0 ;
  assign n8607 = n6376 & ~n8606 ;
  assign n8610 = n8609 ^ n8607 ^ 1'b0 ;
  assign n8611 = n2931 & n2948 ;
  assign n8612 = n8611 ^ n4655 ^ 1'b0 ;
  assign n8613 = n2093 | n8612 ;
  assign n8614 = ( ~x39 & n2107 ) | ( ~x39 & n2681 ) | ( n2107 & n2681 ) ;
  assign n8615 = ~n4721 & n7360 ;
  assign n8616 = n1957 ^ n992 ^ 1'b0 ;
  assign n8617 = n307 & ~n8616 ;
  assign n8618 = n8617 ^ n1527 ^ 1'b0 ;
  assign n8619 = n1554 | n8618 ;
  assign n8620 = n2811 | n8619 ;
  assign n8621 = n8620 ^ n468 ^ 1'b0 ;
  assign n8622 = n8615 | n8621 ;
  assign n8623 = n8614 | n8622 ;
  assign n8624 = n6480 ^ n5413 ^ 1'b0 ;
  assign n8625 = n3622 ^ n1092 ^ 1'b0 ;
  assign n8626 = n2957 & n5990 ;
  assign n8627 = n8626 ^ n325 ^ 1'b0 ;
  assign n8628 = n8625 | n8627 ;
  assign n8631 = ~n173 & n6176 ;
  assign n8632 = ~n5666 & n8631 ;
  assign n8629 = n4316 ^ x119 ^ 1'b0 ;
  assign n8630 = ~n390 & n8629 ;
  assign n8633 = n8632 ^ n8630 ^ 1'b0 ;
  assign n8634 = n1737 & ~n3083 ;
  assign n8635 = n1571 & n8634 ;
  assign n8637 = n3415 & n7875 ;
  assign n8636 = n418 & n7101 ;
  assign n8638 = n8637 ^ n8636 ^ 1'b0 ;
  assign n8639 = n4814 ^ n2578 ^ 1'b0 ;
  assign n8640 = n902 ^ n571 ^ 1'b0 ;
  assign n8641 = ~n6102 & n8640 ;
  assign n8642 = ~n8639 & n8641 ;
  assign n8643 = n847 & n5142 ;
  assign n8644 = n2907 & n4227 ;
  assign n8645 = n307 & n4970 ;
  assign n8646 = n8645 ^ n6282 ^ 1'b0 ;
  assign n8647 = n5257 ^ n3926 ^ 1'b0 ;
  assign n8648 = n701 & n8647 ;
  assign n8649 = n2496 & n8648 ;
  assign n8650 = n2543 | n3107 ;
  assign n8651 = n7823 | n8650 ;
  assign n8652 = n6116 | n8651 ;
  assign n8653 = n8652 ^ n2948 ^ 1'b0 ;
  assign n8654 = n3371 ^ n1651 ^ 1'b0 ;
  assign n8655 = n2708 ^ n1498 ^ 1'b0 ;
  assign n8656 = n8655 ^ n7904 ^ 1'b0 ;
  assign n8657 = ~n8654 & n8656 ;
  assign n8658 = n942 & ~n2546 ;
  assign n8659 = n4954 ^ n2606 ^ 1'b0 ;
  assign n8660 = n2139 & n8659 ;
  assign n8661 = n3813 ^ n961 ^ 1'b0 ;
  assign n8662 = n8660 & ~n8661 ;
  assign n8663 = n8662 ^ n3509 ^ 1'b0 ;
  assign n8664 = n8658 & n8663 ;
  assign n8665 = n8101 ^ n3751 ^ 1'b0 ;
  assign n8666 = n356 | n3740 ;
  assign n8667 = n270 & ~n8344 ;
  assign n8668 = n400 & n1037 ;
  assign n8669 = n5020 & ~n8668 ;
  assign n8670 = ~n3157 & n8669 ;
  assign n8671 = n5067 & ~n8670 ;
  assign n8672 = x66 & ~n865 ;
  assign n8673 = ~n3256 & n8672 ;
  assign n8674 = n8673 ^ n5440 ^ 1'b0 ;
  assign n8675 = n3987 | n8674 ;
  assign n8676 = ~n980 & n1534 ;
  assign n8677 = n8676 ^ x81 ^ 1'b0 ;
  assign n8678 = n845 & ~n8677 ;
  assign n8679 = n788 & n8678 ;
  assign n8680 = n8679 ^ n5649 ^ 1'b0 ;
  assign n8681 = n5090 & ~n8680 ;
  assign n8682 = n6948 ^ n5806 ^ 1'b0 ;
  assign n8683 = n5594 & n8682 ;
  assign n8684 = n7855 ^ n4569 ^ 1'b0 ;
  assign n8685 = n359 & n5263 ;
  assign n8686 = ~n768 & n8685 ;
  assign n8687 = n8686 ^ n4310 ^ n2093 ;
  assign n8688 = n2322 ^ n708 ^ 1'b0 ;
  assign n8689 = n492 & n8688 ;
  assign n8690 = n1510 & n8689 ;
  assign n8691 = n1167 & n8690 ;
  assign n8692 = n8691 ^ n5687 ^ 1'b0 ;
  assign n8693 = n1495 & n8692 ;
  assign n8694 = n5168 & ~n8693 ;
  assign n8695 = n1914 ^ n394 ^ 1'b0 ;
  assign n8696 = n8695 ^ n4415 ^ 1'b0 ;
  assign n8697 = ~n1267 & n8696 ;
  assign n8698 = n4006 & ~n8697 ;
  assign n8699 = ~x77 & n5617 ;
  assign n8700 = n8699 ^ n8170 ^ 1'b0 ;
  assign n8701 = ~n6398 & n8700 ;
  assign n8703 = n237 & ~n2983 ;
  assign n8704 = ~n2468 & n8703 ;
  assign n8705 = n8704 ^ n6699 ^ 1'b0 ;
  assign n8706 = n4995 & n8705 ;
  assign n8707 = n4106 & n8706 ;
  assign n8702 = n1316 & ~n3607 ;
  assign n8708 = n8707 ^ n8702 ^ 1'b0 ;
  assign n8709 = ( n1109 & n2290 ) | ( n1109 & n5354 ) | ( n2290 & n5354 ) ;
  assign n8710 = n5107 & ~n8709 ;
  assign n8711 = n985 & n3417 ;
  assign n8712 = n1015 | n6022 ;
  assign n8713 = n8533 | n8712 ;
  assign n8714 = n146 & n5358 ;
  assign n8715 = n5168 & ~n8714 ;
  assign n8716 = ~n6766 & n8715 ;
  assign n8719 = n6251 ^ n3587 ^ 1'b0 ;
  assign n8720 = ~n6418 & n8719 ;
  assign n8717 = n2512 & ~n7025 ;
  assign n8718 = n1472 | n8717 ;
  assign n8721 = n8720 ^ n8718 ^ 1'b0 ;
  assign n8722 = n5582 | n5754 ;
  assign n8723 = n704 & ~n8722 ;
  assign n8724 = n1708 ^ n1700 ^ n880 ;
  assign n8725 = n3458 & ~n7274 ;
  assign n8726 = n4901 ^ n485 ^ 1'b0 ;
  assign n8727 = n3774 ^ n3090 ^ 1'b0 ;
  assign n8728 = n5802 & n8727 ;
  assign n8729 = n1789 | n1990 ;
  assign n8730 = n8729 ^ n3682 ^ 1'b0 ;
  assign n8732 = n1839 & ~n5488 ;
  assign n8733 = n4003 & n8732 ;
  assign n8731 = ~n4047 & n5289 ;
  assign n8734 = n8733 ^ n8731 ^ 1'b0 ;
  assign n8735 = n8730 | n8734 ;
  assign n8736 = n7616 ^ n5161 ^ 1'b0 ;
  assign n8737 = n8735 | n8736 ;
  assign n8738 = n1496 | n6266 ;
  assign n8739 = n2422 & n8738 ;
  assign n8740 = n967 & n8739 ;
  assign n8741 = n2693 | n3029 ;
  assign n8742 = n8741 ^ n5418 ^ 1'b0 ;
  assign n8743 = ~n2824 & n8742 ;
  assign n8744 = n6482 ^ n6465 ^ 1'b0 ;
  assign n8745 = n8239 ^ n2354 ^ 1'b0 ;
  assign n8746 = n1241 & ~n8745 ;
  assign n8747 = n7066 ^ n2469 ^ 1'b0 ;
  assign n8748 = n2079 & n8747 ;
  assign n8749 = n5144 & n8748 ;
  assign n8750 = n8749 ^ n2315 ^ 1'b0 ;
  assign n8751 = n8180 & ~n8750 ;
  assign n8752 = n246 & ~n3062 ;
  assign n8753 = n1653 & n8752 ;
  assign n8754 = n8753 ^ n5064 ^ n3498 ;
  assign n8757 = n583 & ~n6367 ;
  assign n8758 = n8757 ^ n5976 ^ n5237 ;
  assign n8755 = n3377 ^ n262 ^ 1'b0 ;
  assign n8756 = n1142 & ~n8755 ;
  assign n8759 = n8758 ^ n8756 ^ 1'b0 ;
  assign n8765 = ~n3584 & n7158 ;
  assign n8766 = n8765 ^ n3056 ^ 1'b0 ;
  assign n8767 = x67 & ~n8766 ;
  assign n8768 = x3 & ~n3293 ;
  assign n8769 = ~n8767 & n8768 ;
  assign n8760 = n7981 ^ n960 ^ 1'b0 ;
  assign n8761 = ~n3204 & n8760 ;
  assign n8762 = n8761 ^ n7038 ^ 1'b0 ;
  assign n8763 = n2702 & n8762 ;
  assign n8764 = n4062 & ~n8763 ;
  assign n8770 = n8769 ^ n8764 ^ 1'b0 ;
  assign n8771 = n3667 | n5689 ;
  assign n8772 = n4212 & ~n8771 ;
  assign n8773 = n238 & n1870 ;
  assign n8774 = n6499 | n8773 ;
  assign n8775 = n3875 | n8774 ;
  assign n8776 = ~n7564 & n8775 ;
  assign n8777 = n7202 | n8577 ;
  assign n8778 = n704 | n3296 ;
  assign n8779 = n8778 ^ n2802 ^ 1'b0 ;
  assign n8780 = n3120 | n8779 ;
  assign n8781 = ( n5229 & n5689 ) | ( n5229 & ~n8780 ) | ( n5689 & ~n8780 ) ;
  assign n8782 = n4002 ^ n436 ^ 1'b0 ;
  assign n8783 = n4251 ^ n3904 ^ n2857 ;
  assign n8784 = n4306 | n8783 ;
  assign n8785 = n8782 | n8784 ;
  assign n8786 = ~n262 & n4162 ;
  assign n8787 = ~n3090 & n8786 ;
  assign n8788 = n2614 & ~n8787 ;
  assign n8789 = n8788 ^ n1551 ^ 1'b0 ;
  assign n8790 = n750 & ~n8789 ;
  assign n8791 = n5500 & n8790 ;
  assign n8792 = n5998 | n8791 ;
  assign n8793 = n8785 | n8792 ;
  assign n8794 = n8599 ^ x122 ^ 1'b0 ;
  assign n8795 = n7116 | n8512 ;
  assign n8796 = ~n3474 & n5731 ;
  assign n8797 = n558 & ~n3563 ;
  assign n8798 = n8797 ^ n1550 ^ 1'b0 ;
  assign n8799 = ~n3104 & n8798 ;
  assign n8800 = n1937 | n8799 ;
  assign n8801 = n722 ^ n634 ^ 1'b0 ;
  assign n8802 = ~n457 & n8801 ;
  assign n8803 = ~n8800 & n8802 ;
  assign n8804 = n8266 ^ n221 ^ 1'b0 ;
  assign n8805 = n3369 ^ n1534 ^ 1'b0 ;
  assign n8806 = n914 | n8805 ;
  assign n8807 = n6967 | n8806 ;
  assign n8808 = n558 | n1979 ;
  assign n8809 = ~n4408 & n8808 ;
  assign n8810 = n8809 ^ n1201 ^ 1'b0 ;
  assign n8811 = n8810 ^ n7259 ^ n243 ;
  assign n8813 = ~n1469 & n5317 ;
  assign n8812 = n5556 & n5940 ;
  assign n8814 = n8813 ^ n8812 ^ 1'b0 ;
  assign n8815 = n5320 ^ n3163 ^ 1'b0 ;
  assign n8816 = n5451 & ~n8815 ;
  assign n8817 = ~n2389 & n5146 ;
  assign n8818 = n8817 ^ n5130 ^ 1'b0 ;
  assign n8819 = ~n1290 & n4579 ;
  assign n8820 = n6077 & n8819 ;
  assign n8824 = n3189 ^ n650 ^ 1'b0 ;
  assign n8825 = n2713 & n8824 ;
  assign n8826 = n879 | n8825 ;
  assign n8827 = n8826 ^ n3629 ^ 1'b0 ;
  assign n8828 = n1374 | n8827 ;
  assign n8821 = n5224 ^ n1212 ^ n618 ;
  assign n8822 = ~n2173 & n8821 ;
  assign n8823 = n4325 & n8822 ;
  assign n8829 = n8828 ^ n8823 ^ n1958 ;
  assign n8830 = n482 | n4459 ;
  assign n8831 = n1397 | n8830 ;
  assign n8832 = n2099 & ~n8831 ;
  assign n8833 = n1141 & ~n4002 ;
  assign n8834 = ~n1667 & n4802 ;
  assign n8835 = n8834 ^ n647 ^ 1'b0 ;
  assign n8836 = n4621 | n8835 ;
  assign n8837 = n8836 ^ n7009 ^ 1'b0 ;
  assign n8838 = n2958 & ~n4501 ;
  assign n8839 = n504 & n8838 ;
  assign n8840 = ~x105 & n8839 ;
  assign n8841 = n2660 & n3103 ;
  assign n8842 = n851 & n1997 ;
  assign n8843 = ~n8841 & n8842 ;
  assign n8844 = n2574 ^ n938 ^ 1'b0 ;
  assign n8845 = n8844 ^ n4079 ^ 1'b0 ;
  assign n8846 = n8315 | n8845 ;
  assign n8847 = ~n2091 & n4655 ;
  assign n8848 = n8847 ^ n1067 ^ 1'b0 ;
  assign n8849 = n8848 ^ n5974 ^ 1'b0 ;
  assign n8850 = n3272 ^ n1010 ^ n221 ;
  assign n8851 = n1172 | n8850 ;
  assign n8852 = n571 | n7735 ;
  assign n8853 = n4244 ^ n2579 ^ 1'b0 ;
  assign n8854 = n6348 | n8853 ;
  assign n8855 = n141 | n3917 ;
  assign n8856 = n707 & ~n8855 ;
  assign n8857 = n8856 ^ n4204 ^ 1'b0 ;
  assign n8859 = ~n663 & n3981 ;
  assign n8860 = n2879 & n8859 ;
  assign n8861 = n8018 & n8860 ;
  assign n8858 = n4847 & n7360 ;
  assign n8862 = n8861 ^ n8858 ^ 1'b0 ;
  assign n8863 = n4324 | n8157 ;
  assign n8864 = n167 & ~n1253 ;
  assign n8865 = n8864 ^ n1979 ^ 1'b0 ;
  assign n8866 = n5385 & ~n8865 ;
  assign n8867 = n8866 ^ n3584 ^ 1'b0 ;
  assign n8868 = n7891 ^ n1041 ^ 1'b0 ;
  assign n8869 = n972 & ~n8868 ;
  assign n8870 = n595 & ~n7437 ;
  assign n8871 = n8870 ^ n4472 ^ 1'b0 ;
  assign n8872 = n851 | n4962 ;
  assign n8873 = n8872 ^ n4413 ^ 1'b0 ;
  assign n8874 = n5140 ^ n1415 ^ 1'b0 ;
  assign n8875 = n2177 & ~n8874 ;
  assign n8876 = n1020 & ~n4608 ;
  assign n8877 = n8876 ^ n3229 ^ 1'b0 ;
  assign n8878 = n2073 ^ n1564 ^ 1'b0 ;
  assign n8879 = n8877 & ~n8878 ;
  assign n8880 = n8142 ^ n6078 ^ 1'b0 ;
  assign n8881 = n1663 | n2533 ;
  assign n8882 = n8881 ^ n2996 ^ 1'b0 ;
  assign n8883 = n213 & ~n8882 ;
  assign n8884 = n129 | n889 ;
  assign n8885 = n4071 & ~n8884 ;
  assign n8886 = n1599 & ~n8885 ;
  assign n8887 = n6994 & n8886 ;
  assign n8888 = n1432 ^ n167 ^ 1'b0 ;
  assign n8889 = n8888 ^ n7887 ^ 1'b0 ;
  assign n8890 = n4610 | n7023 ;
  assign n8891 = n8890 ^ n1158 ^ 1'b0 ;
  assign n8892 = ( n221 & ~n1292 ) | ( n221 & n1989 ) | ( ~n1292 & n1989 ) ;
  assign n8893 = n6901 & n8892 ;
  assign n8894 = n3812 & n8893 ;
  assign n8898 = n1366 & ~n6536 ;
  assign n8899 = n8898 ^ n4817 ^ 1'b0 ;
  assign n8895 = ~n1563 & n7146 ;
  assign n8896 = n656 & n8895 ;
  assign n8897 = n7694 | n8896 ;
  assign n8900 = n8899 ^ n8897 ^ 1'b0 ;
  assign n8901 = n3031 | n3644 ;
  assign n8902 = n8901 ^ n1793 ^ 1'b0 ;
  assign n8903 = n4020 ^ n1344 ^ 1'b0 ;
  assign n8904 = n5913 ^ n4218 ^ 1'b0 ;
  assign n8905 = ~n851 & n8904 ;
  assign n8906 = n1333 ^ n558 ^ 1'b0 ;
  assign n8907 = n1753 | n8906 ;
  assign n8908 = n1419 | n7235 ;
  assign n8909 = n5469 ^ n1569 ^ 1'b0 ;
  assign n8910 = n8908 & n8909 ;
  assign n8911 = ~x106 & n4230 ;
  assign n8912 = n8911 ^ n558 ^ 1'b0 ;
  assign n8913 = n1329 & ~n8912 ;
  assign n8914 = ~n2232 & n8913 ;
  assign n8915 = ~n1808 & n6684 ;
  assign n8916 = n3691 & n8915 ;
  assign n8917 = ~n259 & n1470 ;
  assign n8918 = n8917 ^ n7821 ^ 1'b0 ;
  assign n8920 = ~n1645 & n6894 ;
  assign n8921 = n5064 & n8920 ;
  assign n8919 = n4974 & n6671 ;
  assign n8922 = n8921 ^ n8919 ^ 1'b0 ;
  assign n8926 = n4501 ^ n2318 ^ 1'b0 ;
  assign n8927 = n4009 & n8926 ;
  assign n8923 = n4162 & n5688 ;
  assign n8924 = n245 & n8923 ;
  assign n8925 = n1354 & ~n8924 ;
  assign n8928 = n8927 ^ n8925 ^ 1'b0 ;
  assign n8929 = n8928 ^ n5715 ^ 1'b0 ;
  assign n8930 = x56 & ~n8929 ;
  assign n8931 = x73 & n1663 ;
  assign n8932 = ~n1663 & n2261 ;
  assign n8933 = n8932 ^ x39 ^ 1'b0 ;
  assign n8934 = n8933 ^ x94 ^ 1'b0 ;
  assign n8935 = x89 & n8934 ;
  assign n8936 = n8935 ^ n8209 ^ 1'b0 ;
  assign n8937 = ~n473 & n866 ;
  assign n8938 = ( n6259 & ~n7530 ) | ( n6259 & n8937 ) | ( ~n7530 & n8937 ) ;
  assign n8939 = ~x11 & n3846 ;
  assign n8940 = n8939 ^ n1991 ^ 1'b0 ;
  assign n8941 = ~n7996 & n8940 ;
  assign n8942 = ~n868 & n2178 ;
  assign n8947 = n634 & n6567 ;
  assign n8948 = ~n6053 & n8947 ;
  assign n8944 = n273 | n7462 ;
  assign n8945 = n8944 ^ n950 ^ 1'b0 ;
  assign n8946 = n5202 & ~n8945 ;
  assign n8949 = n8948 ^ n8946 ^ 1'b0 ;
  assign n8950 = ~n134 & n8949 ;
  assign n8943 = x95 & n4415 ;
  assign n8951 = n8950 ^ n8943 ^ 1'b0 ;
  assign n8952 = n3382 & ~n8779 ;
  assign n8953 = n2935 ^ n360 ^ 1'b0 ;
  assign n8954 = n2231 & n8953 ;
  assign n8955 = ~n2831 & n7182 ;
  assign n8956 = n8954 & ~n8955 ;
  assign n8957 = n8582 ^ n6832 ^ 1'b0 ;
  assign n8958 = n4571 & ~n8957 ;
  assign n8959 = ( ~n770 & n4100 ) | ( ~n770 & n8286 ) | ( n4100 & n8286 ) ;
  assign n8960 = ~n1010 & n2425 ;
  assign n8961 = n8960 ^ n353 ^ 1'b0 ;
  assign n8962 = n4314 & ~n8961 ;
  assign n8963 = n8962 ^ n660 ^ 1'b0 ;
  assign n8964 = n6024 ^ n2456 ^ 1'b0 ;
  assign n8965 = n6448 & ~n8964 ;
  assign n8966 = n2238 | n8965 ;
  assign n8967 = n482 & ~n2911 ;
  assign n8968 = n8966 & n8967 ;
  assign n8969 = n6057 & ~n7643 ;
  assign n8970 = n8969 ^ n394 ^ 1'b0 ;
  assign n8971 = n8392 ^ n6640 ^ 1'b0 ;
  assign n8972 = n5350 | n8971 ;
  assign n8973 = n5249 ^ n336 ^ 1'b0 ;
  assign n8974 = n7915 ^ n2374 ^ 1'b0 ;
  assign n8975 = n8067 & ~n8974 ;
  assign n8976 = n2212 ^ n786 ^ 1'b0 ;
  assign n8977 = n2649 & ~n8976 ;
  assign n8978 = ~n1945 & n8977 ;
  assign n8979 = n547 & n2993 ;
  assign n8980 = n8979 ^ n4196 ^ 1'b0 ;
  assign n8981 = n7732 | n8427 ;
  assign n8982 = n8980 & ~n8981 ;
  assign n8983 = n8840 | n8982 ;
  assign n8984 = n6088 ^ n5986 ^ n2651 ;
  assign n8985 = n444 | n5977 ;
  assign n8986 = n4279 ^ n1899 ^ 1'b0 ;
  assign n8987 = n5096 | n7781 ;
  assign n8988 = n3244 & n7339 ;
  assign n8989 = ~n7272 & n8988 ;
  assign n8990 = n3966 ^ x31 ^ 1'b0 ;
  assign n8991 = ~n3280 & n8990 ;
  assign n8992 = n283 & n8991 ;
  assign n8993 = n6557 ^ n4013 ^ 1'b0 ;
  assign n8994 = x54 & ~n1046 ;
  assign n8995 = n5018 & ~n8994 ;
  assign n8996 = n4218 & n8995 ;
  assign n8997 = n8996 ^ n420 ^ 1'b0 ;
  assign n8998 = n3840 & n5938 ;
  assign n8999 = n8998 ^ n3114 ^ 1'b0 ;
  assign n9000 = n2253 | n6378 ;
  assign n9001 = n5432 | n9000 ;
  assign n9002 = n4056 ^ n571 ^ 1'b0 ;
  assign n9003 = ~n1532 & n9002 ;
  assign n9004 = n215 & ~n2240 ;
  assign n9005 = n3126 & ~n9004 ;
  assign n9006 = n4282 ^ n1046 ^ 1'b0 ;
  assign n9007 = n9005 & ~n9006 ;
  assign n9008 = n9007 ^ n5006 ^ 1'b0 ;
  assign n9009 = n4730 | n9008 ;
  assign n9010 = n9003 & ~n9009 ;
  assign n9011 = n9010 ^ n6401 ^ 1'b0 ;
  assign n9012 = n4580 & n8892 ;
  assign n9013 = n9012 ^ n7057 ^ 1'b0 ;
  assign n9014 = x8 | n323 ;
  assign n9015 = n1706 & n8937 ;
  assign n9016 = n3156 & n4300 ;
  assign n9017 = n610 & ~n5749 ;
  assign n9018 = n5273 & n9017 ;
  assign n9019 = n9018 ^ n4579 ^ 1'b0 ;
  assign n9020 = ~n2194 & n9019 ;
  assign n9021 = n3587 & n9020 ;
  assign n9022 = n5230 & n8651 ;
  assign n9023 = x127 & ~n1588 ;
  assign n9024 = n9023 ^ x55 ^ 1'b0 ;
  assign n9025 = ~n1034 & n4416 ;
  assign n9026 = n9025 ^ n4406 ^ 1'b0 ;
  assign n9027 = n9026 ^ n3488 ^ 1'b0 ;
  assign n9028 = ~n8258 & n9027 ;
  assign n9029 = n2019 & n5970 ;
  assign n9030 = n9029 ^ n1420 ^ 1'b0 ;
  assign n9031 = ~n516 & n2566 ;
  assign n9032 = n3614 ^ n3468 ^ 1'b0 ;
  assign n9033 = ~n4513 & n9032 ;
  assign n9034 = ~n9031 & n9033 ;
  assign n9035 = n5965 ^ n1770 ^ 1'b0 ;
  assign n9036 = n8047 ^ n1994 ^ 1'b0 ;
  assign n9037 = n6433 | n8343 ;
  assign n9038 = n5403 & ~n9037 ;
  assign n9039 = n1899 & ~n7547 ;
  assign n9040 = n9039 ^ n5485 ^ 1'b0 ;
  assign n9044 = n4332 ^ n2530 ^ 1'b0 ;
  assign n9045 = n2191 & n9044 ;
  assign n9046 = n3700 & ~n4029 ;
  assign n9047 = n9046 ^ n1126 ^ 1'b0 ;
  assign n9048 = n4564 & n9047 ;
  assign n9049 = ~n9045 & n9048 ;
  assign n9041 = n2266 & ~n5893 ;
  assign n9042 = n9041 ^ n8499 ^ 1'b0 ;
  assign n9043 = n2385 & ~n9042 ;
  assign n9050 = n9049 ^ n9043 ^ 1'b0 ;
  assign n9051 = n3633 | n6580 ;
  assign n9052 = n5586 ^ n1877 ^ 1'b0 ;
  assign n9053 = ~n2885 & n9052 ;
  assign n9054 = ~n1149 & n3340 ;
  assign n9055 = n9054 ^ n5865 ^ 1'b0 ;
  assign n9056 = n3602 & n9055 ;
  assign n9057 = n3132 ^ n811 ^ 1'b0 ;
  assign n9058 = n9057 ^ n1135 ^ 1'b0 ;
  assign n9059 = n4117 & ~n4144 ;
  assign n9060 = n6376 ^ n4658 ^ 1'b0 ;
  assign n9061 = x126 & ~n5335 ;
  assign n9062 = n9061 ^ n3201 ^ 1'b0 ;
  assign n9063 = n9062 ^ n2528 ^ 1'b0 ;
  assign n9064 = n6782 | n9063 ;
  assign n9065 = n229 & ~n5233 ;
  assign n9066 = ~n7954 & n9065 ;
  assign n9067 = n358 & ~n3477 ;
  assign n9068 = n9067 ^ n3320 ^ 1'b0 ;
  assign n9069 = n1186 ^ n707 ^ 1'b0 ;
  assign n9070 = n9069 ^ n7231 ^ 1'b0 ;
  assign n9071 = n2532 & n6470 ;
  assign n9072 = ~n1558 & n7295 ;
  assign n9073 = n8827 ^ n5732 ^ 1'b0 ;
  assign n9074 = n3492 | n9073 ;
  assign n9075 = n1880 | n9074 ;
  assign n9076 = ~n9072 & n9075 ;
  assign n9077 = n794 & ~n2107 ;
  assign n9078 = n8079 & n9077 ;
  assign n9079 = n9078 ^ n5338 ^ 1'b0 ;
  assign n9082 = ~n4939 & n5091 ;
  assign n9081 = n4567 ^ n361 ^ 1'b0 ;
  assign n9080 = n1609 & ~n6285 ;
  assign n9083 = n9082 ^ n9081 ^ n9080 ;
  assign n9084 = ~n1437 & n5956 ;
  assign n9085 = n3322 & n9084 ;
  assign n9086 = n1102 & n9085 ;
  assign n9087 = n9086 ^ x60 ^ 1'b0 ;
  assign n9088 = n2479 & n7118 ;
  assign n9089 = n696 | n2635 ;
  assign n9090 = ~n2515 & n4790 ;
  assign n9091 = ~n6024 & n9090 ;
  assign n9092 = n9091 ^ n4323 ^ 1'b0 ;
  assign n9093 = ~n3622 & n9092 ;
  assign n9095 = n2694 & ~n8589 ;
  assign n9094 = n616 & ~n5833 ;
  assign n9096 = n9095 ^ n9094 ^ 1'b0 ;
  assign n9097 = n6064 & ~n9096 ;
  assign n9098 = n9097 ^ n5806 ^ 1'b0 ;
  assign n9106 = n5582 ^ n988 ^ 1'b0 ;
  assign n9107 = ~n4224 & n9106 ;
  assign n9100 = n1501 | n6203 ;
  assign n9101 = n5094 | n9100 ;
  assign n9099 = n1144 | n4150 ;
  assign n9102 = n9101 ^ n9099 ^ 1'b0 ;
  assign n9103 = n1808 & ~n9102 ;
  assign n9104 = n1800 | n8722 ;
  assign n9105 = n9103 & ~n9104 ;
  assign n9108 = n9107 ^ n9105 ^ 1'b0 ;
  assign n9109 = n300 | n1197 ;
  assign n9110 = n3797 & n7172 ;
  assign n9111 = n7210 & n9110 ;
  assign n9112 = n1057 & ~n7364 ;
  assign n9113 = n9112 ^ n6083 ^ 1'b0 ;
  assign n9114 = n8765 ^ n2390 ^ 1'b0 ;
  assign n9115 = n9114 ^ n3632 ^ 1'b0 ;
  assign n9116 = n9113 & ~n9115 ;
  assign n9117 = n3554 | n5579 ;
  assign n9118 = n4322 | n9117 ;
  assign n9119 = n7004 ^ n3208 ^ 1'b0 ;
  assign n9120 = ( n3070 & ~n5257 ) | ( n3070 & n8590 ) | ( ~n5257 & n8590 ) ;
  assign n9121 = n9120 ^ n555 ^ 1'b0 ;
  assign n9122 = n7421 | n9121 ;
  assign n9123 = n1895 | n4513 ;
  assign n9124 = n9123 ^ n6544 ^ 1'b0 ;
  assign n9125 = n570 & ~n4394 ;
  assign n9126 = n9124 & n9125 ;
  assign n9127 = n8947 ^ n930 ^ 1'b0 ;
  assign n9128 = n870 | n9127 ;
  assign n9129 = n3108 ^ n830 ^ 1'b0 ;
  assign n9130 = n367 & ~n529 ;
  assign n9131 = n3286 ^ n3149 ^ 1'b0 ;
  assign n9132 = ~n3428 & n9131 ;
  assign n9133 = ~n4713 & n9132 ;
  assign n9134 = n9133 ^ n1793 ^ 1'b0 ;
  assign n9135 = ~n9130 & n9134 ;
  assign n9136 = ~n2638 & n5974 ;
  assign n9138 = ~n3363 & n3466 ;
  assign n9137 = n6280 | n6298 ;
  assign n9139 = n9138 ^ n9137 ^ 1'b0 ;
  assign n9140 = ~n928 & n1292 ;
  assign n9141 = n9140 ^ x47 ^ 1'b0 ;
  assign n9142 = ~x12 & n9141 ;
  assign n9143 = ~n812 & n5564 ;
  assign n9144 = n9143 ^ n2827 ^ 1'b0 ;
  assign n9145 = ~n8896 & n9144 ;
  assign n9146 = n2293 ^ n1414 ^ 1'b0 ;
  assign n9147 = n1513 | n3983 ;
  assign n9148 = n1146 | n9147 ;
  assign n9149 = n9148 ^ n3547 ^ 1'b0 ;
  assign n9150 = n3826 ^ n3552 ^ 1'b0 ;
  assign n9151 = n3060 ^ x22 ^ 1'b0 ;
  assign n9152 = n4216 & ~n9151 ;
  assign n9153 = n7539 ^ n3223 ^ 1'b0 ;
  assign n9154 = n4304 & ~n9153 ;
  assign n9155 = n5252 & n9154 ;
  assign n9156 = ~n3246 & n9155 ;
  assign n9157 = n4084 ^ n2711 ^ n252 ;
  assign n9158 = n2526 | n9157 ;
  assign n9159 = n2533 ^ n1324 ^ 1'b0 ;
  assign n9160 = n9159 ^ n2691 ^ 1'b0 ;
  assign n9161 = n623 & n9160 ;
  assign n9162 = ~n5487 & n7982 ;
  assign n9163 = n5590 ^ n217 ^ 1'b0 ;
  assign n9164 = n9162 | n9163 ;
  assign n9165 = ~n4853 & n9164 ;
  assign n9166 = n375 | n6722 ;
  assign n9167 = n502 | n7004 ;
  assign n9168 = n179 & ~n9167 ;
  assign n9169 = n4112 & n7938 ;
  assign n9170 = n6528 ^ n1899 ^ 1'b0 ;
  assign n9171 = n1880 & n9170 ;
  assign n9172 = n9171 ^ n3618 ^ 1'b0 ;
  assign n9173 = n4208 ^ n2978 ^ n1515 ;
  assign n9175 = n3082 & ~n3672 ;
  assign n9174 = n1625 | n7875 ;
  assign n9176 = n9175 ^ n9174 ^ 1'b0 ;
  assign n9177 = n6499 | n9176 ;
  assign n9178 = n9173 & ~n9177 ;
  assign n9179 = n1644 & n3608 ;
  assign n9180 = ~n1147 & n4486 ;
  assign n9181 = n4023 & n9180 ;
  assign n9182 = n9181 ^ n1769 ^ n1284 ;
  assign n9183 = ( n2937 & n3087 ) | ( n2937 & ~n9182 ) | ( n3087 & ~n9182 ) ;
  assign n9184 = n5692 ^ n1395 ^ 1'b0 ;
  assign n9185 = n2608 | n9184 ;
  assign n9186 = ~n1487 & n3090 ;
  assign n9187 = ~n549 & n6419 ;
  assign n9188 = ~n7338 & n8514 ;
  assign n9189 = n6902 & n9188 ;
  assign n9190 = n9189 ^ n7848 ^ 1'b0 ;
  assign n9191 = n1854 | n4303 ;
  assign n9192 = n2520 & ~n9191 ;
  assign n9193 = ~n1361 & n2009 ;
  assign n9194 = n9192 & n9193 ;
  assign n9195 = n4745 ^ n1870 ^ 1'b0 ;
  assign n9196 = n9194 | n9195 ;
  assign n9197 = n9196 ^ n6239 ^ 1'b0 ;
  assign n9198 = n3594 | n4521 ;
  assign n9199 = n1453 & ~n2677 ;
  assign n9200 = n9199 ^ n391 ^ 1'b0 ;
  assign n9201 = ~n4253 & n9200 ;
  assign n9202 = n5282 | n9201 ;
  assign n9203 = n353 & ~n9202 ;
  assign n9204 = n1323 & ~n9203 ;
  assign n9205 = n9204 ^ n2171 ^ 1'b0 ;
  assign n9206 = n7094 ^ n2271 ^ 1'b0 ;
  assign n9207 = ~n886 & n9206 ;
  assign n9208 = n1765 & n4098 ;
  assign n9209 = n3983 ^ n2306 ^ 1'b0 ;
  assign n9210 = n4924 & ~n9209 ;
  assign n9211 = n9210 ^ n5488 ^ 1'b0 ;
  assign n9212 = n1625 | n9211 ;
  assign n9213 = n3053 & ~n9212 ;
  assign n9214 = ~n8297 & n8637 ;
  assign n9215 = n7121 & n8190 ;
  assign n9219 = n307 | n1212 ;
  assign n9216 = n2168 ^ n1858 ^ 1'b0 ;
  assign n9217 = n4162 & n9216 ;
  assign n9218 = n9217 ^ n3021 ^ 1'b0 ;
  assign n9220 = n9219 ^ n9218 ^ n3193 ;
  assign n9221 = n6073 & ~n6115 ;
  assign n9222 = n9221 ^ n1506 ^ 1'b0 ;
  assign n9223 = n9222 ^ n1743 ^ 1'b0 ;
  assign n9224 = x120 & ~n9223 ;
  assign n9225 = n4824 ^ n4674 ^ 1'b0 ;
  assign n9226 = ~n200 & n9225 ;
  assign n9227 = n6991 ^ n3824 ^ 1'b0 ;
  assign n9228 = n412 | n2987 ;
  assign n9229 = n9228 ^ n9102 ^ 1'b0 ;
  assign n9230 = x47 & n9229 ;
  assign n9231 = n2623 ^ n1510 ^ 1'b0 ;
  assign n9232 = n3124 | n9231 ;
  assign n9233 = n3446 | n9232 ;
  assign n9234 = n1361 & ~n9233 ;
  assign n9235 = n1817 & n9234 ;
  assign n9236 = n2467 & n9235 ;
  assign n9237 = n9230 & n9236 ;
  assign n9238 = n660 | n1022 ;
  assign n9239 = n5682 & n9238 ;
  assign n9244 = n2091 ^ n375 ^ n279 ;
  assign n9240 = n921 ^ n392 ^ 1'b0 ;
  assign n9241 = ~n889 & n9240 ;
  assign n9242 = n9241 ^ n5235 ^ 1'b0 ;
  assign n9243 = ~n983 & n9242 ;
  assign n9245 = n9244 ^ n9243 ^ 1'b0 ;
  assign n9246 = n8738 ^ n3926 ^ 1'b0 ;
  assign n9247 = n8529 & n9246 ;
  assign n9248 = n1087 & n4277 ;
  assign n9249 = ~n3706 & n9248 ;
  assign n9250 = ~n3310 & n9249 ;
  assign n9251 = n7175 ^ n4842 ^ 1'b0 ;
  assign n9252 = n1628 ^ x54 ^ 1'b0 ;
  assign n9253 = n4188 & ~n4240 ;
  assign n9254 = ~n9252 & n9253 ;
  assign n9255 = n493 & ~n6663 ;
  assign n9256 = n9255 ^ n1534 ^ 1'b0 ;
  assign n9257 = n1624 ^ n391 ^ 1'b0 ;
  assign n9258 = n2058 ^ n444 ^ 1'b0 ;
  assign n9259 = n2486 & n3998 ;
  assign n9260 = n7887 & ~n8188 ;
  assign n9261 = n9260 ^ n2601 ^ 1'b0 ;
  assign n9262 = x37 & n9261 ;
  assign n9263 = n6156 | n6550 ;
  assign n9264 = n5287 | n9263 ;
  assign n9265 = n9264 ^ n4809 ^ 1'b0 ;
  assign n9266 = n5243 ^ n4244 ^ 1'b0 ;
  assign n9267 = n931 & ~n8058 ;
  assign n9268 = ~n1329 & n4687 ;
  assign n9269 = n2792 ^ n1779 ^ 1'b0 ;
  assign n9270 = n4185 & ~n9269 ;
  assign n9271 = n9031 ^ n4102 ^ 1'b0 ;
  assign n9272 = ~n5855 & n9271 ;
  assign n9273 = n9272 ^ n5501 ^ 1'b0 ;
  assign n9274 = n7177 ^ n4791 ^ 1'b0 ;
  assign n9275 = n9274 ^ n2073 ^ 1'b0 ;
  assign n9276 = ~n2743 & n4736 ;
  assign n9277 = ~n7506 & n9276 ;
  assign n9278 = n4681 & n8307 ;
  assign n9279 = n406 & n9278 ;
  assign n9280 = n492 & n6271 ;
  assign n9281 = n8206 ^ n2291 ^ 1'b0 ;
  assign n9282 = n5429 ^ n3072 ^ 1'b0 ;
  assign n9283 = n5522 | n9282 ;
  assign n9284 = n7061 & ~n9283 ;
  assign n9285 = n2451 & n9284 ;
  assign n9286 = n3999 | n9285 ;
  assign n9287 = n6746 ^ n2958 ^ 1'b0 ;
  assign n9288 = n7244 | n9287 ;
  assign n9289 = ~n1394 & n1710 ;
  assign n9290 = n5068 & ~n9289 ;
  assign n9291 = n868 | n9290 ;
  assign n9292 = n7061 | n9291 ;
  assign n9293 = n507 & ~n4965 ;
  assign n9294 = n9203 & n9293 ;
  assign n9295 = n2393 & ~n3906 ;
  assign n9296 = n2600 ^ n1478 ^ 1'b0 ;
  assign n9297 = n3629 & n9296 ;
  assign n9298 = x23 & n9297 ;
  assign n9299 = n9295 & n9298 ;
  assign n9300 = ~n2997 & n3504 ;
  assign n9301 = ~n276 & n763 ;
  assign n9302 = n9301 ^ n6371 ^ 1'b0 ;
  assign n9303 = ~n245 & n6805 ;
  assign n9304 = n9303 ^ n3474 ^ 1'b0 ;
  assign n9305 = ~x53 & n9304 ;
  assign n9308 = n3090 ^ n259 ^ 1'b0 ;
  assign n9306 = n739 & ~n1491 ;
  assign n9307 = n5447 & n9306 ;
  assign n9309 = n9308 ^ n9307 ^ 1'b0 ;
  assign n9310 = n1381 & n9309 ;
  assign n9311 = n1080 ^ n698 ^ 1'b0 ;
  assign n9312 = n1483 | n7784 ;
  assign n9313 = n1247 | n1361 ;
  assign n9314 = n7354 ^ n2243 ^ 1'b0 ;
  assign n9315 = ~n5809 & n9314 ;
  assign n9316 = n9315 ^ n3544 ^ 1'b0 ;
  assign n9317 = n3401 ^ n823 ^ 1'b0 ;
  assign n9318 = ~n1487 & n9317 ;
  assign n9319 = n9316 & n9318 ;
  assign n9320 = n9319 ^ n6874 ^ 1'b0 ;
  assign n9321 = n9320 ^ n1069 ^ 1'b0 ;
  assign n9322 = ( n1170 & ~n5038 ) | ( n1170 & n5961 ) | ( ~n5038 & n5961 ) ;
  assign n9323 = n5859 ^ n2070 ^ 1'b0 ;
  assign n9324 = n9323 ^ n6644 ^ n450 ;
  assign n9325 = n3262 ^ n3201 ^ 1'b0 ;
  assign n9326 = n2360 | n9325 ;
  assign n9327 = n3756 ^ n885 ^ 1'b0 ;
  assign n9328 = n2002 | n9327 ;
  assign n9329 = n978 | n6028 ;
  assign n9330 = n9328 & ~n9329 ;
  assign n9331 = n7114 | n9330 ;
  assign n9332 = n9331 ^ n6634 ^ 1'b0 ;
  assign n9335 = n1579 & ~n2503 ;
  assign n9336 = ~n360 & n9335 ;
  assign n9337 = n7422 & n9336 ;
  assign n9333 = n1530 & n4196 ;
  assign n9334 = ~n6151 & n9333 ;
  assign n9338 = n9337 ^ n9334 ^ 1'b0 ;
  assign n9339 = n4198 & ~n7735 ;
  assign n9340 = n9339 ^ n346 ^ 1'b0 ;
  assign n9341 = n9340 ^ n5913 ^ 1'b0 ;
  assign n9342 = n2658 | n6705 ;
  assign n9343 = n9342 ^ n8210 ^ 1'b0 ;
  assign n9344 = n335 ^ x67 ^ 1'b0 ;
  assign n9345 = ~n2166 & n3675 ;
  assign n9346 = ~n1548 & n9345 ;
  assign n9347 = n9346 ^ n5527 ^ 1'b0 ;
  assign n9348 = ~n1033 & n5816 ;
  assign n9349 = n9348 ^ x15 ^ 1'b0 ;
  assign n9350 = n3381 ^ n1208 ^ 1'b0 ;
  assign n9351 = ( x95 & x105 ) | ( x95 & n238 ) | ( x105 & n238 ) ;
  assign n9352 = n7404 & n9351 ;
  assign n9353 = n9350 & n9352 ;
  assign n9354 = n8757 ^ n610 ^ 1'b0 ;
  assign n9355 = n4385 | n7640 ;
  assign n9356 = ~n5388 & n6278 ;
  assign n9357 = ~n2319 & n4345 ;
  assign n9358 = ~n1498 & n5118 ;
  assign n9359 = ~n1444 & n9358 ;
  assign n9360 = n3629 | n9359 ;
  assign n9361 = n6729 | n9360 ;
  assign n9362 = n6038 | n9361 ;
  assign n9363 = ~n9357 & n9362 ;
  assign n9364 = n9363 ^ n3613 ^ 1'b0 ;
  assign n9365 = ~n1151 & n8817 ;
  assign n9373 = n924 | n4053 ;
  assign n9367 = ~n1243 & n2512 ;
  assign n9368 = n4194 & ~n9367 ;
  assign n9366 = ~n3333 & n4280 ;
  assign n9369 = n9368 ^ n9366 ^ 1'b0 ;
  assign n9370 = ~n5132 & n9369 ;
  assign n9371 = n4873 ^ n250 ^ 1'b0 ;
  assign n9372 = n9370 & ~n9371 ;
  assign n9374 = n9373 ^ n9372 ^ 1'b0 ;
  assign n9375 = n435 | n2198 ;
  assign n9376 = n9375 ^ n3262 ^ 1'b0 ;
  assign n9377 = ~n677 & n7076 ;
  assign n9378 = n9377 ^ n252 ^ 1'b0 ;
  assign n9379 = n3453 ^ n2310 ^ 1'b0 ;
  assign n9380 = n5025 & n9379 ;
  assign n9384 = ~n428 & n2554 ;
  assign n9385 = ~n1035 & n9384 ;
  assign n9381 = n984 & n3504 ;
  assign n9382 = n9381 ^ n6850 ^ 1'b0 ;
  assign n9383 = ~n9381 & n9382 ;
  assign n9386 = n9385 ^ n9383 ^ 1'b0 ;
  assign n9387 = n1099 & ~n6177 ;
  assign n9388 = ~n530 & n1299 ;
  assign n9389 = n9388 ^ n2604 ^ 1'b0 ;
  assign n9390 = n8101 ^ n3091 ^ 1'b0 ;
  assign n9391 = n9389 | n9390 ;
  assign n9392 = n7574 & ~n9391 ;
  assign n9393 = n1060 & n9392 ;
  assign n9394 = n4882 & ~n8808 ;
  assign n9395 = ~n1204 & n9394 ;
  assign n9396 = n986 ^ n799 ^ 1'b0 ;
  assign n9397 = ~n9395 & n9396 ;
  assign n9398 = n6519 ^ n4307 ^ n3512 ;
  assign n9399 = n6166 | n9398 ;
  assign n9405 = n571 | n1467 ;
  assign n9406 = n9405 ^ n1990 ^ 1'b0 ;
  assign n9407 = n1848 & ~n1903 ;
  assign n9408 = n9406 & n9407 ;
  assign n9400 = ~x42 & n3788 ;
  assign n9401 = n9400 ^ n4602 ^ 1'b0 ;
  assign n9402 = n1849 | n9401 ;
  assign n9403 = n9402 ^ n4414 ^ 1'b0 ;
  assign n9404 = n6638 & n9403 ;
  assign n9409 = n9408 ^ n9404 ^ 1'b0 ;
  assign n9410 = ~n1784 & n8086 ;
  assign n9411 = n9409 & ~n9410 ;
  assign n9412 = ~n4414 & n5416 ;
  assign n9413 = n2707 | n2911 ;
  assign n9414 = n201 & n482 ;
  assign n9415 = n3229 ^ n1133 ^ 1'b0 ;
  assign n9416 = n1333 & ~n2173 ;
  assign n9417 = n9416 ^ n2146 ^ 1'b0 ;
  assign n9418 = ~n7153 & n9417 ;
  assign n9419 = n882 & n1290 ;
  assign n9420 = ~n1724 & n4710 ;
  assign n9421 = n5741 & n9420 ;
  assign n9422 = n8094 & n9421 ;
  assign n9423 = n9275 ^ n3462 ^ n354 ;
  assign n9424 = ~n3465 & n8270 ;
  assign n9425 = n6453 ^ n4126 ^ 1'b0 ;
  assign n9426 = n5817 & n6958 ;
  assign n9427 = n9425 & n9426 ;
  assign n9428 = n6309 ^ n6085 ^ 1'b0 ;
  assign n9429 = n9427 & ~n9428 ;
  assign n9430 = n6469 ^ n724 ^ 1'b0 ;
  assign n9431 = n307 | n9430 ;
  assign n9432 = n5519 & ~n9431 ;
  assign n9433 = n4321 & n9432 ;
  assign n9434 = n3074 & n9433 ;
  assign n9435 = n8993 & n9434 ;
  assign n9436 = n3354 | n9435 ;
  assign n9437 = n1846 | n9436 ;
  assign n9438 = n2838 | n4814 ;
  assign n9439 = n6561 & ~n9438 ;
  assign n9440 = ~n1054 & n2198 ;
  assign n9441 = n9350 & n9440 ;
  assign n9442 = n9441 ^ n4027 ^ 1'b0 ;
  assign n9443 = n2016 | n3428 ;
  assign n9444 = n1201 & ~n9443 ;
  assign n9445 = n2677 & ~n6930 ;
  assign n9446 = n4875 & ~n9445 ;
  assign n9447 = n8664 ^ n5254 ^ 1'b0 ;
  assign n9448 = n1325 ^ n507 ^ 1'b0 ;
  assign n9449 = n7261 ^ n6194 ^ n528 ;
  assign n9450 = n1270 | n5816 ;
  assign n9451 = n642 & ~n7922 ;
  assign n9452 = n300 & n9451 ;
  assign n9453 = n363 & n3968 ;
  assign n9454 = n9453 ^ n514 ^ 1'b0 ;
  assign n9455 = n9454 ^ n4578 ^ 1'b0 ;
  assign n9456 = n2533 ^ n227 ^ 1'b0 ;
  assign n9457 = n844 & ~n3737 ;
  assign n9458 = ~n9456 & n9457 ;
  assign n9459 = n1540 ^ n1346 ^ 1'b0 ;
  assign n9460 = n9459 ^ n1996 ^ 1'b0 ;
  assign n9461 = n9458 | n9460 ;
  assign n9462 = n7670 & n8093 ;
  assign n9463 = n6483 ^ n3450 ^ 1'b0 ;
  assign n9464 = n5237 & n9463 ;
  assign n9465 = n1042 | n9464 ;
  assign n9467 = n2226 & ~n4417 ;
  assign n9468 = n1069 & n9467 ;
  assign n9466 = ~n5883 & n8140 ;
  assign n9469 = n9468 ^ n9466 ^ 1'b0 ;
  assign n9470 = ( n5064 & n9465 ) | ( n5064 & ~n9469 ) | ( n9465 & ~n9469 ) ;
  assign n9471 = ( n503 & ~n4458 ) | ( n503 & n8315 ) | ( ~n4458 & n8315 ) ;
  assign n9472 = n9471 ^ n8064 ^ 1'b0 ;
  assign n9473 = ~n4177 & n9472 ;
  assign n9474 = n1513 & n9362 ;
  assign n9475 = n192 | n4291 ;
  assign n9476 = n1890 & n2355 ;
  assign n9477 = ~n528 & n9476 ;
  assign n9478 = n7172 & ~n9477 ;
  assign n9479 = n9478 ^ n6488 ^ 1'b0 ;
  assign n9480 = x126 & ~n7231 ;
  assign n9481 = ( ~n1268 & n3929 ) | ( ~n1268 & n9480 ) | ( n3929 & n9480 ) ;
  assign n9482 = n2653 ^ n2026 ^ 1'b0 ;
  assign n9483 = n482 & ~n3258 ;
  assign n9484 = n335 & n2037 ;
  assign n9485 = n9483 & ~n9484 ;
  assign n9486 = n7101 & n9485 ;
  assign n9487 = n3986 & n9486 ;
  assign n9491 = n1792 ^ n287 ^ 1'b0 ;
  assign n9492 = n4525 & ~n9491 ;
  assign n9488 = n963 ^ n311 ^ 1'b0 ;
  assign n9489 = n9488 ^ n834 ^ 1'b0 ;
  assign n9490 = n2182 & n9489 ;
  assign n9493 = n9492 ^ n9490 ^ 1'b0 ;
  assign n9494 = ~n4056 & n9493 ;
  assign n9495 = n6873 & n7444 ;
  assign n9496 = n3353 & n6225 ;
  assign n9497 = n4376 & n9496 ;
  assign n9498 = n3023 & ~n3289 ;
  assign n9499 = n6456 ^ n4287 ^ 1'b0 ;
  assign n9500 = ~n9498 & n9499 ;
  assign n9501 = n9497 | n9500 ;
  assign n9502 = n3369 ^ n2331 ^ 1'b0 ;
  assign n9503 = n1172 & ~n7463 ;
  assign n9504 = n717 & n1618 ;
  assign n9505 = n1262 & n9504 ;
  assign n9506 = ~n1895 & n9505 ;
  assign n9507 = n9351 ^ n6857 ^ 1'b0 ;
  assign n9508 = n9507 ^ n8179 ^ 1'b0 ;
  assign n9510 = ( n792 & ~n1833 ) | ( n792 & n7462 ) | ( ~n1833 & n7462 ) ;
  assign n9509 = n570 & ~n4871 ;
  assign n9511 = n9510 ^ n9509 ^ 1'b0 ;
  assign n9512 = ~n3475 & n5014 ;
  assign n9513 = n7278 ^ n2980 ^ n1477 ;
  assign n9514 = ~n8714 & n9513 ;
  assign n9515 = x60 & ~n4679 ;
  assign n9516 = ~n4423 & n9515 ;
  assign n9517 = n9516 ^ n5243 ^ 1'b0 ;
  assign n9518 = n3699 | n6685 ;
  assign n9519 = n1695 & ~n9518 ;
  assign n9520 = n530 | n7191 ;
  assign n9522 = n7456 & ~n8590 ;
  assign n9521 = n7001 ^ n707 ^ 1'b0 ;
  assign n9523 = n9522 ^ n9521 ^ 1'b0 ;
  assign n9524 = n1329 | n1398 ;
  assign n9525 = n9524 ^ x34 ^ 1'b0 ;
  assign n9526 = ~n4658 & n9525 ;
  assign n9527 = ~n593 & n1777 ;
  assign n9528 = ~n1908 & n9527 ;
  assign n9529 = n9528 ^ n2948 ^ 1'b0 ;
  assign n9530 = ~n1898 & n9529 ;
  assign n9531 = ~n857 & n1072 ;
  assign n9532 = x50 & ~n3628 ;
  assign n9533 = ~n5351 & n9532 ;
  assign n9534 = ~n6496 & n8731 ;
  assign n9535 = n6437 ^ n5938 ^ 1'b0 ;
  assign n9536 = n6515 & ~n9535 ;
  assign n9538 = x17 & n9483 ;
  assign n9539 = n9538 ^ n5202 ^ 1'b0 ;
  assign n9540 = n2651 & ~n3615 ;
  assign n9541 = ~n9539 & n9540 ;
  assign n9537 = n2826 | n7832 ;
  assign n9542 = n9541 ^ n9537 ^ 1'b0 ;
  assign n9543 = n4611 ^ n2245 ^ 1'b0 ;
  assign n9544 = n4759 & ~n9543 ;
  assign n9546 = n6996 ^ n1849 ^ 1'b0 ;
  assign n9545 = n1207 | n6173 ;
  assign n9547 = n9546 ^ n9545 ^ 1'b0 ;
  assign n9548 = n1912 & n3759 ;
  assign n9549 = n3826 | n9462 ;
  assign n9550 = n450 & n6522 ;
  assign n9551 = n9550 ^ n161 ^ 1'b0 ;
  assign n9552 = n4181 | n9551 ;
  assign n9553 = n1761 | n9552 ;
  assign n9554 = n3354 ^ n2478 ^ 1'b0 ;
  assign n9555 = n3619 ^ x37 ^ 1'b0 ;
  assign n9556 = ~n6423 & n9555 ;
  assign n9557 = n5324 & n6919 ;
  assign n9558 = n1716 & n3934 ;
  assign n9559 = ~n9557 & n9558 ;
  assign n9560 = n5235 & n7954 ;
  assign n9568 = n1784 ^ n1235 ^ 1'b0 ;
  assign n9561 = n5618 ^ n794 ^ 1'b0 ;
  assign n9562 = n1118 | n9561 ;
  assign n9563 = n5839 & ~n9562 ;
  assign n9564 = ~n876 & n9563 ;
  assign n9565 = n9564 ^ n3230 ^ 1'b0 ;
  assign n9566 = n687 & ~n9565 ;
  assign n9567 = n4455 & n9566 ;
  assign n9569 = n9568 ^ n9567 ^ 1'b0 ;
  assign n9570 = n3123 ^ n1616 ^ 1'b0 ;
  assign n9571 = n7399 | n9570 ;
  assign n9572 = n9525 ^ n2261 ^ 1'b0 ;
  assign n9573 = n6610 ^ n5735 ^ 1'b0 ;
  assign n9574 = n9573 ^ n1235 ^ 1'b0 ;
  assign n9575 = n3034 & n6338 ;
  assign n9576 = n4727 | n9445 ;
  assign n9577 = n420 & ~n922 ;
  assign n9578 = n6749 & n9577 ;
  assign n9579 = ~n356 & n9578 ;
  assign n9580 = ~n200 & n4472 ;
  assign n9581 = ~n4472 & n9580 ;
  assign n9582 = n5483 & n5562 ;
  assign n9583 = ~n5562 & n9582 ;
  assign n9584 = n9581 | n9583 ;
  assign n9585 = n9579 | n9584 ;
  assign n9586 = n1493 & ~n6932 ;
  assign n9587 = n2389 | n3537 ;
  assign n9588 = n9587 ^ n1393 ^ 1'b0 ;
  assign n9589 = n4723 & ~n9588 ;
  assign n9590 = n9589 ^ n5442 ^ 1'b0 ;
  assign n9591 = n266 & n4918 ;
  assign n9592 = ~n5519 & n9591 ;
  assign n9593 = n1012 | n3386 ;
  assign n9594 = n4334 | n9593 ;
  assign n9595 = n889 ^ n616 ^ 1'b0 ;
  assign n9596 = n6711 | n9595 ;
  assign n9599 = n636 | n3570 ;
  assign n9600 = n1025 & ~n9599 ;
  assign n9601 = n8767 & ~n9600 ;
  assign n9602 = ~n1064 & n9601 ;
  assign n9597 = n6239 ^ n5096 ^ 1'b0 ;
  assign n9598 = ~n4106 & n9597 ;
  assign n9603 = n9602 ^ n9598 ^ 1'b0 ;
  assign n9604 = n862 | n9603 ;
  assign n9605 = ~n285 & n3336 ;
  assign n9606 = n8289 & ~n9605 ;
  assign n9607 = n4657 & n7698 ;
  assign n9608 = n1387 & ~n9607 ;
  assign n9609 = ~n1341 & n8192 ;
  assign n9610 = n2496 & ~n2763 ;
  assign n9611 = n9610 ^ n330 ^ 1'b0 ;
  assign n9612 = ~n5025 & n9611 ;
  assign n9613 = x52 & ~n9103 ;
  assign n9614 = n9613 ^ n2067 ^ 1'b0 ;
  assign n9615 = n6583 ^ n725 ^ 1'b0 ;
  assign n9616 = n1122 ^ n831 ^ 1'b0 ;
  assign n9617 = n2159 | n9616 ;
  assign n9618 = ~n5966 & n7093 ;
  assign n9619 = ~n6203 & n6344 ;
  assign n9620 = ~x73 & n9619 ;
  assign n9621 = n3358 ^ n3101 ^ 1'b0 ;
  assign n9622 = ~n5249 & n9621 ;
  assign n9623 = ~n242 & n9622 ;
  assign n9624 = n3789 ^ n1542 ^ 1'b0 ;
  assign n9625 = n7476 ^ n2024 ^ 1'b0 ;
  assign n9626 = n9625 ^ n8985 ^ 1'b0 ;
  assign n9627 = n2729 ^ n1833 ^ 1'b0 ;
  assign n9628 = ~n3607 & n9627 ;
  assign n9629 = n6258 & ~n6847 ;
  assign n9630 = x108 & n4333 ;
  assign n9631 = n1146 & n7981 ;
  assign n9632 = n9631 ^ n1874 ^ 1'b0 ;
  assign n9633 = n1191 & ~n9632 ;
  assign n9634 = ~n4254 & n9633 ;
  assign n9635 = n1082 | n2785 ;
  assign n9636 = n1025 | n2722 ;
  assign n9637 = n516 | n8707 ;
  assign n9638 = n9636 | n9637 ;
  assign n9639 = n3415 & ~n9638 ;
  assign n9640 = n9635 & ~n9639 ;
  assign n9641 = n9634 | n9640 ;
  assign n9644 = ( n2974 & n4640 ) | ( n2974 & n9217 ) | ( n4640 & n9217 ) ;
  assign n9645 = n3765 & n9644 ;
  assign n9646 = ~n5904 & n9645 ;
  assign n9647 = n9646 ^ n4212 ^ 1'b0 ;
  assign n9642 = n3565 ^ n830 ^ 1'b0 ;
  assign n9643 = n6078 | n9642 ;
  assign n9648 = n9647 ^ n9643 ^ 1'b0 ;
  assign n9649 = ~n259 & n3144 ;
  assign n9650 = n9649 ^ n2827 ^ 1'b0 ;
  assign n9651 = n9650 ^ n2957 ^ 1'b0 ;
  assign n9652 = n9651 ^ n9302 ^ 1'b0 ;
  assign n9653 = x95 & n9652 ;
  assign n9654 = n1434 & n2099 ;
  assign n9655 = n8122 ^ n1020 ^ 1'b0 ;
  assign n9656 = n9654 & ~n9655 ;
  assign n9657 = n2423 & ~n9656 ;
  assign n9658 = n650 ^ n446 ^ 1'b0 ;
  assign n9659 = ~n4812 & n5090 ;
  assign n9660 = n9659 ^ n5989 ^ 1'b0 ;
  assign n9661 = n1457 ^ x57 ^ 1'b0 ;
  assign n9662 = ~n2168 & n9661 ;
  assign n9663 = n2911 | n7849 ;
  assign n9664 = n3687 & n4194 ;
  assign n9665 = ~n9663 & n9664 ;
  assign n9666 = n9662 & ~n9665 ;
  assign n9667 = n9666 ^ n5178 ^ 1'b0 ;
  assign n9668 = n1480 & ~n9667 ;
  assign n9669 = n7299 ^ n823 ^ 1'b0 ;
  assign n9670 = ~n1609 & n9669 ;
  assign n9671 = n6474 ^ x118 ^ 1'b0 ;
  assign n9672 = n1777 & ~n5638 ;
  assign n9673 = n3385 ^ n2491 ^ n1240 ;
  assign n9674 = n8725 ^ n8426 ^ 1'b0 ;
  assign n9675 = ~n9673 & n9674 ;
  assign n9676 = n5361 & ~n6590 ;
  assign n9677 = n3369 | n9492 ;
  assign n9678 = n328 | n640 ;
  assign n9679 = n2360 & ~n9678 ;
  assign n9680 = n2557 | n9679 ;
  assign n9681 = n7096 ^ n3925 ^ 1'b0 ;
  assign n9682 = n1226 ^ n604 ^ 1'b0 ;
  assign n9683 = n5962 & ~n9682 ;
  assign n9684 = n1057 & ~n4711 ;
  assign n9685 = n992 ^ n616 ^ 1'b0 ;
  assign n9686 = n4265 & ~n9685 ;
  assign n9687 = ~n1161 & n9686 ;
  assign n9688 = n7177 | n9687 ;
  assign n9689 = n3947 & ~n9688 ;
  assign n9690 = n8987 | n9689 ;
  assign n9691 = n165 & ~n6022 ;
  assign n9693 = ~n8191 & n9367 ;
  assign n9692 = n6907 ^ n2934 ^ 1'b0 ;
  assign n9694 = n9693 ^ n9692 ^ 1'b0 ;
  assign n9695 = n9691 & ~n9694 ;
  assign n9696 = ~n177 & n1139 ;
  assign n9697 = n1980 & ~n9696 ;
  assign n9698 = n1082 & ~n2325 ;
  assign n9699 = ~n5430 & n9698 ;
  assign n9700 = ~n6118 & n9699 ;
  assign n9701 = n704 | n3664 ;
  assign n9702 = n9701 ^ n2145 ^ 1'b0 ;
  assign n9703 = n9702 ^ n8581 ^ 1'b0 ;
  assign n9704 = n9700 | n9703 ;
  assign n9705 = n928 & n3911 ;
  assign n9706 = n8888 & n9705 ;
  assign n9707 = n4363 ^ n538 ^ 1'b0 ;
  assign n9708 = n446 | n9707 ;
  assign n9709 = n3813 & n5400 ;
  assign n9710 = ~n837 & n1645 ;
  assign n9711 = n9069 ^ n809 ^ 1'b0 ;
  assign n9712 = n926 | n4013 ;
  assign n9713 = n2237 | n6077 ;
  assign n9714 = n3150 & ~n9713 ;
  assign n9715 = ~n9712 & n9714 ;
  assign n9716 = n3874 | n9715 ;
  assign n9717 = n5941 ^ n5661 ^ n1444 ;
  assign n9718 = n8536 | n9250 ;
  assign n9719 = n5035 | n7421 ;
  assign n9721 = ~n1664 & n2647 ;
  assign n9722 = n9721 ^ n662 ^ 1'b0 ;
  assign n9723 = n6401 & n9722 ;
  assign n9724 = n8278 & n9723 ;
  assign n9720 = n5378 & ~n6908 ;
  assign n9725 = n9724 ^ n9720 ^ 1'b0 ;
  assign n9726 = n926 & n1751 ;
  assign n9727 = n1947 ^ n1355 ^ 1'b0 ;
  assign n9728 = n9726 & ~n9727 ;
  assign n9729 = n9728 ^ n669 ^ 1'b0 ;
  assign n9730 = n9729 ^ n6432 ^ 1'b0 ;
  assign n9731 = n3994 ^ n2361 ^ 1'b0 ;
  assign n9732 = ~n9730 & n9731 ;
  assign n9733 = n1901 ^ n430 ^ 1'b0 ;
  assign n9734 = ~n1636 & n9733 ;
  assign n9735 = x66 & n9734 ;
  assign n9736 = ~n2667 & n9735 ;
  assign n9737 = n8179 & ~n8791 ;
  assign n9738 = x54 & n7508 ;
  assign n9739 = n5637 & n9738 ;
  assign n9740 = ~n737 & n1920 ;
  assign n9741 = n9740 ^ n7020 ^ 1'b0 ;
  assign n9742 = n2481 & ~n7155 ;
  assign n9743 = n9742 ^ n2806 ^ 1'b0 ;
  assign n9744 = ( n9739 & ~n9741 ) | ( n9739 & n9743 ) | ( ~n9741 & n9743 ) ;
  assign n9745 = n8963 & n9744 ;
  assign n9746 = n8409 ^ n4089 ^ 1'b0 ;
  assign n9747 = n1541 ^ n552 ^ 1'b0 ;
  assign n9748 = ~n6301 & n9747 ;
  assign n9749 = n9748 ^ n590 ^ n297 ;
  assign n9750 = n5038 | n9588 ;
  assign n9751 = n9750 ^ n5227 ^ 1'b0 ;
  assign n9752 = n8456 ^ n4625 ^ 1'b0 ;
  assign n9753 = n183 & ~n9752 ;
  assign n9759 = n3947 | n5183 ;
  assign n9760 = x12 & ~n9759 ;
  assign n9754 = n5888 | n7718 ;
  assign n9755 = n2453 & ~n9754 ;
  assign n9756 = n2689 | n9755 ;
  assign n9757 = n1329 & n1539 ;
  assign n9758 = n9756 & n9757 ;
  assign n9761 = n9760 ^ n9758 ^ 1'b0 ;
  assign n9762 = n1306 & ~n5033 ;
  assign n9763 = n1895 & n9762 ;
  assign n9764 = ( x83 & n2704 ) | ( x83 & ~n9763 ) | ( n2704 & ~n9763 ) ;
  assign n9765 = n9764 ^ n8282 ^ n4107 ;
  assign n9766 = n1616 | n9765 ;
  assign n9774 = ~n482 & n972 ;
  assign n9770 = n2653 ^ n2279 ^ 1'b0 ;
  assign n9771 = n394 & ~n9770 ;
  assign n9772 = n8948 ^ n5202 ^ 1'b0 ;
  assign n9773 = n9771 & ~n9772 ;
  assign n9767 = ~n1314 & n4761 ;
  assign n9768 = n9767 ^ n6550 ^ 1'b0 ;
  assign n9769 = n2934 & ~n9768 ;
  assign n9775 = n9774 ^ n9773 ^ n9769 ;
  assign n9776 = n6730 ^ n4806 ^ 1'b0 ;
  assign n9777 = ~n8153 & n9776 ;
  assign n9778 = ~n425 & n6034 ;
  assign n9779 = ~n6328 & n9778 ;
  assign n9780 = n2687 | n4908 ;
  assign n9781 = n9016 & n9780 ;
  assign n9782 = n834 & n9781 ;
  assign n9784 = n3319 ^ n262 ^ 1'b0 ;
  assign n9783 = ~n3544 & n3634 ;
  assign n9785 = n9784 ^ n9783 ^ 1'b0 ;
  assign n9786 = n2800 ^ n1393 ^ 1'b0 ;
  assign n9787 = n1360 & n3554 ;
  assign n9788 = n9787 ^ n1170 ^ 1'b0 ;
  assign n9789 = n9786 & ~n9788 ;
  assign n9794 = n1919 & ~n6817 ;
  assign n9790 = n1491 ^ n566 ^ 1'b0 ;
  assign n9791 = n230 | n9790 ;
  assign n9792 = n9791 ^ n2518 ^ 1'b0 ;
  assign n9793 = n9792 ^ n5388 ^ n3037 ;
  assign n9795 = n9794 ^ n9793 ^ 1'b0 ;
  assign n9796 = n1070 & n3144 ;
  assign n9797 = n9796 ^ n2186 ^ 1'b0 ;
  assign n9798 = n9797 ^ n4267 ^ 1'b0 ;
  assign n9799 = n1846 & ~n7285 ;
  assign n9800 = n7360 ^ n2198 ^ 1'b0 ;
  assign n9803 = n1714 & ~n2776 ;
  assign n9801 = ~n250 & n1645 ;
  assign n9802 = ~n4825 & n9801 ;
  assign n9804 = n9803 ^ n9802 ^ 1'b0 ;
  assign n9805 = n9804 ^ n9287 ^ 1'b0 ;
  assign n9806 = n5560 | n9250 ;
  assign n9807 = ~n575 & n1178 ;
  assign n9808 = ~n8224 & n9807 ;
  assign n9809 = n1616 & n2070 ;
  assign n9810 = n9809 ^ n6099 ^ 1'b0 ;
  assign n9811 = n8203 | n9810 ;
  assign n9815 = ~n6282 & n6311 ;
  assign n9812 = n6565 ^ n749 ^ 1'b0 ;
  assign n9813 = x70 & n9812 ;
  assign n9814 = ~n2981 & n9813 ;
  assign n9816 = n9815 ^ n9814 ^ 1'b0 ;
  assign n9817 = x22 & ~n3240 ;
  assign n9818 = n3204 & n9817 ;
  assign n9819 = n9818 ^ n2386 ^ 1'b0 ;
  assign n9820 = n4482 | n9819 ;
  assign n9821 = n9820 ^ n1469 ^ 1'b0 ;
  assign n9822 = n2604 & ~n9821 ;
  assign n9823 = n1491 | n4844 ;
  assign n9824 = x94 & ~n4557 ;
  assign n9825 = n9824 ^ n5878 ^ 1'b0 ;
  assign n9826 = n2583 & n9825 ;
  assign n9827 = n8576 ^ x9 ^ 1'b0 ;
  assign n9828 = n3504 & n4112 ;
  assign n9830 = n1249 & n5617 ;
  assign n9829 = ~n2132 & n6247 ;
  assign n9831 = n9830 ^ n9829 ^ 1'b0 ;
  assign n9832 = n2887 & n6640 ;
  assign n9833 = ~n6360 & n9832 ;
  assign n9834 = n806 | n2730 ;
  assign n9835 = n1026 | n9834 ;
  assign n9836 = ~n4954 & n9835 ;
  assign n9837 = n8030 & ~n9197 ;
  assign n9838 = n9837 ^ n866 ^ 1'b0 ;
  assign n9839 = n3596 & n3897 ;
  assign n9840 = n6512 ^ n5727 ^ 1'b0 ;
  assign n9842 = n8760 ^ n4048 ^ 1'b0 ;
  assign n9843 = n5666 & ~n9842 ;
  assign n9841 = ~n4204 & n4916 ;
  assign n9844 = n9843 ^ n9841 ^ 1'b0 ;
  assign n9845 = n5596 & ~n9844 ;
  assign n9846 = n4910 ^ n1664 ^ 1'b0 ;
  assign n9847 = n141 & ~n2177 ;
  assign n9848 = n9847 ^ x61 ^ 1'b0 ;
  assign n9849 = ~n6419 & n7900 ;
  assign n9850 = n9849 ^ n7047 ^ 1'b0 ;
  assign n9851 = n1067 ^ n276 ^ 1'b0 ;
  assign n9852 = n9683 & n9835 ;
  assign n9853 = n1838 ^ n1795 ^ 1'b0 ;
  assign n9854 = n6445 ^ n5746 ^ n2906 ;
  assign n9855 = n9431 ^ n7241 ^ 1'b0 ;
  assign n9856 = n9815 & n9855 ;
  assign n9857 = n3066 | n6034 ;
  assign n9858 = n1685 | n9857 ;
  assign n9859 = n9858 ^ n7078 ^ 1'b0 ;
  assign n9860 = n1898 & ~n6461 ;
  assign n9861 = n6038 & n6112 ;
  assign n9862 = n9861 ^ n3675 ^ 1'b0 ;
  assign n9863 = ( n2978 & ~n9860 ) | ( n2978 & n9862 ) | ( ~n9860 & n9862 ) ;
  assign n9864 = n2710 ^ n954 ^ n338 ;
  assign n9865 = n9864 ^ n4443 ^ 1'b0 ;
  assign n9866 = n4847 & n6694 ;
  assign n9867 = ~n1153 & n5003 ;
  assign n9868 = n3472 ^ n790 ^ 1'b0 ;
  assign n9869 = n9868 ^ n4371 ^ 1'b0 ;
  assign n9870 = n8526 ^ n2392 ^ 1'b0 ;
  assign n9871 = ~n8450 & n9524 ;
  assign n9872 = n9871 ^ n806 ^ 1'b0 ;
  assign n9873 = n7190 & n9872 ;
  assign n9874 = ~n1635 & n9873 ;
  assign n9875 = n5006 ^ n2875 ^ 1'b0 ;
  assign n9876 = n5548 & n9875 ;
  assign n9877 = n3062 | n9876 ;
  assign n9878 = n6434 & n6727 ;
  assign n9879 = ~n725 & n9878 ;
  assign n9880 = n9879 ^ n4129 ^ 1'b0 ;
  assign n9881 = n508 | n9880 ;
  assign n9882 = n2153 | n9881 ;
  assign n9883 = n9882 ^ n4847 ^ 1'b0 ;
  assign n9884 = n9883 ^ n2815 ^ 1'b0 ;
  assign n9885 = n741 | n9884 ;
  assign n9886 = n1959 | n9885 ;
  assign n9887 = n7471 & ~n9886 ;
  assign n9888 = n5430 | n6874 ;
  assign n9889 = n1914 & ~n9888 ;
  assign n9890 = n2165 | n9818 ;
  assign n9891 = n9889 & ~n9890 ;
  assign n9892 = ~n328 & n9159 ;
  assign n9893 = n7668 ^ n5950 ^ 1'b0 ;
  assign n9894 = n9893 ^ n8016 ^ 1'b0 ;
  assign n9895 = n3537 ^ x124 ^ 1'b0 ;
  assign n9896 = n3509 ^ n2414 ^ 1'b0 ;
  assign n9897 = n1751 & n2749 ;
  assign n9898 = n548 | n630 ;
  assign n9899 = x49 | n9898 ;
  assign n9900 = n763 & n9899 ;
  assign n9901 = n1277 & n9900 ;
  assign n9902 = n2344 ^ n648 ^ 1'b0 ;
  assign n9903 = n9902 ^ n3422 ^ 1'b0 ;
  assign n9904 = n3862 & ~n7798 ;
  assign n9905 = n2804 & ~n9904 ;
  assign n9906 = n2423 & n9905 ;
  assign n9907 = n547 & n5898 ;
  assign n9908 = n4902 & n9907 ;
  assign n9909 = n1685 & ~n3019 ;
  assign n9910 = n5907 & n9909 ;
  assign n9911 = n9908 | n9910 ;
  assign n9912 = ~n3422 & n5061 ;
  assign n9913 = n9912 ^ n2186 ^ 1'b0 ;
  assign n9914 = n9913 ^ n8309 ^ 1'b0 ;
  assign n9915 = ~n6875 & n8229 ;
  assign n9916 = n6467 ^ n408 ^ x52 ;
  assign n9917 = n6310 ^ n5438 ^ 1'b0 ;
  assign n9918 = n3760 & ~n9917 ;
  assign n9919 = n2366 & n9918 ;
  assign n9920 = n3642 ^ n814 ^ 1'b0 ;
  assign n9921 = n2331 | n9920 ;
  assign n9922 = n3994 & ~n5086 ;
  assign n9923 = n9921 & n9922 ;
  assign n9924 = n8157 & n9923 ;
  assign n9925 = n1236 & n4082 ;
  assign n9926 = ~n3646 & n9925 ;
  assign n9927 = n7731 & n8531 ;
  assign n9928 = n9926 & n9927 ;
  assign n9929 = n3809 ^ n1984 ^ 1'b0 ;
  assign n9930 = ~n1734 & n1827 ;
  assign n9931 = n9929 & n9930 ;
  assign n9932 = n2623 | n9931 ;
  assign n9933 = n2623 & ~n9932 ;
  assign n9934 = n839 | n8614 ;
  assign n9935 = n5211 & ~n9934 ;
  assign n9936 = ~n5211 & n9935 ;
  assign n9937 = n5940 | n9936 ;
  assign n9938 = n9933 & ~n9937 ;
  assign n9939 = n4107 | n6626 ;
  assign n9940 = n9939 ^ n5410 ^ 1'b0 ;
  assign n9944 = ~n3699 & n6549 ;
  assign n9945 = n4565 & n9944 ;
  assign n9941 = n5136 ^ n2979 ^ 1'b0 ;
  assign n9942 = n1321 & ~n9941 ;
  assign n9943 = n2592 & n9942 ;
  assign n9946 = n9945 ^ n9943 ^ 1'b0 ;
  assign n9947 = n5067 ^ n4619 ^ n3662 ;
  assign n9948 = n3417 ^ n1216 ^ 1'b0 ;
  assign n9949 = n9948 ^ n1530 ^ 1'b0 ;
  assign n9950 = n1001 & n9949 ;
  assign n9951 = n9247 & n9950 ;
  assign n9952 = n9951 ^ n520 ^ 1'b0 ;
  assign n9953 = n634 & n788 ;
  assign n9954 = ~n822 & n9953 ;
  assign n9955 = n243 | n9539 ;
  assign n9956 = n2664 & n9955 ;
  assign n9957 = ~n2478 & n9956 ;
  assign n9958 = n9957 ^ n2776 ^ 1'b0 ;
  assign n9959 = n8514 & n9958 ;
  assign n9960 = ~n681 & n4129 ;
  assign n9961 = n9960 ^ n7114 ^ 1'b0 ;
  assign n9962 = n3354 & n5143 ;
  assign n9963 = ~n1423 & n4230 ;
  assign n9964 = n9963 ^ n2919 ^ 1'b0 ;
  assign n9965 = n2122 & ~n9964 ;
  assign n9966 = n9964 & n9965 ;
  assign n9967 = x71 & n1129 ;
  assign n9968 = n9967 ^ n9413 ^ 1'b0 ;
  assign n9969 = n428 | n9968 ;
  assign n9970 = n9966 & ~n9969 ;
  assign n9971 = n899 | n1925 ;
  assign n9972 = n1925 & ~n9971 ;
  assign n9973 = x45 & n5496 ;
  assign n9974 = n3249 & n9973 ;
  assign n9975 = ~n1222 & n9974 ;
  assign n9976 = n7418 | n9975 ;
  assign n9977 = n7418 & ~n9976 ;
  assign n9978 = n9972 | n9977 ;
  assign n9979 = n9970 | n9978 ;
  assign n9980 = n6353 ^ x52 ^ 1'b0 ;
  assign n9981 = n8269 | n9980 ;
  assign n9985 = ~n1176 & n4102 ;
  assign n9986 = n1781 & n9985 ;
  assign n9982 = n731 | n2165 ;
  assign n9983 = n5715 | n9982 ;
  assign n9984 = ~n1571 & n9983 ;
  assign n9987 = n9986 ^ n9984 ^ 1'b0 ;
  assign n9988 = ~n6727 & n9987 ;
  assign n9989 = n6780 ^ n2623 ^ 1'b0 ;
  assign n9990 = n9136 & n9989 ;
  assign n9991 = n811 & n1025 ;
  assign n9992 = n9991 ^ n185 ^ 1'b0 ;
  assign n9994 = n335 & ~n459 ;
  assign n9995 = n459 & n9994 ;
  assign n9993 = n7317 ^ n1203 ^ 1'b0 ;
  assign n9996 = n9995 ^ n9993 ^ 1'b0 ;
  assign n9997 = n3414 & ~n9996 ;
  assign n9999 = n1829 ^ n1569 ^ 1'b0 ;
  assign n10000 = ~n132 & n9999 ;
  assign n10001 = ~n1616 & n10000 ;
  assign n10002 = n7736 & n10001 ;
  assign n10003 = ( n1854 & n3245 ) | ( n1854 & n10002 ) | ( n3245 & n10002 ) ;
  assign n10004 = n3509 & ~n10003 ;
  assign n10005 = n10004 ^ n4998 ^ 1'b0 ;
  assign n9998 = n1319 | n3264 ;
  assign n10006 = n10005 ^ n9998 ^ n2896 ;
  assign n10007 = x93 & ~n1270 ;
  assign n10008 = n10007 ^ n5413 ^ n4832 ;
  assign n10009 = n3538 ^ n2418 ^ 1'b0 ;
  assign n10010 = n948 | n10009 ;
  assign n10011 = n10008 & n10010 ;
  assign n10013 = n2384 | n3844 ;
  assign n10014 = n2573 | n10013 ;
  assign n10012 = n9315 & ~n9679 ;
  assign n10015 = n10014 ^ n10012 ^ 1'b0 ;
  assign n10016 = n5528 ^ n2584 ^ 1'b0 ;
  assign n10017 = n1187 ^ n538 ^ 1'b0 ;
  assign n10018 = ~n717 & n10017 ;
  assign n10019 = ~n6286 & n10018 ;
  assign n10020 = n10019 ^ n9409 ^ 1'b0 ;
  assign n10021 = n6195 | n6335 ;
  assign n10022 = n2313 & n9244 ;
  assign n10023 = ~x119 & n5364 ;
  assign n10024 = n10023 ^ n2649 ^ 1'b0 ;
  assign n10025 = n3500 & n6325 ;
  assign n10026 = n1201 & n10025 ;
  assign n10027 = n2083 & ~n6114 ;
  assign n10028 = n5229 ^ n5223 ^ 1'b0 ;
  assign n10029 = ~n642 & n10028 ;
  assign n10030 = n5413 & n6921 ;
  assign n10031 = n10030 ^ x38 ^ 1'b0 ;
  assign n10032 = n1006 | n3075 ;
  assign n10033 = n2673 | n10032 ;
  assign n10034 = ~x4 & n10033 ;
  assign n10035 = n10034 ^ n1576 ^ 1'b0 ;
  assign n10036 = n10035 ^ n4602 ^ 1'b0 ;
  assign n10037 = n4882 & n10036 ;
  assign n10038 = ~n3153 & n3381 ;
  assign n10039 = n3153 & n10038 ;
  assign n10040 = n588 | n1177 ;
  assign n10041 = n10039 | n10040 ;
  assign n10042 = n10037 | n10041 ;
  assign n10043 = n857 & n6304 ;
  assign n10044 = ~n453 & n10043 ;
  assign n10045 = n10044 ^ n4310 ^ 1'b0 ;
  assign n10046 = n833 | n4806 ;
  assign n10047 = ~n946 & n2394 ;
  assign n10048 = n8952 ^ n6471 ^ 1'b0 ;
  assign n10049 = n1634 & ~n8206 ;
  assign n10050 = ~n3330 & n6522 ;
  assign n10051 = n10050 ^ n1541 ^ 1'b0 ;
  assign n10052 = ( n786 & n812 ) | ( n786 & ~n3010 ) | ( n812 & ~n3010 ) ;
  assign n10053 = n1057 & ~n10052 ;
  assign n10054 = n10053 ^ n1226 ^ n1063 ;
  assign n10055 = n1693 & n3697 ;
  assign n10056 = n3969 ^ n2395 ^ 1'b0 ;
  assign n10057 = n3789 | n10056 ;
  assign n10058 = n8635 & ~n10057 ;
  assign n10059 = n8215 ^ n4580 ^ 1'b0 ;
  assign n10060 = ~n4279 & n10059 ;
  assign n10061 = n192 & ~n5141 ;
  assign n10062 = n10061 ^ n9586 ^ 1'b0 ;
  assign n10063 = n10060 & n10062 ;
  assign n10064 = n3213 ^ n1783 ^ 1'b0 ;
  assign n10065 = n7139 | n10064 ;
  assign n10066 = n4232 & n8059 ;
  assign n10067 = n10066 ^ n2924 ^ 1'b0 ;
  assign n10068 = x106 | n10067 ;
  assign n10069 = n8705 ^ n330 ^ 1'b0 ;
  assign n10070 = x72 | n3667 ;
  assign n10071 = n4602 ^ x41 ^ 1'b0 ;
  assign n10072 = ~n10070 & n10071 ;
  assign n10073 = n7870 ^ n5445 ^ n819 ;
  assign n10074 = ~n5492 & n10073 ;
  assign n10075 = ~n516 & n962 ;
  assign n10076 = ~n8637 & n10075 ;
  assign n10077 = n5926 ^ n205 ^ 1'b0 ;
  assign n10078 = n5313 & n6621 ;
  assign n10079 = n7120 ^ n3716 ^ 1'b0 ;
  assign n10080 = ~n4842 & n8339 ;
  assign n10081 = n2436 ^ x125 ^ 1'b0 ;
  assign n10082 = n586 & n1095 ;
  assign n10083 = ~n9766 & n10082 ;
  assign n10084 = n1361 & n1534 ;
  assign n10085 = n1156 & ~n9285 ;
  assign n10086 = n10084 & ~n10085 ;
  assign n10087 = n7980 ^ n3082 ^ 1'b0 ;
  assign n10088 = n1167 & n10087 ;
  assign n10089 = ~n9534 & n10088 ;
  assign n10090 = n4490 ^ n475 ^ 1'b0 ;
  assign n10091 = n6195 & ~n10090 ;
  assign n10092 = n1974 & n3170 ;
  assign n10093 = ~n2376 & n10092 ;
  assign n10094 = ~n1110 & n10093 ;
  assign n10095 = n3680 & ~n10094 ;
  assign n10096 = n8982 ^ n2992 ^ 1'b0 ;
  assign n10097 = n9106 ^ n4289 ^ 1'b0 ;
  assign n10098 = n1103 & ~n10097 ;
  assign n10099 = n8223 ^ n1714 ^ 1'b0 ;
  assign n10116 = ~n6669 & n7239 ;
  assign n10117 = n6669 & n10116 ;
  assign n10100 = n407 & n4664 ;
  assign n10101 = ~n407 & n10100 ;
  assign n10102 = n809 | n1622 ;
  assign n10103 = n1622 & ~n10102 ;
  assign n10104 = n2010 & ~n5139 ;
  assign n10105 = n10103 & n10104 ;
  assign n10106 = n660 | n10105 ;
  assign n10107 = n10105 & ~n10106 ;
  assign n10110 = ~n741 & n984 ;
  assign n10111 = ~n984 & n10110 ;
  assign n10112 = x55 & n10111 ;
  assign n10108 = n846 & n8229 ;
  assign n10109 = ~n8229 & n10108 ;
  assign n10113 = n10112 ^ n10109 ^ 1'b0 ;
  assign n10114 = n10107 | n10113 ;
  assign n10115 = n10101 | n10114 ;
  assign n10118 = n10117 ^ n10115 ^ 1'b0 ;
  assign n10119 = ~n4553 & n8508 ;
  assign n10120 = n10119 ^ n407 ^ 1'b0 ;
  assign n10121 = n1699 ^ n545 ^ 1'b0 ;
  assign n10122 = n5611 ^ n2427 ^ 1'b0 ;
  assign n10123 = ~n1827 & n10122 ;
  assign n10124 = ~n6736 & n8804 ;
  assign n10125 = ~n10123 & n10124 ;
  assign n10126 = n7712 | n8764 ;
  assign n10127 = n5196 | n7369 ;
  assign n10128 = n921 & ~n10127 ;
  assign n10129 = n7736 & n7802 ;
  assign n10130 = n1741 ^ n1192 ^ 1'b0 ;
  assign n10131 = n1909 & n10130 ;
  assign n10132 = ~n10129 & n10131 ;
  assign n10133 = n1191 & n5367 ;
  assign n10134 = n245 & n10133 ;
  assign n10135 = ~n5302 & n8039 ;
  assign n10136 = n10135 ^ n8848 ^ 1'b0 ;
  assign n10137 = ~n3695 & n5887 ;
  assign n10138 = n9679 | n10137 ;
  assign n10139 = n2291 & ~n10138 ;
  assign n10140 = n2385 & n3272 ;
  assign n10141 = ~n2925 & n10140 ;
  assign n10142 = n2307 & n3369 ;
  assign n10143 = n9684 ^ n409 ^ 1'b0 ;
  assign n10144 = ~n3072 & n10143 ;
  assign n10145 = n8385 ^ n7210 ^ 1'b0 ;
  assign n10146 = ~n5804 & n10145 ;
  assign n10147 = n10146 ^ n7114 ^ 1'b0 ;
  assign n10148 = ~n5622 & n10147 ;
  assign n10149 = n10148 ^ n8900 ^ 1'b0 ;
  assign n10150 = n6536 | n9386 ;
  assign n10151 = n3064 | n10150 ;
  assign n10152 = x64 & n3973 ;
  assign n10153 = n722 & ~n10152 ;
  assign n10154 = n3753 & n9644 ;
  assign n10155 = ~n6835 & n10154 ;
  assign n10156 = n10155 ^ n4341 ^ 1'b0 ;
  assign n10157 = n1226 & n7614 ;
  assign n10158 = n6061 ^ n4007 ^ 1'b0 ;
  assign n10159 = n8217 | n8791 ;
  assign n10160 = n10159 ^ n4666 ^ 1'b0 ;
  assign n10161 = n2109 & ~n7041 ;
  assign n10162 = n7590 & n10161 ;
  assign n10163 = n4662 & ~n8117 ;
  assign n10164 = ~n10162 & n10163 ;
  assign n10165 = n9859 & n10164 ;
  assign n10166 = n553 & n8933 ;
  assign n10167 = n3919 ^ n315 ^ 1'b0 ;
  assign n10168 = n4639 | n10167 ;
  assign n10169 = n4551 ^ n4056 ^ 1'b0 ;
  assign n10170 = n10168 | n10169 ;
  assign n10171 = ~n6037 & n6283 ;
  assign n10172 = n10171 ^ n1393 ^ 1'b0 ;
  assign n10173 = n2232 | n9646 ;
  assign n10174 = x49 & ~n7594 ;
  assign n10175 = n10174 ^ n262 ^ 1'b0 ;
  assign n10176 = n10175 ^ n5369 ^ 1'b0 ;
  assign n10177 = n10173 & ~n10176 ;
  assign n10178 = n8205 ^ n2074 ^ 1'b0 ;
  assign n10179 = n3030 ^ n2226 ^ 1'b0 ;
  assign n10181 = n2392 | n3760 ;
  assign n10180 = n4354 & n5801 ;
  assign n10182 = n10181 ^ n10180 ^ 1'b0 ;
  assign n10183 = ~n5458 & n10182 ;
  assign n10184 = n3812 ^ n3632 ^ 1'b0 ;
  assign n10186 = n3126 ^ n2878 ^ 1'b0 ;
  assign n10185 = ~n446 & n10014 ;
  assign n10187 = n10186 ^ n10185 ^ 1'b0 ;
  assign n10188 = n9190 ^ n9006 ^ 1'b0 ;
  assign n10189 = ~n7624 & n10188 ;
  assign n10190 = ~n2446 & n9795 ;
  assign n10191 = n2313 & n4282 ;
  assign n10192 = n2732 ^ n1723 ^ 1'b0 ;
  assign n10193 = n1135 | n2079 ;
  assign n10194 = n10193 ^ n2833 ^ 1'b0 ;
  assign n10195 = n4037 | n10194 ;
  assign n10196 = n4438 ^ n1602 ^ 1'b0 ;
  assign n10197 = n10196 ^ n3097 ^ 1'b0 ;
  assign n10198 = ~n2771 & n5242 ;
  assign n10199 = n10198 ^ n4461 ^ 1'b0 ;
  assign n10200 = n8093 ^ n3298 ^ 1'b0 ;
  assign n10201 = n3049 & ~n10200 ;
  assign n10202 = ~n4404 & n10201 ;
  assign n10203 = n10202 ^ n358 ^ 1'b0 ;
  assign n10204 = n2155 & ~n2677 ;
  assign n10205 = n227 & n10204 ;
  assign n10206 = n4267 & ~n10205 ;
  assign n10207 = n10206 ^ n6965 ^ 1'b0 ;
  assign n10208 = ~n2923 & n10207 ;
  assign n10209 = ~n195 & n10208 ;
  assign n10210 = n10209 ^ n5885 ^ 1'b0 ;
  assign n10211 = n2749 & n10210 ;
  assign n10212 = n10211 ^ n5679 ^ 1'b0 ;
  assign n10213 = n806 | n8917 ;
  assign n10214 = n2376 ^ n717 ^ 1'b0 ;
  assign n10215 = n8052 | n10214 ;
  assign n10216 = ~n277 & n10215 ;
  assign n10217 = n9736 ^ n6987 ^ n450 ;
  assign n10219 = ~n4014 & n4230 ;
  assign n10220 = n4404 & n10219 ;
  assign n10221 = n8055 | n10220 ;
  assign n10222 = n9218 | n10221 ;
  assign n10218 = ~n3466 & n6266 ;
  assign n10223 = n10222 ^ n10218 ^ 1'b0 ;
  assign n10224 = ~n2204 & n3049 ;
  assign n10225 = n10223 & n10224 ;
  assign n10226 = n3651 & ~n8263 ;
  assign n10227 = n6677 & n10226 ;
  assign n10228 = n9883 ^ n3049 ^ 1'b0 ;
  assign n10229 = n6687 ^ n3401 ^ 1'b0 ;
  assign n10230 = n10228 & n10229 ;
  assign n10231 = n825 & ~n6523 ;
  assign n10232 = n6353 ^ n547 ^ 1'b0 ;
  assign n10233 = n5485 & ~n10232 ;
  assign n10234 = n5695 ^ n185 ^ 1'b0 ;
  assign n10235 = n3746 & ~n10234 ;
  assign n10236 = n10235 ^ n9494 ^ 1'b0 ;
  assign n10237 = n10233 & ~n10236 ;
  assign n10240 = x127 | n1691 ;
  assign n10238 = x11 & ~n7821 ;
  assign n10239 = n4643 & ~n10238 ;
  assign n10241 = n10240 ^ n10239 ^ 1'b0 ;
  assign n10242 = n5852 ^ n5258 ^ 1'b0 ;
  assign n10243 = n2508 & n7898 ;
  assign n10244 = n595 & n6590 ;
  assign n10245 = ~n3673 & n10244 ;
  assign n10246 = ~n5534 & n6085 ;
  assign n10247 = ~n2396 & n10246 ;
  assign n10248 = n3012 | n3165 ;
  assign n10249 = ~n6735 & n10248 ;
  assign n10250 = n10249 ^ n7610 ^ 1'b0 ;
  assign n10251 = ~n161 & n745 ;
  assign n10252 = n161 & n10251 ;
  assign n10253 = ~n560 & n10252 ;
  assign n10254 = ~n2224 & n10253 ;
  assign n10255 = n10254 ^ n7959 ^ 1'b0 ;
  assign n10256 = n7127 ^ n6104 ^ 1'b0 ;
  assign n10257 = n5470 & ~n10256 ;
  assign n10258 = n5150 & ~n7426 ;
  assign n10259 = ~n766 & n10258 ;
  assign n10260 = n10027 | n10259 ;
  assign n10261 = n7449 | n10260 ;
  assign n10262 = n6439 ^ n6296 ^ 1'b0 ;
  assign n10263 = n2245 ^ n1786 ^ 1'b0 ;
  assign n10264 = n1483 | n10263 ;
  assign n10265 = n1012 | n10264 ;
  assign n10266 = n6873 | n8286 ;
  assign n10267 = ~n1979 & n6825 ;
  assign n10268 = n6114 & n10267 ;
  assign n10269 = n3280 ^ n749 ^ x70 ;
  assign n10270 = n1975 | n5265 ;
  assign n10271 = n5265 & ~n10270 ;
  assign n10272 = n4486 ^ n325 ^ 1'b0 ;
  assign n10273 = n3518 & n10272 ;
  assign n10274 = ~n7424 & n10273 ;
  assign n10275 = ~n10273 & n10274 ;
  assign n10276 = n10271 | n10275 ;
  assign n10277 = n10269 & ~n10276 ;
  assign n10278 = ~n1107 & n4632 ;
  assign n10279 = n2598 | n8800 ;
  assign n10280 = n10279 ^ n1470 ^ 1'b0 ;
  assign n10281 = n10280 ^ n9084 ^ 1'b0 ;
  assign n10282 = n1527 | n4882 ;
  assign n10283 = n2575 | n3428 ;
  assign n10284 = n6208 & n9143 ;
  assign n10285 = n3403 & ~n6333 ;
  assign n10286 = n3087 & ~n8580 ;
  assign n10287 = ~n1828 & n10286 ;
  assign n10288 = n984 ^ n904 ^ 1'b0 ;
  assign n10289 = x40 | n10288 ;
  assign n10290 = n10289 ^ n6258 ^ 1'b0 ;
  assign n10291 = ~n851 & n10290 ;
  assign n10292 = ~n7747 & n10291 ;
  assign n10293 = n2198 & n2938 ;
  assign n10294 = n424 & ~n4926 ;
  assign n10295 = n3128 & n10294 ;
  assign n10296 = n5664 | n5720 ;
  assign n10297 = ~n4169 & n7977 ;
  assign n10298 = n6494 & ~n9700 ;
  assign n10299 = n10298 ^ n6260 ^ 1'b0 ;
  assign n10300 = ~n5392 & n10299 ;
  assign n10301 = ~n595 & n10300 ;
  assign n10302 = n6497 ^ n3177 ^ 1'b0 ;
  assign n10303 = n835 ^ n528 ^ 1'b0 ;
  assign n10304 = n5685 & ~n7339 ;
  assign n10305 = n5039 ^ n3027 ^ 1'b0 ;
  assign n10306 = x77 ^ x50 ^ 1'b0 ;
  assign n10307 = ~n2002 & n10306 ;
  assign n10308 = n10307 ^ n3283 ^ 1'b0 ;
  assign n10309 = n7023 ^ n330 ^ 1'b0 ;
  assign n10310 = n512 & n10309 ;
  assign n10311 = ~n5090 & n10310 ;
  assign n10312 = n1290 ^ n504 ^ 1'b0 ;
  assign n10313 = n10312 ^ n510 ^ 1'b0 ;
  assign n10314 = ~n510 & n10313 ;
  assign n10315 = n5595 & ~n10314 ;
  assign n10316 = n2718 & n5418 ;
  assign n10317 = n10316 ^ n2236 ^ 1'b0 ;
  assign n10318 = n10317 ^ n6215 ^ 1'b0 ;
  assign n10319 = ~n9429 & n10230 ;
  assign n10320 = n3079 & n6425 ;
  assign n10321 = n10320 ^ n8007 ^ 1'b0 ;
  assign n10322 = n7349 ^ n7210 ^ 1'b0 ;
  assign n10323 = ~n10321 & n10322 ;
  assign n10324 = n9034 ^ n3027 ^ 1'b0 ;
  assign n10325 = ~n3267 & n8742 ;
  assign n10326 = x7 & n10325 ;
  assign n10327 = n5189 | n10326 ;
  assign n10328 = n10327 ^ n1399 ^ 1'b0 ;
  assign n10329 = n3762 | n9868 ;
  assign n10330 = n811 & ~n10329 ;
  assign n10331 = n10314 & n10330 ;
  assign n10332 = n1816 ^ n1776 ^ 1'b0 ;
  assign n10333 = ~n5603 & n10332 ;
  assign n10334 = n2933 | n10333 ;
  assign n10335 = n10334 ^ n1161 ^ 1'b0 ;
  assign n10336 = n5137 & ~n10335 ;
  assign n10341 = n3819 ^ n1919 ^ 1'b0 ;
  assign n10337 = n3158 ^ n564 ^ 1'b0 ;
  assign n10338 = n4875 & ~n10337 ;
  assign n10339 = n3622 ^ n1998 ^ 1'b0 ;
  assign n10340 = n10338 & ~n10339 ;
  assign n10342 = n10341 ^ n10340 ^ 1'b0 ;
  assign n10343 = ~n1714 & n10342 ;
  assign n10346 = n2255 | n4908 ;
  assign n10347 = n2255 & ~n10346 ;
  assign n10348 = n3120 | n10347 ;
  assign n10349 = n3120 & ~n10348 ;
  assign n10344 = n5008 & n7802 ;
  assign n10345 = n8810 & ~n10344 ;
  assign n10350 = n10349 ^ n10345 ^ 1'b0 ;
  assign n10351 = n502 | n3944 ;
  assign n10352 = n2785 & n10351 ;
  assign n10353 = n10352 ^ n3367 ^ 1'b0 ;
  assign n10354 = n2068 & ~n10353 ;
  assign n10355 = n7709 ^ n7423 ^ 1'b0 ;
  assign n10356 = n7763 | n10355 ;
  assign n10357 = n1728 & n3383 ;
  assign n10358 = n1749 & n7362 ;
  assign n10359 = n7194 | n10358 ;
  assign n10360 = ~n503 & n5243 ;
  assign n10361 = n3739 & n10360 ;
  assign n10362 = n4350 ^ n911 ^ 1'b0 ;
  assign n10363 = n5861 & ~n10362 ;
  assign n10364 = n3140 ^ n1628 ^ 1'b0 ;
  assign n10365 = n7427 | n10364 ;
  assign n10366 = n10365 ^ n3296 ^ 1'b0 ;
  assign n10367 = n10363 & n10366 ;
  assign n10371 = ~n2608 & n8093 ;
  assign n10372 = ~n8093 & n10371 ;
  assign n10368 = n1201 | n2905 ;
  assign n10369 = n2905 & ~n10368 ;
  assign n10370 = n4819 & ~n10369 ;
  assign n10373 = n10372 ^ n10370 ^ 1'b0 ;
  assign n10374 = ~n1089 & n10373 ;
  assign n10375 = ~n10373 & n10374 ;
  assign n10376 = n7253 ^ n304 ^ 1'b0 ;
  assign n10377 = n9159 & ~n10376 ;
  assign n10378 = x22 | n2243 ;
  assign n10379 = n516 ^ x77 ^ 1'b0 ;
  assign n10380 = n7128 & n10379 ;
  assign n10381 = n10380 ^ n9588 ^ 1'b0 ;
  assign n10382 = n1744 & n9641 ;
  assign n10386 = n5038 ^ n716 ^ 1'b0 ;
  assign n10383 = n8494 ^ n3655 ^ n768 ;
  assign n10384 = n507 | n10383 ;
  assign n10385 = n10384 ^ n8571 ^ 1'b0 ;
  assign n10387 = n10386 ^ n10385 ^ 1'b0 ;
  assign n10388 = x59 | n4597 ;
  assign n10389 = n10388 ^ n6434 ^ n2461 ;
  assign n10390 = n3503 & n10389 ;
  assign n10391 = n10390 ^ n7942 ^ 1'b0 ;
  assign n10392 = n10391 ^ n134 ^ 1'b0 ;
  assign n10395 = n5705 ^ n4148 ^ n2959 ;
  assign n10396 = n6877 ^ x7 ^ 1'b0 ;
  assign n10397 = n10395 | n10396 ;
  assign n10393 = n9707 ^ n2537 ^ 1'b0 ;
  assign n10394 = n7460 | n10393 ;
  assign n10398 = n10397 ^ n10394 ^ 1'b0 ;
  assign n10399 = n2012 ^ n571 ^ 1'b0 ;
  assign n10400 = n7739 | n10399 ;
  assign n10401 = n2761 | n8689 ;
  assign n10402 = n5550 & n10401 ;
  assign n10403 = n707 & n1658 ;
  assign n10404 = n10403 ^ n2434 ^ 1'b0 ;
  assign n10405 = ~n10402 & n10404 ;
  assign n10406 = n3763 & n4202 ;
  assign n10407 = n10406 ^ n1497 ^ 1'b0 ;
  assign n10408 = n7727 & ~n10407 ;
  assign n10410 = n2569 & n2850 ;
  assign n10409 = n6747 & n10011 ;
  assign n10411 = n10410 ^ n10409 ^ 1'b0 ;
  assign n10412 = n5489 & ~n7688 ;
  assign n10413 = ~n2980 & n3149 ;
  assign n10414 = n3805 & n10413 ;
  assign n10415 = ~n1685 & n4224 ;
  assign n10416 = n10415 ^ n5019 ^ 1'b0 ;
  assign n10417 = n7672 & ~n10416 ;
  assign n10418 = n3934 | n6417 ;
  assign n10419 = n9305 & ~n10418 ;
  assign n10420 = n1498 | n6096 ;
  assign n10421 = n3014 & ~n3380 ;
  assign n10422 = n2002 & n10421 ;
  assign n10423 = ( n4173 & ~n4388 ) | ( n4173 & n5974 ) | ( ~n4388 & n5974 ) ;
  assign n10424 = n1711 & ~n10285 ;
  assign n10425 = n990 | n3090 ;
  assign n10426 = n2376 | n2732 ;
  assign n10427 = n10426 ^ n7971 ^ 1'b0 ;
  assign n10428 = n10425 & n10427 ;
  assign n10429 = n7898 & n10428 ;
  assign n10430 = n10077 ^ n4419 ^ 1'b0 ;
  assign n10431 = n7395 & ~n10430 ;
  assign n10432 = n8921 ^ n2839 ^ 1'b0 ;
  assign n10433 = ~n2827 & n7355 ;
  assign n10434 = ~n1756 & n10433 ;
  assign n10435 = n7574 & n10434 ;
  assign n10436 = n918 | n2227 ;
  assign n10437 = n6675 | n7365 ;
  assign n10438 = n1115 & ~n10437 ;
  assign n10439 = n153 & n7017 ;
  assign n10440 = ~n305 & n610 ;
  assign n10441 = n10439 | n10440 ;
  assign n10442 = n996 & ~n3149 ;
  assign n10443 = ~n475 & n795 ;
  assign n10444 = n1031 ^ x74 ^ 1'b0 ;
  assign n10445 = n10443 & ~n10444 ;
  assign n10446 = n10445 ^ n9081 ^ 1'b0 ;
  assign n10447 = n922 | n9355 ;
  assign n10448 = n10447 ^ n8473 ^ 1'b0 ;
  assign n10451 = n1315 & ~n6213 ;
  assign n10452 = n10451 ^ n6454 ^ 1'b0 ;
  assign n10449 = ~n6877 & n7135 ;
  assign n10450 = n4648 | n10449 ;
  assign n10453 = n10452 ^ n10450 ^ 1'b0 ;
  assign n10454 = ~n2161 & n3454 ;
  assign n10455 = n7146 & n7955 ;
  assign n10456 = n10454 & n10455 ;
  assign n10457 = n7689 ^ n4363 ^ 1'b0 ;
  assign n10458 = n1031 & n10457 ;
  assign n10459 = n962 & n10458 ;
  assign n10460 = ~n962 & n10459 ;
  assign n10461 = ( n194 & ~n8142 ) | ( n194 & n10460 ) | ( ~n8142 & n10460 ) ;
  assign n10462 = n3353 ^ n2830 ^ 1'b0 ;
  assign n10463 = x2 & ~n4729 ;
  assign n10464 = ~n1839 & n5154 ;
  assign n10465 = n10464 ^ n10190 ^ 1'b0 ;
  assign n10466 = n9566 & ~n10465 ;
  assign n10467 = n6853 ^ n6251 ^ 1'b0 ;
  assign n10468 = ~n6051 & n10467 ;
  assign n10469 = n432 & ~n1900 ;
  assign n10470 = n6423 & n10469 ;
  assign n10471 = n1706 | n6352 ;
  assign n10472 = n574 | n7981 ;
  assign n10473 = n6687 & ~n10472 ;
  assign n10474 = n1623 & n10473 ;
  assign n10475 = ~n704 & n7402 ;
  assign n10476 = n10475 ^ n5792 ^ 1'b0 ;
  assign n10477 = x52 & ~n10476 ;
  assign n10478 = n10477 ^ n3849 ^ 1'b0 ;
  assign n10479 = n4882 & ~n4885 ;
  assign n10480 = n1948 ^ n430 ^ 1'b0 ;
  assign n10481 = n4916 & n10480 ;
  assign n10482 = ~n5861 & n10481 ;
  assign n10483 = n7569 ^ n349 ^ 1'b0 ;
  assign n10484 = n5005 ^ n3632 ^ 1'b0 ;
  assign n10485 = x54 & ~n10484 ;
  assign n10486 = n10485 ^ n3547 ^ n445 ;
  assign n10487 = ~n954 & n1924 ;
  assign n10488 = n5364 | n10487 ;
  assign n10489 = n1114 & ~n10488 ;
  assign n10490 = n1004 | n1935 ;
  assign n10491 = n4898 & n7876 ;
  assign n10492 = ~n10490 & n10491 ;
  assign n10493 = n10005 ^ n613 ^ 1'b0 ;
  assign n10494 = n1254 & n6915 ;
  assign n10495 = n10494 ^ n430 ^ 1'b0 ;
  assign n10496 = n718 | n10495 ;
  assign n10497 = ~n2771 & n6698 ;
  assign n10498 = n2347 | n6579 ;
  assign n10499 = n854 | n4165 ;
  assign n10500 = n1365 ^ n884 ^ 1'b0 ;
  assign n10501 = n1135 ^ n849 ^ 1'b0 ;
  assign n10503 = n5797 ^ n4529 ^ 1'b0 ;
  assign n10502 = n6739 & ~n8382 ;
  assign n10504 = n10503 ^ n10502 ^ 1'b0 ;
  assign n10505 = n10504 ^ n4265 ^ 1'b0 ;
  assign n10506 = n10501 | n10505 ;
  assign n10507 = ~n3350 & n10506 ;
  assign n10508 = n8753 ^ n2388 ^ 1'b0 ;
  assign n10509 = ~n194 & n3748 ;
  assign n10510 = n10509 ^ n595 ^ 1'b0 ;
  assign n10511 = n10510 ^ n3094 ^ 1'b0 ;
  assign n10512 = n3468 | n10511 ;
  assign n10513 = n10508 | n10512 ;
  assign n10514 = n4775 | n7522 ;
  assign n10515 = x54 & ~n394 ;
  assign n10516 = n10515 ^ n2789 ^ 1'b0 ;
  assign n10517 = n549 | n10516 ;
  assign n10518 = n10517 ^ n6335 ^ 1'b0 ;
  assign n10519 = n5500 & n10123 ;
  assign n10520 = n612 & n9017 ;
  assign n10521 = n10520 ^ n9768 ^ 1'b0 ;
  assign n10522 = n2755 ^ n1060 ^ 1'b0 ;
  assign n10523 = n9764 & n10522 ;
  assign n10524 = n8899 ^ n8337 ^ n3702 ;
  assign n10525 = n2019 & n5397 ;
  assign n10526 = n10525 ^ n3215 ^ 1'b0 ;
  assign n10527 = n10526 ^ n3607 ^ 1'b0 ;
  assign n10528 = n1020 & ~n8861 ;
  assign n10529 = n10528 ^ n1035 ^ 1'b0 ;
  assign n10530 = n6553 ^ n1857 ^ 1'b0 ;
  assign n10531 = n221 & n10530 ;
  assign n10532 = n10531 ^ n3969 ^ 1'b0 ;
  assign n10533 = ~n3314 & n10532 ;
  assign n10534 = n10533 ^ n531 ^ 1'b0 ;
  assign n10535 = n4608 & ~n9057 ;
  assign n10536 = n6575 & ~n10535 ;
  assign n10537 = n10536 ^ n394 ^ 1'b0 ;
  assign n10538 = n1107 ^ n131 ^ 1'b0 ;
  assign n10539 = n293 & ~n10538 ;
  assign n10540 = ~n1171 & n10539 ;
  assign n10541 = n10540 ^ n5649 ^ 1'b0 ;
  assign n10542 = n1830 & n9016 ;
  assign n10543 = n10541 & n10542 ;
  assign n10546 = n873 | n4853 ;
  assign n10547 = n3482 | n10546 ;
  assign n10548 = n10547 ^ n6469 ^ 1'b0 ;
  assign n10549 = n10548 ^ n1623 ^ 1'b0 ;
  assign n10550 = n5204 & ~n10549 ;
  assign n10544 = n6766 & ~n7739 ;
  assign n10545 = n4109 & ~n10544 ;
  assign n10551 = n10550 ^ n10545 ^ 1'b0 ;
  assign n10552 = n4227 & n8091 ;
  assign n10553 = n1545 & n6572 ;
  assign n10554 = n7917 ^ n1226 ^ 1'b0 ;
  assign n10555 = n7007 ^ n3477 ^ 1'b0 ;
  assign n10556 = n3788 | n10352 ;
  assign n10557 = n392 & n1948 ;
  assign n10558 = n10557 ^ n3500 ^ 1'b0 ;
  assign n10559 = ~n870 & n5038 ;
  assign n10560 = n7186 & ~n7245 ;
  assign n10561 = n7057 ^ n3790 ^ n1843 ;
  assign n10562 = n608 | n2564 ;
  assign n10563 = ( n2067 & n2413 ) | ( n2067 & n10562 ) | ( n2413 & n10562 ) ;
  assign n10564 = n10561 & ~n10563 ;
  assign n10565 = ~n8387 & n10564 ;
  assign n10566 = n4346 & ~n4413 ;
  assign n10567 = n2174 ^ n1704 ^ 1'b0 ;
  assign n10568 = n10567 ^ n6919 ^ 1'b0 ;
  assign n10569 = n1597 | n4218 ;
  assign n10570 = n2568 | n10569 ;
  assign n10571 = n8720 | n10570 ;
  assign n10572 = ~n3803 & n4205 ;
  assign n10573 = x58 & ~n5113 ;
  assign n10574 = n4193 ^ n3221 ^ 1'b0 ;
  assign n10575 = n10573 & n10574 ;
  assign n10576 = n8113 & n10575 ;
  assign n10588 = n512 & n3301 ;
  assign n10577 = x52 & ~n430 ;
  assign n10578 = n10577 ^ n10517 ^ 1'b0 ;
  assign n10579 = n4336 ^ n3395 ^ 1'b0 ;
  assign n10580 = n2596 ^ n1543 ^ 1'b0 ;
  assign n10581 = ~n2653 & n10580 ;
  assign n10582 = n570 | n10581 ;
  assign n10583 = n10579 & ~n10582 ;
  assign n10584 = n1782 & n7393 ;
  assign n10585 = n10584 ^ n8283 ^ 1'b0 ;
  assign n10586 = n10583 | n10585 ;
  assign n10587 = ~n10578 & n10586 ;
  assign n10589 = n10588 ^ n10587 ^ n2035 ;
  assign n10590 = n2154 ^ n2034 ^ 1'b0 ;
  assign n10591 = n1162 & ~n10590 ;
  assign n10592 = ~n7656 & n10591 ;
  assign n10593 = n4133 ^ n1035 ^ 1'b0 ;
  assign n10594 = n10592 & ~n10593 ;
  assign n10595 = ~n1964 & n10594 ;
  assign n10596 = n8590 ^ n8279 ^ 1'b0 ;
  assign n10597 = n7749 & n10596 ;
  assign n10598 = n2656 | n10500 ;
  assign n10599 = n7498 ^ n1325 ^ 1'b0 ;
  assign n10600 = ~n2241 & n5125 ;
  assign n10601 = ~n3762 & n5854 ;
  assign n10602 = n10601 ^ n8305 ^ 1'b0 ;
  assign n10603 = n5621 ^ n2769 ^ 1'b0 ;
  assign n10604 = n10602 & n10603 ;
  assign n10605 = n6705 ^ n784 ^ 1'b0 ;
  assign n10611 = ( ~n335 & n2390 ) | ( ~n335 & n5181 ) | ( n2390 & n5181 ) ;
  assign n10612 = n10611 ^ n9622 ^ 1'b0 ;
  assign n10606 = n266 & n1883 ;
  assign n10607 = n10606 ^ n2565 ^ 1'b0 ;
  assign n10608 = ~n2650 & n3687 ;
  assign n10609 = n4296 & n10608 ;
  assign n10610 = n10607 & ~n10609 ;
  assign n10613 = n10612 ^ n10610 ^ 1'b0 ;
  assign n10614 = n7112 | n9622 ;
  assign n10615 = n10614 ^ n8518 ^ 1'b0 ;
  assign n10616 = n10613 | n10615 ;
  assign n10617 = n508 | n10586 ;
  assign n10618 = n10217 ^ n7025 ^ n4019 ;
  assign n10619 = n4786 | n6228 ;
  assign n10620 = n3640 | n4313 ;
  assign n10621 = n10620 ^ n277 ^ 1'b0 ;
  assign n10622 = n3573 ^ n945 ^ 1'b0 ;
  assign n10623 = n6824 & n10622 ;
  assign n10624 = n10623 ^ n3774 ^ 1'b0 ;
  assign n10625 = ~n5105 & n9835 ;
  assign n10626 = n4298 & n10625 ;
  assign n10627 = n4715 & ~n10626 ;
  assign n10628 = n10627 ^ n430 ^ 1'b0 ;
  assign n10629 = n2709 ^ n2210 ^ 1'b0 ;
  assign n10630 = n512 & ~n10629 ;
  assign n10631 = ~n735 & n6436 ;
  assign n10632 = n1380 & ~n2171 ;
  assign n10633 = n2037 | n10632 ;
  assign n10634 = n2907 & n10633 ;
  assign n10635 = ~n10631 & n10634 ;
  assign n10636 = n4197 ^ n2650 ^ 1'b0 ;
  assign n10638 = n1945 | n2465 ;
  assign n10639 = n2972 | n10638 ;
  assign n10637 = ~n132 & n4113 ;
  assign n10640 = n10639 ^ n10637 ^ 1'b0 ;
  assign n10641 = n994 | n10640 ;
  assign n10642 = n2608 & ~n6407 ;
  assign n10643 = ~n877 & n3135 ;
  assign n10644 = n10643 ^ n9660 ^ n4038 ;
  assign n10645 = n747 | n834 ;
  assign n10646 = n834 & ~n10645 ;
  assign n10647 = ~n1060 & n10646 ;
  assign n10648 = n4025 & n10647 ;
  assign n10649 = n10648 ^ n1401 ^ 1'b0 ;
  assign n10650 = n2391 | n9307 ;
  assign n10651 = n10649 & n10650 ;
  assign n10652 = ~n10649 & n10651 ;
  assign n10653 = n181 & n2157 ;
  assign n10654 = n7139 ^ n7014 ^ 1'b0 ;
  assign n10655 = ~n3999 & n10654 ;
  assign n10656 = ~n9744 & n10655 ;
  assign n10657 = n9744 & n10656 ;
  assign n10658 = n10653 & ~n10657 ;
  assign n10659 = n10652 & n10658 ;
  assign n10660 = n1867 ^ n1281 ^ 1'b0 ;
  assign n10661 = n2945 & n8722 ;
  assign n10662 = n3692 & ~n10661 ;
  assign n10663 = n1228 & ~n9713 ;
  assign n10664 = n660 | n5790 ;
  assign n10665 = n10664 ^ n8018 ^ 1'b0 ;
  assign n10666 = n2393 | n4600 ;
  assign n10667 = ~n1067 & n7402 ;
  assign n10668 = n10667 ^ n1391 ^ 1'b0 ;
  assign n10669 = n1819 & ~n10668 ;
  assign n10670 = n2563 ^ n1882 ^ 1'b0 ;
  assign n10671 = x36 & n10670 ;
  assign n10672 = n2078 & n3899 ;
  assign n10673 = n10672 ^ n3220 ^ 1'b0 ;
  assign n10674 = n8015 & ~n10673 ;
  assign n10675 = n10674 ^ n4230 ^ n466 ;
  assign n10676 = ~n9441 & n10675 ;
  assign n10677 = ~n9362 & n10676 ;
  assign n10678 = n9275 ^ n5753 ^ 1'b0 ;
  assign n10679 = ~n10677 & n10678 ;
  assign n10680 = n5723 & ~n6834 ;
  assign n10681 = n10680 ^ n294 ^ 1'b0 ;
  assign n10682 = n8352 & n8395 ;
  assign n10683 = n3267 ^ n1412 ^ 1'b0 ;
  assign n10684 = n3413 & ~n10683 ;
  assign n10685 = ~x77 & n9490 ;
  assign n10686 = n10685 ^ n4186 ^ 1'b0 ;
  assign n10687 = n1671 | n5734 ;
  assign n10688 = n10687 ^ n4334 ^ 1'b0 ;
  assign n10689 = ~n3191 & n10688 ;
  assign n10690 = n10689 ^ n6445 ^ 1'b0 ;
  assign n10691 = ( n830 & n1336 ) | ( n830 & ~n5406 ) | ( n1336 & ~n5406 ) ;
  assign n10692 = n6019 | n10691 ;
  assign n10693 = n4859 ^ n584 ^ 1'b0 ;
  assign n10694 = n4515 & ~n10693 ;
  assign n10695 = n3052 & n10694 ;
  assign n10696 = n10692 & ~n10695 ;
  assign n10697 = n884 & n1414 ;
  assign n10698 = n10697 ^ n1548 ^ 1'b0 ;
  assign n10699 = n3145 ^ n478 ^ 1'b0 ;
  assign n10700 = n6442 | n9130 ;
  assign n10701 = n10700 ^ n1368 ^ 1'b0 ;
  assign n10702 = n1939 & n3002 ;
  assign n10703 = ~n10701 & n10702 ;
  assign n10704 = n5990 ^ n1291 ^ 1'b0 ;
  assign n10705 = n1191 & n3596 ;
  assign n10706 = n1550 & n10705 ;
  assign n10707 = n10706 ^ n7887 ^ n6520 ;
  assign n10708 = n10550 ^ n8655 ^ 1'b0 ;
  assign n10709 = x17 & n2885 ;
  assign n10710 = n7818 ^ n7172 ^ n2314 ;
  assign n10711 = x87 & n5090 ;
  assign n10712 = ~n2099 & n10711 ;
  assign n10713 = n2741 ^ n1254 ^ 1'b0 ;
  assign n10714 = n2604 & ~n10713 ;
  assign n10715 = n6244 | n10714 ;
  assign n10716 = n4521 | n9425 ;
  assign n10717 = n2312 & ~n3199 ;
  assign n10718 = n10717 ^ n7554 ^ 1'b0 ;
  assign n10720 = n2366 & n2906 ;
  assign n10719 = n1228 & n8731 ;
  assign n10721 = n10720 ^ n10719 ^ 1'b0 ;
  assign n10723 = n7876 ^ n3350 ^ 1'b0 ;
  assign n10724 = n1241 & ~n10723 ;
  assign n10722 = n3802 & ~n4430 ;
  assign n10725 = n10724 ^ n10722 ^ 1'b0 ;
  assign n10726 = n1206 | n6716 ;
  assign n10727 = n8324 | n10726 ;
  assign n10728 = n10727 ^ n3549 ^ 1'b0 ;
  assign n10729 = n1165 & ~n4746 ;
  assign n10730 = n4746 & n10729 ;
  assign n10731 = n10730 ^ n1909 ^ 1'b0 ;
  assign n10732 = n358 | n427 ;
  assign n10733 = n358 & ~n10732 ;
  assign n10734 = ~n1055 & n10733 ;
  assign n10735 = n616 & n1449 ;
  assign n10736 = n10734 & n10735 ;
  assign n10737 = n1489 & ~n10736 ;
  assign n10738 = ~n1489 & n10737 ;
  assign n10739 = n9524 & n10738 ;
  assign n10740 = ~n10731 & n10739 ;
  assign n10741 = n381 & ~n1067 ;
  assign n10742 = ~n381 & n10741 ;
  assign n10743 = n955 & ~n3191 ;
  assign n10744 = n10742 & n10743 ;
  assign n10745 = n4429 & ~n10744 ;
  assign n10746 = ~n4429 & n10745 ;
  assign n10747 = ( n618 & ~n10740 ) | ( n618 & n10746 ) | ( ~n10740 & n10746 ) ;
  assign n10748 = ~n343 & n4128 ;
  assign n10749 = n942 & ~n6626 ;
  assign n10750 = ~n1467 & n10749 ;
  assign n10751 = n2420 & n2521 ;
  assign n10752 = n10751 ^ n5702 ^ 1'b0 ;
  assign n10753 = ~n10708 & n10752 ;
  assign n10754 = n10753 ^ n1171 ^ 1'b0 ;
  assign n10755 = n1572 ^ n332 ^ 1'b0 ;
  assign n10756 = n2347 & ~n10755 ;
  assign n10757 = ~n624 & n10756 ;
  assign n10758 = ~n10756 & n10757 ;
  assign n10759 = n4579 ^ n1953 ^ 1'b0 ;
  assign n10760 = n7006 ^ n3715 ^ 1'b0 ;
  assign n10761 = n9486 ^ n5595 ^ n5123 ;
  assign n10762 = n311 & n620 ;
  assign n10763 = n10762 ^ n3790 ^ 1'b0 ;
  assign n10764 = n10763 ^ n4775 ^ 1'b0 ;
  assign n10765 = ~n459 & n10764 ;
  assign n10767 = ~n2911 & n5234 ;
  assign n10768 = n10767 ^ n7941 ^ 1'b0 ;
  assign n10766 = n1662 & ~n7835 ;
  assign n10769 = n10768 ^ n10766 ^ 1'b0 ;
  assign n10770 = n2608 ^ n1664 ^ 1'b0 ;
  assign n10771 = n9660 & n10770 ;
  assign n10772 = n7792 ^ n7439 ^ 1'b0 ;
  assign n10773 = n5013 & n10772 ;
  assign n10774 = ~n7597 & n10773 ;
  assign n10775 = n1648 | n4631 ;
  assign n10776 = n3366 & ~n10775 ;
  assign n10777 = x32 & n980 ;
  assign n10778 = n8249 ^ n4061 ^ 1'b0 ;
  assign n10779 = n10777 & n10778 ;
  assign n10780 = n4336 & n10779 ;
  assign n10783 = n3157 ^ n998 ^ n902 ;
  assign n10784 = ~n4296 & n10783 ;
  assign n10785 = n10784 ^ n2655 ^ 1'b0 ;
  assign n10781 = n5243 ^ n5132 ^ 1'b0 ;
  assign n10782 = ~n6158 & n10781 ;
  assign n10786 = n10785 ^ n10782 ^ 1'b0 ;
  assign n10787 = x53 & n10786 ;
  assign n10788 = ~n10780 & n10787 ;
  assign n10789 = n10096 ^ n7211 ^ 1'b0 ;
  assign n10790 = n6992 ^ n4506 ^ 1'b0 ;
  assign n10793 = n4032 ^ n3245 ^ 1'b0 ;
  assign n10791 = n4175 ^ n1180 ^ 1'b0 ;
  assign n10792 = ~n435 & n10791 ;
  assign n10794 = n10793 ^ n10792 ^ 1'b0 ;
  assign n10795 = ~n9727 & n10794 ;
  assign n10796 = n5306 | n10764 ;
  assign n10797 = n10796 ^ n4117 ^ 1'b0 ;
  assign n10798 = n6940 | n9608 ;
  assign n10799 = n10798 ^ n10153 ^ 1'b0 ;
  assign n10800 = n2600 & ~n10537 ;
  assign n10801 = n3895 ^ n3821 ^ 1'b0 ;
  assign n10802 = n7941 & ~n10801 ;
  assign n10803 = n6488 ^ n560 ^ 1'b0 ;
  assign n10804 = n1070 & ~n1759 ;
  assign n10805 = n10804 ^ n8538 ^ 1'b0 ;
  assign n10806 = n6176 ^ n627 ^ 1'b0 ;
  assign n10808 = n6712 ^ n6194 ^ 1'b0 ;
  assign n10807 = x23 & n219 ;
  assign n10809 = n10808 ^ n10807 ^ 1'b0 ;
  assign n10810 = n3163 | n10809 ;
  assign n10811 = n2621 & n6616 ;
  assign n10812 = n10040 & n10811 ;
  assign n10813 = n10812 ^ n8644 ^ 1'b0 ;
  assign n10814 = ~n4014 & n7522 ;
  assign n10815 = n10814 ^ n8965 ^ 1'b0 ;
  assign n10816 = n5741 & n7468 ;
  assign n10817 = n5941 ^ n747 ^ 1'b0 ;
  assign n10818 = n10817 ^ n1059 ^ 1'b0 ;
  assign n10819 = n10816 | n10818 ;
  assign n10820 = n10819 ^ n1041 ^ 1'b0 ;
  assign n10822 = n1502 & ~n2198 ;
  assign n10821 = n1497 & ~n2278 ;
  assign n10823 = n10822 ^ n10821 ^ 1'b0 ;
  assign n10824 = n766 & n10823 ;
  assign n10825 = n10824 ^ n6853 ^ 1'b0 ;
  assign n10826 = n4356 ^ n2091 ^ 1'b0 ;
  assign n10827 = ~n1336 & n10826 ;
  assign n10830 = n6592 & n6935 ;
  assign n10828 = ~n3300 & n7601 ;
  assign n10829 = n7915 & n10828 ;
  assign n10831 = n10830 ^ n10829 ^ 1'b0 ;
  assign n10832 = n10831 ^ n9315 ^ 1'b0 ;
  assign n10833 = n4227 ^ n695 ^ x52 ;
  assign n10834 = n10833 ^ n7427 ^ 1'b0 ;
  assign n10835 = ( n4344 & n7807 ) | ( n4344 & ~n10834 ) | ( n7807 & ~n10834 ) ;
  assign n10836 = ~n931 & n4213 ;
  assign n10837 = n457 | n3760 ;
  assign n10838 = n481 & ~n10837 ;
  assign n10839 = n2948 | n9350 ;
  assign n10840 = x84 | n10839 ;
  assign n10841 = ~n10838 & n10840 ;
  assign n10842 = n5317 ^ x127 ^ 1'b0 ;
  assign n10843 = ~n8621 & n10842 ;
  assign n10845 = n3027 | n3085 ;
  assign n10846 = n10845 ^ n700 ^ 1'b0 ;
  assign n10844 = n190 & ~n7984 ;
  assign n10847 = n10846 ^ n10844 ^ 1'b0 ;
  assign n10848 = n8224 ^ n2139 ^ 1'b0 ;
  assign n10849 = n5119 ^ n371 ^ 1'b0 ;
  assign n10850 = x59 & ~n1508 ;
  assign n10851 = n2786 & n10850 ;
  assign n10852 = n10706 ^ n8319 ^ 1'b0 ;
  assign n10853 = n10851 | n10852 ;
  assign n10854 = n1842 & n3046 ;
  assign n10855 = n10854 ^ n8227 ^ 1'b0 ;
  assign n10856 = n5907 & ~n10855 ;
  assign n10857 = n10553 ^ n5689 ^ 1'b0 ;
  assign n10858 = n2160 & n7237 ;
  assign n10859 = ~n1227 & n3695 ;
  assign n10860 = n6226 ^ n4775 ^ 1'b0 ;
  assign n10861 = n3696 & n6590 ;
  assign n10862 = n9566 ^ n7529 ^ 1'b0 ;
  assign n10863 = n10862 ^ n4623 ^ 1'b0 ;
  assign n10864 = n9588 ^ n3807 ^ 1'b0 ;
  assign n10865 = n10864 ^ n3874 ^ 1'b0 ;
  assign n10866 = ~x58 & n10865 ;
  assign n10867 = n10129 ^ n895 ^ 1'b0 ;
  assign n10868 = n4312 & ~n7548 ;
  assign n10869 = n4790 & ~n5289 ;
  assign n10872 = n3580 ^ n538 ^ 1'b0 ;
  assign n10873 = n7690 & n10872 ;
  assign n10870 = n6407 & n7374 ;
  assign n10871 = n3926 | n10870 ;
  assign n10874 = n10873 ^ n10871 ^ 1'b0 ;
  assign n10875 = n4736 & ~n5469 ;
  assign n10876 = n10875 ^ n2961 ^ 1'b0 ;
  assign n10877 = n1905 & n2374 ;
  assign n10878 = n153 & n10877 ;
  assign n10879 = n3661 | n10878 ;
  assign n10880 = n10879 ^ n5061 ^ 1'b0 ;
  assign n10881 = n5378 & ~n10880 ;
  assign n10882 = ~n1667 & n4217 ;
  assign n10883 = n10882 ^ n749 ^ 1'b0 ;
  assign n10884 = n10883 ^ n2932 ^ 1'b0 ;
  assign n10885 = n9730 ^ n984 ^ 1'b0 ;
  assign n10886 = n10884 & ~n10885 ;
  assign n10887 = n716 & ~n2115 ;
  assign n10888 = n4898 & ~n10887 ;
  assign n10889 = n10888 ^ n9210 ^ 1'b0 ;
  assign n10890 = n363 | n1052 ;
  assign n10891 = ~n4129 & n6444 ;
  assign n10892 = n7033 ^ n1315 ^ 1'b0 ;
  assign n10893 = n6365 & ~n10892 ;
  assign n10894 = ~n4150 & n10893 ;
  assign n10895 = n10894 ^ n562 ^ 1'b0 ;
  assign n10896 = n1013 ^ n325 ^ 1'b0 ;
  assign n10897 = n7092 ^ n4499 ^ 1'b0 ;
  assign n10898 = ~n7827 & n7942 ;
  assign n10899 = n10897 & n10898 ;
  assign n10900 = x106 & n3721 ;
  assign n10901 = n5814 & n10900 ;
  assign n10902 = n5923 ^ n482 ^ 1'b0 ;
  assign n10903 = ~n8260 & n10902 ;
  assign n10904 = n5399 ^ n2601 ^ 1'b0 ;
  assign n10905 = n5595 & ~n10904 ;
  assign n10906 = n3145 & ~n5050 ;
  assign n10907 = n302 & n2313 ;
  assign n10908 = n10906 & n10907 ;
  assign n10909 = ( n200 & n7335 ) | ( n200 & n10908 ) | ( n7335 & n10908 ) ;
  assign n10910 = n4918 ^ n4563 ^ 1'b0 ;
  assign n10911 = ~n5458 & n10910 ;
  assign n10912 = n4124 & ~n10911 ;
  assign n10913 = n3299 ^ n3094 ^ 1'b0 ;
  assign n10914 = x57 | n4847 ;
  assign n10915 = n2452 & n4393 ;
  assign n10916 = n10915 ^ n7972 ^ 1'b0 ;
  assign n10917 = n1994 & ~n2656 ;
  assign n10918 = n10917 ^ n1008 ^ 1'b0 ;
  assign n10919 = n2439 & n10918 ;
  assign n10920 = n4793 & n10919 ;
  assign n10921 = n3525 | n10920 ;
  assign n10922 = n10132 & ~n10921 ;
  assign n10923 = ~n2315 & n4673 ;
  assign n10924 = n10923 ^ x64 ^ 1'b0 ;
  assign n10925 = n261 & n10924 ;
  assign n10926 = n248 & n3509 ;
  assign n10927 = ~n7574 & n10926 ;
  assign n10928 = ~n1764 & n6451 ;
  assign n10929 = n10928 ^ n5832 ^ 1'b0 ;
  assign n10931 = n1786 ^ n342 ^ 1'b0 ;
  assign n10930 = ~n2038 & n5354 ;
  assign n10932 = n10931 ^ n10930 ^ 1'b0 ;
  assign n10933 = n10550 & ~n10932 ;
  assign n10934 = n1079 & n10933 ;
  assign n10935 = n7836 ^ n1552 ^ 1'b0 ;
  assign n10936 = n6694 ^ x119 ^ 1'b0 ;
  assign n10937 = n810 & ~n3015 ;
  assign n10938 = ~n2516 & n6211 ;
  assign n10939 = n932 & n10938 ;
  assign n10940 = n4995 | n10939 ;
  assign n10941 = n10940 ^ n819 ^ 1'b0 ;
  assign n10942 = n9713 | n10941 ;
  assign n10943 = n10937 | n10942 ;
  assign n10944 = n4117 ^ n2775 ^ 1'b0 ;
  assign n10945 = n6128 ^ n451 ^ 1'b0 ;
  assign n10946 = ~n4450 & n10945 ;
  assign n10947 = n1149 | n10946 ;
  assign n10948 = n7991 ^ n5580 ^ 1'b0 ;
  assign n10949 = n9333 ^ n7650 ^ n3558 ;
  assign n10950 = n2732 & n4681 ;
  assign n10951 = n3293 & n10950 ;
  assign n10952 = n323 & ~n590 ;
  assign n10953 = n3552 | n4511 ;
  assign n10954 = n10953 ^ n1397 ^ 1'b0 ;
  assign n10955 = n3149 & n7350 ;
  assign n10956 = n7190 ^ n1602 ^ 1'b0 ;
  assign n10957 = n6177 & n9605 ;
  assign n10958 = n1147 & n7848 ;
  assign n10959 = n8537 & ~n10958 ;
  assign n10960 = n10959 ^ n3838 ^ 1'b0 ;
  assign n10961 = n9560 & ~n10960 ;
  assign n10964 = n4232 & ~n5132 ;
  assign n10965 = ~n400 & n10964 ;
  assign n10966 = n10965 ^ n2144 ^ 1'b0 ;
  assign n10962 = n6430 ^ n5685 ^ 1'b0 ;
  assign n10963 = n439 | n10962 ;
  assign n10967 = n10966 ^ n10963 ^ 1'b0 ;
  assign n10968 = ~n3046 & n7129 ;
  assign n10969 = n6239 ^ n4505 ^ 1'b0 ;
  assign n10970 = n1656 | n10969 ;
  assign n10971 = ~n3064 & n5381 ;
  assign n10972 = ~n1219 & n1713 ;
  assign n10973 = n6461 | n8444 ;
  assign n10974 = n10973 ^ n9290 ^ 1'b0 ;
  assign n10975 = ~n1973 & n4391 ;
  assign n10976 = n9181 ^ n1762 ^ n837 ;
  assign n10977 = ~n10975 & n10976 ;
  assign n10978 = n10974 & n10977 ;
  assign n10979 = n6378 ^ n909 ^ 1'b0 ;
  assign n10980 = n336 & n10979 ;
  assign n10981 = n5635 ^ n5517 ^ 1'b0 ;
  assign n10982 = n3754 & n5110 ;
  assign n10983 = ~n3818 & n10982 ;
  assign n10984 = n10983 ^ n1694 ^ 1'b0 ;
  assign n10985 = ~n10981 & n10984 ;
  assign n10986 = n5769 | n6239 ;
  assign n10994 = n4117 ^ n2566 ^ 1'b0 ;
  assign n10987 = n642 | n1532 ;
  assign n10991 = n1495 ^ n992 ^ 1'b0 ;
  assign n10988 = n5019 ^ n4306 ^ 1'b0 ;
  assign n10989 = ~n1513 & n10988 ;
  assign n10990 = ~n5246 & n10989 ;
  assign n10992 = n10991 ^ n10990 ^ 1'b0 ;
  assign n10993 = n10987 | n10992 ;
  assign n10995 = n10994 ^ n10993 ^ 1'b0 ;
  assign n10996 = n2113 & n2924 ;
  assign n10997 = n10996 ^ n6478 ^ 1'b0 ;
  assign n10998 = n2176 | n9554 ;
  assign n10999 = n8527 ^ n1530 ^ 1'b0 ;
  assign n11000 = n1833 & n9060 ;
  assign n11001 = n11000 ^ n2585 ^ 1'b0 ;
  assign n11002 = n1808 & n2866 ;
  assign n11003 = n11002 ^ n2151 ^ 1'b0 ;
  assign n11005 = n3134 | n3142 ;
  assign n11006 = n11005 ^ n2253 ^ 1'b0 ;
  assign n11004 = n1854 | n3553 ;
  assign n11007 = n11006 ^ n11004 ^ 1'b0 ;
  assign n11008 = n11003 | n11007 ;
  assign n11009 = n2533 & ~n8912 ;
  assign n11010 = ~n806 & n2055 ;
  assign n11011 = ~n6373 & n10986 ;
  assign n11012 = n3195 & n11011 ;
  assign n11013 = n4254 & n9611 ;
  assign n11014 = n11013 ^ n639 ^ 1'b0 ;
  assign n11015 = n11014 ^ n6014 ^ 1'b0 ;
  assign n11016 = ~n7009 & n11015 ;
  assign n11017 = ~n5430 & n6369 ;
  assign n11018 = n7847 ^ n7090 ^ 1'b0 ;
  assign n11019 = n3091 | n11018 ;
  assign n11020 = n5792 ^ n1895 ^ 1'b0 ;
  assign n11021 = n4050 | n11020 ;
  assign n11022 = n5557 & ~n5793 ;
  assign n11023 = n11022 ^ n7870 ^ 1'b0 ;
  assign n11024 = n3371 & n4959 ;
  assign n11025 = n11024 ^ n5783 ^ 1'b0 ;
  assign n11026 = n1185 ^ n604 ^ 1'b0 ;
  assign n11027 = n3669 | n11026 ;
  assign n11028 = n4988 & n6236 ;
  assign n11029 = n2627 & n11028 ;
  assign n11030 = n11027 & ~n11029 ;
  assign n11031 = ~n5141 & n5959 ;
  assign n11032 = n5782 | n7104 ;
  assign n11033 = n6959 & n11032 ;
  assign n11034 = n11033 ^ n5417 ^ 1'b0 ;
  assign n11035 = ~n2512 & n4158 ;
  assign n11036 = ~n216 & n609 ;
  assign n11037 = ~n11035 & n11036 ;
  assign n11038 = n613 & n5354 ;
  assign n11039 = n3230 & n5442 ;
  assign n11040 = n6369 | n11039 ;
  assign n11041 = n10818 ^ n7382 ^ 1'b0 ;
  assign n11042 = n7231 ^ n2585 ^ 1'b0 ;
  assign n11043 = n6421 | n11042 ;
  assign n11044 = ~n7046 & n7259 ;
  assign n11045 = n1786 & ~n6355 ;
  assign n11046 = n744 | n1601 ;
  assign n11047 = n11046 ^ n221 ^ 1'b0 ;
  assign n11048 = ~n6669 & n7118 ;
  assign n11049 = ~n11047 & n11048 ;
  assign n11050 = n11045 | n11049 ;
  assign n11051 = n11050 ^ n2711 ^ 1'b0 ;
  assign n11052 = ~n3510 & n8511 ;
  assign n11053 = x124 & n6549 ;
  assign n11054 = n9277 ^ n9238 ^ 1'b0 ;
  assign n11055 = ( n3302 & n3608 ) | ( n3302 & n4740 ) | ( n3608 & n4740 ) ;
  assign n11056 = n4616 & n5899 ;
  assign n11057 = ~n3461 & n5166 ;
  assign n11058 = n11057 ^ n8615 ^ 1'b0 ;
  assign n11059 = ~n11056 & n11058 ;
  assign n11060 = n11055 & n11059 ;
  assign n11061 = n5632 ^ n4177 ^ 1'b0 ;
  assign n11062 = n11061 ^ n1724 ^ 1'b0 ;
  assign n11063 = n5716 ^ n705 ^ 1'b0 ;
  assign n11064 = ~n11062 & n11063 ;
  assign n11065 = n7781 & n11064 ;
  assign n11066 = n11060 & n11065 ;
  assign n11067 = n6805 | n9713 ;
  assign n11068 = ( ~n771 & n2062 ) | ( ~n771 & n7269 ) | ( n2062 & n7269 ) ;
  assign n11069 = n1903 | n5540 ;
  assign n11070 = n7232 | n10567 ;
  assign n11071 = n3074 | n10129 ;
  assign n11072 = n2650 ^ n1663 ^ 1'b0 ;
  assign n11073 = n6526 & ~n11072 ;
  assign n11074 = n6572 & n9656 ;
  assign n11075 = n11074 ^ n8389 ^ 1'b0 ;
  assign n11076 = n430 & ~n3547 ;
  assign n11077 = n11075 & n11076 ;
  assign n11078 = n3371 | n4701 ;
  assign n11079 = n11078 ^ n1325 ^ 1'b0 ;
  assign n11080 = n2803 & n11079 ;
  assign n11081 = n11080 ^ n3987 ^ 1'b0 ;
  assign n11082 = ~n2705 & n5418 ;
  assign n11083 = n11082 ^ n3559 ^ 1'b0 ;
  assign n11084 = n11081 & ~n11083 ;
  assign n11085 = n3646 & n9300 ;
  assign n11086 = n8052 ^ n5181 ^ 1'b0 ;
  assign n11087 = n1747 & n11086 ;
  assign n11088 = n11087 ^ n1899 ^ 1'b0 ;
  assign n11089 = n8881 ^ n3964 ^ 1'b0 ;
  assign n11090 = n11089 ^ n8382 ^ 1'b0 ;
  assign n11091 = ~n10968 & n11090 ;
  assign n11092 = ~n549 & n728 ;
  assign n11093 = n2759 | n11092 ;
  assign n11094 = x27 | n11093 ;
  assign n11095 = n11094 ^ n8902 ^ 1'b0 ;
  assign n11096 = ~n1885 & n11095 ;
  assign n11097 = n2166 & ~n4731 ;
  assign n11098 = n5602 & n11097 ;
  assign n11099 = n6313 & n11098 ;
  assign n11100 = ~n2171 & n10344 ;
  assign n11101 = n4623 & n4647 ;
  assign n11102 = ~n7158 & n11101 ;
  assign n11104 = ~n1781 & n5343 ;
  assign n11103 = n1188 & ~n8775 ;
  assign n11105 = n11104 ^ n11103 ^ 1'b0 ;
  assign n11106 = ~n9774 & n11105 ;
  assign n11107 = ( x35 & n2090 ) | ( x35 & n2471 ) | ( n2090 & n2471 ) ;
  assign n11108 = n1013 & n7337 ;
  assign n11109 = ~n4823 & n8190 ;
  assign n11110 = n11109 ^ n5656 ^ 1'b0 ;
  assign n11111 = n446 & ~n2867 ;
  assign n11112 = n5098 ^ n2523 ^ 1'b0 ;
  assign n11113 = n11111 | n11112 ;
  assign n11114 = n11113 ^ n4190 ^ 1'b0 ;
  assign n11115 = n2621 & ~n3116 ;
  assign n11116 = n3946 ^ n2767 ^ 1'b0 ;
  assign n11117 = n3428 | n4418 ;
  assign n11118 = ~n11116 & n11117 ;
  assign n11119 = n571 | n945 ;
  assign n11120 = n261 | n10683 ;
  assign n11121 = n4584 & ~n11120 ;
  assign n11122 = n1487 & ~n10846 ;
  assign n11123 = n3970 | n4177 ;
  assign n11124 = n1118 & ~n3764 ;
  assign n11125 = ~n831 & n1439 ;
  assign n11126 = ~n586 & n11125 ;
  assign n11127 = n11124 | n11126 ;
  assign n11128 = n5240 ^ n866 ^ 1'b0 ;
  assign n11129 = n7786 ^ n5373 ^ n3551 ;
  assign n11130 = n3296 & n11129 ;
  assign n11131 = n5885 & ~n11130 ;
  assign n11132 = n832 & n4254 ;
  assign n11133 = ~n865 & n11132 ;
  assign n11134 = n11133 ^ n5821 ^ 1'b0 ;
  assign n11135 = n9333 ^ n2307 ^ 1'b0 ;
  assign n11136 = n11135 ^ n8444 ^ 1'b0 ;
  assign n11137 = ~n1808 & n11136 ;
  assign n11138 = n8046 & n11137 ;
  assign n11139 = ~n8022 & n11138 ;
  assign n11140 = ~n806 & n10403 ;
  assign n11141 = ~n6987 & n11140 ;
  assign n11142 = n8345 ^ n530 ^ 1'b0 ;
  assign n11143 = n177 & n1221 ;
  assign n11144 = ~n4883 & n11143 ;
  assign n11145 = ~n757 & n11144 ;
  assign n11146 = ~n3640 & n11145 ;
  assign n11147 = n1882 ^ n171 ^ 1'b0 ;
  assign n11148 = n5194 & n11147 ;
  assign n11149 = n11148 ^ n3413 ^ 1'b0 ;
  assign n11150 = x19 & n804 ;
  assign n11151 = ~x23 & n3465 ;
  assign n11152 = n5403 | n11151 ;
  assign n11153 = n11152 ^ n2650 ^ 1'b0 ;
  assign n11154 = n7162 & ~n7511 ;
  assign n11155 = n11154 ^ n7360 ^ 1'b0 ;
  assign n11156 = n11155 ^ n4679 ^ 1'b0 ;
  assign n11157 = n1181 & ~n6501 ;
  assign n11158 = n8444 | n10177 ;
  assign n11159 = n2815 | n7624 ;
  assign n11160 = n11159 ^ n1862 ^ 1'b0 ;
  assign n11161 = n11160 ^ n3268 ^ x44 ;
  assign n11162 = n2638 & ~n3635 ;
  assign n11163 = n4095 & n11162 ;
  assign n11164 = n7077 & ~n11163 ;
  assign n11165 = n11164 ^ n7723 ^ 1'b0 ;
  assign n11166 = n7128 ^ n4499 ^ 1'b0 ;
  assign n11167 = n10702 ^ n6632 ^ 1'b0 ;
  assign n11168 = ~n4616 & n11167 ;
  assign n11169 = ~n4417 & n8035 ;
  assign n11170 = ~n8623 & n11169 ;
  assign n11171 = n10283 ^ n8905 ^ 1'b0 ;
  assign n11172 = n11171 ^ n2398 ^ 1'b0 ;
  assign n11173 = ~n3706 & n11172 ;
  assign n11174 = n6251 ^ n5958 ^ 1'b0 ;
  assign n11175 = n6598 ^ n3064 ^ 1'b0 ;
  assign n11176 = n3898 ^ n1529 ^ 1'b0 ;
  assign n11177 = n9419 & n11176 ;
  assign n11178 = ~n4001 & n11177 ;
  assign n11179 = ~n2490 & n6638 ;
  assign n11180 = n2490 & n11179 ;
  assign n11181 = n2136 | n11180 ;
  assign n11182 = n4322 ^ n4296 ^ 1'b0 ;
  assign n11183 = n4835 & ~n11182 ;
  assign n11184 = n2222 & ~n9133 ;
  assign n11185 = n11184 ^ x40 ^ 1'b0 ;
  assign n11186 = n3279 ^ n2691 ^ 1'b0 ;
  assign n11187 = ( n2269 & n2475 ) | ( n2269 & n2986 ) | ( n2475 & n2986 ) ;
  assign n11188 = n11186 & ~n11187 ;
  assign n11189 = ~n2083 & n11188 ;
  assign n11190 = n11189 ^ n9916 ^ 1'b0 ;
  assign n11191 = n5264 ^ n764 ^ 1'b0 ;
  assign n11192 = n5144 ^ n1281 ^ 1'b0 ;
  assign n11193 = n11191 | n11192 ;
  assign n11194 = ~n757 & n1733 ;
  assign n11195 = n11194 ^ n4438 ^ 1'b0 ;
  assign n11196 = n6539 | n11195 ;
  assign n11197 = n4568 & ~n11196 ;
  assign n11198 = n1543 & n1920 ;
  assign n11199 = n650 | n3760 ;
  assign n11200 = n4351 | n11199 ;
  assign n11201 = n7683 | n11200 ;
  assign n11202 = n11201 ^ n7001 ^ 1'b0 ;
  assign n11203 = n7246 ^ x73 ^ 1'b0 ;
  assign n11204 = n6766 & n11203 ;
  assign n11205 = ~n3659 & n11204 ;
  assign n11206 = n3336 | n5874 ;
  assign n11207 = n11206 ^ n10931 ^ 1'b0 ;
  assign n11208 = ( ~n5329 & n8325 ) | ( ~n5329 & n11061 ) | ( n8325 & n11061 ) ;
  assign n11209 = n7676 ^ n5649 ^ 1'b0 ;
  assign n11210 = n1352 ^ n859 ^ 1'b0 ;
  assign n11211 = ~n1986 & n8683 ;
  assign n11212 = n7854 & n11211 ;
  assign n11213 = n196 | n1106 ;
  assign n11214 = n1631 & ~n11213 ;
  assign n11215 = n1349 & ~n11214 ;
  assign n11216 = n11215 ^ n6519 ^ 1'b0 ;
  assign n11219 = n1747 ^ n1137 ^ 1'b0 ;
  assign n11220 = n179 & n11219 ;
  assign n11217 = n373 | n1525 ;
  assign n11218 = n11217 ^ n7203 ^ 1'b0 ;
  assign n11221 = n11220 ^ n11218 ^ 1'b0 ;
  assign n11222 = n11216 & n11221 ;
  assign n11223 = n3672 ^ n3354 ^ 1'b0 ;
  assign n11224 = n2858 ^ n359 ^ 1'b0 ;
  assign n11225 = n356 & n11224 ;
  assign n11226 = ( n1601 & ~n5451 ) | ( n1601 & n11225 ) | ( ~n5451 & n11225 ) ;
  assign n11231 = n7401 ^ x84 ^ 1'b0 ;
  assign n11230 = n4679 | n6358 ;
  assign n11232 = n11231 ^ n11230 ^ 1'b0 ;
  assign n11227 = n6770 ^ n4029 ^ 1'b0 ;
  assign n11228 = n11227 ^ n4636 ^ 1'b0 ;
  assign n11229 = ~n911 & n11228 ;
  assign n11233 = n11232 ^ n11229 ^ 1'b0 ;
  assign n11235 = n8821 ^ n733 ^ 1'b0 ;
  assign n11234 = n4364 | n10026 ;
  assign n11236 = n11235 ^ n11234 ^ 1'b0 ;
  assign n11237 = n1586 | n5596 ;
  assign n11239 = n4279 ^ n1489 ^ 1'b0 ;
  assign n11240 = n5087 & ~n11239 ;
  assign n11238 = n5663 & n6094 ;
  assign n11241 = n11240 ^ n11238 ^ 1'b0 ;
  assign n11242 = n3740 ^ n2064 ^ n1868 ;
  assign n11243 = n11242 ^ n7349 ^ 1'b0 ;
  assign n11244 = n8977 ^ n519 ^ 1'b0 ;
  assign n11245 = n4846 & ~n4985 ;
  assign n11246 = n5019 ^ n985 ^ 1'b0 ;
  assign n11247 = n11245 | n11246 ;
  assign n11248 = n5413 & ~n11238 ;
  assign n11253 = ~n1673 & n3224 ;
  assign n11249 = n4853 ^ n519 ^ 1'b0 ;
  assign n11250 = n221 & ~n482 ;
  assign n11251 = ~n7044 & n11250 ;
  assign n11252 = ( n4310 & ~n11249 ) | ( n4310 & n11251 ) | ( ~n11249 & n11251 ) ;
  assign n11254 = n11253 ^ n11252 ^ n9093 ;
  assign n11257 = n1139 ^ n806 ^ 1'b0 ;
  assign n11258 = ~n1832 & n11257 ;
  assign n11255 = n1909 & n9072 ;
  assign n11256 = n1689 | n11255 ;
  assign n11259 = n11258 ^ n11256 ^ 1'b0 ;
  assign n11260 = n3956 & n7878 ;
  assign n11261 = ~n555 & n2385 ;
  assign n11262 = n8232 & n11261 ;
  assign n11263 = n11262 ^ n6644 ^ 1'b0 ;
  assign n11264 = n8749 ^ n6809 ^ 1'b0 ;
  assign n11265 = n790 & n11264 ;
  assign n11266 = ~n11263 & n11265 ;
  assign n11267 = n877 | n5720 ;
  assign n11268 = n11267 ^ n3268 ^ 1'b0 ;
  assign n11269 = x51 ^ x11 ^ 1'b0 ;
  assign n11270 = n8319 ^ n8024 ^ 1'b0 ;
  assign n11271 = n11269 | n11270 ;
  assign n11272 = n1409 ^ n1403 ^ n131 ;
  assign n11273 = n11272 ^ n6736 ^ 1'b0 ;
  assign n11274 = n4517 & n6781 ;
  assign n11275 = n11274 ^ n221 ^ 1'b0 ;
  assign n11276 = n2136 ^ n1479 ^ 1'b0 ;
  assign n11277 = n1374 & ~n11276 ;
  assign n11278 = n3599 & ~n11277 ;
  assign n11279 = ~x107 & n11278 ;
  assign n11280 = n3809 & ~n9713 ;
  assign n11281 = n3474 & n4676 ;
  assign n11282 = n733 & n11281 ;
  assign n11283 = n3189 & n11282 ;
  assign n11284 = n4701 ^ n2313 ^ 1'b0 ;
  assign n11285 = n5418 & ~n7617 ;
  assign n11286 = n5105 & n11285 ;
  assign n11287 = n2967 & ~n7498 ;
  assign n11288 = n4645 & n11287 ;
  assign n11289 = n539 | n11288 ;
  assign n11290 = n1634 | n11289 ;
  assign n11291 = n7180 ^ n5935 ^ 1'b0 ;
  assign n11292 = ~n566 & n731 ;
  assign n11293 = n1013 & n11292 ;
  assign n11294 = n189 & ~n11293 ;
  assign n11295 = n11294 ^ n3067 ^ 1'b0 ;
  assign n11296 = n11295 ^ n5327 ^ n2930 ;
  assign n11297 = n11293 ^ n1572 ^ 1'b0 ;
  assign n11298 = n1993 & n11297 ;
  assign n11299 = n6378 ^ n5859 ^ 1'b0 ;
  assign n11300 = n4300 | n11299 ;
  assign n11301 = n1777 ^ n1351 ^ 1'b0 ;
  assign n11302 = n11301 ^ n8249 ^ 1'b0 ;
  assign n11303 = n8021 & n11302 ;
  assign n11304 = n4648 ^ n3772 ^ 1'b0 ;
  assign n11305 = n11220 & n11304 ;
  assign n11306 = x28 & ~n9818 ;
  assign n11307 = ~n3734 & n11306 ;
  assign n11308 = n1833 & n3847 ;
  assign n11309 = n894 & n11308 ;
  assign n11310 = n11309 ^ n3793 ^ 1'b0 ;
  assign n11311 = n7543 ^ n528 ^ 1'b0 ;
  assign n11312 = n11310 & ~n11311 ;
  assign n11313 = n10931 ^ n6494 ^ 1'b0 ;
  assign n11314 = n4093 & n11313 ;
  assign n11315 = n811 | n6037 ;
  assign n11316 = ~n5719 & n10015 ;
  assign n11317 = n2649 ^ n2458 ^ 1'b0 ;
  assign n11318 = n3956 | n11317 ;
  assign n11319 = n2884 & n11318 ;
  assign n11322 = n7605 ^ n5254 ^ n2260 ;
  assign n11323 = n6679 | n11322 ;
  assign n11320 = n5429 & n6585 ;
  assign n11321 = n8535 | n11320 ;
  assign n11324 = n11323 ^ n11321 ^ 1'b0 ;
  assign n11325 = n10295 ^ n6519 ^ 1'b0 ;
  assign n11326 = n808 & n5842 ;
  assign n11327 = n11326 ^ n6606 ^ 1'b0 ;
  assign n11329 = n2656 & n11274 ;
  assign n11330 = ( n243 & n568 ) | ( n243 & ~n11329 ) | ( n568 & ~n11329 ) ;
  assign n11328 = n876 & ~n5059 ;
  assign n11331 = n11330 ^ n11328 ^ 1'b0 ;
  assign n11332 = ~n3688 & n5721 ;
  assign n11333 = n1540 | n3195 ;
  assign n11334 = n4234 & ~n11333 ;
  assign n11335 = n11334 ^ n5312 ^ 1'b0 ;
  assign n11336 = n1049 | n11335 ;
  assign n11337 = n1386 | n11336 ;
  assign n11338 = ~n1087 & n11337 ;
  assign n11339 = n11338 ^ n1203 ^ 1'b0 ;
  assign n11340 = ~n2144 & n4459 ;
  assign n11341 = n11340 ^ n3192 ^ 1'b0 ;
  assign n11342 = n2887 | n11089 ;
  assign n11343 = n6408 ^ n1260 ^ 1'b0 ;
  assign n11344 = n757 | n11343 ;
  assign n11345 = n10232 & ~n11344 ;
  assign n11346 = n11345 ^ n1302 ^ 1'b0 ;
  assign n11347 = n4398 ^ n2702 ^ 1'b0 ;
  assign n11348 = n1122 & ~n4627 ;
  assign n11349 = n11348 ^ n4410 ^ 1'b0 ;
  assign n11350 = n5341 ^ n4404 ^ 1'b0 ;
  assign n11351 = n11350 ^ n5959 ^ n3853 ;
  assign n11352 = ( n4244 & ~n5642 ) | ( n4244 & n8737 ) | ( ~n5642 & n8737 ) ;
  assign n11353 = ~n10312 & n11352 ;
  assign n11354 = n1812 & n11353 ;
  assign n11355 = n5744 & n5862 ;
  assign n11356 = n5907 ^ n531 ^ 1'b0 ;
  assign n11357 = n8064 ^ n1526 ^ 1'b0 ;
  assign n11358 = ~n1053 & n5708 ;
  assign n11359 = n8371 ^ n5004 ^ 1'b0 ;
  assign n11360 = n10129 & ~n11359 ;
  assign n11361 = n1015 | n5380 ;
  assign n11362 = n6640 & ~n11361 ;
  assign n11363 = n8035 ^ n4673 ^ n2694 ;
  assign n11365 = n4871 | n5863 ;
  assign n11364 = n934 & n2115 ;
  assign n11366 = n11365 ^ n11364 ^ 1'b0 ;
  assign n11367 = ~n5487 & n11366 ;
  assign n11368 = n9181 ^ n3494 ^ 1'b0 ;
  assign n11369 = n5985 & n8095 ;
  assign n11370 = n6994 ^ n361 ^ 1'b0 ;
  assign n11371 = n1909 & ~n11370 ;
  assign n11372 = n10691 | n11371 ;
  assign n11373 = n1918 & ~n8511 ;
  assign n11374 = n10152 ^ n3073 ^ n305 ;
  assign n11375 = ~n996 & n1880 ;
  assign n11376 = ~n1056 & n2614 ;
  assign n11377 = n8535 ^ n5564 ^ 1'b0 ;
  assign n11378 = n11376 & ~n11377 ;
  assign n11379 = n413 | n1487 ;
  assign n11380 = n962 | n11379 ;
  assign n11381 = ~n11163 & n11380 ;
  assign n11382 = ~n420 & n11381 ;
  assign n11383 = n6792 & ~n8937 ;
  assign n11384 = n11382 & n11383 ;
  assign n11385 = ~n6333 & n7614 ;
  assign n11386 = n5431 ^ n1858 ^ 1'b0 ;
  assign n11387 = n5393 & n11386 ;
  assign n11388 = n11387 ^ n335 ^ 1'b0 ;
  assign n11389 = n1521 & n11388 ;
  assign n11390 = ~n4692 & n10391 ;
  assign n11391 = n1982 & n11390 ;
  assign n11392 = n9234 ^ n2123 ^ 1'b0 ;
  assign n11393 = n1205 & ~n1561 ;
  assign n11394 = n782 ^ x98 ^ 1'b0 ;
  assign n11395 = n5736 ^ n4532 ^ 1'b0 ;
  assign n11396 = n11394 & n11395 ;
  assign n11397 = n6756 ^ n4681 ^ 1'b0 ;
  assign n11398 = n831 & ~n11397 ;
  assign n11399 = n11398 ^ n9662 ^ 1'b0 ;
  assign n11400 = n1815 | n11399 ;
  assign n11401 = n6965 ^ n4387 ^ 1'b0 ;
  assign n11402 = n3076 & n11401 ;
  assign n11403 = n6030 ^ n5146 ^ 1'b0 ;
  assign n11404 = n11402 | n11403 ;
  assign n11405 = n886 & n3070 ;
  assign n11406 = n11405 ^ n7784 ^ 1'b0 ;
  assign n11407 = n2978 & ~n3120 ;
  assign n11408 = n8713 & ~n11407 ;
  assign n11409 = n343 & n11408 ;
  assign n11410 = n6420 & ~n9459 ;
  assign n11411 = n11410 ^ n7019 ^ 1'b0 ;
  assign n11412 = n10568 | n11411 ;
  assign n11413 = n220 & ~n1232 ;
  assign n11414 = n11413 ^ n1540 ^ 1'b0 ;
  assign n11415 = n11414 ^ n2885 ^ 1'b0 ;
  assign n11416 = n4569 & n5735 ;
  assign n11417 = n11416 ^ n7460 ^ 1'b0 ;
  assign n11418 = n11417 ^ n6212 ^ n5940 ;
  assign n11419 = n1983 ^ n938 ^ 1'b0 ;
  assign n11420 = n5097 | n11419 ;
  assign n11421 = n6499 & ~n11420 ;
  assign n11422 = n330 & n9573 ;
  assign n11423 = n5222 & n11422 ;
  assign n11424 = ~n7543 & n11423 ;
  assign n11425 = n11424 ^ n10043 ^ 1'b0 ;
  assign n11426 = ~n9673 & n11425 ;
  assign n11427 = n7416 | n11426 ;
  assign n11428 = n529 | n11427 ;
  assign n11429 = n4558 & n7244 ;
  assign n11430 = ~n11428 & n11429 ;
  assign n11431 = n11430 ^ n3083 ^ 1'b0 ;
  assign n11432 = ~n11421 & n11431 ;
  assign n11433 = n6406 ^ n4384 ^ 1'b0 ;
  assign n11434 = n11433 ^ n3784 ^ 1'b0 ;
  assign n11435 = n1194 | n11434 ;
  assign n11436 = n6458 ^ n2358 ^ 1'b0 ;
  assign n11437 = n689 & n1759 ;
  assign n11438 = n6330 & ~n11334 ;
  assign n11439 = n3066 & ~n3135 ;
  assign n11440 = n8861 & n11439 ;
  assign n11443 = n287 | n4443 ;
  assign n11441 = n5525 & n6240 ;
  assign n11442 = n11441 ^ n1812 ^ 1'b0 ;
  assign n11444 = n11443 ^ n11442 ^ n428 ;
  assign n11445 = n2481 & ~n2828 ;
  assign n11446 = n9009 & ~n11445 ;
  assign n11447 = n1409 & ~n2533 ;
  assign n11448 = n2533 & n11447 ;
  assign n11449 = n1334 & ~n11448 ;
  assign n11450 = ~n1334 & n11449 ;
  assign n11451 = n159 & n11450 ;
  assign n11452 = n11451 ^ n8335 ^ 1'b0 ;
  assign n11453 = n786 | n4384 ;
  assign n11454 = n786 & ~n11453 ;
  assign n11455 = n8942 & ~n11454 ;
  assign n11456 = ~n8942 & n11455 ;
  assign n11457 = n11452 | n11456 ;
  assign n11458 = n11452 & ~n11457 ;
  assign n11459 = n4976 | n6979 ;
  assign n11460 = n11285 & ~n11459 ;
  assign n11461 = n11460 ^ n2119 ^ 1'b0 ;
  assign n11462 = n5274 ^ n2028 ^ 1'b0 ;
  assign n11463 = n911 | n11462 ;
  assign n11464 = n6149 & ~n11463 ;
  assign n11465 = n8365 | n11464 ;
  assign n11466 = n11465 ^ n9928 ^ 1'b0 ;
  assign n11467 = n6832 ^ n5680 ^ 1'b0 ;
  assign n11468 = n11467 ^ n7411 ^ n457 ;
  assign n11469 = ~n300 & n9302 ;
  assign n11470 = ~n4996 & n10980 ;
  assign n11471 = n378 & n11470 ;
  assign n11472 = n9133 ^ n4804 ^ n4041 ;
  assign n11473 = ~n259 & n6645 ;
  assign n11474 = n11473 ^ n5434 ^ 1'b0 ;
  assign n11475 = n225 | n1107 ;
  assign n11476 = n11475 ^ n2328 ^ 1'b0 ;
  assign n11477 = n3958 & n11476 ;
  assign n11478 = n8942 & n11477 ;
  assign n11479 = n707 & n11478 ;
  assign n11480 = n11479 ^ n10238 ^ 1'b0 ;
  assign n11481 = ~n11474 & n11480 ;
  assign n11482 = n2112 | n11481 ;
  assign n11483 = n876 & n3358 ;
  assign n11484 = ~n1539 & n11483 ;
  assign n11485 = n3339 | n11484 ;
  assign n11486 = n3283 | n11485 ;
  assign n11487 = ~n7110 & n11486 ;
  assign n11488 = n11487 ^ n8258 ^ 1'b0 ;
  assign n11489 = n1602 & n11488 ;
  assign n11490 = n3353 & n10391 ;
  assign n11491 = n9286 & n11490 ;
  assign n11492 = n1304 & ~n7352 ;
  assign n11493 = n7352 & n11492 ;
  assign n11494 = n639 & n1905 ;
  assign n11495 = n11493 & n11494 ;
  assign n11496 = n2245 & ~n3947 ;
  assign n11497 = ~n7226 & n11496 ;
  assign n11498 = ( n863 & ~n11495 ) | ( n863 & n11497 ) | ( ~n11495 & n11497 ) ;
  assign n11499 = n1827 & ~n6982 ;
  assign n11500 = n5052 & n11499 ;
  assign n11501 = n11500 ^ n9205 ^ 1'b0 ;
  assign n11502 = x58 & x77 ;
  assign n11503 = n11502 ^ n6219 ^ 1'b0 ;
  assign n11504 = n2232 ^ n866 ^ 1'b0 ;
  assign n11505 = n3974 & ~n11504 ;
  assign n11506 = ~n3403 & n11505 ;
  assign n11507 = n11506 ^ n5488 ^ 1'b0 ;
  assign n11508 = n1571 & ~n7432 ;
  assign n11509 = n830 ^ n268 ^ 1'b0 ;
  assign n11510 = ~n677 & n11509 ;
  assign n11511 = n1618 & ~n11510 ;
  assign n11512 = n8179 ^ x88 ^ 1'b0 ;
  assign n11513 = n11512 ^ n2662 ^ 1'b0 ;
  assign n11515 = x111 & ~n4180 ;
  assign n11514 = n1927 | n4280 ;
  assign n11516 = n11515 ^ n11514 ^ 1'b0 ;
  assign n11517 = n2883 | n11516 ;
  assign n11518 = n6801 ^ n4736 ^ 1'b0 ;
  assign n11519 = n436 & ~n11518 ;
  assign n11520 = n5924 ^ n870 ^ 1'b0 ;
  assign n11521 = n9604 ^ n3019 ^ 1'b0 ;
  assign n11522 = n2115 & ~n11521 ;
  assign n11523 = n10969 ^ n7383 ^ 1'b0 ;
  assign n11530 = x68 & ~n1588 ;
  assign n11531 = ~n9948 & n11530 ;
  assign n11532 = ~n2636 & n3105 ;
  assign n11533 = ~n2090 & n11532 ;
  assign n11534 = ~n11531 & n11533 ;
  assign n11535 = n4579 & n11534 ;
  assign n11524 = n7139 ^ n825 ^ 1'b0 ;
  assign n11525 = n1240 & ~n11524 ;
  assign n11526 = x13 & ~n2839 ;
  assign n11527 = ~n8420 & n11526 ;
  assign n11528 = n11527 ^ n7262 ^ 1'b0 ;
  assign n11529 = n11525 & ~n11528 ;
  assign n11536 = n11535 ^ n11529 ^ 1'b0 ;
  assign n11537 = n1273 & ~n11536 ;
  assign n11538 = n10975 ^ n5661 ^ x75 ;
  assign n11539 = n11538 ^ n9679 ^ 1'b0 ;
  assign n11540 = n785 | n7816 ;
  assign n11541 = n11540 ^ n6536 ^ 1'b0 ;
  assign n11542 = n6975 ^ n5613 ^ 1'b0 ;
  assign n11543 = n2123 ^ n1620 ^ 1'b0 ;
  assign n11544 = n277 & n8247 ;
  assign n11545 = ~n8282 & n11544 ;
  assign n11546 = ( n512 & n6069 ) | ( n512 & ~n11545 ) | ( n6069 & ~n11545 ) ;
  assign n11547 = n10688 ^ n7341 ^ 1'b0 ;
  assign n11548 = n4388 & n4631 ;
  assign n11549 = n9818 ^ n5364 ^ 1'b0 ;
  assign n11550 = ~n2516 & n11549 ;
  assign n11551 = n3678 | n5989 ;
  assign n11552 = n10438 ^ n6352 ^ 1'b0 ;
  assign n11553 = n11551 | n11552 ;
  assign n11554 = n2759 | n9244 ;
  assign n11555 = n8161 | n11554 ;
  assign n11556 = ~n5152 & n11555 ;
  assign n11557 = n1864 & ~n2398 ;
  assign n11558 = n1548 & n4666 ;
  assign n11559 = n11558 ^ n8811 ^ n5144 ;
  assign n11560 = n9760 & n10696 ;
  assign n11561 = ~n1551 & n7116 ;
  assign n11562 = n2604 & n6844 ;
  assign n11563 = n4638 & n11562 ;
  assign n11564 = n11563 ^ n11346 ^ 1'b0 ;
  assign n11565 = ~n1153 & n1328 ;
  assign n11566 = n11565 ^ n4462 ^ 1'b0 ;
  assign n11567 = n6880 ^ n3925 ^ 1'b0 ;
  assign n11568 = n5461 & ~n11567 ;
  assign n11569 = n11568 ^ n8769 ^ 1'b0 ;
  assign n11570 = n7963 & ~n11569 ;
  assign n11572 = n2948 ^ n2310 ^ 1'b0 ;
  assign n11573 = ~n8016 & n11572 ;
  assign n11574 = n11573 ^ n3776 ^ 1'b0 ;
  assign n11575 = n1209 & n11574 ;
  assign n11571 = n137 & ~n397 ;
  assign n11576 = n11575 ^ n11571 ^ 1'b0 ;
  assign n11577 = ( n1574 & ~n2073 ) | ( n1574 & n9823 ) | ( ~n2073 & n9823 ) ;
  assign n11578 = n7547 & ~n8874 ;
  assign n11579 = n11578 ^ n10040 ^ 1'b0 ;
  assign n11580 = n11579 ^ n6480 ^ 1'b0 ;
  assign n11581 = n6837 & n7502 ;
  assign n11582 = n11581 ^ n9562 ^ 1'b0 ;
  assign n11583 = n3789 | n9074 ;
  assign n11584 = n11583 ^ n1980 ^ 1'b0 ;
  assign n11585 = ~n1574 & n10466 ;
  assign n11586 = n11585 ^ n250 ^ 1'b0 ;
  assign n11587 = ~n667 & n2800 ;
  assign n11588 = n3740 ^ n2260 ^ 1'b0 ;
  assign n11589 = n696 | n2673 ;
  assign n11590 = x22 & ~n11240 ;
  assign n11596 = n4240 ^ n2013 ^ 1'b0 ;
  assign n11597 = n456 & ~n11596 ;
  assign n11591 = n1733 ^ n213 ^ 1'b0 ;
  assign n11592 = n4287 & n11591 ;
  assign n11593 = n3336 | n3482 ;
  assign n11594 = n11592 | n11593 ;
  assign n11595 = n11594 ^ n1270 ^ 1'b0 ;
  assign n11598 = n11597 ^ n11595 ^ 1'b0 ;
  assign n11599 = n9343 ^ n6821 ^ 1'b0 ;
  assign n11600 = n600 ^ x109 ^ 1'b0 ;
  assign n11601 = n538 & ~n11600 ;
  assign n11602 = ~n2898 & n11601 ;
  assign n11603 = n11602 ^ n5885 ^ 1'b0 ;
  assign n11604 = n5230 & n6961 ;
  assign n11605 = n11604 ^ n11334 ^ 1'b0 ;
  assign n11606 = n3076 & n6362 ;
  assign n11607 = n11606 ^ n6018 ^ 1'b0 ;
  assign n11608 = n2738 & n11607 ;
  assign n11609 = n2367 ^ x37 ^ 1'b0 ;
  assign n11610 = n874 ^ x87 ^ 1'b0 ;
  assign n11611 = n4578 & n11610 ;
  assign n11612 = n8496 & n11611 ;
  assign n11613 = n5747 & n11612 ;
  assign n11614 = n2481 & ~n11613 ;
  assign n11615 = n5977 & ~n11241 ;
  assign n11616 = n9217 ^ n6881 ^ 1'b0 ;
  assign n11620 = n8787 | n9897 ;
  assign n11621 = n11620 ^ n3678 ^ 1'b0 ;
  assign n11617 = n1124 & ~n8760 ;
  assign n11618 = n11617 ^ n6274 ^ n3018 ;
  assign n11619 = n6546 & ~n11618 ;
  assign n11622 = n11621 ^ n11619 ^ 1'b0 ;
  assign n11624 = n5148 ^ n1444 ^ 1'b0 ;
  assign n11623 = n9719 ^ n8512 ^ 1'b0 ;
  assign n11625 = n11624 ^ n11623 ^ 1'b0 ;
  assign n11626 = n8496 & n11625 ;
  assign n11627 = n456 & ~n1540 ;
  assign n11628 = n2165 & n11627 ;
  assign n11629 = ~n1128 & n10880 ;
  assign n11630 = ~n2618 & n11629 ;
  assign n11631 = n1277 ^ x109 ^ 1'b0 ;
  assign n11632 = n1668 & ~n11631 ;
  assign n11633 = n11632 ^ n7681 ^ 1'b0 ;
  assign n11634 = n3673 & n11633 ;
  assign n11635 = n6511 ^ n1656 ^ 1'b0 ;
  assign n11636 = n2721 & n7755 ;
  assign n11637 = n9045 & ~n11392 ;
  assign n11638 = n7715 ^ n328 ^ 1'b0 ;
  assign n11639 = n1321 & n2468 ;
  assign n11640 = ~n11638 & n11639 ;
  assign n11649 = n7068 | n11240 ;
  assign n11647 = n3073 & n3760 ;
  assign n11643 = n724 & n1628 ;
  assign n11644 = n11643 ^ n1042 ^ 1'b0 ;
  assign n11645 = n3554 | n11644 ;
  assign n11646 = ~n3366 & n11645 ;
  assign n11641 = n4600 & n9691 ;
  assign n11642 = n11641 ^ x88 ^ 1'b0 ;
  assign n11648 = n11647 ^ n11646 ^ n11642 ;
  assign n11650 = n11649 ^ n11648 ^ 1'b0 ;
  assign n11651 = n11640 | n11650 ;
  assign n11652 = n8363 & ~n11651 ;
  assign n11653 = n2481 & ~n9417 ;
  assign n11654 = n2709 | n6777 ;
  assign n11658 = n256 & ~n404 ;
  assign n11659 = n11658 ^ n2182 ^ 1'b0 ;
  assign n11655 = n778 | n2892 ;
  assign n11656 = n5224 | n11655 ;
  assign n11657 = ~n5019 & n11656 ;
  assign n11660 = n11659 ^ n11657 ^ 1'b0 ;
  assign n11661 = n1334 & ~n11660 ;
  assign n11662 = n2222 & ~n11597 ;
  assign n11663 = n10572 & n11662 ;
  assign n11664 = n571 & ~n2414 ;
  assign n11665 = n11664 ^ n638 ^ 1'b0 ;
  assign n11666 = ~n3453 & n11665 ;
  assign n11667 = ( x104 & n2818 ) | ( x104 & ~n11666 ) | ( n2818 & ~n11666 ) ;
  assign n11668 = n11667 ^ n8256 ^ 1'b0 ;
  assign n11669 = n5606 ^ n5000 ^ 1'b0 ;
  assign n11670 = x3 & ~n876 ;
  assign n11671 = n967 | n11670 ;
  assign n11672 = n11671 ^ n2584 ^ 1'b0 ;
  assign n11673 = n11672 ^ n1695 ^ 1'b0 ;
  assign n11674 = n1312 | n6934 ;
  assign n11675 = n5871 ^ n3717 ^ 1'b0 ;
  assign n11676 = n529 & ~n11675 ;
  assign n11677 = n11676 ^ n3271 ^ 1'b0 ;
  assign n11678 = n11677 ^ n10352 ^ n7688 ;
  assign n11679 = ~n4706 & n9512 ;
  assign n11680 = ~n6901 & n11679 ;
  assign n11681 = n11680 ^ n5907 ^ 1'b0 ;
  assign n11682 = n283 & ~n11681 ;
  assign n11683 = ~n5705 & n11682 ;
  assign n11684 = n1734 | n5953 ;
  assign n11685 = ~n1574 & n3038 ;
  assign n11686 = n6699 & n11685 ;
  assign n11687 = n6219 | n8384 ;
  assign n11688 = n3267 & ~n11687 ;
  assign n11689 = n1578 | n11688 ;
  assign n11690 = n5749 & ~n11689 ;
  assign n11691 = n11690 ^ n6325 ^ n1279 ;
  assign n11692 = n2660 & n3362 ;
  assign n11693 = n11692 ^ n2687 ^ 1'b0 ;
  assign n11694 = n822 & ~n6362 ;
  assign n11695 = n11694 ^ x46 ^ 1'b0 ;
  assign n11696 = n11693 | n11695 ;
  assign n11697 = n4692 ^ n2456 ^ 1'b0 ;
  assign n11698 = ~n4683 & n11697 ;
  assign n11699 = n8877 ^ n8848 ^ 1'b0 ;
  assign n11700 = ~n6266 & n11699 ;
  assign n11701 = n1693 & ~n1841 ;
  assign n11702 = n297 & n5466 ;
  assign n11703 = n11702 ^ n3032 ^ 1'b0 ;
  assign n11704 = ~n548 & n3403 ;
  assign n11705 = n2256 & ~n3518 ;
  assign n11706 = n7223 & ~n10017 ;
  assign n11707 = n6766 & ~n11706 ;
  assign n11708 = n1663 | n3840 ;
  assign n11709 = n2505 | n11708 ;
  assign n11710 = n4647 & ~n8628 ;
  assign n11711 = ( n10791 & n11709 ) | ( n10791 & ~n11710 ) | ( n11709 & ~n11710 ) ;
  assign n11712 = n2813 & n4494 ;
  assign n11713 = n7835 ^ n6188 ^ 1'b0 ;
  assign n11714 = n1957 ^ n1908 ^ 1'b0 ;
  assign n11715 = n11714 ^ n3078 ^ 1'b0 ;
  assign n11716 = n4434 ^ n595 ^ 1'b0 ;
  assign n11717 = n9729 & n11716 ;
  assign n11718 = x122 & ~n270 ;
  assign n11719 = n3420 & ~n11718 ;
  assign n11720 = n11719 ^ n10602 ^ 1'b0 ;
  assign n11722 = n1849 ^ n333 ^ 1'b0 ;
  assign n11721 = n4215 & n7644 ;
  assign n11723 = n11722 ^ n11721 ^ 1'b0 ;
  assign n11725 = ~n512 & n10562 ;
  assign n11724 = n3875 | n5664 ;
  assign n11726 = n11725 ^ n11724 ^ 1'b0 ;
  assign n11727 = n422 & ~n571 ;
  assign n11728 = n571 & n11727 ;
  assign n11729 = n11728 ^ n1049 ^ 1'b0 ;
  assign n11730 = n2729 & ~n11729 ;
  assign n11731 = ~n2729 & n11730 ;
  assign n11732 = n134 | n10787 ;
  assign n11733 = x17 & n11666 ;
  assign n11734 = n1547 & n8821 ;
  assign n11735 = x62 & n11734 ;
  assign n11736 = n8946 & ~n11735 ;
  assign n11737 = ~n620 & n11736 ;
  assign n11738 = n2091 & n6671 ;
  assign n11739 = n6985 & n11738 ;
  assign n11740 = n4493 & ~n9357 ;
  assign n11741 = ~n3826 & n5318 ;
  assign n11742 = ~n4095 & n8340 ;
  assign n11743 = n4095 & n11742 ;
  assign n11744 = n5648 ^ n1515 ^ n835 ;
  assign n11745 = n11407 ^ n7015 ^ 1'b0 ;
  assign n11746 = n4380 | n11745 ;
  assign n11747 = ~n1666 & n4198 ;
  assign n11748 = n1534 & ~n1789 ;
  assign n11749 = ~n11747 & n11748 ;
  assign n11750 = n11749 ^ n2136 ^ 1'b0 ;
  assign n11753 = n1768 | n2987 ;
  assign n11754 = n1768 & ~n11753 ;
  assign n11752 = n3388 & ~n3774 ;
  assign n11755 = n11754 ^ n11752 ^ 1'b0 ;
  assign n11751 = ~n2817 & n3359 ;
  assign n11756 = n11755 ^ n11751 ^ 1'b0 ;
  assign n11757 = n724 & n8905 ;
  assign n11758 = ~n2604 & n11757 ;
  assign n11759 = n11569 ^ n9459 ^ 1'b0 ;
  assign n11760 = x57 & n5477 ;
  assign n11761 = n2340 & n11760 ;
  assign n11762 = n1476 ^ n315 ^ 1'b0 ;
  assign n11763 = n776 & n4173 ;
  assign n11764 = n5927 | n9632 ;
  assign n11765 = n11764 ^ n1951 ^ 1'b0 ;
  assign n11766 = n11765 ^ n8511 ^ 1'b0 ;
  assign n11767 = n9868 | n11766 ;
  assign n11768 = n834 | n1129 ;
  assign n11769 = n672 | n11768 ;
  assign n11770 = n11769 ^ n5981 ^ 1'b0 ;
  assign n11771 = ~n2122 & n4606 ;
  assign n11772 = n2969 | n3862 ;
  assign n11773 = n11772 ^ n6890 ^ 1'b0 ;
  assign n11774 = n11773 ^ n1053 ^ 1'b0 ;
  assign n11775 = n10848 ^ n3731 ^ 1'b0 ;
  assign n11776 = n9267 ^ n4067 ^ 1'b0 ;
  assign n11777 = n7481 & ~n11776 ;
  assign n11778 = n3393 | n9766 ;
  assign n11779 = n7211 ^ n5182 ^ 1'b0 ;
  assign n11780 = n1416 | n6842 ;
  assign n11781 = ~n809 & n6883 ;
  assign n11782 = n11781 ^ n392 ^ 1'b0 ;
  assign n11783 = n1714 ^ n1335 ^ 1'b0 ;
  assign n11784 = ~n8874 & n11783 ;
  assign n11785 = n3347 & n10147 ;
  assign n11786 = ~n6427 & n11785 ;
  assign n11787 = n5298 ^ n4749 ^ 1'b0 ;
  assign n11788 = n2667 | n11787 ;
  assign n11789 = n1945 | n4153 ;
  assign n11790 = n4153 & ~n11789 ;
  assign n11791 = n1089 | n3352 ;
  assign n11792 = ~n2608 & n11791 ;
  assign n11793 = n1907 & ~n3116 ;
  assign n11794 = n11793 ^ n6910 ^ 1'b0 ;
  assign n11795 = ~n1093 & n5713 ;
  assign n11796 = n1556 | n1759 ;
  assign n11797 = n11796 ^ n7272 ^ 1'b0 ;
  assign n11798 = ~x22 & n10795 ;
  assign n11799 = n5967 ^ n2868 ^ 1'b0 ;
  assign n11800 = n4128 | n10932 ;
  assign n11801 = n11800 ^ n4655 ^ 1'b0 ;
  assign n11802 = n6589 & n11801 ;
  assign n11803 = n8220 ^ n2420 ^ 1'b0 ;
  assign n11804 = n9431 & n11803 ;
  assign n11805 = n1905 ^ n227 ^ 1'b0 ;
  assign n11806 = n4880 ^ n1831 ^ 1'b0 ;
  assign n11807 = ~n11805 & n11806 ;
  assign n11808 = n7141 ^ n1909 ^ 1'b0 ;
  assign n11809 = n11808 ^ n11503 ^ 1'b0 ;
  assign n11810 = n1981 | n5868 ;
  assign n11811 = n11586 ^ n6634 ^ n448 ;
  assign n11812 = n3266 & n8984 ;
  assign n11813 = n10587 & n11812 ;
  assign n11814 = n7295 ^ n6985 ^ 1'b0 ;
  assign n11815 = x127 | n287 ;
  assign n11816 = ( n5417 & ~n6175 ) | ( n5417 & n6832 ) | ( ~n6175 & n6832 ) ;
  assign n11817 = n5054 ^ n741 ^ 1'b0 ;
  assign n11818 = n11412 & ~n11817 ;
  assign n11819 = n802 & n2241 ;
  assign n11820 = n839 & n6528 ;
  assign n11821 = n9793 & n11820 ;
  assign n11822 = n11821 ^ n7172 ^ 1'b0 ;
  assign n11823 = n9418 & n11822 ;
  assign n11824 = n4530 ^ n1227 ^ 1'b0 ;
  assign n11826 = n4230 ^ n2253 ^ 1'b0 ;
  assign n11825 = n1875 | n5349 ;
  assign n11827 = n11826 ^ n11825 ^ 1'b0 ;
  assign n11828 = n11827 ^ n5907 ^ n1991 ;
  assign n11829 = ~n926 & n5642 ;
  assign n11830 = n2975 & ~n7855 ;
  assign n11831 = n11830 ^ x29 ^ 1'b0 ;
  assign n11832 = n4034 & ~n8651 ;
  assign n11833 = n11832 ^ n10846 ^ 1'b0 ;
  assign n11834 = n2726 | n3572 ;
  assign n11835 = n11277 ^ n7679 ^ 1'b0 ;
  assign n11836 = n11834 | n11835 ;
  assign n11837 = n2440 ^ n231 ^ 1'b0 ;
  assign n11838 = n5152 ^ n4153 ^ 1'b0 ;
  assign n11839 = n11838 ^ n5242 ^ 1'b0 ;
  assign n11840 = n7606 & n11839 ;
  assign n11841 = n1880 & n3866 ;
  assign n11842 = n9687 & n11841 ;
  assign n11843 = ~n4900 & n11842 ;
  assign n11844 = n4933 | n10978 ;
  assign n11845 = n1782 ^ n1637 ^ 1'b0 ;
  assign n11846 = n830 & n11845 ;
  assign n11847 = n11823 & n11846 ;
  assign n11848 = n11847 ^ n2828 ^ 1'b0 ;
  assign n11850 = n690 ^ x100 ^ 1'b0 ;
  assign n11849 = n1116 & n5475 ;
  assign n11851 = n11850 ^ n11849 ^ 1'b0 ;
  assign n11852 = ~n1669 & n3998 ;
  assign n11853 = n11852 ^ n8742 ^ 1'b0 ;
  assign n11854 = n4043 & ~n11853 ;
  assign n11855 = n3956 ^ n2321 ^ 1'b0 ;
  assign n11856 = n7276 | n11855 ;
  assign n11857 = n6214 & n11856 ;
  assign n11858 = ~n6565 & n9323 ;
  assign n11859 = n2630 | n8163 ;
  assign n11860 = n2697 & n5821 ;
  assign n11861 = n11859 & n11860 ;
  assign n11862 = n1890 & n5739 ;
  assign n11863 = n7057 & n7626 ;
  assign n11864 = ~n3169 & n10630 ;
  assign n11865 = n4731 ^ n1724 ^ 1'b0 ;
  assign n11866 = n956 ^ n529 ^ 1'b0 ;
  assign n11867 = n8390 ^ n4133 ^ 1'b0 ;
  assign n11868 = n3480 & n11867 ;
  assign n11871 = n4558 ^ n2337 ^ 1'b0 ;
  assign n11872 = n722 & n11871 ;
  assign n11873 = ~n344 & n11872 ;
  assign n11870 = n1623 | n3050 ;
  assign n11869 = n8570 ^ n6958 ^ 1'b0 ;
  assign n11874 = n11873 ^ n11870 ^ n11869 ;
  assign n11875 = n9656 ^ n1574 ^ 1'b0 ;
  assign n11876 = n11875 ^ n2255 ^ 1'b0 ;
  assign n11877 = n11874 & ~n11876 ;
  assign n11878 = n1868 ^ n806 ^ 1'b0 ;
  assign n11879 = ~n4751 & n11878 ;
  assign n11880 = n2639 & ~n11879 ;
  assign n11881 = n7268 ^ n1681 ^ 1'b0 ;
  assign n11882 = n3624 | n5920 ;
  assign n11883 = n5564 ^ n5134 ^ 1'b0 ;
  assign n11884 = n4706 | n5019 ;
  assign n11885 = n11883 | n11884 ;
  assign n11886 = n9049 ^ x124 ^ 1'b0 ;
  assign n11887 = n3646 & ~n11886 ;
  assign n11888 = n549 | n806 ;
  assign n11889 = n4282 & ~n11888 ;
  assign n11890 = n3765 & ~n11889 ;
  assign n11891 = n11890 ^ n1898 ^ 1'b0 ;
  assign n11892 = n11891 ^ n2550 ^ n1444 ;
  assign n11893 = n535 & n11892 ;
  assign n11894 = n11893 ^ n10351 ^ 1'b0 ;
  assign n11895 = n1064 & ~n6782 ;
  assign n11896 = n11895 ^ n9441 ^ 1'b0 ;
  assign n11897 = n8343 | n9445 ;
  assign n11898 = n11897 ^ n6293 ^ 1'b0 ;
  assign n11899 = n7619 ^ n3358 ^ 1'b0 ;
  assign n11900 = n6631 & ~n11899 ;
  assign n11901 = n671 | n8609 ;
  assign n11902 = n4429 & ~n11901 ;
  assign n11903 = n831 & n9618 ;
  assign n11904 = n11903 ^ n7123 ^ 1'b0 ;
  assign n11905 = ~n1493 & n6818 ;
  assign n11906 = n11905 ^ n652 ^ 1'b0 ;
  assign n11907 = n2925 ^ n2847 ^ 1'b0 ;
  assign n11908 = n741 | n11907 ;
  assign n11909 = n8648 | n11908 ;
  assign n11910 = n5232 ^ n2748 ^ 1'b0 ;
  assign n11911 = n250 & ~n11910 ;
  assign n11912 = n1887 & n11911 ;
  assign n11913 = n11912 ^ n4528 ^ 1'b0 ;
  assign n11914 = n2755 & ~n3341 ;
  assign n11915 = x56 | n307 ;
  assign n11916 = n7160 ^ n5195 ^ 1'b0 ;
  assign n11917 = ~n11915 & n11916 ;
  assign n11918 = n566 & ~n6221 ;
  assign n11919 = n9337 ^ n2257 ^ 1'b0 ;
  assign n11920 = n2637 & ~n11919 ;
  assign n11921 = n2748 & n5014 ;
  assign n11922 = n1356 & ~n6638 ;
  assign n11923 = n2308 & ~n4146 ;
  assign n11924 = n11923 ^ n7539 ^ 1'b0 ;
  assign n11925 = n11924 ^ n6328 ^ 1'b0 ;
  assign n11926 = n5664 | n7511 ;
  assign n11927 = n4848 & ~n11926 ;
  assign n11928 = n629 | n11927 ;
  assign n11929 = n3843 ^ n3385 ^ 1'b0 ;
  assign n11930 = n11929 ^ n1527 ^ 1'b0 ;
  assign n11931 = n9983 & n11930 ;
  assign n11932 = n1656 & n8844 ;
  assign n11933 = n11932 ^ n6923 ^ 1'b0 ;
  assign n11934 = n6296 ^ n5866 ^ n2423 ;
  assign n11935 = ~n8179 & n11393 ;
  assign n11936 = n11934 & n11935 ;
  assign n11937 = n6261 ^ n1946 ^ 1'b0 ;
  assign n11938 = ( n10154 & n11688 ) | ( n10154 & n11937 ) | ( n11688 & n11937 ) ;
  assign n11939 = n2385 & n5704 ;
  assign n11940 = n5392 | n11939 ;
  assign n11941 = n7905 & ~n11940 ;
  assign n11942 = n819 ^ x114 ^ 1'b0 ;
  assign n11943 = n6921 & ~n11942 ;
  assign n11945 = n8086 ^ n2675 ^ 1'b0 ;
  assign n11946 = n6570 | n11945 ;
  assign n11944 = ~n1116 & n4970 ;
  assign n11947 = n11946 ^ n11944 ^ 1'b0 ;
  assign n11948 = n1087 & ~n2602 ;
  assign n11949 = n1754 | n5043 ;
  assign n11950 = n11949 ^ n221 ^ 1'b0 ;
  assign n11951 = n11950 ^ n8476 ^ 1'b0 ;
  assign n11952 = n9696 | n11951 ;
  assign n11956 = n11137 ^ n3580 ^ 1'b0 ;
  assign n11957 = ~n2014 & n11956 ;
  assign n11953 = n6056 ^ n2624 ^ n1842 ;
  assign n11954 = n8903 ^ n1192 ^ 1'b0 ;
  assign n11955 = n11953 | n11954 ;
  assign n11958 = n11957 ^ n11955 ^ 1'b0 ;
  assign n11959 = n11022 & ~n11958 ;
  assign n11960 = n9471 ^ n783 ^ 1'b0 ;
  assign n11961 = n2409 ^ n869 ^ 1'b0 ;
  assign n11962 = n3492 & ~n6037 ;
  assign n11963 = n3899 ^ n1749 ^ 1'b0 ;
  assign n11964 = n2809 & n11963 ;
  assign n11965 = n3070 & n8367 ;
  assign n11966 = ~n7177 & n11236 ;
  assign n11967 = n11966 ^ n424 ^ 1'b0 ;
  assign n11968 = n8245 | n8335 ;
  assign n11969 = n733 | n5170 ;
  assign n11970 = n3348 ^ n942 ^ 1'b0 ;
  assign n11971 = n11969 | n11970 ;
  assign n11972 = n1079 | n11971 ;
  assign n11973 = n8352 ^ n3278 ^ 1'b0 ;
  assign n11974 = ~n4947 & n11973 ;
  assign n11976 = ~n2557 & n3363 ;
  assign n11975 = ~n6851 & n9504 ;
  assign n11977 = n11976 ^ n11975 ^ 1'b0 ;
  assign n11978 = n2907 & n4846 ;
  assign n11979 = n3391 ^ n632 ^ 1'b0 ;
  assign n11982 = ~n4359 & n10777 ;
  assign n11983 = n11982 ^ n10622 ^ 1'b0 ;
  assign n11980 = ~n2591 & n4476 ;
  assign n11981 = n10965 | n11980 ;
  assign n11984 = n11983 ^ n11981 ^ 1'b0 ;
  assign n11985 = n3770 ^ n2915 ^ 1'b0 ;
  assign n11986 = n10121 ^ n3140 ^ 1'b0 ;
  assign n11987 = n11985 & ~n11986 ;
  assign n11988 = n8691 ^ n4817 ^ 1'b0 ;
  assign n11989 = ~n568 & n8256 ;
  assign n11990 = n11989 ^ n1283 ^ 1'b0 ;
  assign n11991 = ~n7383 & n7473 ;
  assign n11992 = n11991 ^ n9806 ^ 1'b0 ;
  assign n11995 = n1065 & n2710 ;
  assign n11993 = n9986 ^ n3872 ^ 1'b0 ;
  assign n11994 = n4891 | n11993 ;
  assign n11996 = n11995 ^ n11994 ^ 1'b0 ;
  assign n11997 = n5814 ^ n4805 ^ 1'b0 ;
  assign n11998 = n5967 & n11997 ;
  assign n11999 = n11998 ^ x15 ^ 1'b0 ;
  assign n12000 = n2381 & ~n4158 ;
  assign n12001 = n12000 ^ n2555 ^ 1'b0 ;
  assign n12002 = x23 & n6064 ;
  assign n12003 = n10831 & n12002 ;
  assign n12004 = n7362 ^ n4551 ^ 1'b0 ;
  assign n12005 = n2946 & ~n5865 ;
  assign n12006 = n12005 ^ n1387 ^ 1'b0 ;
  assign n12007 = n2478 & ~n6451 ;
  assign n12008 = ~n219 & n8787 ;
  assign n12009 = n7256 | n8840 ;
  assign n12010 = n12008 | n12009 ;
  assign n12011 = ~n10157 & n11077 ;
  assign n12012 = x112 & ~n1930 ;
  assign n12013 = n468 & n12012 ;
  assign n12014 = n911 | n2868 ;
  assign n12015 = ~n639 & n4724 ;
  assign n12016 = n12015 ^ n1474 ^ 1'b0 ;
  assign n12017 = n9060 & n12016 ;
  assign n12018 = ~n1059 & n6170 ;
  assign n12019 = n6361 & ~n12018 ;
  assign n12020 = n3305 & n12019 ;
  assign n12021 = n877 & ~n1646 ;
  assign n12022 = n1493 | n8537 ;
  assign n12023 = n1587 | n12022 ;
  assign n12024 = n3834 | n6258 ;
  assign n12025 = n9632 & ~n12024 ;
  assign n12026 = n9143 | n12025 ;
  assign n12027 = n12026 ^ n10668 ^ 1'b0 ;
  assign n12028 = n996 & ~n12027 ;
  assign n12029 = ~n11787 & n12028 ;
  assign n12030 = n6934 ^ n2041 ^ 1'b0 ;
  assign n12031 = n747 | n12030 ;
  assign n12032 = n932 & ~n12031 ;
  assign n12033 = n1883 ^ n417 ^ 1'b0 ;
  assign n12036 = n11145 ^ n7087 ^ 1'b0 ;
  assign n12037 = n391 | n12036 ;
  assign n12034 = n5907 ^ n3018 ^ 1'b0 ;
  assign n12035 = n9660 & ~n12034 ;
  assign n12038 = n12037 ^ n12035 ^ 1'b0 ;
  assign n12039 = n4953 | n12038 ;
  assign n12040 = n1103 & n12039 ;
  assign n12041 = n6626 & ~n8382 ;
  assign n12042 = n1327 & n12041 ;
  assign n12043 = n12042 ^ n5847 ^ 1'b0 ;
  assign n12044 = n9038 ^ n7029 ^ 1'b0 ;
  assign n12045 = n2089 ^ n1935 ^ 1'b0 ;
  assign n12046 = n1475 & ~n12045 ;
  assign n12047 = n1315 & n12046 ;
  assign n12048 = n3298 | n12047 ;
  assign n12049 = n7948 | n12048 ;
  assign n12050 = n1761 & ~n12049 ;
  assign n12051 = n2091 | n4976 ;
  assign n12052 = x109 | n12051 ;
  assign n12053 = n12052 ^ n7806 ^ 1'b0 ;
  assign n12054 = ( n639 & ~n942 ) | ( n639 & n9200 ) | ( ~n942 & n9200 ) ;
  assign n12055 = n4373 & n12054 ;
  assign n12056 = n11934 & n12055 ;
  assign n12057 = n12053 | n12056 ;
  assign n12058 = n1467 ^ n200 ^ 1'b0 ;
  assign n12059 = ~n6182 & n12058 ;
  assign n12060 = ~n972 & n12059 ;
  assign n12061 = n1327 & ~n9185 ;
  assign n12062 = n2752 & n12061 ;
  assign n12063 = n12062 ^ n6257 ^ 1'b0 ;
  assign n12064 = n811 ^ n722 ^ 1'b0 ;
  assign n12065 = n2641 ^ n747 ^ 1'b0 ;
  assign n12066 = ( ~n696 & n6110 ) | ( ~n696 & n12065 ) | ( n6110 & n12065 ) ;
  assign n12067 = n2708 & n5723 ;
  assign n12068 = n12067 ^ n2951 ^ 1'b0 ;
  assign n12069 = ~n7617 & n12068 ;
  assign n12070 = n12069 ^ n1163 ^ 1'b0 ;
  assign n12071 = ~n7948 & n12070 ;
  assign n12072 = n7001 ^ n6562 ^ 1'b0 ;
  assign n12073 = n8168 ^ n1789 ^ x0 ;
  assign n12074 = n2930 & ~n7822 ;
  assign n12075 = n6651 & n12074 ;
  assign n12076 = n7618 & ~n12075 ;
  assign n12077 = n1761 & n3322 ;
  assign n12078 = n2369 & n12077 ;
  assign n12079 = n1329 | n12078 ;
  assign n12080 = n12079 ^ n992 ^ 1'b0 ;
  assign n12081 = n540 & n12080 ;
  assign n12082 = ~n2269 & n12081 ;
  assign n12083 = n2808 | n4274 ;
  assign n12084 = n12083 ^ n10777 ^ 1'b0 ;
  assign n12085 = n7055 ^ n879 ^ 1'b0 ;
  assign n12086 = ~n1344 & n12085 ;
  assign n12087 = n3005 & ~n6774 ;
  assign n12088 = ~n12086 & n12087 ;
  assign n12089 = n233 & n5139 ;
  assign n12090 = n12089 ^ n3935 ^ 1'b0 ;
  assign n12091 = ~n7619 & n12090 ;
  assign n12092 = n636 | n12091 ;
  assign n12093 = n12092 ^ n3251 ^ 1'b0 ;
  assign n12094 = n2215 & ~n4505 ;
  assign n12095 = n12094 ^ n2369 ^ 1'b0 ;
  assign n12096 = n4636 ^ n3935 ^ 1'b0 ;
  assign n12097 = ~n5512 & n11086 ;
  assign n12098 = n12096 & n12097 ;
  assign n12099 = n6373 ^ n4019 ^ 1'b0 ;
  assign n12100 = n2090 | n12099 ;
  assign n12101 = n6017 ^ n949 ^ x105 ;
  assign n12102 = n891 & n2058 ;
  assign n12103 = n277 & ~n11020 ;
  assign n12104 = ~n12102 & n12103 ;
  assign n12105 = n1688 & ~n3564 ;
  assign n12106 = n2732 & ~n12105 ;
  assign n12107 = ~n2643 & n12106 ;
  assign n12108 = ~n1704 & n12107 ;
  assign n12109 = n6304 & n6638 ;
  assign n12110 = n12109 ^ n1786 ^ 1'b0 ;
  assign n12111 = n8324 ^ n4056 ^ 1'b0 ;
  assign n12112 = ~n931 & n12111 ;
  assign n12113 = n10222 & ~n12112 ;
  assign n12114 = ~n10969 & n12113 ;
  assign n12115 = n12110 & n12114 ;
  assign n12116 = ~n2951 & n9636 ;
  assign n12117 = ~n1732 & n12116 ;
  assign n12118 = n7626 ^ n6587 ^ n5541 ;
  assign n12119 = n3721 ^ n1216 ^ 1'b0 ;
  assign n12120 = n996 & n12119 ;
  assign n12121 = ~n12001 & n12120 ;
  assign n12122 = n6964 & n12121 ;
  assign n12123 = n3005 ^ n956 ^ 1'b0 ;
  assign n12124 = n2156 & n12123 ;
  assign n12125 = n539 & ~n11079 ;
  assign n12126 = ~n5008 & n7462 ;
  assign n12127 = ~n5959 & n12126 ;
  assign n12128 = ~n8927 & n12127 ;
  assign n12129 = n4674 ^ n2325 ^ 1'b0 ;
  assign n12130 = n8030 & ~n12129 ;
  assign n12131 = n1618 & ~n11029 ;
  assign n12132 = ~n12130 & n12131 ;
  assign n12133 = n7668 | n8951 ;
  assign n12134 = n12133 ^ n6203 ^ 1'b0 ;
  assign n12135 = ~n1414 & n1816 ;
  assign n12136 = n12135 ^ n409 ^ 1'b0 ;
  assign n12137 = n1324 & n10823 ;
  assign n12138 = n12136 & n12137 ;
  assign n12139 = n11073 ^ n3120 ^ 1'b0 ;
  assign n12140 = n6596 ^ n2827 ^ 1'b0 ;
  assign n12141 = n5360 & n6590 ;
  assign n12142 = n12141 ^ n9665 ^ 1'b0 ;
  assign n12143 = n5520 ^ n926 ^ 1'b0 ;
  assign n12144 = n801 | n2445 ;
  assign n12145 = n12143 & ~n12144 ;
  assign n12146 = x75 & ~n409 ;
  assign n12147 = ( n1062 & n5160 ) | ( n1062 & n12146 ) | ( n5160 & n12146 ) ;
  assign n12148 = n5112 | n11699 ;
  assign n12149 = n3312 ^ n1508 ^ 1'b0 ;
  assign n12150 = ~n5403 & n10621 ;
  assign n12151 = ~n425 & n12150 ;
  assign n12152 = n553 | n2470 ;
  assign n12153 = x124 | n12152 ;
  assign n12154 = ~n7402 & n12153 ;
  assign n12155 = n12154 ^ n7262 ^ 1'b0 ;
  assign n12156 = n9124 | n12155 ;
  assign n12157 = n11126 ^ n8176 ^ 1'b0 ;
  assign n12158 = n8641 & ~n9230 ;
  assign n12159 = ~n9101 & n12158 ;
  assign n12160 = n1191 | n2028 ;
  assign n12161 = n7040 & n12160 ;
  assign n12162 = n11004 ^ n3587 ^ 1'b0 ;
  assign n12163 = n1177 & n8832 ;
  assign n12164 = ~n12162 & n12163 ;
  assign n12165 = n2030 & n9456 ;
  assign n12166 = n12165 ^ n10528 ^ 1'b0 ;
  assign n12167 = n4189 ^ n3023 ^ 1'b0 ;
  assign n12168 = ~n1808 & n12167 ;
  assign n12169 = ~n4139 & n12168 ;
  assign n12170 = n12169 ^ n1498 ^ 1'b0 ;
  assign n12171 = n8171 & ~n12170 ;
  assign n12172 = ~n1147 & n3956 ;
  assign n12173 = n3381 & ~n12172 ;
  assign n12174 = n12173 ^ n9448 ^ 1'b0 ;
  assign n12175 = n836 | n5929 ;
  assign n12176 = n12175 ^ n1137 ^ 1'b0 ;
  assign n12177 = n3211 & ~n12176 ;
  assign n12178 = n12177 ^ n344 ^ 1'b0 ;
  assign n12179 = n12178 ^ n11472 ^ n6371 ;
  assign n12180 = n311 & n2013 ;
  assign n12181 = n4701 | n12180 ;
  assign n12182 = n5395 & n10641 ;
  assign n12183 = n1290 & ~n11869 ;
  assign n12184 = n5059 & ~n5196 ;
  assign n12185 = n3274 ^ n1328 ^ 1'b0 ;
  assign n12186 = n4111 & ~n12185 ;
  assign n12187 = n2592 | n2602 ;
  assign n12188 = n2961 ^ n1376 ^ 1'b0 ;
  assign n12189 = n1194 | n12188 ;
  assign n12190 = n1973 ^ n1395 ^ 1'b0 ;
  assign n12191 = n11670 & ~n12190 ;
  assign n12192 = n1770 ^ n634 ^ 1'b0 ;
  assign n12193 = n2016 | n12192 ;
  assign n12194 = ( n775 & n7719 ) | ( n775 & n12193 ) | ( n7719 & n12193 ) ;
  assign n12195 = n1545 ^ n1020 ^ 1'b0 ;
  assign n12196 = n1057 & n3320 ;
  assign n12197 = n1128 & n11394 ;
  assign n12198 = n11141 ^ n6019 ^ 1'b0 ;
  assign n12200 = ~n857 & n3833 ;
  assign n12201 = n12200 ^ n533 ^ 1'b0 ;
  assign n12199 = x73 & ~n954 ;
  assign n12202 = n12201 ^ n12199 ^ 1'b0 ;
  assign n12203 = n1990 ^ n1128 ^ 1'b0 ;
  assign n12204 = ~n1028 & n12203 ;
  assign n12205 = n12204 ^ n2535 ^ 1'b0 ;
  assign n12206 = n8982 | n12205 ;
  assign n12207 = n6525 & ~n10655 ;
  assign n12208 = ~n1279 & n4167 ;
  assign n12209 = n12207 & n12208 ;
  assign n12210 = n3521 ^ n1950 ^ 1'b0 ;
  assign n12211 = n1502 & ~n12210 ;
  assign n12212 = n1819 & ~n2324 ;
  assign n12213 = n6915 & n12212 ;
  assign n12214 = n1487 & n12213 ;
  assign n12215 = n12211 & ~n12214 ;
  assign n12216 = ~n287 & n12215 ;
  assign n12217 = ~n5018 & n12216 ;
  assign n12218 = n7184 ^ n3714 ^ 1'b0 ;
  assign n12219 = n1279 & ~n2159 ;
  assign n12220 = ( ~n4137 & n8191 ) | ( ~n4137 & n12219 ) | ( n8191 & n12219 ) ;
  assign n12221 = n8921 ^ n6044 ^ 1'b0 ;
  assign n12222 = n10222 & ~n12221 ;
  assign n12223 = n12221 & n12222 ;
  assign n12224 = n12069 | n12223 ;
  assign n12225 = n12220 | n12224 ;
  assign n12227 = n480 & n4993 ;
  assign n12226 = n3449 & n9462 ;
  assign n12228 = n12227 ^ n12226 ^ 1'b0 ;
  assign n12229 = ( ~n2826 & n5812 ) | ( ~n2826 & n12045 ) | ( n5812 & n12045 ) ;
  assign n12230 = ~n920 & n10554 ;
  assign n12231 = n4731 & ~n12230 ;
  assign n12232 = n12231 ^ n10578 ^ 1'b0 ;
  assign n12235 = n6640 ^ n5168 ^ n872 ;
  assign n12233 = n1569 ^ n544 ^ 1'b0 ;
  assign n12234 = ~n6019 & n12233 ;
  assign n12236 = n12235 ^ n12234 ^ 1'b0 ;
  assign n12237 = n8831 & ~n12236 ;
  assign n12238 = n12237 ^ n11858 ^ 1'b0 ;
  assign n12239 = n9088 ^ n3338 ^ 1'b0 ;
  assign n12240 = n1052 | n12239 ;
  assign n12241 = n3505 & ~n9001 ;
  assign n12242 = n3573 & n4217 ;
  assign n12243 = ~n2015 & n12242 ;
  assign n12244 = n12243 ^ n1064 ^ 1'b0 ;
  assign n12245 = n3002 & ~n12244 ;
  assign n12246 = ~n2231 & n7769 ;
  assign n12247 = ~n12245 & n12246 ;
  assign n12248 = n4364 ^ n4128 ^ n1180 ;
  assign n12249 = n9741 ^ n6541 ^ 1'b0 ;
  assign n12250 = n12056 ^ n6074 ^ 1'b0 ;
  assign n12251 = ( n2930 & ~n6731 ) | ( n2930 & n11801 ) | ( ~n6731 & n11801 ) ;
  assign n12252 = n12251 ^ n8757 ^ 1'b0 ;
  assign n12255 = x107 & ~n11092 ;
  assign n12256 = n12255 ^ x100 ^ 1'b0 ;
  assign n12253 = n4444 & n11597 ;
  assign n12254 = n4419 & ~n12253 ;
  assign n12257 = n12256 ^ n12254 ^ 1'b0 ;
  assign n12258 = n5004 | n9428 ;
  assign n12259 = n2310 & ~n8395 ;
  assign n12260 = n3356 & n12259 ;
  assign n12261 = n7454 ^ n4998 ^ 1'b0 ;
  assign n12262 = n1843 | n2307 ;
  assign n12263 = ~n3083 & n4185 ;
  assign n12264 = ~n8802 & n12263 ;
  assign n12265 = n11893 ^ n11375 ^ 1'b0 ;
  assign n12266 = n1910 & ~n12265 ;
  assign n12267 = n2009 | n4621 ;
  assign n12268 = n12267 ^ n11364 ^ 1'b0 ;
  assign n12269 = n7247 | n12105 ;
  assign n12271 = ~n514 & n3622 ;
  assign n12270 = n4558 ^ n1706 ^ 1'b0 ;
  assign n12272 = n12271 ^ n12270 ^ 1'b0 ;
  assign n12273 = n931 | n4602 ;
  assign n12274 = n323 & ~n12273 ;
  assign n12275 = n12274 ^ n1499 ^ 1'b0 ;
  assign n12276 = n5735 & n12275 ;
  assign n12277 = n12276 ^ n6416 ^ 1'b0 ;
  assign n12278 = n5758 ^ n2000 ^ 1'b0 ;
  assign n12279 = n12256 & ~n12278 ;
  assign n12280 = n9356 ^ n9103 ^ 1'b0 ;
  assign n12281 = n5769 | n12280 ;
  assign n12282 = n9312 ^ n5031 ^ 1'b0 ;
  assign n12283 = n3700 & ~n12282 ;
  assign n12284 = n8565 ^ n3764 ^ n1055 ;
  assign n12285 = n12284 ^ n10863 ^ 1'b0 ;
  assign n12286 = ~n7206 & n12285 ;
  assign n12287 = n12286 ^ n5118 ^ 1'b0 ;
  assign n12288 = n3545 & n6826 ;
  assign n12289 = n3673 & n4966 ;
  assign n12290 = n4189 ^ n558 ^ 1'b0 ;
  assign n12291 = n3753 & ~n12290 ;
  assign n12292 = n12291 ^ n2373 ^ 1'b0 ;
  assign n12293 = n3658 & n12292 ;
  assign n12294 = n2882 & ~n12293 ;
  assign n12295 = n12294 ^ n1551 ^ 1'b0 ;
  assign n12296 = n12295 ^ n6632 ^ 1'b0 ;
  assign n12297 = n12289 | n12296 ;
  assign n12298 = n1551 | n12297 ;
  assign n12300 = n3760 | n5566 ;
  assign n12301 = n433 & ~n12300 ;
  assign n12299 = n446 & n841 ;
  assign n12302 = n12301 ^ n12299 ^ 1'b0 ;
  assign n12303 = n8138 ^ n1744 ^ 1'b0 ;
  assign n12304 = n8658 & n12303 ;
  assign n12305 = n4296 | n6698 ;
  assign n12306 = n12305 ^ n2683 ^ 1'b0 ;
  assign n12307 = n5341 & ~n9889 ;
  assign n12308 = n12307 ^ n2013 ^ 1'b0 ;
  assign n12309 = n5037 & ~n12308 ;
  assign n12310 = n909 | n1748 ;
  assign n12311 = n12310 ^ n173 ^ 1'b0 ;
  assign n12312 = n12311 ^ n8142 ^ 1'b0 ;
  assign n12313 = n3892 & n5793 ;
  assign n12314 = ~n8635 & n9832 ;
  assign n12315 = n12314 ^ n9813 ^ 1'b0 ;
  assign n12316 = n9780 & ~n12315 ;
  assign n12317 = ~n12313 & n12316 ;
  assign n12318 = n1173 & ~n3121 ;
  assign n12319 = n7639 & n12318 ;
  assign n12320 = n10584 ^ n2176 ^ 1'b0 ;
  assign n12321 = n12320 ^ x47 ^ 1'b0 ;
  assign n12322 = ( n1035 & n2967 ) | ( n1035 & n8260 ) | ( n2967 & n8260 ) ;
  assign n12323 = n2708 & n12322 ;
  assign n12324 = n4459 | n11463 ;
  assign n12325 = n12324 ^ n737 ^ 1'b0 ;
  assign n12326 = n2385 & ~n12325 ;
  assign n12327 = ( n1955 & ~n2961 ) | ( n1955 & n4521 ) | ( ~n2961 & n4521 ) ;
  assign n12328 = x10 & x43 ;
  assign n12329 = ~x10 & n12328 ;
  assign n12330 = n450 & ~n12329 ;
  assign n12331 = ~n450 & n12330 ;
  assign n12332 = n237 & ~n12331 ;
  assign n12333 = n12331 & n12332 ;
  assign n12334 = n1872 & ~n12333 ;
  assign n12335 = x44 & n12334 ;
  assign n12336 = n12335 ^ n11830 ^ 1'b0 ;
  assign n12337 = n7059 & ~n8306 ;
  assign n12338 = n4908 & n8648 ;
  assign n12339 = n2633 & n3086 ;
  assign n12340 = ~n786 & n12339 ;
  assign n12341 = n146 & ~n9519 ;
  assign n12342 = n6447 | n12341 ;
  assign n12343 = x77 & ~n1608 ;
  assign n12344 = n12343 ^ n2392 ^ 1'b0 ;
  assign n12345 = n6445 & n10644 ;
  assign n12346 = n11393 ^ n10817 ^ 1'b0 ;
  assign n12347 = n237 & n4126 ;
  assign n12348 = ~n1069 & n6122 ;
  assign n12349 = n12348 ^ n11804 ^ 1'b0 ;
  assign n12350 = n5687 ^ n1833 ^ 1'b0 ;
  assign n12351 = n4272 & n12350 ;
  assign n12352 = n12351 ^ n270 ^ 1'b0 ;
  assign n12353 = n9501 & n12352 ;
  assign n12354 = n2885 ^ n2183 ^ n1905 ;
  assign n12355 = n173 | n11505 ;
  assign n12356 = n766 & n835 ;
  assign n12357 = ~x79 & n12356 ;
  assign n12358 = n6788 ^ n6266 ^ 1'b0 ;
  assign n12359 = n4878 & ~n12358 ;
  assign n12360 = n12359 ^ n3970 ^ 1'b0 ;
  assign n12361 = n3038 ^ n2227 ^ 1'b0 ;
  assign n12362 = n1831 | n2776 ;
  assign n12363 = n12362 ^ n5255 ^ 1'b0 ;
  assign n12367 = n12243 ^ n8093 ^ 1'b0 ;
  assign n12364 = n1228 & n2360 ;
  assign n12365 = n8765 ^ n6361 ^ 1'b0 ;
  assign n12366 = ~n12364 & n12365 ;
  assign n12368 = n12367 ^ n12366 ^ 1'b0 ;
  assign n12369 = x97 & ~n453 ;
  assign n12370 = n12369 ^ n4775 ^ 1'b0 ;
  assign n12371 = n8464 | n11440 ;
  assign n12372 = n11680 ^ n6972 ^ 1'b0 ;
  assign n12373 = n2664 ^ n353 ^ 1'b0 ;
  assign n12374 = n5308 & ~n12373 ;
  assign n12375 = n12374 ^ n9307 ^ 1'b0 ;
  assign n12376 = n2255 | n11937 ;
  assign n12377 = n1116 & ~n12376 ;
  assign n12378 = ~n3834 & n10144 ;
  assign n12379 = ~n9244 & n12378 ;
  assign n12380 = ~x7 & n12379 ;
  assign n12381 = n9242 | n10483 ;
  assign n12382 = n4191 & n7865 ;
  assign n12383 = n12382 ^ n6389 ^ 1'b0 ;
  assign n12384 = ~n4497 & n12383 ;
  assign n12385 = ~n3251 & n12384 ;
  assign n12386 = n584 | n6215 ;
  assign n12387 = n12385 & ~n12386 ;
  assign n12388 = n4388 ^ n1447 ^ 1'b0 ;
  assign n12389 = n6455 & n6540 ;
  assign n12390 = n3140 & n12389 ;
  assign n12391 = n6975 & n12390 ;
  assign n12392 = n5827 ^ n1772 ^ 1'b0 ;
  assign n12393 = ~n1240 & n12392 ;
  assign n12394 = n11606 ^ n7354 ^ n2038 ;
  assign n12395 = n6895 ^ n4377 ^ n3341 ;
  assign n12396 = ( n9172 & ~n9241 ) | ( n9172 & n12395 ) | ( ~n9241 & n12395 ) ;
  assign n12397 = ~n7673 & n8791 ;
  assign n12398 = n2266 & n2420 ;
  assign n12399 = ~n9663 & n12398 ;
  assign n12400 = n10065 & n11061 ;
  assign n12401 = n407 & n1645 ;
  assign n12402 = ~n12083 & n12401 ;
  assign n12403 = n5361 | n12402 ;
  assign n12404 = n12403 ^ n10400 ^ 1'b0 ;
  assign n12405 = n1374 | n4117 ;
  assign n12406 = n6192 ^ n1671 ^ 1'b0 ;
  assign n12407 = n11874 ^ n4916 ^ 1'b0 ;
  assign n12408 = n1204 & ~n2503 ;
  assign n12409 = ~n879 & n12408 ;
  assign n12410 = n11693 & n12409 ;
  assign n12411 = n7179 & n12410 ;
  assign n12412 = n2964 ^ n1554 ^ 1'b0 ;
  assign n12413 = n5450 | n6975 ;
  assign n12414 = n12413 ^ n10994 ^ 1'b0 ;
  assign n12415 = n2136 | n8353 ;
  assign n12416 = n12415 ^ n7153 ^ 1'b0 ;
  assign n12417 = n3196 & n7747 ;
  assign n12418 = n11767 ^ n11126 ^ 1'b0 ;
  assign n12419 = n890 | n5883 ;
  assign n12420 = n5883 & ~n12419 ;
  assign n12421 = n12420 ^ n2469 ^ 1'b0 ;
  assign n12422 = n491 | n880 ;
  assign n12423 = n770 & ~n12422 ;
  assign n12424 = ~n12421 & n12423 ;
  assign n12425 = n12424 ^ n6739 ^ 1'b0 ;
  assign n12426 = n1654 & ~n11569 ;
  assign n12427 = n12425 & n12426 ;
  assign n12428 = ~n7131 & n12427 ;
  assign n12429 = n2260 & n7206 ;
  assign n12430 = n12429 ^ n11959 ^ 1'b0 ;
  assign n12431 = n4087 ^ n2732 ^ 1'b0 ;
  assign n12432 = n876 & n12431 ;
  assign n12433 = n5289 & ~n12432 ;
  assign n12434 = n7129 ^ n5261 ^ 1'b0 ;
  assign n12435 = n2892 ^ n2642 ^ 1'b0 ;
  assign n12436 = n1749 & n12435 ;
  assign n12437 = ~n975 & n2306 ;
  assign n12438 = n2759 & n12437 ;
  assign n12439 = n12438 ^ n1823 ^ 1'b0 ;
  assign n12440 = n211 & n7043 ;
  assign n12441 = n2099 & n9450 ;
  assign n12442 = ~n2264 & n12441 ;
  assign n12443 = ~n1722 & n3356 ;
  assign n12444 = ~n6822 & n10588 ;
  assign n12445 = ~n998 & n1173 ;
  assign n12446 = n9185 | n12445 ;
  assign n12447 = n1561 & ~n1762 ;
  assign n12448 = n11277 & n11911 ;
  assign n12449 = n12448 ^ n5022 ^ 1'b0 ;
  assign n12450 = n8795 | n12449 ;
  assign n12451 = n12450 ^ n11137 ^ 1'b0 ;
  assign n12452 = n9636 & ~n12451 ;
  assign n12453 = n583 & ~n2458 ;
  assign n12454 = ~n3608 & n12453 ;
  assign n12455 = n5417 | n12454 ;
  assign n12456 = n4126 | n4689 ;
  assign n12457 = n2323 & n8975 ;
  assign n12458 = n8673 ^ n195 ^ 1'b0 ;
  assign n12459 = n2112 | n2978 ;
  assign n12460 = n12459 ^ n2990 ^ 1'b0 ;
  assign n12461 = n1738 | n2465 ;
  assign n12462 = n12460 | n12461 ;
  assign n12463 = n8816 ^ n6289 ^ 1'b0 ;
  assign n12464 = n11327 & ~n12463 ;
  assign n12465 = n2385 & ~n7643 ;
  assign n12466 = ~n8215 & n12465 ;
  assign n12467 = n12466 ^ n6916 ^ 1'b0 ;
  assign n12472 = n1855 | n8235 ;
  assign n12473 = n12472 ^ n9115 ^ 1'b0 ;
  assign n12468 = n10777 ^ n1632 ^ 1'b0 ;
  assign n12469 = n12468 ^ n1046 ^ n847 ;
  assign n12470 = n804 | n12469 ;
  assign n12471 = ~n11089 & n12470 ;
  assign n12474 = n12473 ^ n12471 ^ n7195 ;
  assign n12475 = n3266 & n8504 ;
  assign n12476 = n12475 ^ n4576 ^ 1'b0 ;
  assign n12477 = ~n238 & n10556 ;
  assign n12479 = ~n926 & n1737 ;
  assign n12478 = n11805 ^ n1991 ^ 1'b0 ;
  assign n12480 = n12479 ^ n12478 ^ 1'b0 ;
  assign n12481 = n10550 ^ n6718 ^ 1'b0 ;
  assign n12482 = n12480 & ~n12481 ;
  assign n12483 = n5667 ^ x126 ^ 1'b0 ;
  assign n12484 = ~n6151 & n12483 ;
  assign n12485 = x2 & ~n6729 ;
  assign n12486 = n4100 & n12485 ;
  assign n12487 = n1491 | n5535 ;
  assign n12488 = n2900 | n12487 ;
  assign n12489 = n1008 & n8543 ;
  assign n12490 = n6925 & ~n12489 ;
  assign n12491 = n12489 & n12490 ;
  assign n12492 = n7088 | n12491 ;
  assign n12493 = n12491 & ~n12492 ;
  assign n12494 = n10145 & ~n10501 ;
  assign n12495 = n12493 & n12494 ;
  assign n12496 = n7756 | n12495 ;
  assign n12497 = n7756 & ~n12496 ;
  assign n12498 = n463 & n2227 ;
  assign n12499 = ~n7606 & n12498 ;
  assign n12500 = n7082 ^ n6528 ^ 1'b0 ;
  assign n12501 = n11663 & ~n12500 ;
  assign n12502 = n12501 ^ x44 ^ 1'b0 ;
  assign n12503 = n3856 ^ n2030 ^ 1'b0 ;
  assign n12504 = n6234 & ~n7160 ;
  assign n12506 = n4411 ^ n3037 ^ 1'b0 ;
  assign n12507 = n4332 & n12506 ;
  assign n12508 = n4136 ^ n1851 ^ 1'b0 ;
  assign n12509 = n12507 & n12508 ;
  assign n12510 = n3112 & ~n12509 ;
  assign n12505 = ~n2981 & n5152 ;
  assign n12511 = n12510 ^ n12505 ^ n896 ;
  assign n12512 = n3179 | n12511 ;
  assign n12513 = n1810 ^ n595 ^ 1'b0 ;
  assign n12514 = n4648 ^ n4107 ^ 1'b0 ;
  assign n12515 = x40 | n12514 ;
  assign n12516 = ~n1724 & n12357 ;
  assign n12517 = n12516 ^ n211 ^ 1'b0 ;
  assign n12518 = n4902 | n6075 ;
  assign n12519 = n12518 ^ n9507 ^ n6499 ;
  assign n12520 = n4494 ^ n4459 ^ 1'b0 ;
  assign n12521 = n2994 | n12520 ;
  assign n12522 = n12521 ^ n9607 ^ 1'b0 ;
  assign n12523 = n4505 & ~n5365 ;
  assign n12524 = n4467 & ~n12523 ;
  assign n12525 = n12522 & n12524 ;
  assign n12526 = ( ~n1080 & n4706 ) | ( ~n1080 & n5292 ) | ( n4706 & n5292 ) ;
  assign n12527 = n8695 & ~n12526 ;
  assign n12528 = n5749 ^ n845 ^ 1'b0 ;
  assign n12529 = n7723 & ~n12528 ;
  assign n12530 = n2694 & n5907 ;
  assign n12531 = ~n1825 & n12530 ;
  assign n12532 = ~n4654 & n12531 ;
  assign n12534 = n4425 ^ n3862 ^ 1'b0 ;
  assign n12533 = n7011 | n7071 ;
  assign n12535 = n12534 ^ n12533 ^ 1'b0 ;
  assign n12536 = n10387 ^ n6301 ^ 1'b0 ;
  assign n12537 = n9001 & ~n12536 ;
  assign n12538 = x2 & n371 ;
  assign n12539 = ( n1686 & n1772 ) | ( n1686 & n12538 ) | ( n1772 & n12538 ) ;
  assign n12540 = n2760 ^ n824 ^ 1'b0 ;
  assign n12541 = n9640 | n12540 ;
  assign n12542 = n5716 & ~n12541 ;
  assign n12543 = n12542 ^ n10406 ^ 1'b0 ;
  assign n12544 = n3338 ^ n1674 ^ 1'b0 ;
  assign n12545 = n230 & ~n12544 ;
  assign n12546 = ~n2715 & n4227 ;
  assign n12547 = ~n7443 & n12546 ;
  assign n12548 = n12545 & ~n12547 ;
  assign n12549 = n3780 | n8230 ;
  assign n12550 = ( n1880 & ~n9908 ) | ( n1880 & n12153 ) | ( ~n9908 & n12153 ) ;
  assign n12551 = n266 & n12550 ;
  assign n12552 = n3336 | n12122 ;
  assign n12553 = n6212 & ~n12552 ;
  assign n12554 = n1135 & ~n7338 ;
  assign n12555 = n12554 ^ n5866 ^ 1'b0 ;
  assign n12556 = n1221 & ~n12555 ;
  assign n12562 = n5560 ^ n1270 ^ 1'b0 ;
  assign n12563 = n10006 | n12562 ;
  assign n12557 = n533 & n1006 ;
  assign n12558 = n632 & ~n12557 ;
  assign n12559 = n632 & n12558 ;
  assign n12560 = ~n11662 & n12559 ;
  assign n12561 = ~n3276 & n12560 ;
  assign n12564 = n12563 ^ n12561 ^ 1'b0 ;
  assign n12565 = n11571 ^ n1548 ^ 1'b0 ;
  assign n12566 = ~n7411 & n12565 ;
  assign n12568 = n5716 ^ n2171 ^ 1'b0 ;
  assign n12569 = n846 & ~n12568 ;
  assign n12567 = n4716 & ~n9389 ;
  assign n12570 = n12569 ^ n12567 ^ 1'b0 ;
  assign n12571 = n3482 & n12570 ;
  assign n12572 = n1583 | n11644 ;
  assign n12573 = ~x88 & n6234 ;
  assign n12574 = n1005 | n9553 ;
  assign n12575 = n2833 ^ n2085 ^ 1'b0 ;
  assign n12576 = n336 & n5809 ;
  assign n12577 = ~n1031 & n9247 ;
  assign n12578 = ~n12576 & n12577 ;
  assign n12579 = ( n9680 & n12575 ) | ( n9680 & ~n12578 ) | ( n12575 & ~n12578 ) ;
  assign n12580 = ~n1759 & n9864 ;
  assign n12581 = n790 & n3922 ;
  assign n12582 = n946 & ~n5967 ;
  assign n12583 = ~n10000 & n12582 ;
  assign n12584 = n9739 | n12583 ;
  assign n12585 = n12584 ^ n6445 ^ 1'b0 ;
  assign n12586 = n12585 ^ n4590 ^ 1'b0 ;
  assign n12587 = n12586 ^ n8565 ^ 1'b0 ;
  assign n12588 = n1556 ^ n324 ^ 1'b0 ;
  assign n12589 = n12588 ^ n8694 ^ 1'b0 ;
  assign n12590 = n6115 ^ n1996 ^ 1'b0 ;
  assign n12591 = n356 | n2476 ;
  assign n12592 = n12591 ^ n5961 ^ 1'b0 ;
  assign n12593 = n12592 ^ n4921 ^ 1'b0 ;
  assign n12594 = n2525 ^ n911 ^ 1'b0 ;
  assign n12595 = n4871 | n12594 ;
  assign n12596 = x77 & n12595 ;
  assign n12597 = ( n12056 & n12593 ) | ( n12056 & ~n12596 ) | ( n12593 & ~n12596 ) ;
  assign n12598 = n2566 | n6790 ;
  assign n12599 = n12598 ^ n1224 ^ 1'b0 ;
  assign n12600 = n3018 & n10092 ;
  assign n12601 = ~n1265 & n2400 ;
  assign n12602 = ~n2090 & n12601 ;
  assign n12603 = n12602 ^ n8418 ^ 1'b0 ;
  assign n12604 = n3468 ^ n2021 ^ n134 ;
  assign n12605 = n11698 & n12604 ;
  assign n12606 = n2707 & ~n6813 ;
  assign n12607 = n5068 & n12606 ;
  assign n12608 = n5293 | n12607 ;
  assign n12609 = n9222 | n12608 ;
  assign n12610 = n12609 ^ n1665 ^ 1'b0 ;
  assign n12611 = ~n539 & n12610 ;
  assign n12612 = n6456 ^ n835 ^ 1'b0 ;
  assign n12613 = n2771 | n12612 ;
  assign n12614 = n12049 & n12613 ;
  assign n12615 = n1177 & ~n3330 ;
  assign n12616 = ~n9330 & n12615 ;
  assign n12617 = n12616 ^ n5828 ^ 1'b0 ;
  assign n12618 = x20 | n262 ;
  assign n12619 = n12618 ^ n6319 ^ 1'b0 ;
  assign n12620 = n8145 ^ n998 ^ 1'b0 ;
  assign n12621 = n7766 & n12620 ;
  assign n12622 = n4869 & ~n9152 ;
  assign n12623 = n696 & ~n9541 ;
  assign n12624 = n8938 | n12623 ;
  assign n12625 = n1798 & n5909 ;
  assign n12626 = n12625 ^ n11929 ^ 1'b0 ;
  assign n12627 = n250 & n12626 ;
  assign n12628 = n6235 ^ n2085 ^ 1'b0 ;
  assign n12629 = ~n340 & n12628 ;
  assign n12630 = n3688 & ~n3929 ;
  assign n12631 = ~n12629 & n12630 ;
  assign n12632 = n12631 ^ n4259 ^ 1'b0 ;
  assign n12633 = n12627 & n12632 ;
  assign n12634 = n8823 ^ n1285 ^ 1'b0 ;
  assign n12635 = n1707 ^ n1187 ^ 1'b0 ;
  assign n12636 = n3211 & n10000 ;
  assign n12637 = n12636 ^ n6383 ^ 1'b0 ;
  assign n12638 = n3816 ^ x83 ^ 1'b0 ;
  assign n12639 = ~n6228 & n12638 ;
  assign n12640 = n9726 ^ n1344 ^ 1'b0 ;
  assign n12641 = n7949 & ~n12640 ;
  assign n12642 = n6973 & ~n12641 ;
  assign n12643 = n3868 & ~n12642 ;
  assign n12644 = ~n5618 & n12082 ;
  assign n12647 = n11216 ^ n4858 ^ 1'b0 ;
  assign n12645 = n2351 ^ n355 ^ 1'b0 ;
  assign n12646 = n1650 & ~n12645 ;
  assign n12648 = n12647 ^ n12646 ^ 1'b0 ;
  assign n12649 = n11014 ^ n6813 ^ 1'b0 ;
  assign n12650 = n4771 ^ n2213 ^ 1'b0 ;
  assign n12651 = ~n12649 & n12650 ;
  assign n12652 = n5951 | n10630 ;
  assign n12653 = n404 & ~n494 ;
  assign n12654 = x1 & ~n12653 ;
  assign n12655 = ~x59 & n3325 ;
  assign n12656 = n12655 ^ n1267 ^ 1'b0 ;
  assign n12657 = n1116 | n2635 ;
  assign n12658 = n12657 ^ n9217 ^ 1'b0 ;
  assign n12659 = n2637 ^ n1798 ^ 1'b0 ;
  assign n12660 = n2157 | n8260 ;
  assign n12661 = n12660 ^ n995 ^ 1'b0 ;
  assign n12662 = n12659 & n12661 ;
  assign n12663 = n4499 & ~n9151 ;
  assign n12664 = n12663 ^ n11510 ^ 1'b0 ;
  assign n12665 = n12664 ^ n5687 ^ 1'b0 ;
  assign n12666 = n1728 & ~n12235 ;
  assign n12667 = n12666 ^ n6848 ^ 1'b0 ;
  assign n12668 = x75 | n1810 ;
  assign n12669 = n3911 & n12668 ;
  assign n12670 = ~n3018 & n12669 ;
  assign n12671 = ( n737 & ~n6667 ) | ( n737 & n8694 ) | ( ~n6667 & n8694 ) ;
  assign n12672 = n938 ^ n519 ^ 1'b0 ;
  assign n12673 = n7259 ^ n1197 ^ 1'b0 ;
  assign n12674 = n6007 & ~n12673 ;
  assign n12675 = n12674 ^ n4208 ^ 1'b0 ;
  assign n12676 = n8571 & n12675 ;
  assign n12677 = ~n1738 & n5867 ;
  assign n12678 = n4267 ^ n1842 ^ 1'b0 ;
  assign n12679 = n245 & ~n1612 ;
  assign n12680 = n12679 ^ x74 ^ 1'b0 ;
  assign n12681 = n2786 & n5653 ;
  assign n12682 = n12680 & n12681 ;
  assign n12684 = n4895 & ~n6463 ;
  assign n12683 = n7613 & ~n10165 ;
  assign n12685 = n12684 ^ n12683 ^ 1'b0 ;
  assign n12686 = ( ~n6536 & n12682 ) | ( ~n6536 & n12685 ) | ( n12682 & n12685 ) ;
  assign n12687 = ~n672 & n877 ;
  assign n12688 = n7251 ^ n2090 ^ 1'b0 ;
  assign n12689 = ~n4489 & n12688 ;
  assign n12690 = n3865 ^ n1180 ^ 1'b0 ;
  assign n12691 = n12445 & ~n12690 ;
  assign n12692 = n7683 & n12691 ;
  assign n12693 = n11341 ^ n4515 ^ 1'b0 ;
  assign n12694 = n11885 & ~n12693 ;
  assign n12695 = n3659 ^ n1989 ^ 1'b0 ;
  assign n12696 = n240 & n12695 ;
  assign n12697 = n7423 | n9194 ;
  assign n12698 = n12697 ^ n3468 ^ 1'b0 ;
  assign n12699 = ( n5445 & n12696 ) | ( n5445 & n12698 ) | ( n12696 & n12698 ) ;
  assign n12700 = ~n3373 & n4040 ;
  assign n12701 = n3179 ^ n2981 ^ 1'b0 ;
  assign n12702 = n3998 | n12701 ;
  assign n12703 = n3120 & ~n12702 ;
  assign n12704 = n12700 & n12703 ;
  assign n12705 = n12704 ^ n6857 ^ 1'b0 ;
  assign n12706 = n618 & ~n11148 ;
  assign n12707 = ~n3426 & n12706 ;
  assign n12708 = n835 & n1756 ;
  assign n12709 = n1131 | n11227 ;
  assign n12710 = n12709 ^ n11341 ^ n652 ;
  assign n12711 = n2978 | n6098 ;
  assign n12712 = x123 | n12711 ;
  assign n12713 = ~n2148 & n3754 ;
  assign n12714 = n11601 ^ n1837 ^ 1'b0 ;
  assign n12715 = ( n2159 & ~n2585 ) | ( n2159 & n3972 ) | ( ~n2585 & n3972 ) ;
  assign n12716 = n12715 ^ n12053 ^ n3708 ;
  assign n12717 = n4505 ^ n3407 ^ 1'b0 ;
  assign n12718 = n8178 & ~n12717 ;
  assign n12719 = n2545 | n4182 ;
  assign n12720 = n828 & ~n2986 ;
  assign n12721 = n12719 & n12720 ;
  assign n12722 = n12721 ^ n3548 ^ n1251 ;
  assign n12723 = n5968 & ~n12722 ;
  assign n12724 = n2436 | n4723 ;
  assign n12725 = n12724 ^ n428 ^ 1'b0 ;
  assign n12726 = ~n969 & n2994 ;
  assign n12727 = n12726 ^ n7077 ^ 1'b0 ;
  assign n12728 = n12727 ^ n6043 ^ n707 ;
  assign n12729 = n5606 ^ n1116 ^ 1'b0 ;
  assign n12730 = ~n7835 & n12729 ;
  assign n12731 = n2608 | n5220 ;
  assign n12732 = n11474 ^ n3958 ^ 1'b0 ;
  assign n12733 = n8625 | n12732 ;
  assign n12734 = n9046 ^ n1517 ^ 1'b0 ;
  assign n12735 = n10588 & n12734 ;
  assign n12736 = ~n408 & n12735 ;
  assign n12737 = n12736 ^ n1795 ^ 1'b0 ;
  assign n12738 = ~n11782 & n12737 ;
  assign n12739 = n9480 & n11622 ;
  assign n12740 = n12739 ^ n10120 ^ 1'b0 ;
  assign n12742 = n2811 ^ n1240 ^ 1'b0 ;
  assign n12743 = n7195 & n12742 ;
  assign n12741 = n2074 & ~n3264 ;
  assign n12744 = n12743 ^ n12741 ^ 1'b0 ;
  assign n12745 = n482 & n3791 ;
  assign n12746 = n12745 ^ n5973 ^ 1'b0 ;
  assign n12748 = ~n839 & n8991 ;
  assign n12749 = n12748 ^ n5208 ^ 1'b0 ;
  assign n12747 = n7350 ^ n3040 ^ 1'b0 ;
  assign n12750 = n12749 ^ n12747 ^ 1'b0 ;
  assign n12752 = ~n2871 & n5474 ;
  assign n12751 = n12383 ^ n2678 ^ 1'b0 ;
  assign n12753 = n12752 ^ n12751 ^ n8511 ;
  assign n12754 = n409 & ~n5231 ;
  assign n12755 = n12754 ^ n5392 ^ 1'b0 ;
  assign n12756 = n3069 & n12755 ;
  assign n12758 = n1216 | n11079 ;
  assign n12757 = n7202 | n7602 ;
  assign n12759 = n12758 ^ n12757 ^ 1'b0 ;
  assign n12760 = x76 & ~n1973 ;
  assign n12761 = ~n11611 & n12760 ;
  assign n12762 = n12761 ^ n2822 ^ 1'b0 ;
  assign n12763 = n1534 & n12762 ;
  assign n12764 = ~n1419 & n8869 ;
  assign n12765 = n12764 ^ n6652 ^ 1'b0 ;
  assign n12766 = n12763 & ~n12765 ;
  assign n12767 = ~n5962 & n12766 ;
  assign n12768 = n741 & n4091 ;
  assign n12769 = ~n4891 & n12768 ;
  assign n12770 = n7298 & ~n12015 ;
  assign n12771 = ~n6549 & n7484 ;
  assign n12772 = n2446 | n4247 ;
  assign n12773 = n12772 ^ n3577 ^ 1'b0 ;
  assign n12774 = ~n1593 & n12773 ;
  assign n12775 = ~n2178 & n2409 ;
  assign n12776 = ( ~n2585 & n8961 ) | ( ~n2585 & n11186 ) | ( n8961 & n11186 ) ;
  assign n12777 = n11061 ^ n3534 ^ 1'b0 ;
  assign n12778 = n1292 | n12777 ;
  assign n12779 = n12778 ^ n1769 ^ 1'b0 ;
  assign n12780 = n12779 ^ n8833 ^ 1'b0 ;
  assign n12781 = n12776 & n12780 ;
  assign n12782 = n12775 & ~n12781 ;
  assign n12783 = n7298 ^ n5388 ^ 1'b0 ;
  assign n12784 = n5132 ^ n3434 ^ 1'b0 ;
  assign n12785 = n11787 ^ n4190 ^ n2361 ;
  assign n12786 = n1578 ^ n245 ^ 1'b0 ;
  assign n12787 = ~n1609 & n12786 ;
  assign n12788 = n4971 ^ n439 ^ 1'b0 ;
  assign n12789 = n1130 | n12788 ;
  assign n12792 = n2821 | n8109 ;
  assign n12793 = n12792 ^ n1301 ^ 1'b0 ;
  assign n12790 = ( n522 & ~n6095 ) | ( n522 & n10027 ) | ( ~n6095 & n10027 ) ;
  assign n12791 = n5437 & ~n12790 ;
  assign n12794 = n12793 ^ n12791 ^ 1'b0 ;
  assign n12795 = n12789 & ~n12794 ;
  assign n12796 = ~n5573 & n6989 ;
  assign n12797 = ~n4048 & n4904 ;
  assign n12798 = n4885 ^ n2411 ^ 1'b0 ;
  assign n12799 = ~n753 & n12798 ;
  assign n12800 = ~n2969 & n12799 ;
  assign n12801 = n12800 ^ n7986 ^ 1'b0 ;
  assign n12802 = n8821 | n9430 ;
  assign n12803 = n8980 ^ n3488 ^ 1'b0 ;
  assign n12804 = n141 & n5008 ;
  assign n12805 = n12804 ^ n2392 ^ 1'b0 ;
  assign n12806 = n12803 & n12805 ;
  assign n12807 = n9763 | n12806 ;
  assign n12808 = n1067 | n3120 ;
  assign n12809 = x7 | n12808 ;
  assign n12810 = n1176 & n1993 ;
  assign n12811 = n1732 ^ n972 ^ 1'b0 ;
  assign n12812 = ~n2041 & n12811 ;
  assign n12813 = ~n1342 & n2689 ;
  assign n12814 = n4919 & n7111 ;
  assign n12815 = n12814 ^ n4417 ^ 1'b0 ;
  assign n12816 = ~n12557 & n12815 ;
  assign n12817 = ~n3484 & n3740 ;
  assign n12818 = n7688 & ~n12817 ;
  assign n12819 = n12818 ^ n8174 ^ 1'b0 ;
  assign n12820 = ~n770 & n3161 ;
  assign n12821 = n1243 & n12820 ;
  assign n12822 = n3500 & n12821 ;
  assign n12823 = ~n356 & n9281 ;
  assign n12824 = n3977 ^ n1407 ^ 1'b0 ;
  assign n12825 = n6451 & ~n12824 ;
  assign n12826 = n8055 & ~n12825 ;
  assign n12827 = n2094 & n12826 ;
  assign n12828 = ~n642 & n911 ;
  assign n12829 = n9727 & n12828 ;
  assign n12830 = n2566 ^ x76 ^ 1'b0 ;
  assign n12831 = n1221 & ~n12830 ;
  assign n12832 = n12829 & n12831 ;
  assign n12833 = n1443 & n5369 ;
  assign n12834 = n12833 ^ n2990 ^ 1'b0 ;
  assign n12835 = n12834 ^ n870 ^ 1'b0 ;
  assign n12836 = n2378 & ~n12835 ;
  assign n12837 = n5985 & n12836 ;
  assign n12838 = n12837 ^ n642 ^ 1'b0 ;
  assign n12839 = n4505 & ~n5898 ;
  assign n12840 = n1618 & ~n6989 ;
  assign n12841 = n12840 ^ n6381 ^ 1'b0 ;
  assign n12842 = n623 & n12841 ;
  assign n12843 = n12842 ^ n11277 ^ 1'b0 ;
  assign n12844 = ~n2518 & n5867 ;
  assign n12845 = n7407 ^ n5855 ^ 1'b0 ;
  assign n12846 = ~n12844 & n12845 ;
  assign n12848 = n2579 & n3069 ;
  assign n12847 = x47 & ~n3640 ;
  assign n12849 = n12848 ^ n12847 ^ 1'b0 ;
  assign n12850 = ~n5488 & n12849 ;
  assign n12851 = n11334 ^ n2271 ^ 1'b0 ;
  assign n12852 = n8367 ^ n8028 ^ 1'b0 ;
  assign n12853 = n12702 ^ n11497 ^ 1'b0 ;
  assign n12854 = n2422 & ~n4992 ;
  assign n12855 = n12854 ^ n1355 ^ 1'b0 ;
  assign n12856 = ~n1558 & n1880 ;
  assign n12857 = ~n12855 & n12856 ;
  assign n12858 = n10458 & n11632 ;
  assign n12859 = n5002 & n12858 ;
  assign n12860 = n2181 | n10515 ;
  assign n12861 = n12860 ^ n1228 ^ 1'b0 ;
  assign n12862 = n1146 & n12861 ;
  assign n12863 = n12859 | n12862 ;
  assign n12864 = ~n3976 & n4484 ;
  assign n12865 = ~n4282 & n5278 ;
  assign n12867 = n2602 ^ n155 ^ 1'b0 ;
  assign n12868 = n4418 & n12867 ;
  assign n12866 = n171 | n11341 ;
  assign n12869 = n12868 ^ n12866 ^ 1'b0 ;
  assign n12870 = n1948 ^ n891 ^ 1'b0 ;
  assign n12871 = n227 & n6337 ;
  assign n12872 = n2819 | n5388 ;
  assign n12873 = n1937 & ~n12872 ;
  assign n12874 = n963 & n11010 ;
  assign n12876 = n9006 & n9498 ;
  assign n12875 = ~n3231 & n4530 ;
  assign n12877 = n12876 ^ n12875 ^ n3295 ;
  assign n12878 = n519 & n3103 ;
  assign n12879 = n12878 ^ n326 ^ 1'b0 ;
  assign n12880 = n5691 & n12879 ;
  assign n12881 = n8028 ^ n1506 ^ 1'b0 ;
  assign n12882 = ~n11092 & n12881 ;
  assign n12883 = n12882 ^ n3283 ^ 1'b0 ;
  assign n12884 = ~n6557 & n12883 ;
  assign n12885 = ~n6059 & n8956 ;
  assign n12886 = n12885 ^ n11648 ^ 1'b0 ;
  assign n12887 = n4907 | n7222 ;
  assign n12888 = n12887 ^ n11329 ^ 1'b0 ;
  assign n12889 = n12888 ^ n2020 ^ 1'b0 ;
  assign n12890 = ~x1 & n5663 ;
  assign n12891 = n5550 ^ n4022 ^ 1'b0 ;
  assign n12892 = n1226 | n4069 ;
  assign n12893 = n9916 & ~n12892 ;
  assign n12894 = n12893 ^ n4045 ^ 1'b0 ;
  assign n12895 = n12894 ^ n6823 ^ 1'b0 ;
  assign n12896 = n678 & ~n2906 ;
  assign n12897 = n12896 ^ n3458 ^ 1'b0 ;
  assign n12898 = n1103 & n10763 ;
  assign n12899 = n7132 ^ n2602 ^ 1'b0 ;
  assign n12900 = n12898 & ~n12899 ;
  assign n12901 = n1091 & n2744 ;
  assign n12902 = n5378 & ~n7236 ;
  assign n12903 = n12902 ^ n3369 ^ 1'b0 ;
  assign n12904 = n983 | n3539 ;
  assign n12905 = n4777 ^ n482 ^ 1'b0 ;
  assign n12906 = n5603 | n12905 ;
  assign n12907 = n6883 & n12906 ;
  assign n12908 = n2105 ^ n1830 ^ 1'b0 ;
  assign n12909 = n4217 & n12908 ;
  assign n12910 = n12909 ^ n11489 ^ 1'b0 ;
  assign n12911 = n4838 & n6226 ;
  assign n12912 = n1894 ^ n1477 ^ 1'b0 ;
  assign n12913 = n1733 & n12912 ;
  assign n12914 = ~n10887 & n12913 ;
  assign n12915 = n12914 ^ n591 ^ 1'b0 ;
  assign n12916 = n3765 & n6965 ;
  assign n12917 = n516 | n9227 ;
  assign n12918 = n12916 & ~n12917 ;
  assign n12919 = n353 | n2448 ;
  assign n12920 = n353 & ~n12919 ;
  assign n12921 = n5508 ^ n830 ^ 1'b0 ;
  assign n12922 = n12920 & ~n12921 ;
  assign n12923 = ( n880 & ~n3310 ) | ( n880 & n3534 ) | ( ~n3310 & n3534 ) ;
  assign n12924 = n11076 | n12923 ;
  assign n12925 = n12922 | n12924 ;
  assign n12926 = n7911 & n12925 ;
  assign n12927 = ~n12925 & n12926 ;
  assign n12928 = ~n978 & n5575 ;
  assign n12929 = n1310 | n2472 ;
  assign n12930 = n4025 | n11023 ;
  assign n12931 = n9495 ^ n4948 ^ 1'b0 ;
  assign n12932 = ~n9197 & n12931 ;
  assign n12933 = ~n992 & n11330 ;
  assign n12934 = n12933 ^ n2358 ^ 1'b0 ;
  assign n12935 = n12934 ^ n11469 ^ 1'b0 ;
  assign n12936 = n3812 ^ n2041 ^ 1'b0 ;
  assign n12937 = ~n1086 & n1478 ;
  assign n12938 = n2526 | n6757 ;
  assign n12939 = n12937 & ~n12938 ;
  assign n12940 = n12051 & n12939 ;
  assign n12941 = n3049 & ~n6301 ;
  assign n12942 = ~n5898 & n12941 ;
  assign n12943 = n1387 | n5151 ;
  assign n12944 = n7001 | n12943 ;
  assign n12949 = n6688 ^ n2481 ^ 1'b0 ;
  assign n12946 = n2932 & ~n3075 ;
  assign n12947 = n12946 ^ n2008 ^ 1'b0 ;
  assign n12948 = n10860 & n12947 ;
  assign n12950 = n12949 ^ n12948 ^ 1'b0 ;
  assign n12945 = ~n3707 & n7991 ;
  assign n12951 = n12950 ^ n12945 ^ 1'b0 ;
  assign n12952 = n8227 | n12478 ;
  assign n12953 = n11681 ^ n6083 ^ 1'b0 ;
  assign n12954 = n2293 & n12953 ;
  assign n12955 = n8599 ^ n267 ^ 1'b0 ;
  assign n12956 = n12954 & ~n12955 ;
  assign n12957 = n6837 & n8658 ;
  assign n12958 = n12957 ^ n240 ^ 1'b0 ;
  assign n12959 = n3364 & ~n4844 ;
  assign n12960 = n678 & n12959 ;
  assign n12961 = n171 & n6341 ;
  assign n12962 = ~n12960 & n12961 ;
  assign n12963 = n5945 ^ n2958 ^ 1'b0 ;
  assign n12964 = n849 & ~n12963 ;
  assign n12965 = ~n2352 & n12964 ;
  assign n12966 = ~n5868 & n12965 ;
  assign n12967 = n4248 | n6835 ;
  assign n12968 = n8205 & ~n12967 ;
  assign n12970 = n217 & n3047 ;
  assign n12971 = ~n2358 & n12970 ;
  assign n12969 = n4038 ^ n3348 ^ 1'b0 ;
  assign n12972 = n12971 ^ n12969 ^ 1'b0 ;
  assign n12973 = n12972 ^ n8746 ^ 1'b0 ;
  assign n12974 = ~n10142 & n12973 ;
  assign n12975 = n2633 & ~n10058 ;
  assign n12976 = n1057 & n12772 ;
  assign n12977 = n503 & ~n4056 ;
  assign n12978 = n11261 & ~n12977 ;
  assign n12979 = n2773 ^ n501 ^ 1'b0 ;
  assign n12980 = ~n10326 & n12979 ;
  assign n12981 = n1345 & ~n1900 ;
  assign n12982 = n5417 & n12981 ;
  assign n12983 = n2478 & ~n3833 ;
  assign n12985 = n10557 ^ n5810 ^ 1'b0 ;
  assign n12986 = n4662 & ~n12985 ;
  assign n12984 = ~n4118 & n10144 ;
  assign n12987 = n12986 ^ n12984 ^ 1'b0 ;
  assign n12988 = n9712 ^ n242 ^ 1'b0 ;
  assign n12989 = ~n2775 & n12988 ;
  assign n12990 = n11209 ^ n4382 ^ 1'b0 ;
  assign n12991 = n1993 & n2815 ;
  assign n12992 = ~n5175 & n12991 ;
  assign n12993 = n1419 & ~n2864 ;
  assign n12994 = n898 & n1908 ;
  assign n12995 = n1905 & ~n3891 ;
  assign n12996 = n12995 ^ n4769 ^ 1'b0 ;
  assign n12997 = n2123 & n9462 ;
  assign n12998 = n1447 & ~n1484 ;
  assign n12999 = n10285 & ~n12998 ;
  assign n13000 = n861 & ~n6110 ;
  assign n13001 = n13000 ^ n5308 ^ 1'b0 ;
  assign n13003 = n1016 & n1623 ;
  assign n13004 = n13003 ^ n1188 ^ 1'b0 ;
  assign n13002 = n4416 & n11840 ;
  assign n13005 = n13004 ^ n13002 ^ 1'b0 ;
  assign n13006 = n6979 ^ n3695 ^ 1'b0 ;
  assign n13007 = n645 & n13006 ;
  assign n13008 = n11992 & n13007 ;
  assign n13009 = n13008 ^ n10840 ^ 1'b0 ;
  assign n13010 = n2875 & n4146 ;
  assign n13011 = n1002 | n13010 ;
  assign n13012 = n10121 | n13011 ;
  assign n13014 = n2624 | n3470 ;
  assign n13015 = n13014 ^ n484 ^ 1'b0 ;
  assign n13016 = n1167 & ~n13015 ;
  assign n13013 = ~x2 & n7848 ;
  assign n13017 = n13016 ^ n13013 ^ 1'b0 ;
  assign n13018 = n3554 ^ n3290 ^ 1'b0 ;
  assign n13019 = n11060 ^ n5160 ^ 1'b0 ;
  assign n13020 = n13018 & n13019 ;
  assign n13021 = ~n3585 & n10597 ;
  assign n13022 = n1226 | n8902 ;
  assign n13023 = ~n6782 & n13022 ;
  assign n13024 = n13023 ^ n6839 ^ 1'b0 ;
  assign n13025 = n7664 ^ n361 ^ 1'b0 ;
  assign n13026 = n7699 & ~n13025 ;
  assign n13027 = n13026 ^ n7401 ^ 1'b0 ;
  assign n13028 = ~n9157 & n10965 ;
  assign n13029 = n1629 & ~n13028 ;
  assign n13031 = n155 | n1493 ;
  assign n13032 = n2173 & ~n13031 ;
  assign n13033 = n2602 & ~n3341 ;
  assign n13034 = n13032 | n13033 ;
  assign n13035 = n555 | n13034 ;
  assign n13036 = n13035 ^ n5196 ^ 1'b0 ;
  assign n13030 = n763 & ~n6284 ;
  assign n13037 = n13036 ^ n13030 ^ n5451 ;
  assign n13038 = n1057 & n7170 ;
  assign n13039 = n9385 ^ n3034 ^ 1'b0 ;
  assign n13040 = n13039 ^ n2264 ^ 1'b0 ;
  assign n13041 = n2313 & ~n9803 ;
  assign n13042 = n718 | n8174 ;
  assign n13043 = n10695 | n13042 ;
  assign n13044 = n6427 ^ n1560 ^ 1'b0 ;
  assign n13045 = n4146 & ~n13044 ;
  assign n13046 = n8619 ^ n7169 ^ 1'b0 ;
  assign n13047 = ~n7405 & n13046 ;
  assign n13048 = n13047 ^ n5790 ^ 1'b0 ;
  assign n13049 = n3429 & n8872 ;
  assign n13050 = ~n6557 & n13049 ;
  assign n13051 = n996 & n13050 ;
  assign n13053 = n2301 & n8296 ;
  assign n13052 = ~n1163 & n5667 ;
  assign n13054 = n13053 ^ n13052 ^ 1'b0 ;
  assign n13055 = n4417 | n13054 ;
  assign n13056 = n5280 & n13055 ;
  assign n13057 = n13056 ^ n12075 ^ 1'b0 ;
  assign n13058 = n6826 ^ n5757 ^ 1'b0 ;
  assign n13059 = ~n3636 & n13058 ;
  assign n13060 = n4661 & n13059 ;
  assign n13061 = n12829 ^ n3659 ^ 1'b0 ;
  assign n13062 = n12971 | n13061 ;
  assign n13063 = n3094 & ~n13062 ;
  assign n13064 = n5522 & ~n10040 ;
  assign n13065 = n13064 ^ n680 ^ 1'b0 ;
  assign n13066 = n1973 ^ n516 ^ 1'b0 ;
  assign n13067 = n13066 ^ n5160 ^ 1'b0 ;
  assign n13068 = n3285 | n6004 ;
  assign n13069 = n13068 ^ n5110 ^ 1'b0 ;
  assign n13070 = n1226 | n13069 ;
  assign n13072 = n5186 & ~n6271 ;
  assign n13073 = ~n7777 & n13072 ;
  assign n13071 = n307 & n9872 ;
  assign n13074 = n13073 ^ n13071 ^ 1'b0 ;
  assign n13075 = ~n663 & n2878 ;
  assign n13076 = n13075 ^ n2273 ^ 1'b0 ;
  assign n13077 = ~n2198 & n6167 ;
  assign n13078 = n13077 ^ n7567 ^ 1'b0 ;
  assign n13079 = ~n3116 & n4385 ;
  assign n13080 = n2215 | n2683 ;
  assign n13081 = ~n724 & n4873 ;
  assign n13082 = ~n13080 & n13081 ;
  assign n13083 = n408 & n5652 ;
  assign n13084 = n13083 ^ n8382 ^ 1'b0 ;
  assign n13085 = n5132 & n11324 ;
  assign n13086 = n13085 ^ n1760 ^ 1'b0 ;
  assign n13087 = n5653 & n7731 ;
  assign n13088 = n3473 & n13087 ;
  assign n13089 = n12619 ^ n8261 ^ 1'b0 ;
  assign n13090 = n3072 & ~n13089 ;
  assign n13091 = ( n2495 & ~n3041 ) | ( n2495 & n5367 ) | ( ~n3041 & n5367 ) ;
  assign n13092 = n1251 & n10233 ;
  assign n13093 = n2775 | n13092 ;
  assign n13094 = n8103 ^ n5647 ^ 1'b0 ;
  assign n13095 = n1534 & ~n6570 ;
  assign n13096 = n6534 & n13095 ;
  assign n13097 = n7898 ^ n1615 ^ 1'b0 ;
  assign n13098 = n3572 | n6940 ;
  assign n13099 = n221 & ~n13098 ;
  assign n13100 = n8473 | n13099 ;
  assign n13101 = n137 & n13100 ;
  assign n13102 = n13101 ^ n12191 ^ 1'b0 ;
  assign n13103 = n4983 ^ n1037 ^ 1'b0 ;
  assign n13104 = ( n1471 & n2743 ) | ( n1471 & ~n13103 ) | ( n2743 & ~n13103 ) ;
  assign n13105 = n3898 | n13104 ;
  assign n13106 = x66 & ~n7809 ;
  assign n13107 = n315 & n13106 ;
  assign n13108 = n3158 | n7237 ;
  assign n13109 = n10436 ^ n4126 ^ n163 ;
  assign n13110 = n2409 & ~n13109 ;
  assign n13111 = ( x108 & n181 ) | ( x108 & ~n4993 ) | ( n181 & ~n4993 ) ;
  assign n13112 = ~n1456 & n13111 ;
  assign n13113 = n13112 ^ n4707 ^ 1'b0 ;
  assign n13114 = ~n986 & n6026 ;
  assign n13115 = ~n10064 & n13114 ;
  assign n13116 = n7517 ^ n963 ^ 1'b0 ;
  assign n13117 = n1773 ^ n773 ^ 1'b0 ;
  assign n13118 = n1798 & n12347 ;
  assign n13119 = ~n491 & n7138 ;
  assign n13120 = n4496 & n7449 ;
  assign n13121 = n11355 ^ n9697 ^ 1'b0 ;
  assign n13122 = n4911 ^ n1654 ^ 1'b0 ;
  assign n13123 = n7439 ^ n132 ^ 1'b0 ;
  assign n13124 = ~n13122 & n13123 ;
  assign n13125 = ~n9213 & n13124 ;
  assign n13126 = n13125 ^ n12219 ^ 1'b0 ;
  assign n13127 = n1613 & n7989 ;
  assign n13128 = n5971 & ~n13127 ;
  assign n13129 = n2434 & ~n3240 ;
  assign n13130 = ~n4376 & n13129 ;
  assign n13131 = n5324 & n13130 ;
  assign n13132 = ~n1927 & n5464 ;
  assign n13133 = n3897 & ~n7498 ;
  assign n13134 = ~n13132 & n13133 ;
  assign n13135 = n13131 | n13134 ;
  assign n13137 = n1001 & n2651 ;
  assign n13136 = ~n8670 & n10152 ;
  assign n13138 = n13137 ^ n13136 ^ 1'b0 ;
  assign n13139 = n3773 | n13138 ;
  assign n13140 = n8199 & n12609 ;
  assign n13141 = n13140 ^ n8568 ^ 1'b0 ;
  assign n13144 = n6073 ^ n570 ^ 1'b0 ;
  assign n13142 = x77 & ~n7257 ;
  assign n13143 = n2478 & n13142 ;
  assign n13145 = n13144 ^ n13143 ^ 1'b0 ;
  assign n13146 = n2321 | n7446 ;
  assign n13147 = n12273 ^ n6840 ^ 1'b0 ;
  assign n13148 = n9845 ^ n2767 ^ 1'b0 ;
  assign n13149 = n2442 ^ n1860 ^ 1'b0 ;
  assign n13150 = n7128 & ~n8279 ;
  assign n13151 = n576 & n13150 ;
  assign n13152 = n13151 ^ n656 ^ 1'b0 ;
  assign n13153 = n9098 & n10619 ;
  assign n13154 = n5771 & ~n7405 ;
  assign n13155 = n9891 & n13154 ;
  assign n13156 = n2983 | n13155 ;
  assign n13157 = n8249 & ~n13156 ;
  assign n13158 = n1188 & n3447 ;
  assign n13159 = n9787 & n13158 ;
  assign n13160 = n1927 | n13159 ;
  assign n13161 = n2233 & ~n13160 ;
  assign n13162 = x16 & ~n8924 ;
  assign n13163 = ( ~n825 & n4182 ) | ( ~n825 & n10687 ) | ( n4182 & n10687 ) ;
  assign n13164 = n5485 | n7454 ;
  assign n13165 = n324 & ~n13164 ;
  assign n13166 = n9630 & ~n13165 ;
  assign n13167 = n6474 ^ n4554 ^ 1'b0 ;
  assign n13168 = n288 & n6933 ;
  assign n13173 = n3333 ^ n425 ^ 1'b0 ;
  assign n13170 = n3837 ^ x3 ^ 1'b0 ;
  assign n13171 = n2321 & ~n13170 ;
  assign n13169 = n6921 ^ n1830 ^ 1'b0 ;
  assign n13172 = n13171 ^ n13169 ^ 1'b0 ;
  assign n13174 = n13173 ^ n13172 ^ 1'b0 ;
  assign n13175 = ~n1051 & n6901 ;
  assign n13176 = n13175 ^ n6959 ^ 1'b0 ;
  assign n13178 = n5956 & ~n6024 ;
  assign n13179 = n13178 ^ n5898 ^ 1'b0 ;
  assign n13180 = ~n2154 & n13179 ;
  assign n13177 = n339 | n10326 ;
  assign n13181 = n13180 ^ n13177 ^ 1'b0 ;
  assign n13182 = n1878 ^ n737 ^ 1'b0 ;
  assign n13183 = n6176 & ~n13182 ;
  assign n13184 = ~n5798 & n13183 ;
  assign n13185 = n849 | n13184 ;
  assign n13186 = n7272 & ~n9006 ;
  assign n13187 = n13186 ^ n12974 ^ 1'b0 ;
  assign n13188 = n3608 | n3629 ;
  assign n13189 = n13188 ^ n5435 ^ 1'b0 ;
  assign n13190 = n9763 | n13189 ;
  assign n13191 = n3157 & ~n7375 ;
  assign n13192 = n13190 | n13191 ;
  assign n13193 = n7987 ^ n980 ^ 1'b0 ;
  assign n13194 = n129 ^ x81 ^ 1'b0 ;
  assign n13195 = x18 & ~n13194 ;
  assign n13196 = n13195 ^ n8084 ^ 1'b0 ;
  assign n13197 = n1057 & n13196 ;
  assign n13198 = n8316 ^ n7946 ^ 1'b0 ;
  assign n13199 = n10463 ^ n722 ^ 1'b0 ;
  assign n13200 = n3792 & n13199 ;
  assign n13201 = n1028 | n11795 ;
  assign n13202 = ~n5276 & n6652 ;
  assign n13203 = n7852 & n9345 ;
  assign n13204 = ~n1344 & n5659 ;
  assign n13205 = ~n3206 & n13204 ;
  assign n13206 = ~n4746 & n5857 ;
  assign n13207 = n13206 ^ n2555 ^ 1'b0 ;
  assign n13208 = n5822 & ~n13207 ;
  assign n13209 = n13205 & n13208 ;
  assign n13210 = n11397 ^ n9130 ^ 1'b0 ;
  assign n13211 = n8235 & n13210 ;
  assign n13212 = n2755 ^ n1753 ^ 1'b0 ;
  assign n13213 = n13212 ^ n11496 ^ n1120 ;
  assign n13214 = n1526 | n2874 ;
  assign n13215 = n13214 ^ n1534 ^ 1'b0 ;
  assign n13216 = n7372 | n13215 ;
  assign n13217 = n8329 ^ n4461 ^ 1'b0 ;
  assign n13218 = n13217 ^ n1158 ^ 1'b0 ;
  assign n13219 = n3664 | n13218 ;
  assign n13220 = ( n514 & ~n3733 ) | ( n514 & n13219 ) | ( ~n3733 & n13219 ) ;
  assign n13221 = n12445 ^ n5475 ^ 1'b0 ;
  assign n13222 = ~n2992 & n13221 ;
  assign n13223 = ~n823 & n8244 ;
  assign n13227 = ( n144 & ~n5148 ) | ( n144 & n7762 ) | ( ~n5148 & n7762 ) ;
  assign n13224 = n586 & ~n4402 ;
  assign n13225 = n10827 & n13224 ;
  assign n13226 = n13225 ^ n11258 ^ 1'b0 ;
  assign n13228 = n13227 ^ n13226 ^ 1'b0 ;
  assign n13229 = n13223 & n13228 ;
  assign n13230 = ~n7747 & n9871 ;
  assign n13231 = n13230 ^ n1923 ^ 1'b0 ;
  assign n13232 = ~x72 & n4307 ;
  assign n13233 = ~n5649 & n13232 ;
  assign n13234 = n8589 ^ n1720 ^ 1'b0 ;
  assign n13236 = n2467 ^ n922 ^ 1'b0 ;
  assign n13237 = n3166 & n13236 ;
  assign n13235 = n5839 ^ n914 ^ 1'b0 ;
  assign n13238 = n13237 ^ n13235 ^ 1'b0 ;
  assign n13239 = n294 & n13238 ;
  assign n13240 = n1576 & n1581 ;
  assign n13241 = ~n3188 & n3853 ;
  assign n13242 = n7824 ^ n1741 ^ 1'b0 ;
  assign n13243 = n12834 ^ n9351 ^ 1'b0 ;
  assign n13244 = n4708 & ~n11254 ;
  assign n13245 = n3195 ^ n945 ^ 1'b0 ;
  assign n13246 = ~n2743 & n13245 ;
  assign n13247 = ~n12430 & n13246 ;
  assign n13248 = n1599 ^ n721 ^ 1'b0 ;
  assign n13249 = n8526 ^ n2629 ^ 1'b0 ;
  assign n13250 = n2127 & ~n13249 ;
  assign n13251 = n10754 ^ n8955 ^ 1'b0 ;
  assign n13252 = n4948 ^ n2215 ^ 1'b0 ;
  assign n13253 = n7044 & n13252 ;
  assign n13254 = ~n4402 & n13253 ;
  assign n13255 = n782 & ~n1774 ;
  assign n13256 = n2030 | n3952 ;
  assign n13257 = n13256 ^ n2656 ^ 1'b0 ;
  assign n13258 = n2482 ^ n354 ^ 1'b0 ;
  assign n13259 = n4584 & n13258 ;
  assign n13260 = n13259 ^ n4660 ^ 1'b0 ;
  assign n13261 = n5954 & ~n7736 ;
  assign n13262 = n9778 ^ n7226 ^ 1'b0 ;
  assign n13263 = n509 & ~n5794 ;
  assign n13264 = n5018 & ~n13263 ;
  assign n13265 = n3338 & n13264 ;
  assign n13266 = n2478 ^ n2467 ^ 1'b0 ;
  assign n13267 = n1913 & n5504 ;
  assign n13268 = n13267 ^ n4846 ^ 1'b0 ;
  assign n13269 = x119 & n13268 ;
  assign n13270 = n3035 & n13269 ;
  assign n13271 = n13270 ^ n978 ^ 1'b0 ;
  assign n13273 = n1808 | n1867 ;
  assign n13272 = ~n2928 & n7231 ;
  assign n13274 = n13273 ^ n13272 ^ 1'b0 ;
  assign n13275 = n11437 ^ n8675 ^ 1'b0 ;
  assign n13276 = ~n744 & n10554 ;
  assign n13277 = n13276 ^ n11082 ^ 1'b0 ;
  assign n13278 = n2606 & n3759 ;
  assign n13279 = ~n648 & n13278 ;
  assign n13280 = n6987 ^ n4457 ^ n3386 ;
  assign n13281 = n8326 | n11016 ;
  assign n13282 = n13281 ^ n9069 ^ 1'b0 ;
  assign n13285 = n11873 ^ n4814 ^ 1'b0 ;
  assign n13283 = ~n3729 & n5860 ;
  assign n13284 = ~n6850 & n13283 ;
  assign n13286 = n13285 ^ n13284 ^ 1'b0 ;
  assign n13287 = n6435 ^ n5779 ^ 1'b0 ;
  assign n13288 = n3217 & n4882 ;
  assign n13289 = ~n13287 & n13288 ;
  assign n13290 = ~n230 & n5159 ;
  assign n13291 = ~n2048 & n13290 ;
  assign n13292 = n5996 & ~n8596 ;
  assign n13293 = n6504 ^ n766 ^ 1'b0 ;
  assign n13294 = ~n921 & n13293 ;
  assign n13295 = n13294 ^ n6457 ^ 1'b0 ;
  assign n13296 = n3488 ^ n788 ^ 1'b0 ;
  assign n13297 = n13296 ^ n2848 ^ 1'b0 ;
  assign n13298 = n5923 | n13297 ;
  assign n13299 = ~x16 & n595 ;
  assign n13300 = n3482 ^ n1948 ^ 1'b0 ;
  assign n13301 = n6690 & n12969 ;
  assign n13302 = n6488 ^ n6324 ^ 1'b0 ;
  assign n13303 = x37 | n6519 ;
  assign n13304 = n1487 & ~n6324 ;
  assign n13305 = n4002 & n8079 ;
  assign n13306 = n5090 ^ n1414 ^ 1'b0 ;
  assign n13307 = ~n3677 & n13306 ;
  assign n13308 = n1420 & n10945 ;
  assign n13309 = n5278 & n13308 ;
  assign n13310 = n13309 ^ n7266 ^ 1'b0 ;
  assign n13311 = n2854 & ~n7498 ;
  assign n13312 = ~n6170 & n13311 ;
  assign n13313 = n13312 ^ n1122 ^ 1'b0 ;
  assign n13314 = n4218 & ~n6912 ;
  assign n13315 = n11496 | n13314 ;
  assign n13316 = n13315 ^ n8791 ^ 1'b0 ;
  assign n13317 = ~n5530 & n8185 ;
  assign n13318 = n9203 ^ n2978 ^ 1'b0 ;
  assign n13319 = n13317 & n13318 ;
  assign n13320 = n2091 | n5722 ;
  assign n13321 = n5274 | n5578 ;
  assign n13322 = n198 | n1561 ;
  assign n13323 = n13322 ^ n12251 ^ 1'b0 ;
  assign n13324 = ~n1258 & n3816 ;
  assign n13325 = n13324 ^ n1737 ^ 1'b0 ;
  assign n13326 = ~n753 & n13325 ;
  assign n13327 = n5089 & ~n7002 ;
  assign n13328 = n8707 & n13327 ;
  assign n13330 = n6242 ^ n3637 ^ 1'b0 ;
  assign n13329 = n4366 & n9865 ;
  assign n13331 = n13330 ^ n13329 ^ 1'b0 ;
  assign n13332 = n3672 ^ n390 ^ 1'b0 ;
  assign n13333 = n8799 ^ n5067 ^ 1'b0 ;
  assign n13334 = n13333 ^ n6669 ^ 1'b0 ;
  assign n13335 = x5 & x95 ;
  assign n13336 = ~x95 & n13335 ;
  assign n13337 = x25 & ~n13336 ;
  assign n13338 = n13336 & n13337 ;
  assign n13339 = x126 & ~n13338 ;
  assign n13340 = n13338 & n13339 ;
  assign n13341 = n304 & ~n13340 ;
  assign n13342 = ~n304 & n13341 ;
  assign n13343 = ~n134 & n179 ;
  assign n13344 = n134 & n13343 ;
  assign n13345 = n195 & ~n614 ;
  assign n13346 = ~n195 & n13345 ;
  assign n13347 = n338 | n13346 ;
  assign n13348 = n338 & ~n13347 ;
  assign n13349 = n13344 | n13348 ;
  assign n13350 = n13342 & ~n13349 ;
  assign n13351 = n13188 | n13350 ;
  assign n13352 = n13334 | n13351 ;
  assign n13353 = n12715 ^ n1711 ^ 1'b0 ;
  assign n13354 = n11662 | n13353 ;
  assign n13355 = n11474 | n13354 ;
  assign n13356 = n13355 ^ n4677 ^ 1'b0 ;
  assign n13357 = n13356 ^ n13053 ^ 1'b0 ;
  assign n13358 = n2330 & ~n13357 ;
  assign n13359 = n5967 ^ n1395 ^ 1'b0 ;
  assign n13360 = n2391 & ~n13359 ;
  assign n13361 = n5037 ^ n4900 ^ 1'b0 ;
  assign n13362 = n7512 ^ n4904 ^ 1'b0 ;
  assign n13363 = ~x53 & n335 ;
  assign n13364 = ~n164 & n13363 ;
  assign n13365 = n5685 & ~n13364 ;
  assign n13366 = n11499 ^ n4191 ^ n2542 ;
  assign n13367 = n12724 | n13366 ;
  assign n13368 = ~n6716 & n8020 ;
  assign n13369 = ~n914 & n13368 ;
  assign n13370 = n13369 ^ n5943 ^ 1'b0 ;
  assign n13371 = n3140 ^ n2490 ^ 1'b0 ;
  assign n13372 = n8022 & n10142 ;
  assign n13373 = n7162 & n12518 ;
  assign n13374 = n13373 ^ n2850 ^ 1'b0 ;
  assign n13381 = x119 & ~n8353 ;
  assign n13382 = n4931 & n13381 ;
  assign n13377 = n305 & ~n1086 ;
  assign n13378 = n13377 ^ n1054 ^ 1'b0 ;
  assign n13375 = n8806 ^ n2109 ^ 1'b0 ;
  assign n13376 = n822 & ~n13375 ;
  assign n13379 = n13378 ^ n13376 ^ n7153 ;
  assign n13380 = n2030 | n13379 ;
  assign n13383 = n13382 ^ n13380 ^ 1'b0 ;
  assign n13384 = n3764 | n13383 ;
  assign n13385 = n13384 ^ x70 ^ 1'b0 ;
  assign n13389 = n750 & ~n3037 ;
  assign n13386 = ~n344 & n4224 ;
  assign n13387 = n13386 ^ n12143 ^ 1'b0 ;
  assign n13388 = ~n1868 & n13387 ;
  assign n13390 = n13389 ^ n13388 ^ 1'b0 ;
  assign n13391 = n6575 & n7355 ;
  assign n13392 = n299 & ~n13391 ;
  assign n13393 = n7033 ^ n3377 ^ 1'b0 ;
  assign n13394 = n13393 ^ n5364 ^ 1'b0 ;
  assign n13395 = n3602 ^ n1372 ^ 1'b0 ;
  assign n13396 = ~n1194 & n13395 ;
  assign n13397 = ~n3512 & n13396 ;
  assign n13398 = n11775 ^ n7124 ^ 1'b0 ;
  assign n13399 = n9077 & n13398 ;
  assign n13400 = n3465 ^ n2448 ^ 1'b0 ;
  assign n13401 = ~n1563 & n13400 ;
  assign n13402 = ~n8251 & n13401 ;
  assign n13403 = n3800 & ~n7854 ;
  assign n13404 = n4433 & n13403 ;
  assign n13405 = n177 & ~n1363 ;
  assign n13406 = ~n177 & n13405 ;
  assign n13407 = ~n1158 & n2056 ;
  assign n13408 = n1158 & n13407 ;
  assign n13409 = n13406 | n13408 ;
  assign n13410 = n13406 & ~n13409 ;
  assign n13411 = n4554 | n13410 ;
  assign n13412 = n4554 & ~n13411 ;
  assign n13413 = n13412 ^ n10513 ^ 1'b0 ;
  assign n13414 = n13404 | n13413 ;
  assign n13415 = n13404 & ~n13414 ;
  assign n13416 = ~n5346 & n5425 ;
  assign n13417 = n3624 & ~n11135 ;
  assign n13418 = n13417 ^ n2944 ^ 1'b0 ;
  assign n13419 = n2592 & n11516 ;
  assign n13420 = n13419 ^ n6056 ^ 1'b0 ;
  assign n13421 = n13418 & ~n13420 ;
  assign n13422 = ~n4480 & n13421 ;
  assign n13423 = n221 | n6933 ;
  assign n13424 = n3585 & ~n10089 ;
  assign n13425 = n13424 ^ n8082 ^ 1'b0 ;
  assign n13426 = n5090 & ~n7594 ;
  assign n13427 = n13426 ^ n3509 ^ 1'b0 ;
  assign n13428 = ~n1004 & n13427 ;
  assign n13429 = n1837 & n5990 ;
  assign n13430 = n1937 ^ n432 ^ 1'b0 ;
  assign n13431 = n13429 & n13430 ;
  assign n13432 = ~n10932 & n13431 ;
  assign n13433 = n12971 & n13432 ;
  assign n13434 = n8316 ^ n3763 ^ 1'b0 ;
  assign n13435 = ~n6257 & n9120 ;
  assign n13436 = ~x58 & n13435 ;
  assign n13437 = n2079 ^ n1545 ^ 1'b0 ;
  assign n13438 = n2988 & ~n13437 ;
  assign n13439 = n1443 & n3534 ;
  assign n13440 = n13439 ^ n3872 ^ 1'b0 ;
  assign n13441 = n2603 ^ n297 ^ 1'b0 ;
  assign n13442 = n12466 | n13441 ;
  assign n13443 = n10776 ^ n1420 ^ 1'b0 ;
  assign n13444 = n2034 | n13443 ;
  assign n13445 = n2943 | n4806 ;
  assign n13446 = n13445 ^ n11597 ^ 1'b0 ;
  assign n13447 = ~n1487 & n6104 ;
  assign n13448 = n13447 ^ n3434 ^ n2694 ;
  assign n13449 = n3906 & ~n6175 ;
  assign n13450 = n2231 & n4045 ;
  assign n13451 = n13450 ^ n5609 ^ 1'b0 ;
  assign n13452 = n7362 & n9628 ;
  assign n13453 = ~n7063 & n7069 ;
  assign n13454 = ~n1376 & n6667 ;
  assign n13455 = ( n1128 & ~n3504 ) | ( n1128 & n6512 ) | ( ~n3504 & n6512 ) ;
  assign n13456 = n13455 ^ n7955 ^ n5064 ;
  assign n13457 = ~n516 & n13456 ;
  assign n13458 = x127 & n8082 ;
  assign n13459 = n13458 ^ n5702 ^ 1'b0 ;
  assign n13460 = n13459 ^ n2756 ^ 1'b0 ;
  assign n13461 = n9813 & n13460 ;
  assign n13462 = ~n9709 & n13461 ;
  assign n13463 = ~n13457 & n13462 ;
  assign n13464 = n1963 & n5072 ;
  assign n13465 = n482 & n13464 ;
  assign n13466 = n8427 & n13465 ;
  assign n13467 = n12510 & ~n13466 ;
  assign n13468 = n671 & n7777 ;
  assign n13469 = ~n7777 & n13468 ;
  assign n13470 = n6180 & ~n11862 ;
  assign n13471 = n3184 & ~n8670 ;
  assign n13472 = n492 | n3195 ;
  assign n13473 = n13472 ^ n8057 ^ n230 ;
  assign n13474 = x104 & ~n7226 ;
  assign n13475 = n13474 ^ n2666 ^ 1'b0 ;
  assign n13476 = ~n6436 & n13475 ;
  assign n13477 = n13476 ^ n242 ^ 1'b0 ;
  assign n13478 = n4001 & n5378 ;
  assign n13479 = n13478 ^ n11295 ^ 1'b0 ;
  assign n13480 = n10974 ^ n9815 ^ n3869 ;
  assign n13481 = n570 ^ n430 ^ 1'b0 ;
  assign n13482 = n8577 ^ n800 ^ 1'b0 ;
  assign n13483 = n13481 & ~n13482 ;
  assign n13484 = ~n6310 & n13320 ;
  assign n13485 = n1112 | n6570 ;
  assign n13486 = n3987 & ~n13485 ;
  assign n13487 = n3288 & n5724 ;
  assign n13488 = n5208 & n7055 ;
  assign n13489 = n4854 & ~n13488 ;
  assign n13490 = n1675 & n13489 ;
  assign n13491 = n9082 & ~n13490 ;
  assign n13492 = n6098 & n13491 ;
  assign n13493 = n6996 ^ n5227 ^ 1'b0 ;
  assign n13494 = n7926 & ~n11830 ;
  assign n13495 = n13494 ^ n3611 ^ 1'b0 ;
  assign n13496 = ~n7602 & n8827 ;
  assign n13497 = n698 & n10653 ;
  assign n13498 = n3563 & n13497 ;
  assign n13499 = n3917 & n6640 ;
  assign n13500 = n13499 ^ n10687 ^ 1'b0 ;
  assign n13501 = x120 & ~n13500 ;
  assign n13502 = n2921 & n13501 ;
  assign n13503 = n5834 ^ n1146 ^ 1'b0 ;
  assign n13504 = x12 & n13503 ;
  assign n13505 = n294 | n9725 ;
  assign n13506 = n7462 ^ n5349 ^ 1'b0 ;
  assign n13507 = ~n506 & n13506 ;
  assign n13508 = ~n391 & n3132 ;
  assign n13509 = n6979 & n11104 ;
  assign n13510 = ~n9511 & n13509 ;
  assign n13511 = n9964 ^ n6590 ^ n2259 ;
  assign n13512 = n4195 & ~n13511 ;
  assign n13513 = n3009 & n11201 ;
  assign n13514 = n13513 ^ n3275 ^ 1'b0 ;
  assign n13515 = n1052 | n11038 ;
  assign n13516 = n13515 ^ n4412 ^ 1'b0 ;
  assign n13517 = ~n4180 & n5889 ;
  assign n13518 = n747 | n13517 ;
  assign n13519 = n1181 | n1517 ;
  assign n13520 = n10458 ^ n1304 ^ 1'b0 ;
  assign n13521 = n7369 ^ n2271 ^ 1'b0 ;
  assign n13522 = n9846 ^ n2826 ^ 1'b0 ;
  assign n13524 = n245 | n5383 ;
  assign n13523 = ~n3992 & n11415 ;
  assign n13525 = n13524 ^ n13523 ^ 1'b0 ;
  assign n13526 = n5132 & n10998 ;
  assign n13527 = n13526 ^ n2921 ^ 1'b0 ;
  assign n13528 = n2686 ^ x109 ^ 1'b0 ;
  assign n13529 = n3280 | n7736 ;
  assign n13530 = n13529 ^ n6787 ^ 1'b0 ;
  assign n13531 = n684 | n13530 ;
  assign n13532 = n13531 ^ n5967 ^ 1'b0 ;
  assign n13533 = ~n13528 & n13532 ;
  assign n13535 = n5018 ^ n4511 ^ 1'b0 ;
  assign n13539 = x82 & n9045 ;
  assign n13536 = ~n4484 & n4771 ;
  assign n13537 = n13536 ^ n893 ^ 1'b0 ;
  assign n13538 = ~n983 & n13537 ;
  assign n13540 = n13539 ^ n13538 ^ 1'b0 ;
  assign n13541 = ~n13535 & n13540 ;
  assign n13534 = n4918 & n6665 ;
  assign n13542 = n13541 ^ n13534 ^ 1'b0 ;
  assign n13543 = n1952 & ~n4911 ;
  assign n13544 = n13543 ^ n9504 ^ 1'b0 ;
  assign n13545 = n13544 ^ n11651 ^ 1'b0 ;
  assign n13546 = n2199 & n13545 ;
  assign n13547 = n5973 | n9283 ;
  assign n13548 = n13547 ^ n6982 ^ 1'b0 ;
  assign n13549 = n13548 ^ n7760 ^ n2193 ;
  assign n13550 = n4169 & ~n7401 ;
  assign n13551 = n2843 & ~n7391 ;
  assign n13552 = n8245 & n13551 ;
  assign n13553 = n13552 ^ n3557 ^ 1'b0 ;
  assign n13554 = ~n12538 & n13553 ;
  assign n13555 = n5541 & n5837 ;
  assign n13556 = n13555 ^ n5248 ^ 1'b0 ;
  assign n13557 = n13556 ^ n11337 ^ 1'b0 ;
  assign n13558 = n8927 & n11459 ;
  assign n13559 = n1664 & n11310 ;
  assign n13560 = n13559 ^ n1249 ^ 1'b0 ;
  assign n13561 = ~n272 & n13560 ;
  assign n13562 = n1228 & n13561 ;
  assign n13563 = n11642 & n12821 ;
  assign n13564 = n4022 | n13563 ;
  assign n13565 = n5405 ^ n3960 ^ 1'b0 ;
  assign n13566 = n4958 & ~n13565 ;
  assign n13567 = ~n7899 & n13566 ;
  assign n13568 = n1593 ^ n825 ^ 1'b0 ;
  assign n13569 = n8691 ^ n2418 ^ 1'b0 ;
  assign n13570 = ~n292 & n1400 ;
  assign n13571 = ~n1400 & n13570 ;
  assign n13572 = ~n1089 & n1170 ;
  assign n13573 = n1089 & n13572 ;
  assign n13574 = x92 & ~n13573 ;
  assign n13575 = n13573 & n13574 ;
  assign n13576 = n13575 ^ n2203 ^ 1'b0 ;
  assign n13577 = n13576 ^ n6704 ^ 1'b0 ;
  assign n13578 = n13571 | n13577 ;
  assign n13579 = ~n1578 & n13578 ;
  assign n13580 = n4694 ^ n3359 ^ 1'b0 ;
  assign n13581 = ~n1845 & n13580 ;
  assign n13582 = n13581 ^ n8643 ^ 1'b0 ;
  assign n13583 = n167 | n13582 ;
  assign n13584 = n8185 ^ n6423 ^ 1'b0 ;
  assign n13585 = n9333 & n13584 ;
  assign n13587 = n1432 & n3245 ;
  assign n13588 = ~n3255 & n13587 ;
  assign n13586 = ~n2639 & n3695 ;
  assign n13589 = n13588 ^ n13586 ^ 1'b0 ;
  assign n13590 = n1054 & ~n9874 ;
  assign n13591 = n9340 ^ n1622 ^ 1'b0 ;
  assign n13592 = n409 | n13591 ;
  assign n13593 = n1063 ^ n1001 ^ 1'b0 ;
  assign n13594 = ~n287 & n13593 ;
  assign n13595 = n13066 & ~n13594 ;
  assign n13596 = n10223 & n10771 ;
  assign n13597 = ~n4967 & n6250 ;
  assign n13598 = n2453 & n13597 ;
  assign n13599 = n6684 ^ n921 ^ 1'b0 ;
  assign n13600 = n2285 & n13599 ;
  assign n13601 = n8387 ^ n3777 ^ 1'b0 ;
  assign n13602 = n2999 ^ x82 ^ 1'b0 ;
  assign n13603 = n13602 ^ n9512 ^ 1'b0 ;
  assign n13604 = n3045 | n3320 ;
  assign n13605 = n13604 ^ n9066 ^ 1'b0 ;
  assign n13606 = ~n1355 & n13605 ;
  assign n13607 = n4923 ^ n1724 ^ 1'b0 ;
  assign n13608 = n5927 | n13607 ;
  assign n13609 = n5526 & ~n7625 ;
  assign n13610 = ~n701 & n13609 ;
  assign n13611 = ( n4755 & n13608 ) | ( n4755 & ~n13610 ) | ( n13608 & ~n13610 ) ;
  assign n13612 = n13611 ^ n12041 ^ 1'b0 ;
  assign n13613 = n13606 & n13612 ;
  assign n13614 = n5132 & n13613 ;
  assign n13615 = n3126 ^ n2308 ^ 1'b0 ;
  assign n13616 = n4186 & n4311 ;
  assign n13617 = n1181 & n13616 ;
  assign n13618 = n13617 ^ n297 ^ 1'b0 ;
  assign n13619 = n5686 | n13618 ;
  assign n13620 = n13615 | n13619 ;
  assign n13621 = n13620 ^ n13499 ^ 1'b0 ;
  assign n13622 = n7867 ^ n2329 ^ 1'b0 ;
  assign n13623 = n1576 | n13622 ;
  assign n13624 = n1002 | n13623 ;
  assign n13625 = n8780 ^ n542 ^ 1'b0 ;
  assign n13626 = n4079 ^ n2083 ^ 1'b0 ;
  assign n13627 = ~n4847 & n13626 ;
  assign n13628 = n862 | n8506 ;
  assign n13629 = n3152 | n5450 ;
  assign n13630 = n5027 & ~n13629 ;
  assign n13631 = n5187 | n12604 ;
  assign n13632 = n970 | n5364 ;
  assign n13633 = n1728 | n13632 ;
  assign n13634 = ~n1722 & n13633 ;
  assign n13635 = n13634 ^ n8760 ^ 1'b0 ;
  assign n13636 = ~n5327 & n13635 ;
  assign n13637 = n13634 ^ n5068 ^ 1'b0 ;
  assign n13638 = ~n5689 & n7803 ;
  assign n13639 = n13638 ^ x118 ^ 1'b0 ;
  assign n13640 = ~n2440 & n5268 ;
  assign n13641 = n13639 & n13640 ;
  assign n13642 = n3454 ^ n1808 ^ n775 ;
  assign n13643 = n5825 & n13642 ;
  assign n13644 = n13004 ^ n9045 ^ 1'b0 ;
  assign n13645 = n13644 ^ n5943 ^ 1'b0 ;
  assign n13646 = n6223 & ~n12916 ;
  assign n13647 = x84 & n2604 ;
  assign n13648 = n13646 | n13647 ;
  assign n13649 = n5950 | n7672 ;
  assign n13650 = ~n4098 & n13649 ;
  assign n13651 = n13650 ^ n2883 ^ 1'b0 ;
  assign n13652 = n1702 ^ n859 ^ 1'b0 ;
  assign n13653 = n11505 & n13652 ;
  assign n13654 = n1228 & ~n5228 ;
  assign n13655 = n3615 & n13654 ;
  assign n13656 = n5258 & ~n13655 ;
  assign n13657 = ~n5202 & n11004 ;
  assign n13658 = n13543 ^ n8473 ^ n7438 ;
  assign n13659 = n9526 & ~n10023 ;
  assign n13660 = n10691 ^ x94 ^ 1'b0 ;
  assign n13661 = n1864 | n12631 ;
  assign n13662 = n3575 & n6935 ;
  assign n13663 = n1348 | n13662 ;
  assign n13664 = n159 & n6461 ;
  assign n13665 = ~n784 & n4873 ;
  assign n13666 = ~x75 & n13665 ;
  assign n13667 = n4197 | n13666 ;
  assign n13668 = n4081 ^ n2201 ^ 1'b0 ;
  assign n13669 = ~n1770 & n2006 ;
  assign n13670 = n13669 ^ n5096 ^ 1'b0 ;
  assign n13671 = n13670 ^ n3784 ^ 1'b0 ;
  assign n13672 = n11787 ^ n10470 ^ 1'b0 ;
  assign n13673 = ~n6078 & n13672 ;
  assign n13674 = n7037 & ~n10027 ;
  assign n13675 = n10978 & n13674 ;
  assign n13676 = n5442 ^ x29 ^ 1'b0 ;
  assign n13677 = n851 & n13676 ;
  assign n13678 = ~n5562 & n13677 ;
  assign n13679 = n994 & ~n3833 ;
  assign n13680 = n13679 ^ n2634 ^ 1'b0 ;
  assign n13681 = n10932 ^ n3415 ^ 1'b0 ;
  assign n13682 = n7146 ^ n4757 ^ 1'b0 ;
  assign n13683 = ~n11624 & n13682 ;
  assign n13684 = x52 & n1056 ;
  assign n13685 = n8578 & ~n13039 ;
  assign n13686 = n13685 ^ n363 ^ 1'b0 ;
  assign n13687 = n13684 | n13686 ;
  assign n13688 = n13521 & ~n13687 ;
  assign n13689 = n6291 ^ n2741 ^ 1'b0 ;
  assign n13690 = n3994 & ~n13689 ;
  assign n13691 = n1506 & n7530 ;
  assign n13692 = n3458 & ~n6760 ;
  assign n13693 = ~n7280 & n13692 ;
  assign n13694 = n5143 & ~n6578 ;
  assign n13695 = ~n3335 & n13694 ;
  assign n13696 = ~n8048 & n13695 ;
  assign n13697 = n3012 & ~n3526 ;
  assign n13698 = n1918 & n13697 ;
  assign n13699 = n3968 & ~n5265 ;
  assign n13700 = n5731 ^ n1908 ^ 1'b0 ;
  assign n13701 = n13699 | n13700 ;
  assign n13702 = n13701 ^ n950 ^ 1'b0 ;
  assign n13703 = n6855 | n13702 ;
  assign n13704 = n4110 & ~n13703 ;
  assign n13705 = ~n8028 & n12848 ;
  assign n13706 = n13705 ^ n7381 ^ 1'b0 ;
  assign n13707 = ( ~n3393 & n5337 ) | ( ~n3393 & n13503 ) | ( n5337 & n13503 ) ;
  assign n13708 = ~n4350 & n8927 ;
  assign n13709 = n13707 & n13708 ;
  assign n13710 = n2859 ^ n2399 ^ 1'b0 ;
  assign n13711 = n8954 & n13710 ;
  assign n13712 = ~n7137 & n13711 ;
  assign n13713 = ~n4227 & n13712 ;
  assign n13714 = n13713 ^ n1245 ^ 1'b0 ;
  assign n13715 = n8767 ^ n7627 ^ 1'b0 ;
  assign n13716 = n13715 ^ n4248 ^ 1'b0 ;
  assign n13717 = ~n553 & n7089 ;
  assign n13718 = ~n1916 & n13717 ;
  assign n13719 = ( ~n3438 & n13716 ) | ( ~n3438 & n13718 ) | ( n13716 & n13718 ) ;
  assign n13720 = n8861 | n9898 ;
  assign n13721 = n13036 & ~n13720 ;
  assign n13722 = n2159 | n13721 ;
  assign n13723 = n13722 ^ n2288 ^ 1'b0 ;
  assign n13724 = n5880 ^ n5519 ^ 1'b0 ;
  assign n13726 = n6448 ^ n4916 ^ 1'b0 ;
  assign n13727 = n4554 ^ n194 ^ 1'b0 ;
  assign n13728 = ~n1830 & n13727 ;
  assign n13729 = ~n13726 & n13728 ;
  assign n13725 = x60 | n4449 ;
  assign n13730 = n13729 ^ n13725 ^ 1'b0 ;
  assign n13731 = ( ~n930 & n2930 ) | ( ~n930 & n3637 ) | ( n2930 & n3637 ) ;
  assign n13732 = n361 & n4311 ;
  assign n13733 = n13732 ^ n336 ^ 1'b0 ;
  assign n13734 = n1853 & n7523 ;
  assign n13737 = n1202 | n4701 ;
  assign n13735 = ~n1258 & n2087 ;
  assign n13736 = n13049 & n13735 ;
  assign n13738 = n13737 ^ n13736 ^ 1'b0 ;
  assign n13739 = n2637 | n10596 ;
  assign n13740 = n1609 ^ n550 ^ 1'b0 ;
  assign n13741 = n2866 | n13740 ;
  assign n13742 = ~n201 & n7441 ;
  assign n13743 = ~n2369 & n10773 ;
  assign n13744 = n13743 ^ n13455 ^ 1'b0 ;
  assign n13745 = ~n7182 & n9224 ;
  assign n13746 = ~n13246 & n13745 ;
  assign n13747 = n1952 & n13746 ;
  assign n13751 = n514 | n5571 ;
  assign n13748 = n4598 & n4901 ;
  assign n13749 = ~n12178 & n13748 ;
  assign n13750 = n10857 & ~n13749 ;
  assign n13752 = n13751 ^ n13750 ^ 1'b0 ;
  assign n13758 = ~n542 & n3156 ;
  assign n13753 = n4660 ^ n321 ^ 1'b0 ;
  assign n13754 = n3947 & ~n13753 ;
  assign n13755 = n5418 & n13754 ;
  assign n13756 = n13755 ^ x44 ^ 1'b0 ;
  assign n13757 = n6871 & ~n13756 ;
  assign n13759 = n13758 ^ n13757 ^ 1'b0 ;
  assign n13760 = ~n2566 & n8059 ;
  assign n13761 = n696 & n13760 ;
  assign n13762 = n2283 ^ n287 ^ 1'b0 ;
  assign n13763 = n13761 | n13762 ;
  assign n13764 = n264 & ~n3834 ;
  assign n13765 = ~n2354 & n13764 ;
  assign n13766 = n4033 | n13765 ;
  assign n13767 = n9170 | n13766 ;
  assign n13768 = n13767 ^ n8508 ^ 1'b0 ;
  assign n13769 = ~n3737 & n13768 ;
  assign n13770 = n1963 ^ x11 ^ 1'b0 ;
  assign n13771 = n2136 & ~n9143 ;
  assign n13772 = ~n3186 & n13771 ;
  assign n13773 = n13772 ^ n7167 ^ 1'b0 ;
  assign n13774 = n13770 & n13773 ;
  assign n13775 = n6504 ^ n254 ^ 1'b0 ;
  assign n13776 = ~n3019 & n13775 ;
  assign n13777 = n8148 & n13776 ;
  assign n13778 = n11472 ^ n5987 ^ 1'b0 ;
  assign n13779 = n5338 & n13778 ;
  assign n13780 = ~n8079 & n13779 ;
  assign n13781 = n5564 & ~n8775 ;
  assign n13782 = n1101 | n3548 ;
  assign n13783 = n4289 & n13782 ;
  assign n13784 = n12298 ^ n11407 ^ 1'b0 ;
  assign n13785 = n2847 | n13784 ;
  assign n13786 = n6321 ^ n3548 ^ 1'b0 ;
  assign n13787 = n1160 & n13786 ;
  assign n13788 = n1987 & ~n2089 ;
  assign n13789 = n678 & ~n13788 ;
  assign n13790 = n2087 & ~n9382 ;
  assign n13791 = n13790 ^ n11885 ^ 1'b0 ;
  assign n13792 = ~n11354 & n13791 ;
  assign n13793 = ~x74 & n13792 ;
  assign n13794 = ~n13789 & n13793 ;
  assign n13795 = n12408 ^ n516 ^ 1'b0 ;
  assign n13796 = n6607 & ~n13795 ;
  assign n13797 = n13796 ^ n7719 ^ 1'b0 ;
  assign n13798 = n217 & n13797 ;
  assign n13799 = n10240 ^ n1680 ^ 1'b0 ;
  assign n13800 = n13799 ^ n8361 ^ n7251 ;
  assign n13801 = n6599 & ~n11272 ;
  assign n13802 = n13801 ^ n4674 ^ 1'b0 ;
  assign n13803 = n3166 ^ n2682 ^ 1'b0 ;
  assign n13804 = n13803 ^ n2200 ^ 1'b0 ;
  assign n13805 = n13802 | n13804 ;
  assign n13806 = n246 & n6575 ;
  assign n13807 = n13806 ^ n1758 ^ 1'b0 ;
  assign n13808 = n13807 ^ n11348 ^ 1'b0 ;
  assign n13809 = n483 & n13808 ;
  assign n13810 = n237 & n5745 ;
  assign n13811 = ~n6054 & n13810 ;
  assign n13812 = n7057 ^ n6045 ^ 1'b0 ;
  assign n13813 = n13811 | n13812 ;
  assign n13814 = ~n6425 & n8693 ;
  assign n13815 = n10702 & n13814 ;
  assign n13816 = n1996 | n2091 ;
  assign n13817 = n10698 ^ n7407 ^ 1'b0 ;
  assign n13818 = n3278 & ~n13817 ;
  assign n13819 = ~n3855 & n13818 ;
  assign n13820 = n13819 ^ x66 ^ 1'b0 ;
  assign n13821 = n1189 & n13820 ;
  assign n13822 = n1070 | n1277 ;
  assign n13823 = n9349 ^ n5674 ^ 1'b0 ;
  assign n13824 = n2481 | n4363 ;
  assign n13825 = n6883 ^ n896 ^ 1'b0 ;
  assign n13826 = ~n2082 & n13825 ;
  assign n13827 = n672 ^ n516 ^ 1'b0 ;
  assign n13828 = n507 & ~n13827 ;
  assign n13829 = n12375 & ~n13828 ;
  assign n13830 = n3507 ^ n3428 ^ 1'b0 ;
  assign n13831 = n2673 & n13830 ;
  assign n13832 = n9736 | n13321 ;
  assign n13833 = n6181 | n9292 ;
  assign n13834 = n2566 ^ n1235 ^ 1'b0 ;
  assign n13835 = n3482 & ~n13834 ;
  assign n13836 = n753 & ~n5629 ;
  assign n13837 = n13835 & ~n13836 ;
  assign n13838 = n2093 & n4991 ;
  assign n13839 = n13838 ^ n1419 ^ 1'b0 ;
  assign n13840 = n6451 & n7843 ;
  assign n13841 = n5652 ^ n4643 ^ 1'b0 ;
  assign n13842 = n13841 ^ n6059 ^ 1'b0 ;
  assign n13843 = n7052 & ~n13842 ;
  assign n13844 = ~n8024 & n13843 ;
  assign n13845 = n10583 ^ n4873 ^ 1'b0 ;
  assign n13846 = ( ~n3291 & n7489 ) | ( ~n3291 & n13845 ) | ( n7489 & n13845 ) ;
  assign n13847 = n3545 ^ n1973 ^ 1'b0 ;
  assign n13848 = n13847 ^ n6012 ^ 1'b0 ;
  assign n13849 = n2733 | n13848 ;
  assign n13850 = ~n1244 & n11505 ;
  assign n13851 = ~n177 & n13850 ;
  assign n13852 = n3970 & ~n9910 ;
  assign n13853 = n13851 & n13852 ;
  assign n13854 = ~n12319 & n12790 ;
  assign n13855 = n8704 ^ n7247 ^ 1'b0 ;
  assign n13856 = n6610 & n13855 ;
  assign n13858 = n1517 & n3096 ;
  assign n13857 = n3295 | n8777 ;
  assign n13859 = n13858 ^ n13857 ^ 1'b0 ;
  assign n13860 = n5418 & ~n10859 ;
  assign n13861 = n13860 ^ n8217 ^ 1'b0 ;
  assign n13862 = n467 & n4220 ;
  assign n13863 = n466 & n13862 ;
  assign n13864 = n13863 ^ n428 ^ 1'b0 ;
  assign n13866 = n550 & ~n1475 ;
  assign n13865 = n2561 | n2819 ;
  assign n13867 = n13866 ^ n13865 ^ 1'b0 ;
  assign n13868 = n6732 & ~n13867 ;
  assign n13869 = n9895 & n13868 ;
  assign n13870 = n3949 | n13869 ;
  assign n13871 = n13864 & ~n13870 ;
  assign n13872 = n3338 ^ n2438 ^ 1'b0 ;
  assign n13873 = n2395 & n3347 ;
  assign n13875 = n4373 & n9702 ;
  assign n13874 = n4602 & ~n6664 ;
  assign n13876 = n13875 ^ n13874 ^ 1'b0 ;
  assign n13877 = n6423 ^ n4335 ^ 1'b0 ;
  assign n13878 = n13877 ^ n12045 ^ 1'b0 ;
  assign n13879 = ~n129 & n3719 ;
  assign n13880 = n7469 & n13879 ;
  assign n13881 = n7179 ^ n5664 ^ 1'b0 ;
  assign n13882 = n2051 | n13881 ;
  assign n13884 = n1595 & ~n2496 ;
  assign n13885 = n4253 | n13884 ;
  assign n13883 = x75 & ~n2761 ;
  assign n13886 = n13885 ^ n13883 ^ 1'b0 ;
  assign n13887 = n13886 ^ n5395 ^ 1'b0 ;
  assign n13888 = n13882 | n13887 ;
  assign n13889 = n7426 ^ n6154 ^ 1'b0 ;
  assign n13890 = ~n696 & n6232 ;
  assign n13891 = ~n11380 & n13890 ;
  assign n13892 = n7716 & ~n13891 ;
  assign n13893 = n13889 & n13892 ;
  assign n13894 = x41 & n4086 ;
  assign n13895 = ~n2377 & n13894 ;
  assign n13896 = n13877 & ~n13895 ;
  assign n13897 = n4027 ^ n2198 ^ 1'b0 ;
  assign n13898 = n10489 ^ n9161 ^ 1'b0 ;
  assign n13899 = n13898 ^ n11842 ^ n2881 ;
  assign n13900 = n3283 & ~n13899 ;
  assign n13901 = n11512 ^ n2935 ^ 1'b0 ;
  assign n13902 = ~n568 & n2786 ;
  assign n13903 = n12685 & n13902 ;
  assign n13904 = n2427 ^ n171 ^ 1'b0 ;
  assign n13905 = ~n3221 & n13904 ;
  assign n13906 = n12352 ^ n1883 ^ 1'b0 ;
  assign n13907 = n13905 & n13906 ;
  assign n13908 = ~n2936 & n6478 ;
  assign n13909 = n6330 | n11891 ;
  assign n13910 = n9083 ^ n811 ^ 1'b0 ;
  assign n13911 = n4706 & ~n5882 ;
  assign n13912 = n13911 ^ n3658 ^ 1'b0 ;
  assign n13913 = n4056 | n4641 ;
  assign n13914 = n5651 | n13913 ;
  assign n13915 = n13914 ^ n9554 ^ 1'b0 ;
  assign n13916 = ~n8596 & n13915 ;
  assign n13917 = n3651 & n7719 ;
  assign n13918 = ~n13916 & n13917 ;
  assign n13919 = n3063 & ~n12761 ;
  assign n13920 = n4113 & ~n9391 ;
  assign n13921 = n13920 ^ n6206 ^ 1'b0 ;
  assign n13922 = ( n1011 & n7969 ) | ( n1011 & ~n13921 ) | ( n7969 & ~n13921 ) ;
  assign n13923 = n1316 & ~n10132 ;
  assign n13924 = ~x115 & n13923 ;
  assign n13925 = n13924 ^ n6268 ^ 1'b0 ;
  assign n13926 = n6145 & n6239 ;
  assign n13927 = n5927 & n13926 ;
  assign n13928 = n11601 ^ n9368 ^ 1'b0 ;
  assign n13929 = n1001 | n13928 ;
  assign n13930 = n12001 & ~n13929 ;
  assign n13931 = ~n3818 & n13930 ;
  assign n13932 = n1616 & ~n13931 ;
  assign n13933 = n1774 & ~n12936 ;
  assign n13934 = ~n5038 & n13933 ;
  assign n13935 = n13934 ^ n8664 ^ 1'b0 ;
  assign n13936 = n12936 ^ n4206 ^ 1'b0 ;
  assign n13937 = n5470 & n13936 ;
  assign n13938 = n9246 ^ n7898 ^ n6067 ;
  assign n13939 = ~n1395 & n1867 ;
  assign n13940 = n7752 & n11320 ;
  assign n13941 = ~n4935 & n9573 ;
  assign n13942 = n1016 & n13941 ;
  assign n13944 = n3807 ^ n1470 ^ 1'b0 ;
  assign n13943 = n2859 & ~n9103 ;
  assign n13945 = n13944 ^ n13943 ^ 1'b0 ;
  assign n13946 = n5491 & ~n11850 ;
  assign n13947 = n6994 | n13946 ;
  assign n13948 = n10259 ^ n8533 ^ 1'b0 ;
  assign n13949 = n6175 & ~n6829 ;
  assign n13950 = n9526 ^ n6840 ^ 1'b0 ;
  assign n13951 = x22 & n4444 ;
  assign n13952 = n13951 ^ n6321 ^ 1'b0 ;
  assign n13953 = ~x35 & x101 ;
  assign n13954 = n8881 & ~n13953 ;
  assign n13955 = n13954 ^ n1042 ^ 1'b0 ;
  assign n13956 = n2537 | n13955 ;
  assign n13957 = n13952 | n13956 ;
  assign n13958 = n7280 & n13269 ;
  assign n13959 = n8627 | n13958 ;
  assign n13960 = n485 & n520 ;
  assign n13961 = n13960 ^ n1327 ^ 1'b0 ;
  assign n13962 = n5204 ^ n4212 ^ 1'b0 ;
  assign n13963 = n2260 & n13962 ;
  assign n13964 = ~n6201 & n13963 ;
  assign n13965 = n5976 & n8111 ;
  assign n13966 = n13965 ^ n2664 ^ 1'b0 ;
  assign n13967 = n4296 & ~n13966 ;
  assign n13968 = ~n4311 & n13967 ;
  assign n13969 = n9502 ^ n1079 ^ 1'b0 ;
  assign n13970 = n900 & ~n13969 ;
  assign n13971 = n1543 | n5695 ;
  assign n13972 = n643 | n13971 ;
  assign n13973 = n5327 & ~n13972 ;
  assign n13974 = n5388 ^ n1576 ^ 1'b0 ;
  assign n13975 = n922 | n5836 ;
  assign n13976 = n13975 ^ n12682 ^ 1'b0 ;
  assign n13977 = n13974 & ~n13976 ;
  assign n13978 = n13977 ^ n2161 ^ 1'b0 ;
  assign n13979 = n10123 ^ n6675 ^ 1'b0 ;
  assign n13980 = n13049 & ~n13979 ;
  assign n13984 = n571 | n3251 ;
  assign n13985 = n13984 ^ n487 ^ 1'b0 ;
  assign n13981 = n7215 & n11295 ;
  assign n13982 = ~n11137 & n13981 ;
  assign n13983 = n13982 ^ n4025 ^ 1'b0 ;
  assign n13986 = n13985 ^ n13983 ^ 1'b0 ;
  assign n13987 = n6797 | n13986 ;
  assign n13988 = n1226 | n13974 ;
  assign n13989 = n7986 ^ n1899 ^ 1'b0 ;
  assign n13990 = n2289 & n13989 ;
  assign n13991 = n3474 ^ n1101 ^ 1'b0 ;
  assign n13992 = n1026 & ~n7283 ;
  assign n13993 = ~n667 & n13992 ;
  assign n13994 = n7446 & ~n13993 ;
  assign n13995 = n13994 ^ n3919 ^ 1'b0 ;
  assign n13997 = n4341 ^ n2843 ^ 1'b0 ;
  assign n13998 = n1651 | n13997 ;
  assign n13996 = n8590 ^ n3949 ^ 1'b0 ;
  assign n13999 = n13998 ^ n13996 ^ 1'b0 ;
  assign n14000 = n11649 ^ n4602 ^ 1'b0 ;
  assign n14001 = ~n4687 & n7539 ;
  assign n14002 = n351 & n1329 ;
  assign n14003 = n11329 & ~n14002 ;
  assign n14009 = n2094 & n4505 ;
  assign n14004 = n6985 & n12855 ;
  assign n14005 = n4089 & n14004 ;
  assign n14006 = n7453 & ~n8242 ;
  assign n14007 = x3 & n14006 ;
  assign n14008 = n14005 & n14007 ;
  assign n14010 = n14009 ^ n14008 ^ 1'b0 ;
  assign n14011 = n3888 & ~n8972 ;
  assign n14012 = ~n3826 & n14011 ;
  assign n14013 = n1737 & n6240 ;
  assign n14014 = n4545 ^ n302 ^ 1'b0 ;
  assign n14016 = n2091 & ~n4282 ;
  assign n14017 = ~n2091 & n14016 ;
  assign n14018 = n14017 ^ n7193 ^ 1'b0 ;
  assign n14015 = ( ~n6559 & n9454 ) | ( ~n6559 & n12762 ) | ( n9454 & n12762 ) ;
  assign n14019 = n14018 ^ n14015 ^ 1'b0 ;
  assign n14020 = n14014 & n14019 ;
  assign n14021 = ~n3784 & n12841 ;
  assign n14022 = n3045 & ~n8502 ;
  assign n14023 = n5112 & n6945 ;
  assign n14024 = n14023 ^ n7837 ^ 1'b0 ;
  assign n14025 = n14024 ^ n1508 ^ 1'b0 ;
  assign n14026 = n14022 & n14025 ;
  assign n14027 = n12351 ^ n1241 ^ 1'b0 ;
  assign n14028 = n4883 ^ n3542 ^ 1'b0 ;
  assign n14029 = n14028 ^ n11710 ^ 1'b0 ;
  assign n14030 = n7523 | n14029 ;
  assign n14031 = ~x14 & n13285 ;
  assign n14032 = n10086 | n14031 ;
  assign n14033 = n8682 & n14032 ;
  assign n14034 = n978 | n7141 ;
  assign n14035 = n10422 | n14034 ;
  assign n14036 = n5154 ^ n1226 ^ 1'b0 ;
  assign n14037 = n3245 & n10768 ;
  assign n14038 = n14037 ^ n2928 ^ 1'b0 ;
  assign n14039 = n4812 ^ n1106 ^ 1'b0 ;
  assign n14040 = n11164 & n14039 ;
  assign n14041 = ~n14038 & n14040 ;
  assign n14042 = ~n354 & n9539 ;
  assign n14043 = n2667 & n3961 ;
  assign n14044 = ~n231 & n14043 ;
  assign n14045 = n14044 ^ n1110 ^ n1080 ;
  assign n14046 = n7199 & n14045 ;
  assign n14047 = n9433 ^ n962 ^ 1'b0 ;
  assign n14048 = ~n11968 & n14047 ;
  assign n14049 = ~n14046 & n14048 ;
  assign n14050 = n7488 & n7780 ;
  assign n14051 = n14050 ^ n8374 ^ n363 ;
  assign n14052 = n3223 | n13219 ;
  assign n14053 = n10562 | n14052 ;
  assign n14054 = n10963 & n14053 ;
  assign n14055 = ~n2967 & n3098 ;
  assign n14056 = n3760 & n14055 ;
  assign n14058 = n7545 ^ n2309 ^ 1'b0 ;
  assign n14057 = n12364 ^ n1080 ^ 1'b0 ;
  assign n14059 = n14058 ^ n14057 ^ 1'b0 ;
  assign n14060 = ~n14056 & n14059 ;
  assign n14061 = n3105 ^ n2315 ^ 1'b0 ;
  assign n14062 = n14061 ^ n9686 ^ 1'b0 ;
  assign n14063 = n1033 | n14062 ;
  assign n14064 = n6371 & ~n14063 ;
  assign n14065 = n7592 & ~n12013 ;
  assign n14066 = ~n6180 & n14065 ;
  assign n14067 = n3797 & n6718 ;
  assign n14068 = n1993 & n4083 ;
  assign n14069 = n5630 & n14068 ;
  assign n14070 = ~n2966 & n9667 ;
  assign n14071 = ~n1235 & n2602 ;
  assign n14072 = n3152 | n7297 ;
  assign n14073 = n7848 ^ n2208 ^ 1'b0 ;
  assign n14074 = n588 & n7902 ;
  assign n14075 = n14074 ^ n7518 ^ 1'b0 ;
  assign n14076 = n14073 & ~n14075 ;
  assign n14077 = n14076 ^ n2389 ^ 1'b0 ;
  assign n14078 = n444 & n9845 ;
  assign n14079 = n3079 & ~n6495 ;
  assign n14080 = n14079 ^ n6711 ^ 1'b0 ;
  assign n14081 = ~n6064 & n14080 ;
  assign n14082 = n10184 & ~n10263 ;
  assign n14083 = ~n2108 & n6727 ;
  assign n14084 = ~n8760 & n14083 ;
  assign n14085 = n5761 & n5996 ;
  assign n14086 = n8785 ^ n3557 ^ 1'b0 ;
  assign n14087 = n14085 | n14086 ;
  assign n14088 = n5704 ^ n1284 ^ 1'b0 ;
  assign n14089 = n14087 | n14088 ;
  assign n14090 = n1079 & n3696 ;
  assign n14091 = n14090 ^ n7393 ^ 1'b0 ;
  assign n14092 = n4627 | n8056 ;
  assign n14093 = ( n2486 & ~n4623 ) | ( n2486 & n14092 ) | ( ~n4623 & n14092 ) ;
  assign n14094 = n6366 ^ n1781 ^ 1'b0 ;
  assign n14095 = n5990 & ~n12047 ;
  assign n14096 = n3396 & n14095 ;
  assign n14097 = ~x55 & n14096 ;
  assign n14098 = n1203 & n12859 ;
  assign n14099 = n216 | n5773 ;
  assign n14100 = n5773 & ~n14099 ;
  assign n14101 = ~n1025 & n14100 ;
  assign n14102 = n2947 & ~n14101 ;
  assign n14103 = n4534 ^ n707 ^ 1'b0 ;
  assign n14104 = n14103 ^ n2835 ^ 1'b0 ;
  assign n14105 = n14102 | n14104 ;
  assign n14106 = n9340 & n14105 ;
  assign n14107 = n14106 ^ n12579 ^ 1'b0 ;
  assign n14108 = n6719 & n7174 ;
  assign n14109 = n2030 ^ n909 ^ 1'b0 ;
  assign n14110 = n3483 & n14109 ;
  assign n14111 = ~n10756 & n14110 ;
  assign n14112 = n1982 | n4208 ;
  assign n14113 = n10281 & ~n14112 ;
  assign n14114 = n14113 ^ n9056 ^ 1'b0 ;
  assign n14115 = n10069 ^ x73 ^ 1'b0 ;
  assign n14116 = n11145 | n14115 ;
  assign n14117 = n2681 ^ n2040 ^ 1'b0 ;
  assign n14118 = n13788 ^ n8888 ^ 1'b0 ;
  assign n14119 = n304 & n14118 ;
  assign n14120 = n14119 ^ n13882 ^ 1'b0 ;
  assign n14121 = n1854 | n8353 ;
  assign n14122 = ~n346 & n9433 ;
  assign n14123 = n11905 & n14122 ;
  assign n14124 = n6265 | n14123 ;
  assign n14125 = n7002 | n8968 ;
  assign n14126 = n10329 ^ n7078 ^ n6848 ;
  assign n14127 = n2923 & n8762 ;
  assign n14128 = n14127 ^ n10589 ^ 1'b0 ;
  assign n14129 = n501 | n14128 ;
  assign n14130 = x50 | n14129 ;
  assign n14131 = ~n11414 & n12535 ;
  assign n14132 = ~n192 & n7166 ;
  assign n14133 = ~n7143 & n14132 ;
  assign n14134 = n1604 | n1652 ;
  assign n14135 = n14134 ^ n1677 ^ 1'b0 ;
  assign n14136 = n7029 & n13402 ;
  assign n14137 = ~n14135 & n14136 ;
  assign n14138 = n5667 ^ n4032 ^ 1'b0 ;
  assign n14139 = n11064 | n14138 ;
  assign n14140 = n7537 ^ n1880 ^ n1722 ;
  assign n14141 = n2213 & n14140 ;
  assign n14142 = n14141 ^ n6975 ^ 1'b0 ;
  assign n14143 = ~n2557 & n3575 ;
  assign n14144 = n724 & n14143 ;
  assign n14145 = n481 & n8157 ;
  assign n14146 = n6250 | n14145 ;
  assign n14147 = n1948 & n1983 ;
  assign n14148 = n2815 ^ n835 ^ 1'b0 ;
  assign n14149 = n14147 & ~n14148 ;
  assign n14150 = n14149 ^ n9987 ^ 1'b0 ;
  assign n14151 = n5522 & n14150 ;
  assign n14152 = n4436 & ~n6115 ;
  assign n14153 = n1091 & n14152 ;
  assign n14154 = n6197 ^ n870 ^ 1'b0 ;
  assign n14155 = ~n2241 & n7888 ;
  assign n14156 = ~n1841 & n4177 ;
  assign n14157 = n896 | n14156 ;
  assign n14158 = n14157 ^ n5927 ^ 1'b0 ;
  assign n14159 = n6417 ^ n5363 ^ 1'b0 ;
  assign n14160 = n10184 ^ n3128 ^ 1'b0 ;
  assign n14161 = n1937 | n8945 ;
  assign n14162 = n1098 & n10145 ;
  assign n14163 = n2647 & ~n9289 ;
  assign n14164 = n4500 ^ n1446 ^ 1'b0 ;
  assign n14165 = n530 & n14164 ;
  assign n14166 = ~n14163 & n14165 ;
  assign n14167 = n1925 | n6998 ;
  assign n14168 = n360 & ~n14167 ;
  assign n14169 = n4941 ^ x34 ^ 1'b0 ;
  assign n14170 = ~n5982 & n8514 ;
  assign n14171 = n12809 ^ n4671 ^ 1'b0 ;
  assign n14172 = ~n12101 & n14171 ;
  assign n14173 = n1062 | n11921 ;
  assign n14174 = n14173 ^ n4618 ^ 1'b0 ;
  assign n14175 = n13527 ^ n3678 ^ 1'b0 ;
  assign n14176 = ~n8249 & n9265 ;
  assign n14177 = ~n3038 & n14176 ;
  assign n14178 = n12089 ^ n2161 ^ 1'b0 ;
  assign n14179 = n493 & ~n3848 ;
  assign n14180 = n14179 ^ n13395 ^ 1'b0 ;
  assign n14181 = n3754 & n13464 ;
  assign n14182 = n221 & ~n267 ;
  assign n14183 = ~n694 & n955 ;
  assign n14184 = ~n4816 & n14183 ;
  assign n14185 = n14182 & n14184 ;
  assign n14186 = n8731 & ~n10147 ;
  assign n14187 = n4135 & ~n13383 ;
  assign n14188 = ~n673 & n3224 ;
  assign n14189 = n1666 & n14188 ;
  assign n14190 = n14189 ^ n7658 ^ n810 ;
  assign n14191 = n6281 ^ n884 ^ 1'b0 ;
  assign n14192 = ~n5300 & n8838 ;
  assign n14193 = n14192 ^ n13880 ^ 1'b0 ;
  assign n14194 = n1648 | n11505 ;
  assign n14195 = n14194 ^ n879 ^ 1'b0 ;
  assign n14196 = ~n701 & n1380 ;
  assign n14197 = n8773 & n14196 ;
  assign n14198 = n14197 ^ n4415 ^ 1'b0 ;
  assign n14199 = ~n2752 & n7739 ;
  assign n14200 = n14199 ^ n11253 ^ 1'b0 ;
  assign n14201 = ~n300 & n10147 ;
  assign n14202 = n14200 & n14201 ;
  assign n14203 = n2465 ^ n296 ^ 1'b0 ;
  assign n14204 = n2148 & n14203 ;
  assign n14205 = n14202 & n14204 ;
  assign n14206 = n14205 ^ n10435 ^ 1'b0 ;
  assign n14207 = n7087 & ~n14206 ;
  assign n14208 = n870 & ~n4819 ;
  assign n14209 = n14208 ^ n1765 ^ 1'b0 ;
  assign n14210 = n4053 & n7449 ;
  assign n14211 = n14210 ^ n2469 ^ 1'b0 ;
  assign n14212 = ~n2775 & n14211 ;
  assign n14213 = n8492 ^ x82 ^ 1'b0 ;
  assign n14214 = n2267 & n14213 ;
  assign n14215 = n7891 ^ n868 ^ 1'b0 ;
  assign n14216 = n1080 | n14215 ;
  assign n14217 = n2315 & ~n12859 ;
  assign n14218 = n7137 & n14217 ;
  assign n14219 = ~n227 & n1073 ;
  assign n14220 = ~n6044 & n14219 ;
  assign n14221 = n1281 | n1499 ;
  assign n14222 = n12181 ^ n12082 ^ n3096 ;
  assign n14223 = n14221 | n14222 ;
  assign n14229 = n10629 ^ n8695 ^ 1'b0 ;
  assign n14226 = n998 & ~n2041 ;
  assign n14227 = ~n14106 & n14226 ;
  assign n14228 = n7996 & ~n14227 ;
  assign n14224 = n14118 ^ n2565 ^ 1'b0 ;
  assign n14225 = ~n1961 & n14224 ;
  assign n14230 = n14229 ^ n14228 ^ n14225 ;
  assign n14231 = ( n3876 & n4916 ) | ( n3876 & n7830 ) | ( n4916 & n7830 ) ;
  assign n14232 = n7204 | n11535 ;
  assign n14233 = n1226 | n14232 ;
  assign n14234 = n1710 & n2143 ;
  assign n14235 = n14234 ^ x12 ^ 1'b0 ;
  assign n14236 = n9916 ^ n3633 ^ n2165 ;
  assign n14237 = n4227 & ~n14236 ;
  assign n14238 = ( n2176 & n2325 ) | ( n2176 & ~n3615 ) | ( n2325 & ~n3615 ) ;
  assign n14239 = ~n4098 & n9568 ;
  assign n14240 = n14239 ^ n4388 ^ 1'b0 ;
  assign n14241 = n7973 | n14240 ;
  assign n14242 = n14241 ^ n483 ^ 1'b0 ;
  assign n14243 = ~n7276 & n14242 ;
  assign n14244 = n14238 & n14243 ;
  assign n14245 = n4650 | n8765 ;
  assign n14246 = n5718 ^ n4139 ^ 1'b0 ;
  assign n14247 = n14246 ^ n8789 ^ n2579 ;
  assign n14248 = n14247 ^ n4019 ^ 1'b0 ;
  assign n14249 = n4838 & ~n7938 ;
  assign n14250 = n14249 ^ n8686 ^ 1'b0 ;
  assign n14251 = n3217 & n14250 ;
  assign n14252 = n1232 & n14251 ;
  assign n14253 = n14252 ^ n10292 ^ 1'b0 ;
  assign n14254 = n6934 | n13334 ;
  assign n14255 = n9207 & ~n14092 ;
  assign n14256 = n14255 ^ n9347 ^ 1'b0 ;
  assign n14257 = ~n11057 & n13065 ;
  assign n14258 = n3017 & n9138 ;
  assign n14259 = n2060 & n8902 ;
  assign n14260 = n567 & ~n2342 ;
  assign n14261 = n14260 ^ n12361 ^ 1'b0 ;
  assign n14262 = ~n14259 & n14261 ;
  assign n14263 = n359 & ~n1899 ;
  assign n14264 = n9500 ^ n9161 ^ 1'b0 ;
  assign n14265 = n3388 & n14264 ;
  assign n14266 = ~n3699 & n9364 ;
  assign n14267 = n14266 ^ n1060 ^ 1'b0 ;
  assign n14268 = n5613 & ~n12414 ;
  assign n14271 = n3791 | n9809 ;
  assign n14272 = n1467 | n14271 ;
  assign n14269 = n1782 ^ n1401 ^ 1'b0 ;
  assign n14270 = n1753 | n14269 ;
  assign n14273 = n14272 ^ n14270 ^ 1'b0 ;
  assign n14274 = n262 & ~n14273 ;
  assign n14275 = ~n367 & n3267 ;
  assign n14276 = n14275 ^ n2699 ^ 1'b0 ;
  assign n14277 = n3420 & n14276 ;
  assign n14278 = n1648 | n7139 ;
  assign n14279 = n1827 | n14278 ;
  assign n14280 = n14279 ^ n2062 ^ 1'b0 ;
  assign n14281 = n2664 & n14028 ;
  assign n14282 = n7460 ^ n3426 ^ 1'b0 ;
  assign n14283 = n3483 & n13419 ;
  assign n14284 = ~n6145 & n8290 ;
  assign n14285 = n3189 ^ n2614 ^ n2233 ;
  assign n14286 = n10357 & n14285 ;
  assign n14288 = n2313 ^ n1907 ^ 1'b0 ;
  assign n14287 = n7004 | n10800 ;
  assign n14289 = n14288 ^ n14287 ^ 1'b0 ;
  assign n14290 = n3810 | n4117 ;
  assign n14291 = n2354 ^ x106 ^ 1'b0 ;
  assign n14292 = ~n14290 & n14291 ;
  assign n14293 = n14292 ^ n6002 ^ 1'b0 ;
  assign n14294 = n4300 ^ n2809 ^ 1'b0 ;
  assign n14295 = n5317 & ~n14294 ;
  assign n14296 = n14295 ^ n12017 ^ 1'b0 ;
  assign n14297 = ~n9921 & n14296 ;
  assign n14298 = n4378 ^ n3192 ^ 1'b0 ;
  assign n14299 = n2678 & n14298 ;
  assign n14300 = n3688 & n14299 ;
  assign n14301 = n880 & n5611 ;
  assign n14302 = n14301 ^ n13934 ^ 1'b0 ;
  assign n14303 = n13467 | n14302 ;
  assign n14304 = n5840 ^ n2289 ^ 1'b0 ;
  assign n14305 = n2073 | n14304 ;
  assign n14306 = n14305 ^ n11128 ^ 1'b0 ;
  assign n14307 = n1948 & ~n14306 ;
  assign n14308 = n3496 & n7414 ;
  assign n14309 = n14308 ^ n428 ^ 1'b0 ;
  assign n14310 = n14309 ^ n3792 ^ 1'b0 ;
  assign n14311 = n2948 & ~n14310 ;
  assign n14312 = n14311 ^ n7694 ^ 1'b0 ;
  assign n14313 = x72 & ~n14312 ;
  assign n14314 = n1352 & ~n10287 ;
  assign n14315 = n3716 & n14314 ;
  assign n14316 = n3328 ^ n984 ^ 1'b0 ;
  assign n14317 = n945 | n2026 ;
  assign n14318 = n14317 ^ n12272 ^ 1'b0 ;
  assign n14319 = n6473 ^ n4489 ^ n948 ;
  assign n14320 = n7752 & ~n9156 ;
  assign n14321 = n14319 & n14320 ;
  assign n14322 = n4623 & ~n8177 ;
  assign n14323 = n10614 & n14322 ;
  assign n14324 = n10763 ^ n5018 ^ 1'b0 ;
  assign n14327 = ~n1042 & n3462 ;
  assign n14325 = n3268 ^ n2454 ^ 1'b0 ;
  assign n14326 = n1786 & ~n14325 ;
  assign n14328 = n14327 ^ n14326 ^ 1'b0 ;
  assign n14329 = ~n948 & n14328 ;
  assign n14330 = n1928 & n14329 ;
  assign n14331 = n13886 ^ n11030 ^ n8527 ;
  assign n14332 = n4647 & n7789 ;
  assign n14333 = ~n9573 & n14332 ;
  assign n14334 = ~n2171 & n5810 ;
  assign n14335 = ~x71 & n14334 ;
  assign n14336 = n8535 | n8737 ;
  assign n14337 = n4472 | n14336 ;
  assign n14338 = n6793 & ~n12793 ;
  assign n14339 = n13979 ^ n9316 ^ 1'b0 ;
  assign n14340 = n2708 & n14339 ;
  assign n14341 = n1862 ^ n1160 ^ 1'b0 ;
  assign n14342 = ( n5662 & n7063 ) | ( n5662 & n14341 ) | ( n7063 & n14341 ) ;
  assign n14343 = n9611 ^ n5485 ^ 1'b0 ;
  assign n14344 = n10037 ^ n7594 ^ 1'b0 ;
  assign n14345 = n1103 & ~n13108 ;
  assign n14346 = n14345 ^ n10553 ^ 1'b0 ;
  assign n14347 = n1008 & n9691 ;
  assign n14348 = n921 & n2155 ;
  assign n14349 = n1224 & ~n14348 ;
  assign n14350 = n14349 ^ n727 ^ 1'b0 ;
  assign n14351 = n11618 ^ n3955 ^ 1'b0 ;
  assign n14352 = n9274 & ~n14351 ;
  assign n14353 = n14352 ^ n8576 ^ n2240 ;
  assign n14354 = n3772 & ~n4296 ;
  assign n14355 = n1540 & ~n8188 ;
  assign n14356 = n1251 | n14355 ;
  assign n14358 = n995 ^ n586 ^ 1'b0 ;
  assign n14357 = ~n4730 & n5094 ;
  assign n14359 = n14358 ^ n14357 ^ 1'b0 ;
  assign n14360 = n3445 & n7668 ;
  assign n14361 = n10710 ^ n920 ^ 1'b0 ;
  assign n14362 = n4467 ^ n2660 ^ x18 ;
  assign n14363 = ~n2317 & n2830 ;
  assign n14364 = n7513 & n14363 ;
  assign n14365 = n1861 & n14364 ;
  assign n14369 = n972 & ~n4923 ;
  assign n14370 = n5388 & n14369 ;
  assign n14371 = n14370 ^ n339 ^ 1'b0 ;
  assign n14366 = n5562 ^ n2415 ^ 1'b0 ;
  assign n14367 = n4842 | n14366 ;
  assign n14368 = n2819 | n14367 ;
  assign n14372 = n14371 ^ n14368 ^ 1'b0 ;
  assign n14373 = n2673 & ~n4729 ;
  assign n14374 = n3764 & n14373 ;
  assign n14375 = n2034 & ~n14374 ;
  assign n14376 = n14375 ^ n4796 ^ 1'b0 ;
  assign n14377 = n1262 & ~n13332 ;
  assign n14378 = n2828 & n14377 ;
  assign n14379 = n11699 ^ n7242 ^ 1'b0 ;
  assign n14380 = n507 & ~n13816 ;
  assign n14381 = ~n7597 & n14380 ;
  assign n14382 = ~n4916 & n10776 ;
  assign n14383 = n6594 ^ n5313 ^ 1'b0 ;
  assign n14384 = n14383 ^ n2194 ^ n1552 ;
  assign n14385 = ( ~x73 & n1864 ) | ( ~x73 & n14384 ) | ( n1864 & n14384 ) ;
  assign n14386 = n7235 ^ n5536 ^ 1'b0 ;
  assign n14387 = n3712 & ~n14386 ;
  assign n14388 = n1214 & n8007 ;
  assign n14389 = n3158 ^ n877 ^ 1'b0 ;
  assign n14390 = n14388 & n14389 ;
  assign n14391 = n8032 & ~n10932 ;
  assign n14392 = n9385 & n14391 ;
  assign n14393 = n684 ^ n131 ^ 1'b0 ;
  assign n14394 = n2946 | n14393 ;
  assign n14395 = n181 & n14394 ;
  assign n14396 = n7245 & n14395 ;
  assign n14397 = n2667 ^ n642 ^ 1'b0 ;
  assign n14398 = n14396 & ~n14397 ;
  assign n14399 = ~n1833 & n6265 ;
  assign n14400 = x30 & n604 ;
  assign n14401 = ~x30 & n14400 ;
  assign n14402 = ~n328 & n1095 ;
  assign n14403 = n14401 & n14402 ;
  assign n14404 = n1644 & ~n14403 ;
  assign n14405 = n4047 | n14404 ;
  assign n14406 = n14405 ^ n7911 ^ 1'b0 ;
  assign n14407 = n3037 ^ n2974 ^ 1'b0 ;
  assign n14408 = n14406 & n14407 ;
  assign n14409 = n8190 ^ n3973 ^ 1'b0 ;
  assign n14410 = n1414 & n3100 ;
  assign n14411 = n1015 ^ n687 ^ 1'b0 ;
  assign n14412 = n2264 & n11318 ;
  assign n14413 = n1137 ^ n371 ^ 1'b0 ;
  assign n14414 = ~n14412 & n14413 ;
  assign n14415 = ~n4559 & n6853 ;
  assign n14416 = n2264 ^ n2241 ^ n1013 ;
  assign n14417 = ~n8362 & n14416 ;
  assign n14418 = n3655 & ~n5719 ;
  assign n14419 = n2322 ^ n882 ^ 1'b0 ;
  assign n14420 = n1154 & n14419 ;
  assign n14421 = ( n1221 & n1628 ) | ( n1221 & ~n8846 ) | ( n1628 & ~n8846 ) ;
  assign n14422 = n2190 | n5557 ;
  assign n14423 = n14422 ^ n9026 ^ 1'b0 ;
  assign n14424 = n14421 & n14423 ;
  assign n14425 = n6122 & n14424 ;
  assign n14426 = n14246 ^ n11254 ^ 1'b0 ;
  assign n14427 = n2347 & ~n2709 ;
  assign n14428 = n14427 ^ n10082 ^ n9665 ;
  assign n14429 = n3031 ^ n2517 ^ 1'b0 ;
  assign n14430 = n8139 | n14429 ;
  assign n14431 = n9676 & ~n14430 ;
  assign n14432 = n824 & ~n3946 ;
  assign n14435 = n1317 & n9351 ;
  assign n14433 = n3482 & ~n4288 ;
  assign n14434 = n14433 ^ n2438 ^ 1'b0 ;
  assign n14436 = n14435 ^ n14434 ^ 1'b0 ;
  assign n14437 = n7191 ^ n3844 ^ 1'b0 ;
  assign n14438 = n2499 & n14437 ;
  assign n14439 = n2374 ^ n2107 ^ 1'b0 ;
  assign n14440 = n5940 ^ n1086 ^ 1'b0 ;
  assign n14441 = ~n9124 & n14440 ;
  assign n14442 = ~n540 & n14441 ;
  assign n14443 = ( n10811 & ~n12181 ) | ( n10811 & n14341 ) | ( ~n12181 & n14341 ) ;
  assign n14444 = n12446 ^ n1487 ^ 1'b0 ;
  assign n14445 = n12364 | n14444 ;
  assign n14446 = n14445 ^ x17 ^ 1'b0 ;
  assign n14447 = ~n3401 & n13466 ;
  assign n14448 = ~n2626 & n14341 ;
  assign n14449 = n7057 & n14448 ;
  assign n14450 = ~n2499 & n14449 ;
  assign n14456 = n2739 & ~n5336 ;
  assign n14457 = n1456 & n14456 ;
  assign n14458 = ~n14456 & n14457 ;
  assign n14451 = ~n1137 & n7486 ;
  assign n14452 = ~n7486 & n14451 ;
  assign n14453 = ~n2352 & n3204 ;
  assign n14454 = n14452 & n14453 ;
  assign n14455 = n4726 | n14454 ;
  assign n14459 = n14458 ^ n14455 ^ 1'b0 ;
  assign n14460 = n3218 | n14459 ;
  assign n14461 = n14459 & ~n14460 ;
  assign n14462 = n14461 ^ n4144 ^ 1'b0 ;
  assign n14463 = n14450 & n14462 ;
  assign n14464 = n11108 ^ n5397 ^ 1'b0 ;
  assign n14465 = n5598 & n9871 ;
  assign n14466 = n1493 | n14465 ;
  assign n14467 = n2395 & n5068 ;
  assign n14468 = n11176 & n14467 ;
  assign n14469 = n12157 & n14468 ;
  assign n14470 = ( n4833 & n4964 ) | ( n4833 & n6829 ) | ( n4964 & n6829 ) ;
  assign n14471 = n1394 & n8811 ;
  assign n14472 = ~n14470 & n14471 ;
  assign n14473 = n14472 ^ x82 ^ 1'b0 ;
  assign n14474 = ~n9903 & n11144 ;
  assign n14475 = n9353 & ~n14474 ;
  assign n14476 = ~n8899 & n11356 ;
  assign n14477 = n1471 & n14476 ;
  assign n14478 = n590 | n5513 ;
  assign n14479 = ~n4610 & n5227 ;
  assign n14480 = n14478 & n14479 ;
  assign n14481 = n607 & ~n2864 ;
  assign n14482 = ~n607 & n14481 ;
  assign n14483 = n14482 ^ n2399 ^ 1'b0 ;
  assign n14484 = n12112 & n14483 ;
  assign n14485 = n14484 ^ n8588 ^ 1'b0 ;
  assign n14486 = n1414 & n14485 ;
  assign n14487 = n254 & n14486 ;
  assign n14488 = n707 | n14487 ;
  assign n14489 = n14488 ^ n8529 ^ 1'b0 ;
  assign n14490 = n11668 ^ n1758 ^ 1'b0 ;
  assign n14491 = n6124 & n14490 ;
  assign n14493 = n937 ^ x112 ^ 1'b0 ;
  assign n14494 = ~n4370 & n14493 ;
  assign n14495 = n3137 & n14494 ;
  assign n14492 = n7133 & n9636 ;
  assign n14496 = n14495 ^ n14492 ^ 1'b0 ;
  assign n14497 = n2040 ^ n754 ^ 1'b0 ;
  assign n14498 = n14497 ^ n3509 ^ 1'b0 ;
  assign n14499 = n11744 ^ n9200 ^ 1'b0 ;
  assign n14500 = n13502 ^ n1963 ^ 1'b0 ;
  assign n14501 = n12870 ^ n9053 ^ 1'b0 ;
  assign n14502 = n800 | n12738 ;
  assign n14503 = ~n473 & n10493 ;
  assign n14504 = n11130 & n14503 ;
  assign n14505 = n4500 ^ n3360 ^ 1'b0 ;
  assign n14506 = n11512 ^ n9910 ^ 1'b0 ;
  assign n14507 = n5677 & n14506 ;
  assign n14508 = n14505 & n14507 ;
  assign n14509 = n14508 ^ n13144 ^ 1'b0 ;
  assign n14510 = n11781 & ~n14509 ;
  assign n14511 = n6822 ^ n6578 ^ n5008 ;
  assign n14512 = n8094 ^ n132 ^ 1'b0 ;
  assign n14513 = ~n1115 & n6112 ;
  assign n14514 = n11714 & n14513 ;
  assign n14515 = ~n1946 & n11875 ;
  assign n14516 = n2585 & ~n4559 ;
  assign n14517 = n14516 ^ n8639 ^ 1'b0 ;
  assign n14518 = n4148 & n7876 ;
  assign n14519 = ~n7876 & n14518 ;
  assign n14520 = ~n14517 & n14519 ;
  assign n14521 = n14520 ^ n14519 ^ 1'b0 ;
  assign n14525 = ~n1482 & n7043 ;
  assign n14526 = n1335 & n14525 ;
  assign n14527 = n358 | n14526 ;
  assign n14528 = n14527 ^ n5067 ^ 1'b0 ;
  assign n14522 = n3890 & ~n8980 ;
  assign n14523 = ~n6095 & n14522 ;
  assign n14524 = n3083 | n14523 ;
  assign n14529 = n14528 ^ n14524 ^ 1'b0 ;
  assign n14530 = n10510 | n13934 ;
  assign n14531 = n5358 | n14530 ;
  assign n14532 = ( n14521 & n14529 ) | ( n14521 & n14531 ) | ( n14529 & n14531 ) ;
  assign n14533 = n1156 & n1158 ;
  assign n14534 = ~n181 & n10817 ;
  assign n14536 = ~n392 & n623 ;
  assign n14535 = n1718 & n11883 ;
  assign n14537 = n14536 ^ n14535 ^ 1'b0 ;
  assign n14538 = n1351 & n3062 ;
  assign n14539 = n8369 | n11035 ;
  assign n14540 = n12944 ^ n3700 ^ 1'b0 ;
  assign n14541 = n2895 & ~n2898 ;
  assign n14542 = n5491 ^ n1499 ^ 1'b0 ;
  assign n14543 = n8642 ^ n6799 ^ 1'b0 ;
  assign n14544 = ~n14542 & n14543 ;
  assign n14545 = n1508 & ~n11901 ;
  assign n14546 = ~n14544 & n14545 ;
  assign n14547 = n9841 & ~n14546 ;
  assign n14548 = n10699 ^ n5558 ^ n528 ;
  assign n14549 = n14548 ^ n6333 ^ 1'b0 ;
  assign n14550 = n2087 | n11257 ;
  assign n14551 = n7675 ^ n3318 ^ 1'b0 ;
  assign n14552 = n14550 | n14551 ;
  assign n14553 = ~n1850 & n4040 ;
  assign n14554 = n14552 & n14553 ;
  assign n14555 = n3847 | n5961 ;
  assign n14556 = n1839 & n8505 ;
  assign n14557 = n8831 ^ x91 ^ 1'b0 ;
  assign n14558 = n4907 ^ n407 ^ 1'b0 ;
  assign n14559 = n4928 ^ n2119 ^ 1'b0 ;
  assign n14560 = ~n7473 & n14559 ;
  assign n14561 = n11129 & ~n13261 ;
  assign n14562 = n14561 ^ n2854 ^ 1'b0 ;
  assign n14563 = n9279 | n13169 ;
  assign n14564 = n14563 ^ n1051 ^ 1'b0 ;
  assign n14565 = n13131 ^ n11309 ^ 1'b0 ;
  assign n14566 = n3074 & n14565 ;
  assign n14567 = ~n13613 & n14566 ;
  assign n14568 = n6211 & n14567 ;
  assign n14569 = ~n1316 & n14568 ;
  assign n14570 = n7296 ^ n3770 ^ 1'b0 ;
  assign n14571 = n6400 | n14570 ;
  assign n14572 = n6876 | n11098 ;
  assign n14573 = n10070 & ~n14572 ;
  assign n14574 = n707 | n14573 ;
  assign n14575 = n14571 & ~n14574 ;
  assign n14578 = n10220 ^ n5847 ^ 1'b0 ;
  assign n14579 = n7492 & n14578 ;
  assign n14576 = n7785 | n8494 ;
  assign n14577 = ~n10897 & n14576 ;
  assign n14580 = n14579 ^ n14577 ^ 1'b0 ;
  assign n14581 = n5948 ^ n2729 ^ 1'b0 ;
  assign n14582 = ~n625 & n14581 ;
  assign n14583 = n14582 ^ n13845 ^ 1'b0 ;
  assign n14584 = n10866 ^ n9501 ^ 1'b0 ;
  assign n14585 = n724 | n14584 ;
  assign n14586 = n6638 ^ n873 ^ 1'b0 ;
  assign n14587 = n5336 & n14586 ;
  assign n14588 = ~n7677 & n14587 ;
  assign n14589 = n3283 | n7245 ;
  assign n14590 = n14589 ^ n7898 ^ 1'b0 ;
  assign n14591 = n2475 | n14590 ;
  assign n14592 = n7096 ^ n6964 ^ 1'b0 ;
  assign n14593 = n2087 & ~n14592 ;
  assign n14595 = ~n1016 & n1839 ;
  assign n14596 = n7498 | n14595 ;
  assign n14597 = n229 | n14596 ;
  assign n14594 = ~n2107 & n10524 ;
  assign n14598 = n14597 ^ n14594 ^ 1'b0 ;
  assign n14599 = ~n4310 & n4707 ;
  assign n14600 = n4664 | n14599 ;
  assign n14601 = n1891 ^ n509 ^ 1'b0 ;
  assign n14602 = ~n3454 & n14601 ;
  assign n14603 = ~n1487 & n14602 ;
  assign n14604 = n9138 & n9235 ;
  assign n14605 = ( n3698 & n11869 ) | ( n3698 & n13432 ) | ( n11869 & n13432 ) ;
  assign n14606 = ~n1937 & n14605 ;
  assign n14607 = n3725 & n11569 ;
  assign n14608 = ~n3829 & n14607 ;
  assign n14609 = n14608 ^ n14047 ^ 1'b0 ;
  assign n14610 = n2112 ^ n1399 ^ 1'b0 ;
  assign n14611 = n10216 & n14610 ;
  assign n14612 = n7292 | n9362 ;
  assign n14613 = n1875 & n5525 ;
  assign n14617 = n4318 & ~n6970 ;
  assign n14618 = n5127 & n14617 ;
  assign n14614 = n7871 ^ n2328 ^ 1'b0 ;
  assign n14615 = ~n14394 & n14614 ;
  assign n14616 = ~n349 & n14615 ;
  assign n14619 = n14618 ^ n14616 ^ n9839 ;
  assign n14620 = n12731 ^ n2549 ^ 1'b0 ;
  assign n14621 = n3108 & ~n14620 ;
  assign n14622 = n11186 ^ n4471 ^ n1900 ;
  assign n14623 = n14622 ^ n13660 ^ n1355 ;
  assign n14624 = ~n7938 & n14623 ;
  assign n14625 = n14624 ^ n9408 ^ 1'b0 ;
  assign n14626 = x23 & n14625 ;
  assign n14627 = n8900 ^ n4098 ^ 1'b0 ;
  assign n14628 = ( n3353 & n7270 ) | ( n3353 & n14627 ) | ( n7270 & n14627 ) ;
  assign n14629 = n14628 ^ n5383 ^ 1'b0 ;
  assign n14630 = x24 & ~n2134 ;
  assign n14631 = n14630 ^ n2385 ^ 1'b0 ;
  assign n14632 = n7980 | n14631 ;
  assign n14633 = n7129 & n9201 ;
  assign n14634 = n14633 ^ n8694 ^ n7692 ;
  assign n14635 = n14634 ^ n163 ^ 1'b0 ;
  assign n14636 = n13960 & n14635 ;
  assign n14637 = n14180 ^ n6587 ^ 1'b0 ;
  assign n14638 = n1439 & ~n14566 ;
  assign n14639 = n7953 & n9893 ;
  assign n14641 = ~n190 & n2986 ;
  assign n14640 = ~n1079 & n2884 ;
  assign n14642 = n14641 ^ n14640 ^ 1'b0 ;
  assign n14643 = ~x75 & n825 ;
  assign n14644 = n14643 ^ n6483 ^ n3482 ;
  assign n14645 = n10675 ^ n2722 ^ 1'b0 ;
  assign n14646 = n11994 & ~n14645 ;
  assign n14647 = n5028 & ~n6110 ;
  assign n14648 = n8441 & ~n14647 ;
  assign n14649 = ~n2318 & n6244 ;
  assign n14650 = n14649 ^ n6736 ^ 1'b0 ;
  assign n14651 = n7550 & ~n13811 ;
  assign n14652 = n14651 ^ n10785 ^ 1'b0 ;
  assign n14653 = n1932 | n2539 ;
  assign n14654 = n14653 ^ n9607 ^ n487 ;
  assign n14655 = n14654 ^ n9431 ^ 1'b0 ;
  assign n14656 = n886 | n8673 ;
  assign n14657 = n6679 | n14656 ;
  assign n14658 = x13 | n14240 ;
  assign n14659 = ~x40 & n11750 ;
  assign n14660 = ~n11592 & n14659 ;
  assign n14661 = n3496 ^ n790 ^ 1'b0 ;
  assign n14662 = n6214 & n14661 ;
  assign n14663 = ( ~n3897 & n4189 ) | ( ~n3897 & n11551 ) | ( n4189 & n11551 ) ;
  assign n14664 = n12507 & ~n14663 ;
  assign n14665 = n811 & n12732 ;
  assign n14666 = n10470 | n14665 ;
  assign n14667 = ~n399 & n810 ;
  assign n14668 = ~n810 & n14667 ;
  assign n14669 = n1217 & ~n1389 ;
  assign n14670 = n14668 & n14669 ;
  assign n14671 = n3298 & ~n14670 ;
  assign n14672 = n949 & ~n14671 ;
  assign n14673 = n14672 ^ n475 ^ 1'b0 ;
  assign n14674 = ~n6298 & n8313 ;
  assign n14675 = n5195 & n14674 ;
  assign n14676 = n14675 ^ n13807 ^ 1'b0 ;
  assign n14677 = n11693 & n14465 ;
  assign n14678 = n4990 ^ n2851 ^ 1'b0 ;
  assign n14679 = n13777 ^ n12830 ^ 1'b0 ;
  assign n14680 = x50 & n12796 ;
  assign n14681 = ~n5736 & n14680 ;
  assign n14682 = n4005 & ~n12078 ;
  assign n14683 = n14682 ^ n7566 ^ 1'b0 ;
  assign n14684 = n8709 & n14683 ;
  assign n14685 = n4284 | n14684 ;
  assign n14686 = ~n14681 & n14685 ;
  assign n14688 = n3445 & n5093 ;
  assign n14689 = n14688 ^ n5639 ^ 1'b0 ;
  assign n14687 = n4727 & n5603 ;
  assign n14690 = n14689 ^ n14687 ^ 1'b0 ;
  assign n14691 = n7344 & n14690 ;
  assign n14693 = ( n2145 & ~n3791 ) | ( n2145 & n4464 ) | ( ~n3791 & n4464 ) ;
  assign n14692 = n4600 | n8972 ;
  assign n14694 = n14693 ^ n14692 ^ 1'b0 ;
  assign n14695 = n5172 ^ n493 ^ 1'b0 ;
  assign n14696 = n14694 | n14695 ;
  assign n14697 = n3900 ^ n1030 ^ 1'b0 ;
  assign n14698 = n1165 & ~n1183 ;
  assign n14699 = n14698 ^ n1329 ^ 1'b0 ;
  assign n14700 = n8204 | n14699 ;
  assign n14701 = n14700 ^ n1201 ^ 1'b0 ;
  assign n14702 = n14701 ^ n10801 ^ 1'b0 ;
  assign n14703 = ~n13699 & n14702 ;
  assign n14704 = ~x54 & n14703 ;
  assign n14705 = n12408 ^ n6069 ^ 1'b0 ;
  assign n14706 = n2109 & n4330 ;
  assign n14707 = ~n14705 & n14706 ;
  assign n14708 = n14435 ^ n858 ^ 1'b0 ;
  assign n14709 = n4291 | n14708 ;
  assign n14710 = n14709 ^ n7371 ^ 1'b0 ;
  assign n14711 = ~n4885 & n14710 ;
  assign n14712 = ~n2414 & n3498 ;
  assign n14713 = n5163 | n7994 ;
  assign n14714 = n14713 ^ n11129 ^ 1'b0 ;
  assign n14715 = ~n1790 & n5140 ;
  assign n14716 = n389 & ~n14715 ;
  assign n14717 = ~n272 & n7549 ;
  assign n14718 = n7473 & ~n9227 ;
  assign n14719 = n1976 & n14718 ;
  assign n14720 = n14717 & n14719 ;
  assign n14721 = n473 | n13286 ;
  assign n14722 = n14721 ^ n9458 ^ 1'b0 ;
  assign n14723 = ( n4387 & n6652 ) | ( n4387 & ~n8511 ) | ( n6652 & ~n8511 ) ;
  assign n14725 = n7770 & ~n9067 ;
  assign n14724 = n2253 & n6309 ;
  assign n14726 = n14725 ^ n14724 ^ 1'b0 ;
  assign n14727 = x112 & n11634 ;
  assign n14728 = n3280 & n14727 ;
  assign n14729 = n14229 ^ n8702 ^ 1'b0 ;
  assign n14730 = ~n4760 & n6631 ;
  assign n14731 = n539 & n14730 ;
  assign n14732 = ~n537 & n7311 ;
  assign n14733 = n14732 ^ n3570 ^ 1'b0 ;
  assign n14734 = n4112 & n6039 ;
  assign n14735 = n14734 ^ n3188 ^ 1'b0 ;
  assign n14736 = n14733 & n14735 ;
  assign n14737 = n14168 ^ n13383 ^ 1'b0 ;
  assign n14738 = n5691 ^ n1632 ^ 1'b0 ;
  assign n14739 = n2157 | n3195 ;
  assign n14740 = n11565 | n14739 ;
  assign n14741 = n14740 ^ n5067 ^ 1'b0 ;
  assign n14742 = n14738 | n14741 ;
  assign n14743 = n10287 | n11547 ;
  assign n14744 = n14743 ^ n6544 ^ 1'b0 ;
  assign n14745 = ~n1496 & n5448 ;
  assign n14746 = ~n5627 & n6017 ;
  assign n14747 = n14184 | n14746 ;
  assign n14748 = n14745 & ~n14747 ;
  assign n14749 = n14744 & ~n14748 ;
  assign n14750 = ~n7436 & n10439 ;
  assign n14751 = ~n1990 & n14750 ;
  assign n14752 = n6268 | n9827 ;
  assign n14753 = n9142 ^ n4746 ^ 1'b0 ;
  assign n14754 = n1022 ^ n709 ^ 1'b0 ;
  assign n14755 = n8673 | n14754 ;
  assign n14756 = n8821 & ~n14755 ;
  assign n14757 = n11595 & n14756 ;
  assign n14758 = n14757 ^ n6469 ^ 1'b0 ;
  assign n14759 = n13540 & n14758 ;
  assign n14760 = n14274 ^ n5235 ^ 1'b0 ;
  assign n14761 = n359 | n6122 ;
  assign n14762 = ~n4455 & n14761 ;
  assign n14763 = ~n12602 & n14762 ;
  assign n14764 = n1079 & ~n11009 ;
  assign n14765 = x45 & n13632 ;
  assign n14766 = n14765 ^ n11804 ^ 1'b0 ;
  assign n14767 = n5148 | n6718 ;
  assign n14768 = n539 | n1729 ;
  assign n14769 = x81 & ~n14768 ;
  assign n14770 = n7920 | n14769 ;
  assign n14771 = n1189 & ~n8983 ;
  assign n14772 = ~n14770 & n14771 ;
  assign n14773 = n7444 | n8022 ;
  assign n14774 = n14773 ^ n3551 ^ 1'b0 ;
  assign n14780 = ~x12 & n2040 ;
  assign n14781 = x12 & n14780 ;
  assign n14775 = n2383 & n3821 ;
  assign n14776 = n7881 & n14775 ;
  assign n14777 = ~n6374 & n8799 ;
  assign n14778 = ~n14520 & n14777 ;
  assign n14779 = n14776 | n14778 ;
  assign n14782 = n14781 ^ n14779 ^ 1'b0 ;
  assign n14783 = n5882 ^ n1315 ^ 1'b0 ;
  assign n14784 = n448 & n14783 ;
  assign n14785 = n14784 ^ n325 ^ 1'b0 ;
  assign n14786 = n12641 & ~n13124 ;
  assign n14787 = n9168 ^ n8008 ^ 1'b0 ;
  assign n14788 = ~n6271 & n7723 ;
  assign n14789 = n3874 ^ n3784 ^ 1'b0 ;
  assign n14790 = n7550 & n14789 ;
  assign n14791 = n14790 ^ n3652 ^ 1'b0 ;
  assign n14793 = ~n8619 & n9349 ;
  assign n14792 = ~n1463 & n14761 ;
  assign n14794 = n14793 ^ n14792 ^ 1'b0 ;
  assign n14795 = ~n7085 & n14794 ;
  assign n14796 = ~n3267 & n12086 ;
  assign n14797 = n806 & n14796 ;
  assign n14798 = n1020 | n10851 ;
  assign n14799 = n9718 & ~n10235 ;
  assign n14800 = n2198 | n3859 ;
  assign n14801 = ~n980 & n7513 ;
  assign n14803 = n1515 | n3650 ;
  assign n14802 = ~n895 & n2425 ;
  assign n14804 = n14803 ^ n14802 ^ 1'b0 ;
  assign n14805 = n14804 ^ n11651 ^ 1'b0 ;
  assign n14807 = x92 & n1547 ;
  assign n14806 = n6979 & n13427 ;
  assign n14808 = n14807 ^ n14806 ^ 1'b0 ;
  assign n14809 = n14805 | n14808 ;
  assign n14810 = n5448 & ~n9588 ;
  assign n14811 = ~n1764 & n14810 ;
  assign n14812 = n14811 ^ n4277 ^ 1'b0 ;
  assign n14813 = n806 | n6192 ;
  assign n14814 = n14812 & ~n14813 ;
  assign n14815 = n1434 & ~n6501 ;
  assign n14816 = n14815 ^ n4402 ^ 1'b0 ;
  assign n14817 = n12916 ^ n3429 ^ 1'b0 ;
  assign n14818 = n12165 & n14817 ;
  assign n14819 = n8425 ^ n2113 ^ 1'b0 ;
  assign n14820 = n14819 ^ n1487 ^ 1'b0 ;
  assign n14821 = n4835 & n14820 ;
  assign n14822 = n4086 ^ n1224 ^ 1'b0 ;
  assign n14823 = n1002 | n1661 ;
  assign n14824 = n9860 ^ n1118 ^ 1'b0 ;
  assign n14825 = n318 & n10985 ;
  assign n14826 = n6747 | n14631 ;
  assign n14827 = n4597 ^ n739 ^ 1'b0 ;
  assign n14828 = n1870 & n8062 ;
  assign n14829 = n14828 ^ n12125 ^ 1'b0 ;
  assign n14830 = n14827 & ~n14829 ;
  assign n14831 = n7946 ^ n6461 ^ 1'b0 ;
  assign n14832 = n14831 ^ x27 ^ 1'b0 ;
  assign n14833 = n5723 & n14832 ;
  assign n14834 = n14833 ^ n9145 ^ 1'b0 ;
  assign n14835 = n2604 & n14823 ;
  assign n14838 = n2528 | n3030 ;
  assign n14839 = n14838 ^ n14319 ^ 1'b0 ;
  assign n14840 = n8337 | n14839 ;
  assign n14836 = ~n6714 & n10379 ;
  assign n14837 = n14836 ^ n5553 ^ 1'b0 ;
  assign n14841 = n14840 ^ n14837 ^ 1'b0 ;
  assign n14842 = ~n830 & n11614 ;
  assign n14843 = n1588 & ~n7987 ;
  assign n14844 = n7443 | n13393 ;
  assign n14845 = ~n509 & n998 ;
  assign n14846 = ( ~n4361 & n8763 ) | ( ~n4361 & n13737 ) | ( n8763 & n13737 ) ;
  assign n14847 = ~n894 & n14846 ;
  assign n14848 = n6557 ^ n3059 ^ 1'b0 ;
  assign n14849 = n4366 | n14456 ;
  assign n14850 = n4188 & n8449 ;
  assign n14851 = n7543 & n14850 ;
  assign n14852 = n5264 ^ x100 ^ 1'b0 ;
  assign n14853 = n9168 | n14852 ;
  assign n14854 = ( n7359 & n8946 ) | ( n7359 & ~n10840 ) | ( n8946 & ~n10840 ) ;
  assign n14855 = n4296 ^ n1629 ^ 1'b0 ;
  assign n14856 = ~n4660 & n14496 ;
  assign n14857 = n2602 | n2734 ;
  assign n14858 = n14857 ^ n1997 ^ 1'b0 ;
  assign n14859 = ~n10156 & n14858 ;
  assign n14860 = n14859 ^ n10386 ^ 1'b0 ;
  assign n14861 = n4444 ^ n3358 ^ 1'b0 ;
  assign n14862 = n14860 & ~n14861 ;
  assign n14863 = n9308 & n14862 ;
  assign n14864 = n877 & ~n2243 ;
  assign n14865 = ~n5990 & n14864 ;
  assign n14866 = n14865 ^ n11856 ^ 1'b0 ;
  assign n14867 = n3906 ^ n594 ^ 1'b0 ;
  assign n14868 = n1501 | n14867 ;
  assign n14869 = n2638 & n14868 ;
  assign n14870 = n2638 & ~n4377 ;
  assign n14871 = ~n5543 & n14870 ;
  assign n14872 = ~n5345 & n11961 ;
  assign n14873 = n14871 & ~n14872 ;
  assign n14874 = ~n4942 & n5224 ;
  assign n14875 = n1497 & n14299 ;
  assign n14876 = n2618 & n14875 ;
  assign n14877 = n10388 ^ n6042 ^ n1639 ;
  assign n14878 = n14877 ^ n4941 ^ 1'b0 ;
  assign n14879 = n1245 & n3052 ;
  assign n14880 = n14879 ^ n6404 ^ 1'b0 ;
  assign n14881 = n7001 & ~n7124 ;
  assign n14882 = n14881 ^ n7029 ^ 1'b0 ;
  assign n14883 = n10584 & ~n11914 ;
  assign n14884 = ~n1536 & n14883 ;
  assign n14885 = n307 & n7615 ;
  assign n14886 = n14885 ^ n9785 ^ 1'b0 ;
  assign n14888 = n2948 | n9168 ;
  assign n14889 = n14888 ^ n9525 ^ 1'b0 ;
  assign n14887 = n7643 & ~n10633 ;
  assign n14890 = n14889 ^ n14887 ^ 1'b0 ;
  assign n14891 = n14886 | n14890 ;
  assign n14892 = n8021 ^ n745 ^ 1'b0 ;
  assign n14893 = n1188 & n14892 ;
  assign n14894 = n10080 | n14893 ;
  assign n14895 = n14894 ^ n7356 ^ 1'b0 ;
  assign n14896 = n3981 | n4400 ;
  assign n14897 = n5006 ^ x127 ^ 1'b0 ;
  assign n14898 = n8039 & n14897 ;
  assign n14899 = n1395 | n7590 ;
  assign n14900 = n14898 | n14899 ;
  assign n14901 = x57 & ~n4529 ;
  assign n14902 = n14901 ^ n8689 ^ 1'b0 ;
  assign n14903 = n3486 | n14902 ;
  assign n14904 = n14903 ^ n6723 ^ 1'b0 ;
  assign n14905 = ( n10926 & ~n14900 ) | ( n10926 & n14904 ) | ( ~n14900 & n14904 ) ;
  assign n14906 = n13826 ^ n2335 ^ 1'b0 ;
  assign n14907 = ~n8101 & n14906 ;
  assign n14908 = n14905 & ~n14907 ;
  assign n14909 = n784 & ~n11288 ;
  assign n14910 = n9848 & ~n12361 ;
  assign n14911 = n5146 & n14910 ;
  assign n14914 = ~n5982 & n13660 ;
  assign n14915 = n14914 ^ n8387 ^ 1'b0 ;
  assign n14912 = n516 | n10668 ;
  assign n14913 = n14912 ^ n4181 ^ 1'b0 ;
  assign n14916 = n14915 ^ n14913 ^ 1'b0 ;
  assign n14917 = n983 ^ x27 ^ 1'b0 ;
  assign n14918 = n12653 ^ n10398 ^ 1'b0 ;
  assign n14919 = n5152 & ~n14918 ;
  assign n14920 = n8209 ^ n526 ^ 1'b0 ;
  assign n14921 = ~n1758 & n2642 ;
  assign n14922 = n221 & ~n5231 ;
  assign n14923 = n14922 ^ n5622 ^ 1'b0 ;
  assign n14924 = n1882 & ~n2887 ;
  assign n14926 = n1206 ^ n945 ^ 1'b0 ;
  assign n14925 = n7361 & n8079 ;
  assign n14927 = n14926 ^ n14925 ^ 1'b0 ;
  assign n14928 = n6322 | n6541 ;
  assign n14929 = n4175 ^ n782 ^ 1'b0 ;
  assign n14930 = n4507 & ~n14929 ;
  assign n14931 = n14928 & n14930 ;
  assign n14932 = n9378 ^ n6490 ^ 1'b0 ;
  assign n14933 = n6420 & ~n14932 ;
  assign n14934 = n8209 & ~n14933 ;
  assign n14935 = n14934 ^ n4855 ^ 1'b0 ;
  assign n14936 = n4802 | n13974 ;
  assign n14937 = n14936 ^ n806 ^ 1'b0 ;
  assign n14938 = n1561 ^ n998 ^ 1'b0 ;
  assign n14939 = n2636 | n14938 ;
  assign n14940 = n13481 ^ n11112 ^ 1'b0 ;
  assign n14941 = n553 & ~n14940 ;
  assign n14942 = n7701 ^ n4757 ^ n1762 ;
  assign n14943 = n8374 & ~n14942 ;
  assign n14944 = n8179 & n14943 ;
  assign n14945 = n7244 | n14944 ;
  assign n14946 = n14941 | n14945 ;
  assign n14947 = ~n459 & n7679 ;
  assign n14948 = x29 & n10018 ;
  assign n14949 = ~n14947 & n14948 ;
  assign n14950 = n4985 ^ n984 ^ 1'b0 ;
  assign n14951 = n6627 ^ n2091 ^ 1'b0 ;
  assign n14952 = n14950 & n14951 ;
  assign n14953 = ( n4205 & n14652 ) | ( n4205 & ~n14952 ) | ( n14652 & ~n14952 ) ;
  assign n14954 = n6680 & n9341 ;
  assign n14955 = n7837 & ~n9071 ;
  assign n14956 = n12126 ^ n5096 ^ 1'b0 ;
  assign n14957 = n7601 ^ n2909 ^ 1'b0 ;
  assign n14958 = n9551 | n14957 ;
  assign n14959 = n14958 ^ n3270 ^ 1'b0 ;
  assign n14960 = ~n12959 & n14959 ;
  assign n14961 = n1356 ^ n1329 ^ 1'b0 ;
  assign n14962 = n14960 | n14961 ;
  assign n14963 = n12680 ^ n1467 ^ 1'b0 ;
  assign n14964 = n576 | n8232 ;
  assign n14966 = n2473 & ~n12289 ;
  assign n14967 = ~n13972 & n14966 ;
  assign n14965 = ~n4296 & n8198 ;
  assign n14968 = n14967 ^ n14965 ^ 1'b0 ;
  assign n14969 = n2238 & ~n9787 ;
  assign n14970 = n2293 & n3777 ;
  assign n14971 = n14969 & n14970 ;
  assign n14972 = n428 | n4826 ;
  assign n14973 = n12894 & ~n14972 ;
  assign n14974 = n2008 & ~n4216 ;
  assign n14975 = n4303 & n14974 ;
  assign n14976 = ~n4650 & n14975 ;
  assign n14977 = n6932 | n11309 ;
  assign n14978 = n11834 ^ n6259 ^ 1'b0 ;
  assign n14979 = n8283 | n14978 ;
  assign n14980 = n12154 | n14979 ;
  assign n14981 = n6554 & ~n14980 ;
  assign n14982 = n14981 ^ n2456 ^ 1'b0 ;
  assign n14983 = n7397 ^ n1680 ^ 1'b0 ;
  assign n14984 = n10443 & ~n14983 ;
  assign n14985 = n14984 ^ n11407 ^ 1'b0 ;
  assign n14986 = n11705 ^ n4359 ^ 1'b0 ;
  assign n14987 = n4050 ^ n2178 ^ 1'b0 ;
  assign n14988 = n14156 ^ n1202 ^ 1'b0 ;
  assign n14989 = ( ~n7683 & n14987 ) | ( ~n7683 & n14988 ) | ( n14987 & n14988 ) ;
  assign n14990 = n2023 & n10389 ;
  assign n14991 = n13790 & ~n14990 ;
  assign n14992 = n14991 ^ n1186 ^ 1'b0 ;
  assign n14996 = n2377 ^ x66 ^ 1'b0 ;
  assign n14993 = n1042 | n6591 ;
  assign n14994 = n14993 ^ n1723 ^ 1'b0 ;
  assign n14995 = n998 & ~n14994 ;
  assign n14997 = n14996 ^ n14995 ^ 1'b0 ;
  assign n14998 = n496 | n3080 ;
  assign n14999 = ~n1506 & n14998 ;
  assign n15000 = ( ~n1107 & n1930 ) | ( ~n1107 & n9651 ) | ( n1930 & n9651 ) ;
  assign n15001 = n701 & n12168 ;
  assign n15002 = n15001 ^ n14044 ^ 1'b0 ;
  assign n15003 = n15002 ^ n6278 ^ n1109 ;
  assign n15004 = n5301 ^ n508 ^ 1'b0 ;
  assign n15005 = n2364 & ~n15004 ;
  assign n15006 = ~n4310 & n15005 ;
  assign n15007 = n15003 & n15006 ;
  assign n15008 = ~n1115 & n14697 ;
  assign n15009 = ~n4153 & n7547 ;
  assign n15010 = ~n6557 & n8705 ;
  assign n15011 = n15010 ^ n3989 ^ 1'b0 ;
  assign n15012 = n8614 & ~n9586 ;
  assign n15013 = n15011 & n15012 ;
  assign n15014 = ~n5224 & n11330 ;
  assign n15015 = ~n2819 & n4612 ;
  assign n15016 = n15015 ^ n4216 ^ 1'b0 ;
  assign n15017 = n2505 & ~n5096 ;
  assign n15018 = n15017 ^ n548 ^ 1'b0 ;
  assign n15019 = n4826 | n8127 ;
  assign n15020 = n15019 ^ n8606 ^ 1'b0 ;
  assign n15021 = n2664 & ~n6173 ;
  assign n15022 = n15021 ^ n2979 ^ 1'b0 ;
  assign n15023 = ( n2896 & ~n6182 ) | ( n2896 & n10341 ) | ( ~n6182 & n10341 ) ;
  assign n15024 = n797 & ~n3195 ;
  assign n15025 = n15024 ^ n8806 ^ 1'b0 ;
  assign n15026 = n4493 ^ n1491 ^ 1'b0 ;
  assign n15027 = n1628 & n15026 ;
  assign n15028 = ~n2658 & n3691 ;
  assign n15029 = n6603 | n15028 ;
  assign n15030 = n15027 & ~n15029 ;
  assign n15031 = n9530 & n11666 ;
  assign n15032 = n15030 & n15031 ;
  assign n15033 = n15032 ^ n5633 ^ 1'b0 ;
  assign n15035 = n11104 ^ n1260 ^ 1'b0 ;
  assign n15034 = n12269 ^ n7175 ^ 1'b0 ;
  assign n15036 = n15035 ^ n15034 ^ n5895 ;
  assign n15037 = ~n328 & n2345 ;
  assign n15038 = n15037 ^ n14734 ^ 1'b0 ;
  assign n15039 = n3512 & ~n5014 ;
  assign n15040 = ~n11067 & n15039 ;
  assign n15041 = n4569 & ~n6094 ;
  assign n15042 = n1925 | n15041 ;
  assign n15043 = n15040 & ~n15042 ;
  assign n15044 = n6412 & n10850 ;
  assign n15045 = n12426 ^ n1548 ^ 1'b0 ;
  assign n15046 = n5274 & ~n15045 ;
  assign n15047 = n4980 & n15023 ;
  assign n15048 = n9074 | n12190 ;
  assign n15049 = n15048 ^ n7224 ^ 1'b0 ;
  assign n15050 = n10932 ^ n5038 ^ 1'b0 ;
  assign n15051 = n634 & n4538 ;
  assign n15052 = n2385 & n15051 ;
  assign n15053 = ~n339 & n701 ;
  assign n15054 = n339 & n15053 ;
  assign n15055 = ~n482 & n15054 ;
  assign n15056 = n293 & n15055 ;
  assign n15057 = n15052 & n15056 ;
  assign n15058 = ~n7129 & n15057 ;
  assign n15059 = n7129 & n15058 ;
  assign n15060 = n15059 ^ n14454 ^ 1'b0 ;
  assign n15061 = n2980 | n6587 ;
  assign n15062 = n15061 ^ n7498 ^ 1'b0 ;
  assign n15063 = n4809 & ~n15062 ;
  assign n15064 = n8199 ^ n783 ^ 1'b0 ;
  assign n15065 = n4576 | n15064 ;
  assign n15066 = n1469 & ~n2928 ;
  assign n15067 = n287 & n15066 ;
  assign n15068 = n1628 & ~n1723 ;
  assign n15069 = n6016 | n13147 ;
  assign n15070 = n7789 & ~n15069 ;
  assign n15071 = n8166 & ~n15070 ;
  assign n15072 = n9865 & ~n12938 ;
  assign n15073 = n6221 & n15072 ;
  assign n15074 = ( x123 & ~n9431 ) | ( x123 & n15073 ) | ( ~n9431 & n15073 ) ;
  assign n15075 = n3843 & ~n15074 ;
  assign n15076 = n15075 ^ n13863 ^ 1'b0 ;
  assign n15077 = ~n15071 & n15076 ;
  assign n15078 = ~n444 & n10401 ;
  assign n15079 = n15078 ^ n13141 ^ 1'b0 ;
  assign n15080 = n1317 & ~n4113 ;
  assign n15081 = n15080 ^ n2472 ^ 1'b0 ;
  assign n15082 = n10916 | n15081 ;
  assign n15083 = n984 & ~n1351 ;
  assign n15084 = n15083 ^ n2469 ^ 1'b0 ;
  assign n15085 = n13808 & n15084 ;
  assign n15086 = n4339 ^ n1232 ^ 1'b0 ;
  assign n15087 = n15086 ^ n13212 ^ 1'b0 ;
  assign n15088 = ~n10850 & n15087 ;
  assign n15089 = n5611 & n15088 ;
  assign n15090 = n1880 & ~n4258 ;
  assign n15091 = n15090 ^ n2615 ^ 1'b0 ;
  assign n15092 = n7478 ^ n3937 ^ 1'b0 ;
  assign n15093 = n15091 & ~n15092 ;
  assign n15094 = ( n4812 & n11805 ) | ( n4812 & n14998 ) | ( n11805 & n14998 ) ;
  assign n15095 = n1405 ^ n1240 ^ 1'b0 ;
  assign n15096 = n2105 & ~n15095 ;
  assign n15097 = n7718 | n15096 ;
  assign n15098 = n5981 & n15097 ;
  assign n15099 = n809 & ~n2420 ;
  assign n15100 = n1732 | n5958 ;
  assign n15101 = n1016 | n6112 ;
  assign n15102 = n7196 | n15101 ;
  assign n15103 = n836 | n15102 ;
  assign n15104 = n4189 & ~n15103 ;
  assign n15105 = n1191 | n9371 ;
  assign n15106 = ( n2290 & n7378 ) | ( n2290 & ~n10205 ) | ( n7378 & ~n10205 ) ;
  assign n15107 = n10526 ^ n7900 ^ 1'b0 ;
  assign n15108 = n4621 | n15107 ;
  assign n15109 = n15106 | n15108 ;
  assign n15110 = n15109 ^ n13742 ^ 1'b0 ;
  assign n15111 = ~n994 & n4072 ;
  assign n15112 = ~n3837 & n7092 ;
  assign n15113 = ~n10425 & n15112 ;
  assign n15114 = n12349 | n15113 ;
  assign n15115 = n13376 ^ n4871 ^ 1'b0 ;
  assign n15116 = n2285 & ~n2909 ;
  assign n15117 = n14655 ^ n5290 ^ 1'b0 ;
  assign n15118 = n15116 | n15117 ;
  assign n15119 = n794 & ~n3017 ;
  assign n15120 = n2094 & ~n15119 ;
  assign n15121 = n15120 ^ n9360 ^ 1'b0 ;
  assign n15122 = n1031 | n5038 ;
  assign n15123 = n5007 ^ n3230 ^ 1'b0 ;
  assign n15124 = n10617 ^ n2176 ^ 1'b0 ;
  assign n15125 = n3556 | n6414 ;
  assign n15126 = n6667 & ~n9449 ;
  assign n15127 = n15126 ^ n12873 ^ 1'b0 ;
  assign n15128 = n4469 | n12870 ;
  assign n15129 = n5715 | n15128 ;
  assign n15130 = ~n13266 & n14189 ;
  assign n15131 = n1909 & ~n4397 ;
  assign n15132 = n15131 ^ n8673 ^ 1'b0 ;
  assign n15133 = ~n10799 & n15132 ;
  assign n15135 = n1216 & ~n3464 ;
  assign n15136 = ~n1867 & n15135 ;
  assign n15134 = n2945 & ~n6587 ;
  assign n15137 = n15136 ^ n15134 ^ 1'b0 ;
  assign n15138 = n4855 & n7109 ;
  assign n15139 = ~n15137 & n15138 ;
  assign n15140 = n6982 & n7282 ;
  assign n15141 = n15140 ^ n5753 ^ 1'b0 ;
  assign n15142 = n6973 ^ n1934 ^ 1'b0 ;
  assign n15147 = n3716 & ~n6712 ;
  assign n15145 = n3834 | n7631 ;
  assign n15146 = n15145 ^ n15025 ^ 1'b0 ;
  assign n15143 = n1662 ^ n1139 ^ 1'b0 ;
  assign n15144 = ~n3335 & n15143 ;
  assign n15148 = n15147 ^ n15146 ^ n15144 ;
  assign n15149 = n4105 | n10010 ;
  assign n15150 = n3422 | n15149 ;
  assign n15151 = n15150 ^ n4416 ^ 1'b0 ;
  assign n15152 = n4759 & ~n9185 ;
  assign n15153 = n5322 & n15152 ;
  assign n15154 = n4216 & ~n6019 ;
  assign n15155 = n15154 ^ n3138 ^ 1'b0 ;
  assign n15156 = n6043 ^ n1823 ^ 1'b0 ;
  assign n15157 = n1267 & ~n15156 ;
  assign n15158 = ~n8527 & n10639 ;
  assign n15159 = n3725 & n15158 ;
  assign n15160 = n15159 ^ n614 ^ 1'b0 ;
  assign n15161 = n7179 | n7295 ;
  assign n15162 = ~n5271 & n15148 ;
  assign n15163 = ~n2329 & n6437 ;
  assign n15164 = n15163 ^ n6212 ^ 1'b0 ;
  assign n15165 = ~n4037 & n4433 ;
  assign n15166 = n15165 ^ n11943 ^ 1'b0 ;
  assign n15167 = n2958 ^ n1948 ^ 1'b0 ;
  assign n15168 = ~n1115 & n15167 ;
  assign n15169 = n7841 ^ n2602 ^ 1'b0 ;
  assign n15170 = n4753 & n7195 ;
  assign n15171 = n15170 ^ n3407 ^ 1'b0 ;
  assign n15172 = n2681 & ~n10609 ;
  assign n15173 = n15172 ^ n7619 ^ 1'b0 ;
  assign n15174 = n2101 & n5016 ;
  assign n15175 = n3137 & n15174 ;
  assign n15177 = n3842 ^ n1726 ^ 1'b0 ;
  assign n15176 = n5186 & ~n9608 ;
  assign n15178 = n15177 ^ n15176 ^ 1'b0 ;
  assign n15179 = n782 | n1055 ;
  assign n15180 = n15179 ^ n14390 ^ 1'b0 ;
  assign n15181 = n5535 ^ n3526 ^ 1'b0 ;
  assign n15182 = n2242 ^ n945 ^ 1'b0 ;
  assign n15183 = n15181 & n15182 ;
  assign n15184 = n2763 | n5181 ;
  assign n15185 = n365 | n15184 ;
  assign n15186 = n6485 & ~n11148 ;
  assign n15187 = n6310 & ~n13811 ;
  assign n15188 = n15187 ^ n2530 ^ 1'b0 ;
  assign n15189 = n1380 & ~n15188 ;
  assign n15190 = n15189 ^ n3714 ^ 1'b0 ;
  assign n15191 = n8441 ^ n3358 ^ n962 ;
  assign n15193 = n2163 & n2414 ;
  assign n15192 = ~n464 & n10079 ;
  assign n15194 = n15193 ^ n15192 ^ 1'b0 ;
  assign n15195 = n9774 ^ n4296 ^ 1'b0 ;
  assign n15196 = n15195 ^ n6455 ^ 1'b0 ;
  assign n15197 = n4364 ^ n2427 ^ 1'b0 ;
  assign n15198 = n4755 & n15197 ;
  assign n15199 = n10674 & n15198 ;
  assign n15200 = ~n6022 & n15199 ;
  assign n15201 = ~n15199 & n15200 ;
  assign n15202 = n15201 ^ n1017 ^ 1'b0 ;
  assign n15203 = n5886 | n15202 ;
  assign n15204 = ~n5986 & n7830 ;
  assign n15206 = ~n8279 & n13985 ;
  assign n15207 = ~n830 & n15206 ;
  assign n15208 = n15207 ^ n9445 ^ 1'b0 ;
  assign n15205 = ~n708 & n12083 ;
  assign n15209 = n15208 ^ n15205 ^ 1'b0 ;
  assign n15210 = n4929 ^ n1034 ^ 1'b0 ;
  assign n15211 = n5417 & ~n15210 ;
  assign n15212 = n5525 & n9530 ;
  assign n15213 = n8121 & n15212 ;
  assign n15214 = n516 | n4623 ;
  assign n15215 = n4277 & n11703 ;
  assign n15216 = n863 & ~n2905 ;
  assign n15217 = n15216 ^ n1098 ^ 1'b0 ;
  assign n15218 = n3310 ^ n2584 ^ 1'b0 ;
  assign n15219 = n4800 & ~n15218 ;
  assign n15220 = ~n2608 & n8152 ;
  assign n15221 = n15220 ^ n254 ^ 1'b0 ;
  assign n15222 = ~n3780 & n15221 ;
  assign n15223 = ~n15219 & n15222 ;
  assign n15224 = n4960 | n13877 ;
  assign n15225 = n15223 & ~n15224 ;
  assign n15226 = n15225 ^ n749 ^ 1'b0 ;
  assign n15227 = n6454 & ~n15226 ;
  assign n15228 = n7199 & n12569 ;
  assign n15229 = n6587 & n15228 ;
  assign n15230 = ~n692 & n5004 ;
  assign n15231 = n15230 ^ n2081 ^ 1'b0 ;
  assign n15232 = n15231 ^ n3126 ^ 1'b0 ;
  assign n15233 = n15232 ^ n7245 ^ 1'b0 ;
  assign n15234 = n1267 & ~n15233 ;
  assign n15235 = n568 & ~n1069 ;
  assign n15236 = ~n6844 & n15235 ;
  assign n15237 = n9176 | n15236 ;
  assign n15238 = n7899 | n15237 ;
  assign n15240 = n1726 & ~n4204 ;
  assign n15239 = n625 | n4458 ;
  assign n15241 = n15240 ^ n15239 ^ 1'b0 ;
  assign n15242 = n15241 ^ n10922 ^ 1'b0 ;
  assign n15243 = n13108 ^ n10232 ^ 1'b0 ;
  assign n15244 = n1644 & ~n15243 ;
  assign n15245 = n6582 & n15244 ;
  assign n15246 = n775 & ~n14263 ;
  assign n15247 = n15146 ^ n9179 ^ 1'b0 ;
  assign n15248 = ~n14886 & n15247 ;
  assign n15249 = n1537 | n3336 ;
  assign n15250 = n1566 | n15249 ;
  assign n15251 = n1506 & n15250 ;
  assign n15253 = ~n198 & n2649 ;
  assign n15254 = n15253 ^ n7825 ^ 1'b0 ;
  assign n15252 = n8439 | n8473 ;
  assign n15255 = n15254 ^ n15252 ^ 1'b0 ;
  assign n15256 = n7129 & ~n15255 ;
  assign n15257 = n2130 ^ n2107 ^ 1'b0 ;
  assign n15258 = n2067 & ~n15257 ;
  assign n15259 = n4296 ^ n2755 ^ 1'b0 ;
  assign n15260 = n15258 & n15259 ;
  assign n15261 = ~n12890 & n15260 ;
  assign n15262 = n11737 | n14810 ;
  assign n15263 = n7198 | n15262 ;
  assign n15264 = x82 | n15263 ;
  assign n15265 = n14790 ^ n294 ^ 1'b0 ;
  assign n15266 = n2056 & n2598 ;
  assign n15267 = n7736 ^ n6467 ^ 1'b0 ;
  assign n15268 = n3803 | n7250 ;
  assign n15269 = n15268 ^ n8531 ^ 1'b0 ;
  assign n15270 = n15267 | n15269 ;
  assign n15271 = n4028 & ~n13057 ;
  assign n15272 = n3785 & ~n5356 ;
  assign n15273 = n15272 ^ n7928 ^ n2513 ;
  assign n15274 = n6160 & n15273 ;
  assign n15275 = n1656 | n11718 ;
  assign n15276 = n15275 ^ n7305 ^ 1'b0 ;
  assign n15277 = n4267 ^ n4234 ^ 1'b0 ;
  assign n15278 = n2675 & n15277 ;
  assign n15281 = n5921 ^ x82 ^ 1'b0 ;
  assign n15282 = n1342 & n15281 ;
  assign n15279 = x19 | n3536 ;
  assign n15280 = n15279 ^ n283 ^ 1'b0 ;
  assign n15283 = n15282 ^ n15280 ^ n12825 ;
  assign n15284 = n3280 ^ n1317 ^ 1'b0 ;
  assign n15285 = ~n1212 & n5445 ;
  assign n15286 = n4502 | n10895 ;
  assign n15287 = n2980 | n4556 ;
  assign n15288 = n15287 ^ n2592 ^ 1'b0 ;
  assign n15289 = ( n3433 & n9333 ) | ( n3433 & ~n10763 ) | ( n9333 & ~n10763 ) ;
  assign n15290 = n11072 & n15289 ;
  assign n15291 = n15290 ^ n5381 ^ 1'b0 ;
  assign n15292 = ~n1732 & n7093 ;
  assign n15293 = n5104 | n7050 ;
  assign n15294 = n15293 ^ n4224 ^ 1'b0 ;
  assign n15295 = n9116 & ~n10498 ;
  assign n15296 = n9114 & n15295 ;
  assign n15297 = n13066 & ~n15296 ;
  assign n15298 = ~n13828 & n15297 ;
  assign n15299 = n15252 ^ n9096 ^ n5189 ;
  assign n15300 = n3356 | n11725 ;
  assign n15301 = n7378 ^ n5973 ^ 1'b0 ;
  assign n15302 = n1738 | n15301 ;
  assign n15303 = n15302 ^ n6117 ^ 1'b0 ;
  assign n15304 = n1302 & ~n1994 ;
  assign n15305 = ~n181 & n11286 ;
  assign n15306 = n539 & ~n13623 ;
  assign n15307 = n11587 & n15306 ;
  assign n15308 = ~n1950 & n7280 ;
  assign n15309 = n15308 ^ n13127 ^ 1'b0 ;
  assign n15310 = ~n7437 & n15309 ;
  assign n15311 = n15310 ^ n1952 ^ 1'b0 ;
  assign n15313 = n185 | n2188 ;
  assign n15312 = n1103 & ~n2385 ;
  assign n15314 = n15313 ^ n15312 ^ n8573 ;
  assign n15315 = n3438 | n8235 ;
  assign n15316 = x0 | n15315 ;
  assign n15317 = n15314 & n15316 ;
  assign n15318 = n1181 ^ n920 ^ x107 ;
  assign n15319 = n3116 | n3531 ;
  assign n15320 = ~x123 & n15319 ;
  assign n15321 = x27 & ~n4759 ;
  assign n15322 = n15321 ^ n7250 ^ 1'b0 ;
  assign n15323 = n2505 & n11747 ;
  assign n15324 = n15323 ^ n10862 ^ 1'b0 ;
  assign n15325 = n13599 ^ n3282 ^ 1'b0 ;
  assign n15326 = n15325 ^ n11568 ^ 1'b0 ;
  assign n15327 = n4328 ^ n3600 ^ 1'b0 ;
  assign n15328 = ~n3702 & n15327 ;
  assign n15330 = n3728 ^ n1806 ^ 1'b0 ;
  assign n15331 = n11186 & n15330 ;
  assign n15332 = n15331 ^ n9707 ^ 1'b0 ;
  assign n15329 = n1737 & n3445 ;
  assign n15333 = n15332 ^ n15329 ^ 1'b0 ;
  assign n15334 = ~n3334 & n12366 ;
  assign n15335 = n15334 ^ n13625 ^ 1'b0 ;
  assign n15336 = n224 & ~n15335 ;
  assign n15337 = n12468 ^ n7946 ^ 1'b0 ;
  assign n15338 = n7009 | n11712 ;
  assign n15339 = n10939 ^ n7289 ^ 1'b0 ;
  assign n15342 = n5228 | n10505 ;
  assign n15340 = n9381 ^ n6039 ^ 1'b0 ;
  assign n15341 = ~n973 & n15340 ;
  assign n15343 = n15342 ^ n15341 ^ 1'b0 ;
  assign n15344 = n588 | n1731 ;
  assign n15345 = n1280 | n15344 ;
  assign n15346 = n12916 ^ n9421 ^ 1'b0 ;
  assign n15347 = ( n3433 & n15345 ) | ( n3433 & n15346 ) | ( n15345 & n15346 ) ;
  assign n15348 = n4554 | n10000 ;
  assign n15349 = ~n9916 & n15348 ;
  assign n15350 = n825 & n15349 ;
  assign n15351 = n15350 ^ n8042 ^ 1'b0 ;
  assign n15352 = n8773 ^ n5961 ^ 1'b0 ;
  assign n15353 = n526 | n15352 ;
  assign n15354 = ( n307 & n8096 ) | ( n307 & ~n15353 ) | ( n8096 & ~n15353 ) ;
  assign n15355 = n3798 & ~n15354 ;
  assign n15356 = n11365 ^ n2073 ^ 1'b0 ;
  assign n15357 = n6943 & n15356 ;
  assign n15358 = n3128 | n15357 ;
  assign n15359 = n5090 ^ n3833 ^ 1'b0 ;
  assign n15360 = n13279 & ~n14595 ;
  assign n15361 = n14257 ^ n9646 ^ 1'b0 ;
  assign n15362 = n1568 & ~n1980 ;
  assign n15363 = n15362 ^ n14304 ^ 1'b0 ;
  assign n15364 = n10299 & ~n10539 ;
  assign n15365 = n3505 & n15364 ;
  assign n15366 = ~n2800 & n15365 ;
  assign n15367 = n6145 & ~n7857 ;
  assign n15368 = ~n3714 & n8767 ;
  assign n15369 = n15368 ^ n2438 ^ 1'b0 ;
  assign n15370 = n5358 & ~n8986 ;
  assign n15371 = n1270 & n15370 ;
  assign n15372 = n2358 & n7852 ;
  assign n15373 = n13058 & ~n15372 ;
  assign n15374 = n9646 ^ n3300 ^ 1'b0 ;
  assign n15375 = n15373 & n15374 ;
  assign n15376 = n279 & ~n5350 ;
  assign n15377 = n15376 ^ n7204 ^ 1'b0 ;
  assign n15378 = n8755 | n15377 ;
  assign n15379 = n158 & ~n5971 ;
  assign n15380 = n4527 | n7139 ;
  assign n15381 = n15380 ^ n7627 ^ 1'b0 ;
  assign n15382 = ~n12710 & n15381 ;
  assign n15383 = n8127 ^ n812 ^ 1'b0 ;
  assign n15384 = n10482 ^ n6284 ^ 1'b0 ;
  assign n15396 = ~n1455 & n2467 ;
  assign n15397 = n3072 & n15396 ;
  assign n15388 = n4816 ^ n3829 ^ 1'b0 ;
  assign n15385 = ~x46 & n1051 ;
  assign n15386 = ( ~n998 & n1680 ) | ( ~n998 & n15385 ) | ( n1680 & n15385 ) ;
  assign n15387 = n1331 | n15386 ;
  assign n15389 = n15388 ^ n15387 ^ 1'b0 ;
  assign n15390 = n9235 ^ n3549 ^ 1'b0 ;
  assign n15391 = ~n15389 & n15390 ;
  assign n15392 = n297 | n2127 ;
  assign n15393 = n4592 | n15392 ;
  assign n15394 = n15393 ^ n718 ^ 1'b0 ;
  assign n15395 = n15391 & n15394 ;
  assign n15398 = n15397 ^ n15395 ^ 1'b0 ;
  assign n15399 = n355 & ~n10666 ;
  assign n15400 = n15399 ^ n11925 ^ 1'b0 ;
  assign n15401 = n5096 & n8899 ;
  assign n15403 = ~n346 & n3669 ;
  assign n15402 = n3956 | n11108 ;
  assign n15404 = n15403 ^ n15402 ^ 1'b0 ;
  assign n15405 = n2188 | n2767 ;
  assign n15406 = n15405 ^ n4052 ^ 1'b0 ;
  assign n15407 = n8059 & ~n13568 ;
  assign n15408 = n15407 ^ n14260 ^ 1'b0 ;
  assign n15409 = ~n6007 & n10051 ;
  assign n15410 = ~n12575 & n15409 ;
  assign n15411 = n920 & ~n3628 ;
  assign n15412 = n15411 ^ n8459 ^ 1'b0 ;
  assign n15413 = n1841 | n5453 ;
  assign n15414 = n15413 ^ n4212 ^ 1'b0 ;
  assign n15415 = x11 & ~n6309 ;
  assign n15416 = n5301 & n6994 ;
  assign n15417 = n9103 | n11037 ;
  assign n15418 = n15417 ^ n6906 ^ 1'b0 ;
  assign n15419 = ~n2367 & n6594 ;
  assign n15420 = x54 & n13697 ;
  assign n15421 = n15419 & n15420 ;
  assign n15422 = n9734 ^ n3898 ^ 1'b0 ;
  assign n15423 = n1556 & ~n15422 ;
  assign n15424 = ~n2259 & n15423 ;
  assign n15425 = ~n7596 & n15424 ;
  assign n15426 = n2696 & ~n15425 ;
  assign n15427 = n7629 & ~n14061 ;
  assign n15428 = n3472 & ~n5007 ;
  assign n15429 = ~x104 & n15428 ;
  assign n15430 = n12687 ^ n5913 ^ 1'b0 ;
  assign n15431 = n5289 & n5716 ;
  assign n15432 = ~n15430 & n15431 ;
  assign n15433 = n2156 & ~n2636 ;
  assign n15434 = n15433 ^ n1158 ^ 1'b0 ;
  assign n15435 = n15434 ^ n6080 ^ 1'b0 ;
  assign n15436 = ~n10588 & n15435 ;
  assign n15437 = n4489 ^ n1675 ^ 1'b0 ;
  assign n15438 = n15437 ^ n1668 ^ 1'b0 ;
  assign n15439 = n1652 & ~n15438 ;
  assign n15440 = n15439 ^ n7887 ^ 1'b0 ;
  assign n15441 = n15440 ^ n11700 ^ 1'b0 ;
  assign n15442 = n2453 ^ n2210 ^ 1'b0 ;
  assign n15443 = n4457 ^ n510 ^ 1'b0 ;
  assign n15444 = n1048 | n15443 ;
  assign n15445 = n3270 | n15444 ;
  assign n15446 = n15445 ^ n9573 ^ 1'b0 ;
  assign n15447 = ~n3116 & n15446 ;
  assign n15448 = n15442 & n15447 ;
  assign n15449 = n2395 & ~n13721 ;
  assign n15450 = n15448 & n15449 ;
  assign n15451 = n2136 ^ x65 ^ 1'b0 ;
  assign n15452 = ~n6009 & n15451 ;
  assign n15453 = n2824 & ~n9868 ;
  assign n15454 = ~n15452 & n15453 ;
  assign n15462 = ~n8435 & n9650 ;
  assign n15455 = n245 | n2469 ;
  assign n15456 = ~n934 & n15455 ;
  assign n15457 = x85 & ~n7140 ;
  assign n15458 = n15456 & n15457 ;
  assign n15459 = n11035 & ~n11316 ;
  assign n15460 = n15459 ^ n13530 ^ 1'b0 ;
  assign n15461 = ~n15458 & n15460 ;
  assign n15463 = n15462 ^ n15461 ^ 1'b0 ;
  assign n15464 = n6766 ^ n2441 ^ 1'b0 ;
  assign n15465 = n965 & n15464 ;
  assign n15466 = n6705 ^ n5154 ^ 1'b0 ;
  assign n15467 = n15466 ^ n2953 ^ 1'b0 ;
  assign n15468 = n1317 & ~n2928 ;
  assign n15469 = ~n2624 & n7375 ;
  assign n15470 = n2847 ^ n2469 ^ n614 ;
  assign n15471 = n15470 ^ n1449 ^ 1'b0 ;
  assign n15472 = n9340 ^ n9173 ^ 1'b0 ;
  assign n15473 = ~n3949 & n15472 ;
  assign n15474 = n900 & n4336 ;
  assign n15475 = n13885 ^ n3622 ^ 1'b0 ;
  assign n15476 = n15266 & ~n15475 ;
  assign n15477 = ~n5072 & n13543 ;
  assign n15478 = n15477 ^ n11124 ^ 1'b0 ;
  assign n15479 = ~n4296 & n11089 ;
  assign n15480 = ~n3736 & n15479 ;
  assign n15481 = ~n7184 & n13522 ;
  assign n15482 = n15481 ^ n12586 ^ 1'b0 ;
  assign n15483 = n7926 & ~n8679 ;
  assign n15484 = n15483 ^ n7194 ^ 1'b0 ;
  assign n15485 = n3075 | n12308 ;
  assign n15486 = n2515 | n15485 ;
  assign n15487 = n2043 & ~n3134 ;
  assign n15488 = n707 | n15487 ;
  assign n15489 = n15419 ^ n11442 ^ n9133 ;
  assign n15490 = n1599 & ~n6587 ;
  assign n15491 = n3706 & n15490 ;
  assign n15492 = ~n2357 & n5700 ;
  assign n15493 = n15492 ^ n13782 ^ 1'b0 ;
  assign n15494 = n12367 & n15493 ;
  assign n15495 = n2980 & n14198 ;
  assign n15496 = n2009 & n2156 ;
  assign n15497 = ~n2009 & n15496 ;
  assign n15498 = n3813 & ~n15497 ;
  assign n15499 = n8145 ^ n5035 ^ 1'b0 ;
  assign n15500 = n15498 & ~n15499 ;
  assign n15501 = n669 | n1030 ;
  assign n15502 = n1030 & ~n15501 ;
  assign n15503 = n15502 ^ n14006 ^ 1'b0 ;
  assign n15504 = ~n6197 & n15503 ;
  assign n15505 = ~n1315 & n9896 ;
  assign n15506 = ~n15504 & n15505 ;
  assign n15507 = n2091 & n9377 ;
  assign n15508 = n3931 & ~n5290 ;
  assign n15509 = ~n161 & n15508 ;
  assign n15510 = ~n2765 & n12815 ;
  assign n15511 = ~n15509 & n15510 ;
  assign n15512 = ~n15507 & n15511 ;
  assign n15513 = n10237 ^ n2931 ^ 1'b0 ;
  assign n15514 = x107 & n15513 ;
  assign n15515 = n9872 ^ n1543 ^ 1'b0 ;
  assign n15516 = n4213 | n15515 ;
  assign n15517 = n4497 & n9459 ;
  assign n15518 = n15517 ^ n14355 ^ 1'b0 ;
  assign n15519 = n7509 ^ n1644 ^ 1'b0 ;
  assign n15520 = ~n2291 & n11290 ;
  assign n15521 = n15519 & n15520 ;
  assign n15522 = n15521 ^ n307 ^ 1'b0 ;
  assign n15523 = n9410 ^ n439 ^ 1'b0 ;
  assign n15524 = n482 & ~n14960 ;
  assign n15525 = n15524 ^ n3433 ^ 1'b0 ;
  assign n15526 = n14232 & ~n14842 ;
  assign n15527 = ~n1212 & n3057 ;
  assign n15528 = n7613 & n15527 ;
  assign n15529 = n8522 | n15528 ;
  assign n15530 = n5139 | n9910 ;
  assign n15531 = n9910 & ~n15530 ;
  assign n15532 = n7841 & ~n15531 ;
  assign n15545 = n2267 & ~n2811 ;
  assign n15546 = n2811 & n15545 ;
  assign n15533 = x44 & ~n1880 ;
  assign n15534 = ~x44 & n15533 ;
  assign n15535 = x76 & n336 ;
  assign n15536 = ~x76 & n15535 ;
  assign n15537 = n314 & n15536 ;
  assign n15538 = n899 & ~n15537 ;
  assign n15539 = n15534 & ~n15538 ;
  assign n15540 = x112 & ~n3666 ;
  assign n15541 = n15539 & n15540 ;
  assign n15542 = n1951 & n15541 ;
  assign n15543 = n895 | n7186 ;
  assign n15544 = n15542 & ~n15543 ;
  assign n15547 = n15546 ^ n15544 ^ 1'b0 ;
  assign n15548 = n3899 & n15547 ;
  assign n15549 = ~n15532 & n15548 ;
  assign n15550 = n15549 ^ n2792 ^ 1'b0 ;
  assign n15551 = ~n3634 & n6223 ;
  assign n15552 = n1457 | n10089 ;
  assign n15553 = n14157 ^ n3862 ^ 1'b0 ;
  assign n15554 = n14627 ^ n14187 ^ 1'b0 ;
  assign n15555 = ~n10003 & n15554 ;
  assign n15556 = n10191 ^ n2456 ^ 1'b0 ;
  assign n15557 = n4880 & ~n5549 ;
  assign n15558 = n11746 ^ n6402 ^ 1'b0 ;
  assign n15559 = ~n1993 & n15558 ;
  assign n15560 = ~n8127 & n13073 ;
  assign n15561 = n1216 & ~n3009 ;
  assign n15562 = n3483 & ~n15561 ;
  assign n15563 = n15562 ^ n7057 ^ 1'b0 ;
  assign n15564 = n11939 | n15563 ;
  assign n15565 = ~n4656 & n5974 ;
  assign n15566 = n15565 ^ n13715 ^ 1'b0 ;
  assign n15567 = ~n11145 & n15566 ;
  assign n15568 = n8670 ^ n3385 ^ x73 ;
  assign n15569 = n9709 ^ n1983 ^ 1'b0 ;
  assign n15570 = ~n6181 & n15569 ;
  assign n15571 = n15570 ^ n15388 ^ 1'b0 ;
  assign n15572 = n1612 | n7676 ;
  assign n15573 = n5365 ^ n5154 ^ 1'b0 ;
  assign n15574 = n15573 ^ n13542 ^ 1'b0 ;
  assign n15575 = ~n3926 & n5802 ;
  assign n15576 = n12454 | n15575 ;
  assign n15577 = n949 & ~n2091 ;
  assign n15578 = ~n3236 & n15577 ;
  assign n15579 = n7530 ^ n483 ^ 1'b0 ;
  assign n15580 = ~n2480 & n12911 ;
  assign n15581 = n1726 ^ n1645 ^ 1'b0 ;
  assign n15582 = n8763 ^ n5592 ^ n387 ;
  assign n15583 = ~n1810 & n14158 ;
  assign n15584 = ~n15582 & n15583 ;
  assign n15585 = n3091 | n10780 ;
  assign n15586 = n6128 & n6184 ;
  assign n15587 = ~n8901 & n15586 ;
  assign n15588 = n3548 | n5451 ;
  assign n15589 = n1601 & n11176 ;
  assign n15590 = n4726 & ~n15589 ;
  assign n15591 = ~n5240 & n12311 ;
  assign n15592 = n15591 ^ n171 ^ 1'b0 ;
  assign n15593 = n466 | n2673 ;
  assign n15594 = n11209 ^ n7259 ^ n4382 ;
  assign n15595 = n10011 ^ n1385 ^ 1'b0 ;
  assign n15596 = n11911 & ~n15595 ;
  assign n15597 = n8127 & n15367 ;
  assign n15598 = ~n10840 & n15597 ;
  assign n15599 = n2799 & n14674 ;
  assign n15600 = n5526 ^ n2245 ^ 1'b0 ;
  assign n15601 = n2267 & ~n15600 ;
  assign n15602 = n15601 ^ n10698 ^ 1'b0 ;
  assign n15603 = n12590 | n13851 ;
  assign n15604 = n5383 | n9425 ;
  assign n15605 = n15604 ^ n3130 ^ 1'b0 ;
  assign n15606 = n13686 ^ n5763 ^ 1'b0 ;
  assign n15607 = ~n15605 & n15606 ;
  assign n15608 = n6575 | n10499 ;
  assign n15609 = n15608 ^ n1948 ^ 1'b0 ;
  assign n15610 = n10173 & n15609 ;
  assign n15611 = n15610 ^ n5215 ^ 1'b0 ;
  assign n15612 = n15611 ^ n6131 ^ 1'b0 ;
  assign n15613 = ~n1156 & n9196 ;
  assign n15614 = ~n2661 & n10591 ;
  assign n15615 = n15614 ^ n12102 ^ 1'b0 ;
  assign n15616 = n5234 & ~n10359 ;
  assign n15617 = ~n15615 & n15616 ;
  assign n15618 = n14889 ^ n1221 ^ 1'b0 ;
  assign n15619 = n7435 ^ n4570 ^ 1'b0 ;
  assign n15620 = x127 & ~n15619 ;
  assign n15621 = n15620 ^ n8846 ^ 1'b0 ;
  assign n15622 = n144 & n3224 ;
  assign n15623 = ( ~n7622 & n9642 ) | ( ~n7622 & n13378 ) | ( n9642 & n13378 ) ;
  assign n15624 = ~n15622 & n15623 ;
  assign n15625 = ( n2872 & n3415 ) | ( n2872 & ~n4450 ) | ( n3415 & ~n4450 ) ;
  assign n15626 = n7462 | n15625 ;
  assign n15627 = n10641 ^ n1525 ^ 1'b0 ;
  assign n15628 = ~n1930 & n2503 ;
  assign n15629 = n3360 ^ n888 ^ 1'b0 ;
  assign n15630 = ~n3551 & n15629 ;
  assign n15631 = n9502 & ~n12613 ;
  assign n15632 = ~n6722 & n15631 ;
  assign n15633 = n1645 ^ n1126 ^ 1'b0 ;
  assign n15634 = n6992 | n15633 ;
  assign n15635 = n15632 & ~n15634 ;
  assign n15636 = n3688 ^ n2602 ^ 1'b0 ;
  assign n15637 = n3353 & ~n15636 ;
  assign n15638 = n4318 | n7782 ;
  assign n15640 = n6044 & n10040 ;
  assign n15639 = n2347 & n11286 ;
  assign n15641 = n15640 ^ n15639 ^ 1'b0 ;
  assign n15642 = n4871 | n6772 ;
  assign n15643 = n1519 & ~n15642 ;
  assign n15644 = n662 | n6787 ;
  assign n15645 = n8152 | n15644 ;
  assign n15646 = n2811 | n7098 ;
  assign n15647 = n15645 & n15646 ;
  assign n15648 = n8426 ^ n7027 ^ 1'b0 ;
  assign n15649 = n8803 ^ n867 ^ 1'b0 ;
  assign n15650 = n7059 | n15649 ;
  assign n15651 = n1624 ^ n272 ^ 1'b0 ;
  assign n15652 = n5764 & n5839 ;
  assign n15653 = n13551 ^ n5239 ^ 1'b0 ;
  assign n15654 = n15652 | n15653 ;
  assign n15655 = n1273 & ~n11624 ;
  assign n15656 = n1178 & n2550 ;
  assign n15657 = ~n2396 & n15656 ;
  assign n15658 = ~n1580 & n15657 ;
  assign n15659 = x37 & ~n1016 ;
  assign n15660 = n14044 ^ n3929 ^ 1'b0 ;
  assign n15661 = n4110 & ~n15660 ;
  assign n15662 = n450 & n9072 ;
  assign n15663 = n12830 ^ n8713 ^ 1'b0 ;
  assign n15664 = n15663 ^ n3072 ^ 1'b0 ;
  assign n15665 = ~n5294 & n6212 ;
  assign n15666 = n15665 ^ n9469 ^ 1'b0 ;
  assign n15668 = n2932 | n3563 ;
  assign n15667 = n7904 & ~n14184 ;
  assign n15669 = n15668 ^ n15667 ^ 1'b0 ;
  assign n15670 = ~n577 & n15669 ;
  assign n15671 = n15670 ^ n12315 ^ 1'b0 ;
  assign n15672 = n15671 ^ n9913 ^ 1'b0 ;
  assign n15673 = n11474 ^ n5520 ^ 1'b0 ;
  assign n15674 = n2261 & ~n15673 ;
  assign n15675 = n15674 ^ n8571 ^ 1'b0 ;
  assign n15676 = ~n950 & n5704 ;
  assign n15677 = ~n5063 & n14038 ;
  assign n15678 = n15271 ^ n12397 ^ 1'b0 ;
  assign n15679 = n9102 | n9711 ;
  assign n15680 = n13684 ^ n7574 ^ n3793 ;
  assign n15681 = n3759 & ~n11276 ;
  assign n15682 = n15681 ^ n1526 ^ 1'b0 ;
  assign n15683 = x14 & ~n15682 ;
  assign n15684 = n15683 ^ n4980 ^ 1'b0 ;
  assign n15685 = n1711 ^ n828 ^ 1'b0 ;
  assign n15686 = n15685 ^ n5158 ^ 1'b0 ;
  assign n15687 = n15686 ^ n3817 ^ 1'b0 ;
  assign n15688 = ~n6972 & n8954 ;
  assign n15689 = n15688 ^ n5562 ^ 1'b0 ;
  assign n15690 = ~n2632 & n13604 ;
  assign n15691 = ~n5991 & n6030 ;
  assign n15692 = n8263 & n15691 ;
  assign n15693 = n494 | n15692 ;
  assign n15694 = n15693 ^ n5789 ^ 1'b0 ;
  assign n15695 = n15319 ^ n1985 ^ 1'b0 ;
  assign n15696 = n3017 ^ n1059 ^ 1'b0 ;
  assign n15697 = ~n3987 & n15696 ;
  assign n15698 = x22 & ~n2418 ;
  assign n15699 = n1172 | n2465 ;
  assign n15700 = n8137 & ~n15699 ;
  assign n15701 = n15700 ^ n5436 ^ 1'b0 ;
  assign n15702 = ~n1051 & n15701 ;
  assign n15703 = n3872 & n4265 ;
  assign n15704 = ~n1888 & n15703 ;
  assign n15705 = n15704 ^ n5746 ^ 1'b0 ;
  assign n15706 = ( n1861 & n3941 ) | ( n1861 & n7268 ) | ( n3941 & n7268 ) ;
  assign n15707 = n15706 ^ n1268 ^ 1'b0 ;
  assign n15708 = n10151 & n15707 ;
  assign n15709 = n371 | n2615 ;
  assign n15710 = ( n6289 & n7747 ) | ( n6289 & ~n15709 ) | ( n7747 & ~n15709 ) ;
  assign n15713 = n8033 & n8090 ;
  assign n15711 = n3075 & ~n4169 ;
  assign n15712 = n14134 & n15711 ;
  assign n15714 = n15713 ^ n15712 ^ 1'b0 ;
  assign n15715 = n14422 ^ n13296 ^ 1'b0 ;
  assign n15716 = n15714 & n15715 ;
  assign n15717 = n11173 & n12271 ;
  assign n15718 = n3561 ^ n1833 ^ 1'b0 ;
  assign n15719 = n12112 & ~n15718 ;
  assign n15720 = n10688 ^ n1755 ^ 1'b0 ;
  assign n15721 = n15720 ^ n2091 ^ 1'b0 ;
  assign n15722 = n1800 & ~n4056 ;
  assign n15723 = x106 | n4853 ;
  assign n15724 = n3314 & ~n15723 ;
  assign n15725 = n1016 & n15724 ;
  assign n15726 = ~n7776 & n12911 ;
  assign n15727 = ~n5872 & n15726 ;
  assign n15728 = n10351 & n15551 ;
  assign n15729 = n487 | n7884 ;
  assign n15730 = ~n3611 & n7987 ;
  assign n15731 = n3142 & n15730 ;
  assign n15732 = n5870 ^ n1838 ^ 1'b0 ;
  assign n15733 = n731 | n7739 ;
  assign n15734 = n15733 ^ n4180 ^ 1'b0 ;
  assign n15735 = n542 & n15734 ;
  assign n15736 = n2979 ^ n1790 ^ 1'b0 ;
  assign n15737 = n2091 | n15736 ;
  assign n15738 = n2585 & n8354 ;
  assign n15739 = n376 & n15738 ;
  assign n15740 = n15739 ^ n882 ^ 1'b0 ;
  assign n15741 = n9865 & n15740 ;
  assign n15742 = n15737 | n15741 ;
  assign n15743 = ~n3611 & n13641 ;
  assign n15744 = n1686 | n15743 ;
  assign n15745 = n9034 | n12726 ;
  assign n15746 = n3539 | n15745 ;
  assign n15747 = ~n4886 & n6651 ;
  assign n15748 = ~n1238 & n9148 ;
  assign n15749 = ~n2638 & n15748 ;
  assign n15750 = n15749 ^ n2530 ^ 1'b0 ;
  assign n15751 = n11892 ^ n2394 ^ n1901 ;
  assign n15752 = n2194 & ~n15751 ;
  assign n15753 = n15752 ^ n7747 ^ 1'b0 ;
  assign n15754 = n7900 ^ n4617 ^ 1'b0 ;
  assign n15755 = n2222 & n15754 ;
  assign n15756 = n15747 ^ n12569 ^ 1'b0 ;
  assign n15757 = n809 | n4351 ;
  assign n15758 = n3428 & ~n15757 ;
  assign n15759 = ~n13467 & n15758 ;
  assign n15760 = n12661 ^ n2517 ^ 1'b0 ;
  assign n15761 = n741 | n15760 ;
  assign n15762 = n15761 ^ n1894 ^ 1'b0 ;
  assign n15763 = n2067 | n3108 ;
  assign n15764 = x86 | n15763 ;
  assign n15765 = n6587 ^ n1793 ^ 1'b0 ;
  assign n15766 = ~n15764 & n15765 ;
  assign n15767 = ~n12530 & n15766 ;
  assign n15768 = n135 & n15767 ;
  assign n15769 = n7475 ^ n7268 ^ 1'b0 ;
  assign n15770 = n2326 ^ n2142 ^ 1'b0 ;
  assign n15771 = n12317 ^ n673 ^ 1'b0 ;
  assign n15772 = n6811 ^ n6623 ^ 1'b0 ;
  assign n15773 = n2578 & n15484 ;
  assign n15774 = n12147 ^ n9931 ^ 1'b0 ;
  assign n15775 = ~n4303 & n15774 ;
  assign n15776 = n5574 ^ n1930 ^ 1'b0 ;
  assign n15777 = n14740 & n15776 ;
  assign n15778 = n3651 & n6401 ;
  assign n15779 = ~n15777 & n15778 ;
  assign n15780 = n5223 & n13302 ;
  assign n15781 = n8224 | n12655 ;
  assign n15782 = n2653 | n15781 ;
  assign n15783 = x11 & n4674 ;
  assign n15784 = n13395 ^ n9222 ^ n159 ;
  assign n15785 = n7989 & ~n9302 ;
  assign n15786 = n15784 & n15785 ;
  assign n15787 = n2792 & ~n2896 ;
  assign n15788 = n15787 ^ n5720 ^ 1'b0 ;
  assign n15789 = ~n4654 & n12472 ;
  assign n15790 = n1984 ^ n618 ^ 1'b0 ;
  assign n15791 = n4819 & n6438 ;
  assign n15792 = n12315 ^ n390 ^ 1'b0 ;
  assign n15793 = ~n3932 & n15792 ;
  assign n15794 = n15793 ^ n13863 ^ 1'b0 ;
  assign n15795 = n15794 ^ n10901 ^ n4840 ;
  assign n15797 = n2314 & n14852 ;
  assign n15796 = n4234 & n14858 ;
  assign n15798 = n15797 ^ n15796 ^ 1'b0 ;
  assign n15799 = n15798 ^ n10259 ^ 1'b0 ;
  assign n15800 = n1365 ^ n311 ^ 1'b0 ;
  assign n15801 = n12425 & n15800 ;
  assign n15802 = n5960 ^ n1147 ^ 1'b0 ;
  assign n15803 = n15802 ^ n10225 ^ 1'b0 ;
  assign n15804 = n6922 ^ n671 ^ 1'b0 ;
  assign n15805 = ~n3677 & n15804 ;
  assign n15806 = n15803 & ~n15805 ;
  assign n15807 = n6534 | n11491 ;
  assign n15808 = n10443 ^ n7020 ^ 1'b0 ;
  assign n15809 = n211 & ~n10263 ;
  assign n15810 = n15809 ^ n15251 ^ 1'b0 ;
  assign n15811 = ~n3289 & n6283 ;
  assign n15812 = ~n15523 & n15811 ;
  assign n15813 = n7953 & ~n12585 ;
  assign n15814 = n8767 & ~n15813 ;
  assign n15815 = n9019 ^ n2385 ^ 1'b0 ;
  assign n15816 = n1493 & n15815 ;
  assign n15817 = n6470 & n12509 ;
  assign n15818 = n8302 & n15817 ;
  assign n15819 = n15818 ^ n7715 ^ 1'b0 ;
  assign n15820 = ~n15816 & n15819 ;
  assign n15821 = x87 & ~n356 ;
  assign n15822 = ~n2480 & n15821 ;
  assign n15823 = n15822 ^ n7635 ^ 1'b0 ;
  assign n15824 = n288 | n722 ;
  assign n15825 = n270 ^ x97 ^ 1'b0 ;
  assign n15826 = ~n904 & n15825 ;
  assign n15827 = n13132 ^ n12434 ^ 1'b0 ;
  assign n15828 = ~n9517 & n15827 ;
  assign n15829 = ~n4079 & n8991 ;
  assign n15830 = ~n11482 & n15829 ;
  assign n15831 = ~n6495 & n9378 ;
  assign n15832 = n15830 & n15831 ;
  assign n15833 = n4942 & ~n6006 ;
  assign n15834 = n4962 ^ n2839 ^ 1'b0 ;
  assign n15835 = n15833 & n15834 ;
  assign n15836 = n9576 | n15835 ;
  assign n15837 = n3060 & ~n15438 ;
  assign n15838 = n4965 & n15837 ;
  assign n15839 = n15838 ^ n1456 ^ 1'b0 ;
  assign n15840 = n2755 | n9459 ;
  assign n15841 = n15840 ^ n163 ^ 1'b0 ;
  assign n15842 = ~n502 & n3489 ;
  assign n15843 = ~n15841 & n15842 ;
  assign n15844 = ~n15839 & n15843 ;
  assign n15845 = n616 & ~n8921 ;
  assign n15846 = ~n766 & n15845 ;
  assign n15847 = ~n7810 & n14147 ;
  assign n15848 = x74 & n15847 ;
  assign n15849 = n213 & n7847 ;
  assign n15850 = ~n5962 & n15849 ;
  assign n15851 = ~n1572 & n15850 ;
  assign n15852 = n5840 ^ n753 ^ 1'b0 ;
  assign n15853 = ~n1072 & n9082 ;
  assign n15854 = n15853 ^ n7955 ^ 1'b0 ;
  assign n15855 = n15854 ^ n3281 ^ 1'b0 ;
  assign n15856 = n8986 | n11072 ;
  assign n15857 = n15855 & ~n15856 ;
  assign n15858 = n15857 ^ n5941 ^ 1'b0 ;
  assign n15859 = n4817 & n14531 ;
  assign n15860 = n847 & n1655 ;
  assign n15861 = n1519 & n15860 ;
  assign n15862 = n3872 ^ n3486 ^ 1'b0 ;
  assign n15863 = ~n851 & n3426 ;
  assign n15864 = n15862 & ~n15863 ;
  assign n15865 = n3090 & ~n12966 ;
  assign n15866 = ~n15864 & n15865 ;
  assign n15867 = n1037 | n2423 ;
  assign n15868 = n15867 ^ n10629 ^ 1'b0 ;
  assign n15869 = n12499 & n15868 ;
  assign n15870 = n2179 & n14032 ;
  assign n15871 = n13294 ^ n3878 ^ 1'b0 ;
  assign n15872 = n15871 ^ n13743 ^ n10126 ;
  assign n15873 = n2808 | n14900 ;
  assign n15874 = n4364 ^ n4062 ^ 1'b0 ;
  assign n15875 = n6019 | n15874 ;
  assign n15876 = n7299 & ~n15875 ;
  assign n15877 = n15873 & n15876 ;
  assign n15878 = n1782 & n15877 ;
  assign n15879 = n4062 ^ n1181 ^ 1'b0 ;
  assign n15880 = n6092 & ~n15879 ;
  assign n15881 = n7253 | n10157 ;
  assign n15882 = n7920 | n15881 ;
  assign n15883 = n4428 & ~n11863 ;
  assign n15884 = n3290 | n3774 ;
  assign n15885 = x52 & n14986 ;
  assign n15886 = n15885 ^ n15479 ^ 1'b0 ;
  assign n15887 = n198 & n1022 ;
  assign n15888 = n510 & n15887 ;
  assign n15889 = n15888 ^ n3201 ^ 1'b0 ;
  assign n15891 = ~n1691 & n2367 ;
  assign n15890 = n3691 ^ n2953 ^ 1'b0 ;
  assign n15892 = n15891 ^ n15890 ^ 1'b0 ;
  assign n15894 = ~n6473 & n6553 ;
  assign n15893 = ~n4298 & n13027 ;
  assign n15895 = n15894 ^ n15893 ^ n10862 ;
  assign n15896 = ~n507 & n4895 ;
  assign n15897 = n15896 ^ n2399 ^ 1'b0 ;
  assign n15900 = x74 & ~n3262 ;
  assign n15901 = n15900 ^ n10539 ^ 1'b0 ;
  assign n15898 = n5985 ^ n5223 ^ 1'b0 ;
  assign n15899 = n15898 ^ n3132 ^ 1'b0 ;
  assign n15902 = n15901 ^ n15899 ^ 1'b0 ;
  assign n15903 = n14180 ^ n571 ^ 1'b0 ;
  assign n15904 = n6089 & ~n15903 ;
  assign n15905 = n2603 & n10905 ;
  assign n15906 = n13132 & n15905 ;
  assign n15907 = n5937 ^ n3833 ^ 1'b0 ;
  assign n15908 = n7463 & n15907 ;
  assign n15909 = n15908 ^ n3805 ^ 1'b0 ;
  assign n15910 = n8145 & ~n10692 ;
  assign n15911 = ~n916 & n15910 ;
  assign n15912 = n15911 ^ n418 ^ 1'b0 ;
  assign n15913 = n9607 ^ n2826 ^ 1'b0 ;
  assign n15914 = n971 & ~n1414 ;
  assign n15915 = n2165 | n15914 ;
  assign n15916 = n10314 & ~n15915 ;
  assign n15917 = n12415 ^ n3324 ^ 1'b0 ;
  assign n15918 = n15588 ^ n11164 ^ 1'b0 ;
  assign n15919 = ~n15917 & n15918 ;
  assign n15920 = n13127 | n15272 ;
  assign n15921 = n15920 ^ n9133 ^ 1'b0 ;
  assign n15922 = n15830 ^ n6249 ^ 1'b0 ;
  assign n15923 = n1228 | n7273 ;
  assign n15924 = n3496 & n5666 ;
  assign n15925 = ~n3496 & n15924 ;
  assign n15926 = n2479 | n15925 ;
  assign n15927 = n2479 & ~n15926 ;
  assign n15928 = n7468 ^ n5016 ^ 1'b0 ;
  assign n15929 = ~n4316 & n15928 ;
  assign n15930 = ~n6964 & n15929 ;
  assign n15931 = ~n5290 & n15930 ;
  assign n15932 = ~n3428 & n3890 ;
  assign n15933 = n15932 ^ n9770 ^ 1'b0 ;
  assign n15934 = n7001 ^ n1170 ^ 1'b0 ;
  assign n15935 = n9707 | n15934 ;
  assign n15936 = n2787 & ~n11348 ;
  assign n15937 = n1197 & n15936 ;
  assign n15938 = n7132 ^ n831 ^ 1'b0 ;
  assign n15939 = ~n15937 & n15938 ;
  assign n15942 = n2324 ^ n2085 ^ 1'b0 ;
  assign n15943 = n733 & n15942 ;
  assign n15940 = n8518 ^ n4032 ^ 1'b0 ;
  assign n15941 = n10832 & n15940 ;
  assign n15944 = n15943 ^ n15941 ^ 1'b0 ;
  assign n15945 = x111 & ~n4170 ;
  assign n15946 = n15945 ^ n11958 ^ 1'b0 ;
  assign n15947 = n747 | n15946 ;
  assign n15948 = n624 | n2960 ;
  assign n15949 = n9076 & ~n15948 ;
  assign n15950 = ( n4768 & ~n4944 ) | ( n4768 & n7614 ) | ( ~n4944 & n7614 ) ;
  assign n15951 = n11111 ^ n1351 ^ 1'b0 ;
  assign n15952 = n528 & ~n6918 ;
  assign n15953 = ~n11128 & n15952 ;
  assign n15954 = n6214 & ~n7129 ;
  assign n15955 = n15954 ^ n10699 ^ 1'b0 ;
  assign n15956 = n15955 ^ n12412 ^ 1'b0 ;
  assign n15957 = n1993 & ~n3953 ;
  assign n15958 = n5320 & n15957 ;
  assign n15959 = n15958 ^ n6315 ^ 1'b0 ;
  assign n15960 = n1634 & n4662 ;
  assign n15961 = n2735 | n3089 ;
  assign n15962 = n13666 ^ n8241 ^ 1'b0 ;
  assign n15963 = ~n2771 & n15962 ;
  assign n15964 = n12762 & ~n15963 ;
  assign n15965 = n6026 & n10939 ;
  assign n15966 = n12197 | n15965 ;
  assign n15967 = n15966 ^ n2986 ^ 1'b0 ;
  assign n15968 = x47 & ~n13501 ;
  assign n15969 = ~n2478 & n15968 ;
  assign n15970 = x33 & ~n14902 ;
  assign n15971 = n14902 & n15970 ;
  assign n15972 = n2276 & ~n15971 ;
  assign n15973 = ~n2276 & n15972 ;
  assign n15974 = n3978 | n4858 ;
  assign n15975 = n4858 & ~n15974 ;
  assign n15976 = n15514 & ~n15975 ;
  assign n15977 = n15973 & n15976 ;
  assign n15978 = ~n1766 & n10669 ;
  assign n15979 = ~n4060 & n15978 ;
  assign n15980 = ~n11546 & n15979 ;
  assign n15981 = n12741 ^ n12214 ^ 1'b0 ;
  assign n15982 = ~n15980 & n15981 ;
  assign n15983 = n3251 & ~n8769 ;
  assign n15984 = n2409 & ~n11773 ;
  assign n15985 = n7911 ^ n7543 ^ 1'b0 ;
  assign n15986 = n1790 ^ n1770 ^ 1'b0 ;
  assign n15987 = n13633 | n15986 ;
  assign n15988 = n15987 ^ n13925 ^ 1'b0 ;
  assign n15989 = ~n5214 & n15988 ;
  assign n15990 = ~n5611 & n11374 ;
  assign n15991 = n15990 ^ n2330 ^ 1'b0 ;
  assign n15993 = n7767 ^ n2079 ^ 1'b0 ;
  assign n15992 = n6685 | n15761 ;
  assign n15994 = n15993 ^ n15992 ^ 1'b0 ;
  assign n15995 = ~n2838 & n9836 ;
  assign n15996 = n8636 & n15995 ;
  assign n15997 = n4505 ^ n2470 ^ 1'b0 ;
  assign n15998 = n15996 & ~n15997 ;
  assign n15999 = ~n355 & n1280 ;
  assign n16002 = ~n4860 & n5224 ;
  assign n16000 = n155 & n3874 ;
  assign n16001 = ~n5165 & n16000 ;
  assign n16003 = n16002 ^ n16001 ^ 1'b0 ;
  assign n16004 = ( ~n642 & n6232 ) | ( ~n642 & n16003 ) | ( n6232 & n16003 ) ;
  assign n16005 = n15799 ^ n6381 ^ 1'b0 ;
  assign n16006 = n4650 ^ n2423 ^ 1'b0 ;
  assign n16007 = n16006 ^ n15969 ^ 1'b0 ;
  assign n16008 = ~n338 & n4081 ;
  assign n16009 = n1756 ^ n831 ^ 1'b0 ;
  assign n16010 = n16009 ^ n7573 ^ 1'b0 ;
  assign n16011 = n16008 & n16010 ;
  assign n16012 = n5358 & n14257 ;
  assign n16013 = n2892 & n9082 ;
  assign n16014 = n695 | n819 ;
  assign n16015 = n16014 ^ n302 ^ 1'b0 ;
  assign n16016 = n14621 ^ n549 ^ 1'b0 ;
  assign n16017 = n2785 | n16016 ;
  assign n16018 = n16017 ^ n11291 ^ 1'b0 ;
  assign n16019 = n150 & ~n3314 ;
  assign n16020 = n3722 & n16019 ;
  assign n16021 = n16020 ^ n4214 ^ 1'b0 ;
  assign n16022 = n15957 & ~n16021 ;
  assign n16023 = n13236 ^ n10132 ^ 1'b0 ;
  assign n16024 = n1133 & n2308 ;
  assign n16025 = n12743 & ~n13670 ;
  assign n16026 = n2299 & ~n12013 ;
  assign n16027 = ( ~n4999 & n8763 ) | ( ~n4999 & n16026 ) | ( n8763 & n16026 ) ;
  assign n16028 = ~n15705 & n16027 ;
  assign n16029 = ( n8127 & n10544 ) | ( n8127 & n11380 ) | ( n10544 & n11380 ) ;
  assign n16030 = ~n10198 & n12351 ;
  assign n16031 = n14631 ^ n9030 ^ n8735 ;
  assign n16032 = n441 | n16031 ;
  assign n16033 = n6504 & ~n16032 ;
  assign n16034 = n3556 & n6180 ;
  assign n16035 = ~n3765 & n7681 ;
  assign n16036 = ~n428 & n2979 ;
  assign n16037 = ~n1255 & n10473 ;
  assign n16038 = ~n11782 & n16037 ;
  assign n16039 = n3632 ^ n3434 ^ 1'b0 ;
  assign n16040 = n7093 & ~n16039 ;
  assign n16041 = n2602 & n16040 ;
  assign n16042 = ~n7088 & n16041 ;
  assign n16043 = n806 & ~n13224 ;
  assign n16045 = n8783 ^ n3707 ^ 1'b0 ;
  assign n16046 = x76 | n16045 ;
  assign n16047 = n9217 & ~n16046 ;
  assign n16044 = n2009 & ~n9220 ;
  assign n16048 = n16047 ^ n16044 ^ 1'b0 ;
  assign n16049 = ~n16043 & n16048 ;
  assign n16050 = n10691 ^ n2649 ^ 1'b0 ;
  assign n16051 = ~n7259 & n16050 ;
  assign n16052 = ~n5985 & n16051 ;
  assign n16053 = n3450 & n3658 ;
  assign n16054 = n16053 ^ n6352 ^ 1'b0 ;
  assign n16055 = n11858 ^ n10831 ^ 1'b0 ;
  assign n16056 = ~n934 & n12635 ;
  assign n16057 = ~n3706 & n6954 ;
  assign n16058 = n16057 ^ n3930 ^ 1'b0 ;
  assign n16061 = n5590 | n9389 ;
  assign n16062 = n16061 ^ n2932 ^ 1'b0 ;
  assign n16059 = n1425 & ~n12817 ;
  assign n16060 = n10220 & n16059 ;
  assign n16063 = n16062 ^ n16060 ^ 1'b0 ;
  assign n16064 = x99 & ~n4147 ;
  assign n16065 = ~n3592 & n16064 ;
  assign n16066 = n5819 | n16065 ;
  assign n16067 = n2215 & n3589 ;
  assign n16068 = ~n1861 & n8220 ;
  assign n16069 = n2835 & n9456 ;
  assign n16070 = ~n15945 & n16069 ;
  assign n16071 = n354 & ~n15096 ;
  assign n16072 = n5652 & ~n14166 ;
  assign n16073 = n9458 & n16072 ;
  assign n16074 = n549 | n7681 ;
  assign n16075 = ( n11889 & n14731 ) | ( n11889 & n16074 ) | ( n14731 & n16074 ) ;
  assign n16076 = n11496 ^ n9724 ^ 1'b0 ;
  assign n16077 = ~n3965 & n16076 ;
  assign n16078 = n11918 & ~n16077 ;
  assign n16080 = ~n211 & n3786 ;
  assign n16081 = n1222 | n16080 ;
  assign n16079 = x60 | n9604 ;
  assign n16082 = n16081 ^ n16079 ^ 1'b0 ;
  assign n16083 = n1534 | n7339 ;
  assign n16084 = n1331 & ~n3611 ;
  assign n16085 = ~n4310 & n16084 ;
  assign n16086 = n16085 ^ n6445 ^ 1'b0 ;
  assign n16087 = n2633 & ~n16086 ;
  assign n16088 = n12923 & n16087 ;
  assign n16089 = ~n5265 & n6311 ;
  assign n16090 = n16089 ^ n10918 ^ 1'b0 ;
  assign n16091 = n5213 ^ n2355 ^ 1'b0 ;
  assign n16092 = n6926 & ~n16091 ;
  assign n16093 = x59 & ~n4071 ;
  assign n16094 = n13929 & n16093 ;
  assign n16095 = n16094 ^ n6144 ^ 1'b0 ;
  assign n16096 = n9344 & ~n9458 ;
  assign n16098 = n1987 | n8840 ;
  assign n16099 = n13895 & ~n16098 ;
  assign n16097 = x21 | n1105 ;
  assign n16100 = n16099 ^ n16097 ^ 1'b0 ;
  assign n16101 = n16096 & ~n16100 ;
  assign n16102 = ~n8577 & n16101 ;
  assign n16103 = n7855 ^ n6064 ^ 1'b0 ;
  assign n16104 = ~n4778 & n13991 ;
  assign n16105 = n3443 | n15790 ;
  assign n16106 = n16105 ^ n14489 ^ 1'b0 ;
  assign n16107 = n12825 ^ n1640 ^ 1'b0 ;
  assign n16108 = x42 & n10033 ;
  assign n16109 = n16108 ^ n402 ^ 1'b0 ;
  assign n16110 = n16109 ^ n8508 ^ n2191 ;
  assign n16111 = n1480 | n1841 ;
  assign n16112 = n7096 | n16111 ;
  assign n16113 = n3270 | n8577 ;
  assign n16114 = ~n430 & n1842 ;
  assign n16115 = n16114 ^ n3800 ^ 1'b0 ;
  assign n16116 = ~n16113 & n16115 ;
  assign n16117 = n3324 | n15301 ;
  assign n16118 = n16117 ^ n8705 ^ 1'b0 ;
  assign n16119 = ~n1954 & n16118 ;
  assign n16120 = n16119 ^ n11695 ^ 1'b0 ;
  assign n16121 = n16120 ^ n1823 ^ 1'b0 ;
  assign n16122 = n16116 & n16121 ;
  assign n16123 = n15254 ^ n5541 ^ 1'b0 ;
  assign n16124 = n2155 & ~n16123 ;
  assign n16125 = n16124 ^ n16062 ^ 1'b0 ;
  assign n16126 = n3362 ^ n2561 ^ 1'b0 ;
  assign n16127 = n4390 & n11961 ;
  assign n16128 = n15214 & n16127 ;
  assign n16129 = n11347 | n12812 ;
  assign n16130 = n2453 ^ n229 ^ 1'b0 ;
  assign n16131 = n6148 ^ n2660 ^ n1875 ;
  assign n16132 = n16131 ^ n12045 ^ 1'b0 ;
  assign n16133 = n10087 & ~n16132 ;
  assign n16134 = ~n4587 & n6325 ;
  assign n16136 = n9343 ^ n1540 ^ 1'b0 ;
  assign n16137 = ~n2642 & n16136 ;
  assign n16135 = n1147 | n3298 ;
  assign n16138 = n16137 ^ n16135 ^ 1'b0 ;
  assign n16139 = n12432 ^ n3525 ^ 1'b0 ;
  assign n16140 = n6070 & ~n6542 ;
  assign n16141 = n2073 | n8400 ;
  assign n16142 = n16141 ^ n1368 ^ 1'b0 ;
  assign n16143 = n16142 ^ x16 ^ 1'b0 ;
  assign n16144 = n14441 & ~n16143 ;
  assign n16145 = ~n2281 & n2806 ;
  assign n16146 = n1179 ^ n868 ^ 1'b0 ;
  assign n16147 = n16146 ^ n8322 ^ 1'b0 ;
  assign n16148 = n788 & ~n16147 ;
  assign n16149 = ~n238 & n10193 ;
  assign n16150 = n2233 & n16149 ;
  assign n16151 = n5825 & ~n10622 ;
  assign n16152 = ~n3764 & n10866 ;
  assign n16153 = n16152 ^ n13958 ^ 1'b0 ;
  assign n16154 = ~n894 & n10653 ;
  assign n16155 = n16154 ^ n13847 ^ 1'b0 ;
  assign n16156 = n15454 ^ n9143 ^ 1'b0 ;
  assign n16157 = n7585 & n16156 ;
  assign n16158 = n11119 ^ n9568 ^ 1'b0 ;
  assign n16159 = n3373 & ~n4217 ;
  assign n16160 = ~n656 & n2085 ;
  assign n16161 = n12520 & n16160 ;
  assign n16162 = n10273 & n16161 ;
  assign n16163 = n6499 & n16162 ;
  assign n16164 = n10927 | n13666 ;
  assign n16165 = n5986 & ~n16164 ;
  assign n16166 = ~n12911 & n16165 ;
  assign n16167 = ~n7944 & n8660 ;
  assign n16168 = n16167 ^ n3445 ^ 1'b0 ;
  assign n16169 = n3764 ^ n3482 ^ 1'b0 ;
  assign n16170 = n510 | n16169 ;
  assign n16171 = n5814 ^ n5282 ^ 1'b0 ;
  assign n16172 = n13838 ^ n2121 ^ 1'b0 ;
  assign n16173 = ~n13440 & n15038 ;
  assign n16174 = ~n3140 & n9230 ;
  assign n16175 = ~n13053 & n16174 ;
  assign n16176 = n16175 ^ n2961 ^ 1'b0 ;
  assign n16177 = ~n5228 & n11787 ;
  assign n16178 = ~n3504 & n16177 ;
  assign n16179 = n11045 & n16178 ;
  assign n16180 = ~n8369 & n10452 ;
  assign n16182 = n1856 ^ n420 ^ 1'b0 ;
  assign n16181 = n3919 & n5429 ;
  assign n16183 = n16182 ^ n16181 ^ 1'b0 ;
  assign n16184 = n9229 & n10232 ;
  assign n16185 = n16184 ^ n6712 ^ 1'b0 ;
  assign n16186 = n8247 & ~n10517 ;
  assign n16187 = ~n4638 & n16186 ;
  assign n16188 = ~n287 & n4219 ;
  assign n16189 = n1341 | n9745 ;
  assign n16190 = n1795 | n16189 ;
  assign n16191 = ~n3544 & n13364 ;
  assign n16192 = n6042 & ~n10506 ;
  assign n16193 = ~n9803 & n11188 ;
  assign n16194 = n5503 ^ n1162 ^ 1'b0 ;
  assign n16195 = n387 & n689 ;
  assign n16196 = ~n689 & n16195 ;
  assign n16197 = n3628 | n16196 ;
  assign n16198 = n4390 | n16197 ;
  assign n16200 = n1848 & ~n2067 ;
  assign n16201 = n4911 & n16200 ;
  assign n16202 = n4393 & ~n16201 ;
  assign n16203 = ~n5682 & n16202 ;
  assign n16199 = n3343 | n13625 ;
  assign n16204 = n16203 ^ n16199 ^ 1'b0 ;
  assign n16205 = n6218 | n12795 ;
  assign n16206 = n10338 ^ n5215 ^ 1'b0 ;
  assign n16207 = n2608 & n16206 ;
  assign n16208 = n9528 ^ x116 ^ 1'b0 ;
  assign n16209 = ~n7873 & n8290 ;
  assign n16210 = n8825 ^ n1418 ^ 1'b0 ;
  assign n16211 = n16209 & n16210 ;
  assign n16212 = ~n2407 & n2949 ;
  assign n16213 = n16212 ^ n8129 ^ 1'b0 ;
  assign n16214 = n2188 & ~n16213 ;
  assign n16215 = n16214 ^ n2630 ^ 1'b0 ;
  assign n16216 = n1588 | n9571 ;
  assign n16217 = n16215 & ~n16216 ;
  assign n16218 = n1387 & n1711 ;
  assign n16219 = n3078 | n4218 ;
  assign n16220 = n194 & ~n16219 ;
  assign n16221 = ~n632 & n16046 ;
  assign n16222 = n6719 ^ n131 ^ 1'b0 ;
  assign n16223 = n12313 ^ n1499 ^ 1'b0 ;
  assign n16224 = ~n16222 & n16223 ;
  assign n16225 = n9357 ^ n867 ^ n281 ;
  assign n16226 = n16225 ^ n9248 ^ 1'b0 ;
  assign n16227 = n4853 & n16226 ;
  assign n16228 = n16227 ^ n356 ^ 1'b0 ;
  assign n16229 = ~x76 & n6747 ;
  assign n16230 = n9868 ^ n8069 ^ 1'b0 ;
  assign n16231 = ~n4459 & n16230 ;
  assign n16232 = n2265 & n13548 ;
  assign n16233 = ~n16231 & n16232 ;
  assign n16234 = n2815 & n6634 ;
  assign n16235 = n9860 & ~n14216 ;
  assign n16236 = ~n5434 & n16235 ;
  assign n16237 = ~n8799 & n14607 ;
  assign n16238 = ~n1637 & n5338 ;
  assign n16239 = n12503 ^ n7356 ^ 1'b0 ;
  assign n16240 = n3843 & n16239 ;
  assign n16246 = n5045 & ~n8491 ;
  assign n16241 = n8190 & n10890 ;
  assign n16242 = ~n4579 & n16241 ;
  assign n16243 = n8529 ^ n4598 ^ 1'b0 ;
  assign n16244 = x47 | n16243 ;
  assign n16245 = n16242 | n16244 ;
  assign n16247 = n16246 ^ n16245 ^ 1'b0 ;
  assign n16248 = n4655 ^ n2091 ^ 1'b0 ;
  assign n16249 = n8633 & ~n9096 ;
  assign n16250 = n2506 & ~n4921 ;
  assign n16251 = n3648 & ~n6542 ;
  assign n16252 = n8679 | n9798 ;
  assign n16253 = n16251 & ~n16252 ;
  assign n16254 = n14129 ^ n7707 ^ 1'b0 ;
  assign n16255 = ( ~n1329 & n2456 ) | ( ~n1329 & n9252 ) | ( n2456 & n9252 ) ;
  assign n16256 = n8575 & n16255 ;
  assign n16257 = n13395 ^ n3509 ^ 1'b0 ;
  assign n16258 = n4289 | n4765 ;
  assign n16259 = n16258 ^ n7574 ^ 1'b0 ;
  assign n16260 = n1749 & ~n3926 ;
  assign n16261 = n16260 ^ n285 ^ 1'b0 ;
  assign n16262 = n7194 ^ n6921 ^ 1'b0 ;
  assign n16263 = n7752 & ~n16262 ;
  assign n16264 = n985 & n16263 ;
  assign n16265 = n16264 ^ n3380 ^ 1'b0 ;
  assign n16266 = n1206 & n5438 ;
  assign n16267 = n16266 ^ n5159 ^ 1'b0 ;
  assign n16268 = n13296 ^ n3107 ^ 1'b0 ;
  assign n16269 = ~n1226 & n16268 ;
  assign n16270 = n11309 ^ n6220 ^ 1'b0 ;
  assign n16271 = n8273 ^ n4643 ^ 1'b0 ;
  assign n16272 = n4679 | n16271 ;
  assign n16273 = n3722 & n7179 ;
  assign n16274 = ~n13783 & n16273 ;
  assign n16275 = n4298 | n14304 ;
  assign n16276 = n4241 ^ n2119 ^ 1'b0 ;
  assign n16277 = n638 | n1983 ;
  assign n16278 = n16277 ^ n2923 ^ 1'b0 ;
  assign n16279 = n14975 & n16278 ;
  assign n16280 = n16279 ^ n7114 ^ x37 ;
  assign n16281 = n15320 ^ n14956 ^ 1'b0 ;
  assign n16282 = n8465 | n16281 ;
  assign n16283 = n10811 ^ n1851 ^ 1'b0 ;
  assign n16284 = ~n13108 & n16283 ;
  assign n16285 = n12320 ^ n10310 ^ 1'b0 ;
  assign n16286 = n1185 & n16285 ;
  assign n16287 = n9410 & ~n12088 ;
  assign n16288 = n16287 ^ n4615 ^ 1'b0 ;
  assign n16289 = n4567 & ~n16288 ;
  assign n16290 = n10173 & n12525 ;
  assign n16291 = n5789 ^ n928 ^ 1'b0 ;
  assign n16292 = n14902 | n16291 ;
  assign n16293 = ~n700 & n16292 ;
  assign n16294 = n2650 | n5746 ;
  assign n16295 = n16294 ^ x22 ^ 1'b0 ;
  assign n16296 = n16293 & ~n16295 ;
  assign n16297 = n1662 & ~n2883 ;
  assign n16298 = n16297 ^ n1202 ^ 1'b0 ;
  assign n16299 = n4289 | n16298 ;
  assign n16305 = n1004 & n2718 ;
  assign n16306 = n4971 & n8276 ;
  assign n16307 = n16306 ^ n886 ^ 1'b0 ;
  assign n16308 = n16307 ^ x110 ^ 1'b0 ;
  assign n16309 = n16305 & n16308 ;
  assign n16310 = ~n221 & n16309 ;
  assign n16300 = n4705 ^ n1048 ^ 1'b0 ;
  assign n16301 = n12423 ^ n830 ^ 1'b0 ;
  assign n16302 = n3784 & ~n16301 ;
  assign n16303 = n16302 ^ n10848 ^ 1'b0 ;
  assign n16304 = ~n16300 & n16303 ;
  assign n16311 = n16310 ^ n16304 ^ 1'b0 ;
  assign n16312 = n629 & n1103 ;
  assign n16313 = n16312 ^ n1618 ^ 1'b0 ;
  assign n16314 = n13694 & n16313 ;
  assign n16315 = n5810 ^ n5739 ^ 1'b0 ;
  assign n16316 = n926 & ~n2459 ;
  assign n16317 = n16316 ^ n895 ^ 1'b0 ;
  assign n16318 = n6445 & ~n16317 ;
  assign n16319 = n12862 ^ n11274 ^ n931 ;
  assign n16320 = x98 & ~n9359 ;
  assign n16321 = n16320 ^ n1589 ^ 1'b0 ;
  assign n16322 = n16321 ^ n5938 ^ 1'b0 ;
  assign n16323 = n3696 & n16322 ;
  assign n16324 = ~n2389 & n6570 ;
  assign n16325 = ~n10760 & n14581 ;
  assign n16326 = n16325 ^ n945 ^ 1'b0 ;
  assign n16327 = n7017 | n11166 ;
  assign n16328 = ~n5160 & n11684 ;
  assign n16329 = n16328 ^ n2689 ^ 1'b0 ;
  assign n16330 = n134 & n595 ;
  assign n16331 = n16330 ^ n8775 ^ 1'b0 ;
  assign n16332 = n1374 | n3754 ;
  assign n16333 = n888 & ~n16332 ;
  assign n16334 = n9691 ^ n4993 ^ 1'b0 ;
  assign n16335 = n2821 | n3359 ;
  assign n16336 = n4582 & ~n16335 ;
  assign n16337 = n6311 ^ n4117 ^ 1'b0 ;
  assign n16339 = n4749 ^ n4158 ^ 1'b0 ;
  assign n16340 = n7605 & n16339 ;
  assign n16338 = n11301 ^ n5972 ^ 1'b0 ;
  assign n16341 = n16340 ^ n16338 ^ 1'b0 ;
  assign n16342 = ~n1051 & n4276 ;
  assign n16343 = n16342 ^ n4160 ^ 1'b0 ;
  assign n16344 = n16343 ^ n12172 ^ 1'b0 ;
  assign n16345 = n5144 & ~n7000 ;
  assign n16346 = n13682 ^ n1504 ^ n1457 ;
  assign n16347 = n4779 ^ n4605 ^ 1'b0 ;
  assign n16348 = n16347 ^ n15663 ^ n6131 ;
  assign n16349 = n12295 | n14041 ;
  assign n16350 = n16349 ^ n9452 ^ 1'b0 ;
  assign n16351 = n4867 & ~n6645 ;
  assign n16352 = n10622 | n16203 ;
  assign n16353 = n16352 ^ n11547 ^ 1'b0 ;
  assign n16354 = ~n3220 & n16353 ;
  assign n16355 = n3904 ^ n2181 ^ 1'b0 ;
  assign n16356 = n2099 & ~n4413 ;
  assign n16357 = n4413 & n16356 ;
  assign n16358 = n1681 & ~n7917 ;
  assign n16359 = ~n7274 & n16358 ;
  assign n16360 = n10064 & ~n16180 ;
  assign n16361 = n16359 & n16360 ;
  assign n16362 = ~n2876 & n4253 ;
  assign n16363 = n2324 ^ n1423 ^ 1'b0 ;
  assign n16364 = n737 | n13816 ;
  assign n16365 = n13071 & ~n16364 ;
  assign n16366 = n8035 & ~n8439 ;
  assign n16367 = n16366 ^ n9683 ^ 1'b0 ;
  assign n16368 = ~n11592 & n13816 ;
  assign n16369 = n2993 & ~n3166 ;
  assign n16370 = n16369 ^ n3909 ^ 1'b0 ;
  assign n16371 = x2 & ~n16370 ;
  assign n16372 = n15727 ^ n4937 ^ 1'b0 ;
  assign n16373 = n16371 & ~n16372 ;
  assign n16374 = n5072 & n6030 ;
  assign n16375 = n1436 & n3809 ;
  assign n16376 = n3557 ^ n1053 ^ 1'b0 ;
  assign n16377 = n16375 & n16376 ;
  assign n16378 = n16377 ^ n2635 ^ 1'b0 ;
  assign n16379 = n15472 ^ n9864 ^ n5355 ;
  assign n16385 = n1202 & n9000 ;
  assign n16386 = ~n8315 & n16385 ;
  assign n16380 = n433 | n3711 ;
  assign n16381 = n307 & ~n16380 ;
  assign n16382 = n16381 ^ n2023 ^ 1'b0 ;
  assign n16383 = n4804 & ~n16382 ;
  assign n16384 = n6283 & ~n16383 ;
  assign n16387 = n16386 ^ n16384 ^ 1'b0 ;
  assign n16388 = n16387 ^ n11124 ^ 1'b0 ;
  assign n16389 = n7997 & n16388 ;
  assign n16390 = n10954 ^ n2136 ^ 1'b0 ;
  assign n16391 = n16390 ^ n13663 ^ 1'b0 ;
  assign n16392 = ~n2176 & n3080 ;
  assign n16393 = n11202 ^ n2511 ^ 1'b0 ;
  assign n16394 = n13100 ^ n3584 ^ 1'b0 ;
  assign n16395 = ~n14058 & n16394 ;
  assign n16396 = n5676 & n16395 ;
  assign n16397 = n15749 ^ n13993 ^ n3622 ;
  assign n16398 = n11084 ^ n1243 ^ 1'b0 ;
  assign n16399 = n13721 | n16398 ;
  assign n16400 = n4254 & n7547 ;
  assign n16401 = n6370 ^ n4143 ^ 1'b0 ;
  assign n16402 = x59 & n16401 ;
  assign n16403 = ~n5902 & n16402 ;
  assign n16404 = n2000 & n16403 ;
  assign n16405 = n3585 | n6064 ;
  assign n16406 = n13188 & ~n16405 ;
  assign n16407 = n5485 ^ n3452 ^ 1'b0 ;
  assign n16408 = n12369 | n16407 ;
  assign n16409 = n2023 ^ n340 ^ 1'b0 ;
  assign n16410 = n16408 & n16409 ;
  assign n16411 = n8333 ^ n630 ^ 1'b0 ;
  assign n16412 = ( n277 & ~n9722 ) | ( n277 & n16411 ) | ( ~n9722 & n16411 ) ;
  assign n16413 = n9679 ^ x37 ^ 1'b0 ;
  assign n16414 = n4013 & n15290 ;
  assign n16415 = n1808 | n7933 ;
  assign n16416 = n16415 ^ n6480 ^ 1'b0 ;
  assign n16417 = n867 & n16416 ;
  assign n16418 = n5466 ^ n5019 ^ 1'b0 ;
  assign n16419 = n4713 | n16418 ;
  assign n16420 = n14272 & n16419 ;
  assign n16421 = ~n2037 & n13501 ;
  assign n16422 = n9111 & n16421 ;
  assign n16423 = n413 | n15268 ;
  assign n16424 = n1623 | n13895 ;
  assign n16425 = n5704 ^ n4029 ^ 1'b0 ;
  assign n16426 = ~n5708 & n16425 ;
  assign n16427 = n11481 ^ n8993 ^ 1'b0 ;
  assign n16428 = n7129 & ~n11199 ;
  assign n16429 = n16428 ^ n2390 ^ 1'b0 ;
  assign n16430 = n8459 ^ n3135 ^ 1'b0 ;
  assign n16431 = n16429 | n16430 ;
  assign n16432 = n2240 & ~n11762 ;
  assign n16433 = n3584 & n5193 ;
  assign n16434 = n1376 & ~n2847 ;
  assign n16435 = n16434 ^ n3910 ^ 1'b0 ;
  assign n16436 = n12090 & ~n16435 ;
  assign n16437 = n492 | n12230 ;
  assign n16438 = n1708 | n5011 ;
  assign n16439 = x127 & n9075 ;
  assign n16440 = ~n16438 & n16439 ;
  assign n16441 = n4404 & ~n5647 ;
  assign n16442 = n7269 & n14567 ;
  assign n16443 = n2834 & n16442 ;
  assign n16444 = n9911 ^ n7548 ^ 1'b0 ;
  assign n16445 = n13680 & n16444 ;
  assign n16446 = n13446 ^ n10356 ^ 1'b0 ;
  assign n16447 = ~n9848 & n12873 ;
  assign n16448 = n4303 | n4904 ;
  assign n16449 = n4904 & ~n16448 ;
  assign n16450 = n16449 ^ n12836 ^ 1'b0 ;
  assign n16451 = ~n339 & n16450 ;
  assign n16452 = n16451 ^ n5001 ^ 1'b0 ;
  assign n16453 = n5907 ^ n453 ^ 1'b0 ;
  assign n16454 = n4757 | n16453 ;
  assign n16455 = ~n15296 & n16454 ;
  assign n16456 = n1356 & ~n6282 ;
  assign n16457 = n10313 | n16456 ;
  assign n16458 = n478 ^ n153 ^ 1'b0 ;
  assign n16459 = n16457 & ~n16458 ;
  assign n16460 = ~n1996 & n16459 ;
  assign n16461 = n16460 ^ n8505 ^ 1'b0 ;
  assign n16462 = n16461 ^ n4724 ^ 1'b0 ;
  assign n16463 = n8724 & ~n9421 ;
  assign n16464 = n7994 ^ n3403 ^ 1'b0 ;
  assign n16465 = ~n2624 & n8848 ;
  assign n16466 = ~n645 & n16465 ;
  assign n16467 = n11718 ^ x123 ^ 1'b0 ;
  assign n16468 = ~n16466 & n16467 ;
  assign n16469 = n153 & ~n7802 ;
  assign n16470 = n727 & n16469 ;
  assign n16471 = n1724 & n16470 ;
  assign n16472 = n937 & ~n13103 ;
  assign n16473 = n13103 & n16472 ;
  assign n16474 = n4993 & n16473 ;
  assign n16475 = n1170 & ~n4985 ;
  assign n16476 = ~n1170 & n16475 ;
  assign n16477 = n3367 & n16476 ;
  assign n16478 = x38 & ~n1459 ;
  assign n16479 = ~x38 & n16478 ;
  assign n16480 = n16479 ^ n5427 ^ 1'b0 ;
  assign n16481 = n3379 & n16480 ;
  assign n16482 = n16477 & n16481 ;
  assign n16483 = n16482 ^ n610 ^ 1'b0 ;
  assign n16484 = n1080 | n3262 ;
  assign n16485 = n1080 & ~n16484 ;
  assign n16486 = n16485 ^ n14674 ^ 1'b0 ;
  assign n16487 = ~n16483 & n16486 ;
  assign n16488 = n16474 & n16487 ;
  assign n16489 = n13277 & ~n16488 ;
  assign n16490 = n16488 & n16489 ;
  assign n16491 = n5451 & ~n10235 ;
  assign n16492 = n10692 ^ n9175 ^ 1'b0 ;
  assign n16493 = ~n4965 & n16492 ;
  assign n16494 = n16493 ^ n11664 ^ 1'b0 ;
  assign n16495 = n10035 ^ n4805 ^ 1'b0 ;
  assign n16496 = n4761 & n11089 ;
  assign n16497 = ~n12458 & n12551 ;
  assign n16498 = n16497 ^ n14453 ^ 1'b0 ;
  assign n16499 = n5356 ^ n2010 ^ 1'b0 ;
  assign n16500 = n1076 & ~n16499 ;
  assign n16501 = ( ~n1756 & n7905 ) | ( ~n1756 & n8808 ) | ( n7905 & n8808 ) ;
  assign n16502 = n16501 ^ n6234 ^ 1'b0 ;
  assign n16503 = n2638 & ~n16502 ;
  assign n16504 = n4038 & ~n4679 ;
  assign n16505 = n15474 ^ n5243 ^ 1'b0 ;
  assign n16506 = n8179 | n16505 ;
  assign n16507 = n1586 | n6622 ;
  assign n16508 = n4059 ^ n591 ^ 1'b0 ;
  assign n16509 = n6258 | n16508 ;
  assign n16510 = n13132 & n16509 ;
  assign n16511 = n4573 ^ n3667 ^ 1'b0 ;
  assign n16512 = ~n3718 & n16511 ;
  assign n16513 = n3182 & n16512 ;
  assign n16514 = n16513 ^ n2992 ^ 1'b0 ;
  assign n16515 = n5230 & ~n6544 ;
  assign n16516 = n16515 ^ n14788 ^ 1'b0 ;
  assign n16517 = n4076 & n11258 ;
  assign n16518 = n11057 & n16517 ;
  assign n16519 = n12426 ^ n5336 ^ n3547 ;
  assign n16520 = n11802 ^ n305 ^ 1'b0 ;
  assign n16521 = ~n2636 & n5691 ;
  assign n16522 = n16521 ^ n11076 ^ 1'b0 ;
  assign n16523 = n4148 & ~n16522 ;
  assign n16524 = n737 & n11367 ;
  assign n16525 = n6880 | n8333 ;
  assign n16526 = n11872 ^ n132 ^ 1'b0 ;
  assign n16527 = n980 | n16526 ;
  assign n16528 = n11474 ^ n1470 ^ 1'b0 ;
  assign n16529 = n2986 & n16528 ;
  assign n16530 = n16527 | n16529 ;
  assign n16531 = ~n5463 & n8050 ;
  assign n16532 = ~n14705 & n16531 ;
  assign n16533 = n9371 ^ n7404 ^ 1'b0 ;
  assign n16534 = ( n16258 & n16532 ) | ( n16258 & ~n16533 ) | ( n16532 & ~n16533 ) ;
  assign n16535 = n8016 ^ n1456 ^ 1'b0 ;
  assign n16536 = ~n3082 & n14690 ;
  assign n16537 = n11735 ^ n6731 ^ 1'b0 ;
  assign n16538 = n1402 | n16537 ;
  assign n16539 = n1487 | n16538 ;
  assign n16540 = n9525 & ~n16539 ;
  assign n16541 = n3632 | n9887 ;
  assign n16542 = n16541 ^ n898 ^ 1'b0 ;
  assign n16543 = n4072 & ~n16542 ;
  assign n16544 = n16543 ^ n2530 ^ 1'b0 ;
  assign n16545 = ~n673 & n6195 ;
  assign n16546 = n9381 ^ n7712 ^ n7041 ;
  assign n16547 = n5562 ^ n980 ^ 1'b0 ;
  assign n16548 = n3093 & ~n16547 ;
  assign n16549 = n16110 & n16548 ;
  assign n16550 = n1095 | n6272 ;
  assign n16551 = n3369 ^ n895 ^ 1'b0 ;
  assign n16552 = n16550 | n16551 ;
  assign n16553 = n14631 ^ n1991 ^ 1'b0 ;
  assign n16554 = ~n14624 & n16553 ;
  assign n16555 = n6258 & n16554 ;
  assign n16556 = n6570 ^ n2328 ^ 1'b0 ;
  assign n16557 = n3242 & n16556 ;
  assign n16558 = n1441 & n16557 ;
  assign n16559 = ~n14975 & n16558 ;
  assign n16560 = n1578 & ~n7139 ;
  assign n16561 = n6874 | n9769 ;
  assign n16562 = n3262 | n4011 ;
  assign n16563 = n701 | n16562 ;
  assign n16564 = x62 & n2606 ;
  assign n16565 = n2813 & n16564 ;
  assign n16566 = n13663 | n16565 ;
  assign n16567 = n16563 | n16566 ;
  assign n16568 = n2773 ^ n2127 ^ 1'b0 ;
  assign n16569 = n16568 ^ n7683 ^ 1'b0 ;
  assign n16570 = ~n15136 & n16569 ;
  assign n16571 = n16570 ^ n1329 ^ 1'b0 ;
  assign n16572 = n13807 ^ n4587 ^ 1'b0 ;
  assign n16573 = n7675 & ~n16572 ;
  assign n16574 = ~n1042 & n16573 ;
  assign n16575 = n16571 & n16574 ;
  assign n16576 = n7419 ^ n909 ^ 1'b0 ;
  assign n16577 = ~n3986 & n16576 ;
  assign n16578 = n8779 ^ n2153 ^ 1'b0 ;
  assign n16579 = n15824 ^ n1846 ^ 1'b0 ;
  assign n16580 = n12682 | n16579 ;
  assign n16581 = n12156 ^ n5530 ^ 1'b0 ;
  assign n16582 = n2763 & ~n3536 ;
  assign n16583 = n852 & ~n8203 ;
  assign n16584 = n16582 & ~n16583 ;
  assign n16585 = ~n1153 & n6911 ;
  assign n16586 = ~n735 & n16585 ;
  assign n16587 = n5796 & ~n10801 ;
  assign n16588 = n5144 ^ n788 ^ 1'b0 ;
  assign n16589 = n4502 | n16588 ;
  assign n16590 = n16587 & n16589 ;
  assign n16593 = n1924 & ~n6213 ;
  assign n16591 = n3688 & n8505 ;
  assign n16592 = ~n1158 & n16591 ;
  assign n16594 = n16593 ^ n16592 ^ 1'b0 ;
  assign n16595 = n6931 ^ n5810 ^ 1'b0 ;
  assign n16596 = n173 & ~n4321 ;
  assign n16597 = n16596 ^ n3474 ^ 1'b0 ;
  assign n16598 = n16597 ^ x2 ^ 1'b0 ;
  assign n16599 = n972 & n16598 ;
  assign n16600 = n8589 | n12315 ;
  assign n16601 = n2323 & ~n8515 ;
  assign n16602 = n6853 ^ n3837 ^ n2221 ;
  assign n16603 = n16602 ^ n1968 ^ n296 ;
  assign n16604 = n6871 | n16603 ;
  assign n16605 = ( n2245 & ~n9105 ) | ( n2245 & n9214 ) | ( ~n9105 & n9214 ) ;
  assign n16606 = n16605 ^ n2053 ^ 1'b0 ;
  assign n16607 = n2901 ^ n163 ^ 1'b0 ;
  assign n16608 = ~n4423 & n16607 ;
  assign n16609 = ~n851 & n3893 ;
  assign n16610 = n16609 ^ n13678 ^ n4107 ;
  assign n16611 = n4465 | n16610 ;
  assign n16612 = n5470 ^ n4303 ^ 1'b0 ;
  assign n16613 = ( ~n11323 & n13776 ) | ( ~n11323 & n16612 ) | ( n13776 & n16612 ) ;
  assign n16614 = n7092 & n11858 ;
  assign n16615 = n8185 & n16614 ;
  assign n16616 = n7141 ^ n3677 ^ 1'b0 ;
  assign n16617 = n2532 | n16616 ;
  assign n16618 = n8650 & ~n16617 ;
  assign n16619 = n9096 & n11706 ;
  assign n16620 = n1170 | n16619 ;
  assign n16621 = n558 & n1133 ;
  assign n16622 = ~n4011 & n16621 ;
  assign n16623 = n16622 ^ n8668 ^ 1'b0 ;
  assign n16624 = n1651 & ~n11160 ;
  assign n16625 = ( n6427 & ~n16623 ) | ( n6427 & n16624 ) | ( ~n16623 & n16624 ) ;
  assign n16626 = n7621 & ~n12847 ;
  assign n16627 = n16602 ^ n7134 ^ 1'b0 ;
  assign n16628 = n2525 | n16627 ;
  assign n16629 = n8215 & ~n16628 ;
  assign n16630 = n1947 & n3295 ;
  assign n16631 = n12053 & n16630 ;
  assign n16632 = ~n6212 & n16631 ;
  assign n16633 = n934 & n8961 ;
  assign n16634 = ( ~n4564 & n7186 ) | ( ~n4564 & n16633 ) | ( n7186 & n16633 ) ;
  assign n16635 = ~n1843 & n3413 ;
  assign n16636 = n7433 & n16635 ;
  assign n16637 = n5713 & ~n9803 ;
  assign n16638 = n16637 ^ n5074 ^ 1'b0 ;
  assign n16639 = n4619 | n11773 ;
  assign n16640 = x12 | n9964 ;
  assign n16641 = n13841 ^ n13372 ^ 1'b0 ;
  assign n16642 = n11315 ^ n5625 ^ 1'b0 ;
  assign n16643 = n1046 & ~n3618 ;
  assign n16644 = ( n2579 & n3420 ) | ( n2579 & ~n6428 ) | ( n3420 & ~n6428 ) ;
  assign n16645 = ~n16643 & n16644 ;
  assign n16646 = n16645 ^ n5203 ^ 1'b0 ;
  assign n16647 = n6505 & n8247 ;
  assign n16648 = n1018 & n16647 ;
  assign n16649 = n627 ^ n606 ^ 1'b0 ;
  assign n16650 = n10322 ^ n3672 ^ 1'b0 ;
  assign n16651 = n16650 ^ n10232 ^ 1'b0 ;
  assign n16652 = n12556 ^ n1077 ^ 1'b0 ;
  assign n16653 = n11997 ^ n11137 ^ 1'b0 ;
  assign n16654 = n992 & n3114 ;
  assign n16655 = n9246 & ~n16654 ;
  assign n16656 = n12458 | n13065 ;
  assign n16662 = n6428 ^ n2947 ^ 1'b0 ;
  assign n16657 = n1293 | n3003 ;
  assign n16658 = n16657 ^ n4474 ^ 1'b0 ;
  assign n16659 = n16658 ^ n13053 ^ 1'b0 ;
  assign n16660 = n5168 & n16659 ;
  assign n16661 = n1685 & n16660 ;
  assign n16663 = n16662 ^ n16661 ^ 1'b0 ;
  assign n16664 = n16663 ^ n7683 ^ n4623 ;
  assign n16666 = n8193 & n12526 ;
  assign n16665 = n7270 | n12045 ;
  assign n16667 = n16666 ^ n16665 ^ 1'b0 ;
  assign n16668 = n8159 ^ n1226 ^ 1'b0 ;
  assign n16669 = n3876 & ~n16668 ;
  assign n16670 = ( n1837 & n1954 ) | ( n1837 & n16669 ) | ( n1954 & n16669 ) ;
  assign n16671 = ~n2839 & n16670 ;
  assign n16672 = n4861 ^ n662 ^ 1'b0 ;
  assign n16673 = ~n1930 & n16672 ;
  assign n16674 = n16673 ^ n1167 ^ 1'b0 ;
  assign n16675 = ~n1035 & n2882 ;
  assign n16676 = n8260 ^ n5293 ^ 1'b0 ;
  assign n16677 = ~n16675 & n16676 ;
  assign n16678 = n7608 ^ n5028 ^ 1'b0 ;
  assign n16679 = n7040 & n16678 ;
  assign n16680 = n2354 & n3237 ;
  assign n16681 = n16680 ^ n8194 ^ 1'b0 ;
  assign n16682 = n3494 & n4817 ;
  assign n16683 = n7918 & n16682 ;
  assign n16684 = n3434 ^ n916 ^ 1'b0 ;
  assign n16685 = n2833 | n7986 ;
  assign n16686 = ~n5871 & n15706 ;
  assign n16687 = n6456 ^ n3328 ^ 1'b0 ;
  assign n16688 = n2554 & ~n3132 ;
  assign n16689 = n16688 ^ n15119 ^ 1'b0 ;
  assign n16690 = ~n5940 & n16689 ;
  assign n16691 = n8831 ^ n7845 ^ 1'b0 ;
  assign n16692 = n5806 | n16691 ;
  assign n16693 = n7631 | n12785 ;
  assign n16694 = n8921 ^ x59 ^ 1'b0 ;
  assign n16700 = n13701 ^ n12267 ^ 1'b0 ;
  assign n16701 = n4817 & n16700 ;
  assign n16696 = n5156 ^ n4497 ^ 1'b0 ;
  assign n16697 = n1590 & n16696 ;
  assign n16695 = x85 & ~n6698 ;
  assign n16698 = n16697 ^ n16695 ^ 1'b0 ;
  assign n16699 = n4153 & ~n16698 ;
  assign n16702 = n16701 ^ n16699 ^ 1'b0 ;
  assign n16703 = n5491 & ~n16702 ;
  assign n16704 = n14908 & n16703 ;
  assign n16705 = n6091 & n11437 ;
  assign n16706 = n450 & n4576 ;
  assign n16707 = n16706 ^ n4112 ^ 1'b0 ;
  assign n16708 = n13370 & n16707 ;
  assign n16709 = n16708 ^ n3354 ^ 1'b0 ;
  assign n16710 = ~n1634 & n1713 ;
  assign n16711 = n6310 ^ n409 ^ 1'b0 ;
  assign n16712 = n13496 & ~n16711 ;
  assign n16713 = n9713 ^ n2650 ^ 1'b0 ;
  assign n16714 = n4032 ^ x16 ^ 1'b0 ;
  assign n16715 = ~n3905 & n16714 ;
  assign n16716 = n1918 | n7075 ;
  assign n16717 = n11141 ^ n9433 ^ 1'b0 ;
  assign n16718 = n1872 | n16717 ;
  assign n16719 = n6242 ^ n5586 ^ 1'b0 ;
  assign n16720 = ~n684 & n16719 ;
  assign n16721 = ~n1361 & n4532 ;
  assign n16722 = n16721 ^ n3898 ^ 1'b0 ;
  assign n16723 = n4567 & n9676 ;
  assign n16724 = n2917 | n4743 ;
  assign n16725 = n4105 & ~n16724 ;
  assign n16726 = n16725 ^ n4011 ^ 1'b0 ;
  assign n16727 = n7158 ^ n268 ^ 1'b0 ;
  assign n16728 = n3640 | n16727 ;
  assign n16729 = n4747 & ~n6017 ;
  assign n16730 = n12298 & ~n13104 ;
  assign n16731 = ~n13434 & n16730 ;
  assign n16732 = n16731 ^ n16099 ^ 1'b0 ;
  assign n16733 = n3642 & n13363 ;
  assign n16734 = n5186 ^ n882 ^ 1'b0 ;
  assign n16735 = n6199 | n16734 ;
  assign n16736 = n2020 | n16735 ;
  assign n16737 = n11380 & n16736 ;
  assign n16738 = n16737 ^ n3532 ^ 1'b0 ;
  assign n16739 = n2951 | n5485 ;
  assign n16740 = x110 & ~n1402 ;
  assign n16741 = ~n1718 & n16740 ;
  assign n16742 = n16741 ^ n3230 ^ 1'b0 ;
  assign n16743 = n8058 | n16742 ;
  assign n16744 = n10470 ^ n2919 ^ 1'b0 ;
  assign n16745 = n8314 & n16744 ;
  assign n16746 = n1602 & ~n11411 ;
  assign n16747 = n16746 ^ n11767 ^ 1'b0 ;
  assign n16748 = n11081 & n16747 ;
  assign n16749 = n8683 & ~n16748 ;
  assign n16751 = n4406 ^ n4029 ^ n3635 ;
  assign n16752 = n5789 | n16751 ;
  assign n16750 = ~n868 & n1788 ;
  assign n16753 = n16752 ^ n16750 ^ 1'b0 ;
  assign n16754 = n3195 | n8633 ;
  assign n16755 = n2166 | n7469 ;
  assign n16756 = n16538 & ~n16755 ;
  assign n16757 = n9062 ^ n339 ^ 1'b0 ;
  assign n16758 = n15807 | n16757 ;
  assign n16759 = n7635 | n12523 ;
  assign n16760 = n16759 ^ n9676 ^ 1'b0 ;
  assign n16761 = n6780 | n16760 ;
  assign n16762 = n7963 ^ n5898 ^ 1'b0 ;
  assign n16763 = n4636 & ~n14041 ;
  assign n16764 = n16669 ^ n5367 ^ 1'b0 ;
  assign n16765 = ~n3700 & n8499 ;
  assign n16766 = n11187 | n13781 ;
  assign n16767 = n3620 ^ n2037 ^ 1'b0 ;
  assign n16768 = n5453 | n16767 ;
  assign n16769 = n2271 | n16768 ;
  assign n16770 = n10573 & n13528 ;
  assign n16771 = n3158 | n3400 ;
  assign n16772 = n16771 ^ n2718 ^ 1'b0 ;
  assign n16773 = n16772 ^ n4855 ^ 1'b0 ;
  assign n16774 = n9797 ^ n4412 ^ 1'b0 ;
  assign n16775 = n2256 & ~n14127 ;
  assign n16776 = n830 & n981 ;
  assign n16777 = ~x39 & n16776 ;
  assign n16778 = n1177 & ~n4372 ;
  assign n16779 = n16778 ^ n6677 ^ n1477 ;
  assign n16780 = n2873 & n16779 ;
  assign n16781 = n16777 & n16780 ;
  assign n16782 = n926 & n12186 ;
  assign n16783 = n10858 & n16782 ;
  assign n16784 = n16783 ^ n12276 ^ 1'b0 ;
  assign n16785 = n16781 | n16784 ;
  assign n16786 = n5753 & n6203 ;
  assign n16787 = n2493 | n14006 ;
  assign n16788 = n4440 | n16663 ;
  assign n16789 = ~n839 & n2614 ;
  assign n16790 = n9047 & n16789 ;
  assign n16791 = n6823 & n16536 ;
  assign n16793 = n8137 ^ n1087 ^ 1'b0 ;
  assign n16792 = n645 ^ n526 ^ n296 ;
  assign n16794 = n16793 ^ n16792 ^ 1'b0 ;
  assign n16795 = n6259 & n6398 ;
  assign n16796 = n2792 & ~n4096 ;
  assign n16797 = ~n2808 & n16796 ;
  assign n16798 = n6716 & ~n16797 ;
  assign n16799 = n6438 ^ n2499 ^ 1'b0 ;
  assign n16800 = n921 & n2315 ;
  assign n16801 = n165 & n7096 ;
  assign n16802 = n16801 ^ n7096 ^ 1'b0 ;
  assign n16805 = n8146 & n11081 ;
  assign n16806 = n4056 & n16805 ;
  assign n16803 = ~n9095 & n10320 ;
  assign n16804 = ~n9501 & n16803 ;
  assign n16807 = n16806 ^ n16804 ^ 1'b0 ;
  assign n16808 = n6389 ^ n825 ^ 1'b0 ;
  assign n16809 = n1867 | n16808 ;
  assign n16810 = n7236 ^ n1880 ^ 1'b0 ;
  assign n16811 = n16810 ^ n4636 ^ 1'b0 ;
  assign n16812 = n7894 ^ n594 ^ 1'b0 ;
  assign n16813 = n14941 & ~n16812 ;
  assign n16814 = n8538 | n13252 ;
  assign n16815 = n16685 ^ n1899 ^ 1'b0 ;
  assign n16816 = ~x56 & n10207 ;
  assign n16817 = ~x95 & n16816 ;
  assign n16818 = n6907 ^ n412 ^ 1'b0 ;
  assign n16819 = ~n16817 & n16818 ;
  assign n16820 = n1157 & n3046 ;
  assign n16821 = n16820 ^ n2955 ^ 1'b0 ;
  assign n16822 = n1685 & ~n16821 ;
  assign n16823 = ( n2041 & ~n7433 ) | ( n2041 & n12923 ) | ( ~n7433 & n12923 ) ;
  assign n16824 = n16823 ^ n11587 ^ 1'b0 ;
  assign n16826 = ~n7548 & n15258 ;
  assign n16825 = ~n6186 & n10669 ;
  assign n16827 = n16826 ^ n16825 ^ 1'b0 ;
  assign n16828 = n6655 ^ n4991 ^ n801 ;
  assign n16829 = n16062 ^ n786 ^ 1'b0 ;
  assign n16830 = n16828 & n16829 ;
  assign n16831 = n7393 & ~n7991 ;
  assign n16832 = ( n1523 & n10840 ) | ( n1523 & n16831 ) | ( n10840 & n16831 ) ;
  assign n16833 = n10843 & n12560 ;
  assign n16834 = n16833 ^ n6716 ^ 1'b0 ;
  assign n16835 = n5200 ^ n4939 ^ 1'b0 ;
  assign n16836 = n12888 ^ n12857 ^ 1'b0 ;
  assign n16837 = n655 & n7784 ;
  assign n16838 = n7544 & n16837 ;
  assign n16839 = ~n11842 & n13833 ;
  assign n16840 = n16839 ^ n14194 ^ 1'b0 ;
  assign n16841 = n1501 | n5191 ;
  assign n16842 = n16841 ^ n4321 ^ 1'b0 ;
  assign n16843 = n16842 ^ n11516 ^ 1'b0 ;
  assign n16844 = ~n2200 & n16843 ;
  assign n16847 = n5876 ^ n4816 ^ n4280 ;
  assign n16848 = n5273 & n16847 ;
  assign n16845 = ( n339 & n696 ) | ( n339 & ~n8888 ) | ( n696 & ~n8888 ) ;
  assign n16846 = n10675 & ~n16845 ;
  assign n16849 = n16848 ^ n16846 ^ 1'b0 ;
  assign n16850 = n7339 ^ n782 ^ 1'b0 ;
  assign n16851 = ~n12702 & n16850 ;
  assign n16852 = n8958 & ~n16851 ;
  assign n16854 = n6714 ^ n1156 ^ 1'b0 ;
  assign n16855 = ~n12065 & n16854 ;
  assign n16853 = n6268 & n13634 ;
  assign n16856 = n16855 ^ n16853 ^ 1'b0 ;
  assign n16857 = n13333 ^ n13165 ^ 1'b0 ;
  assign n16858 = n16856 | n16857 ;
  assign n16859 = n9286 ^ n7690 ^ 1'b0 ;
  assign n16860 = n2893 & ~n4413 ;
  assign n16861 = n16860 ^ n846 ^ 1'b0 ;
  assign n16862 = n3275 & n9328 ;
  assign n16863 = n14211 & ~n16675 ;
  assign n16864 = ~n16862 & n16863 ;
  assign n16865 = n14623 ^ n12692 ^ 1'b0 ;
  assign n16866 = ( n481 & ~n2854 ) | ( n481 & n5365 ) | ( ~n2854 & n5365 ) ;
  assign n16867 = ~n430 & n16866 ;
  assign n16868 = n1644 | n10400 ;
  assign n16869 = n10415 | n16868 ;
  assign n16870 = n16869 ^ n11022 ^ 1'b0 ;
  assign n16871 = n5477 | n12196 ;
  assign n16872 = n2971 & n16871 ;
  assign n16873 = n9115 | n9954 ;
  assign n16878 = n9859 ^ n8016 ^ 1'b0 ;
  assign n16874 = ~n4635 & n5938 ;
  assign n16875 = n16874 ^ n12062 ^ 1'b0 ;
  assign n16876 = ~n2402 & n16875 ;
  assign n16877 = n4137 | n16876 ;
  assign n16879 = n16878 ^ n16877 ^ 1'b0 ;
  assign n16880 = n1419 | n11714 ;
  assign n16881 = n16880 ^ n1044 ^ 1'b0 ;
  assign n16882 = n12172 ^ n1966 ^ 1'b0 ;
  assign n16883 = n12452 & n16882 ;
  assign n16884 = n15074 & n16883 ;
  assign n16885 = ~n5874 & n16884 ;
  assign n16886 = n6598 ^ n288 ^ 1'b0 ;
  assign n16887 = n13434 ^ n5038 ^ 1'b0 ;
  assign n16888 = n6699 | n10641 ;
  assign n16889 = n8758 & ~n16888 ;
  assign n16890 = ( n555 & n2351 ) | ( n555 & n4280 ) | ( n2351 & n4280 ) ;
  assign n16891 = n3615 | n4079 ;
  assign n16892 = ~n3466 & n16891 ;
  assign n16893 = n14926 ^ n5022 ^ 1'b0 ;
  assign n16894 = n1792 & ~n4661 ;
  assign n16895 = n16894 ^ n5527 ^ 1'b0 ;
  assign n16896 = n7926 ^ x77 ^ 1'b0 ;
  assign n16897 = x60 & n3086 ;
  assign n16898 = ~n11850 & n16897 ;
  assign n16899 = n15843 ^ n14221 ^ n11479 ;
  assign n16900 = ~n4247 & n14955 ;
  assign n16901 = ~n8841 & n16900 ;
  assign n16902 = n16901 ^ n7283 ^ 1'b0 ;
  assign n16903 = n9618 ^ n1008 ^ 1'b0 ;
  assign n16904 = ~n6017 & n16903 ;
  assign n16905 = n6325 & n16904 ;
  assign n16906 = n1958 & n16905 ;
  assign n16907 = n16906 ^ n4195 ^ 1'b0 ;
  assign n16908 = ~n12522 & n16288 ;
  assign n16909 = n12809 ^ n10017 ^ 1'b0 ;
  assign n16910 = x102 & n4344 ;
  assign n16911 = n3666 | n9858 ;
  assign n16912 = n2087 ^ n702 ^ 1'b0 ;
  assign n16913 = n16912 ^ n4212 ^ 1'b0 ;
  assign n16914 = ~n444 & n14674 ;
  assign n16915 = ~n16913 & n16914 ;
  assign n16916 = n16081 ^ n2615 ^ 1'b0 ;
  assign n16917 = n16915 | n16916 ;
  assign n16918 = n6594 & ~n16917 ;
  assign n16919 = n7639 & ~n9254 ;
  assign n16920 = ~n8749 & n14626 ;
  assign n16921 = n16920 ^ n13273 ^ 1'b0 ;
  assign n16922 = n1695 & n10588 ;
  assign n16923 = n5609 | n11316 ;
  assign n16924 = n2176 & ~n16923 ;
  assign n16925 = n2947 ^ n1203 ^ 1'b0 ;
  assign n16926 = n16924 | n16925 ;
  assign n16927 = n6357 | n16926 ;
  assign n16928 = n6230 | n16927 ;
  assign n16929 = n1644 | n10967 ;
  assign n16930 = n1430 & n1436 ;
  assign n16931 = n16930 ^ n7171 ^ 1'b0 ;
  assign n16932 = n702 & n16931 ;
  assign n16933 = ~n2469 & n16932 ;
  assign n16934 = n16933 ^ n8352 ^ 1'b0 ;
  assign n16935 = n3683 | n16934 ;
  assign n16936 = n1482 & ~n16935 ;
  assign n16937 = n296 | n6964 ;
  assign n16938 = n16937 ^ n433 ^ 1'b0 ;
  assign n16939 = n15697 ^ n8823 ^ 1'b0 ;
  assign n16940 = n8857 & ~n10677 ;
  assign n16941 = n16940 ^ n701 ^ 1'b0 ;
  assign n16942 = n1892 & n13324 ;
  assign n16943 = x23 & ~n1325 ;
  assign n16945 = n2887 | n5048 ;
  assign n16946 = n6977 | n16945 ;
  assign n16944 = n6115 ^ n4529 ^ 1'b0 ;
  assign n16947 = n16946 ^ n16944 ^ 1'b0 ;
  assign n16948 = n13530 | n16947 ;
  assign n16949 = n13864 | n14745 ;
  assign n16950 = n16949 ^ n6710 ^ 1'b0 ;
  assign n16951 = n10662 ^ n6893 ^ 1'b0 ;
  assign n16952 = n10551 | n16951 ;
  assign n16953 = n14602 ^ n6208 ^ 1'b0 ;
  assign n16954 = n6026 & n16185 ;
  assign n16955 = ~n2660 & n11518 ;
  assign n16956 = n8506 & n16955 ;
  assign n16957 = ~n2559 & n7236 ;
  assign n16958 = ~n2369 & n5027 ;
  assign n16959 = n7335 & n16958 ;
  assign n16960 = n2792 & n3309 ;
  assign n16961 = n16959 & n16960 ;
  assign n16962 = n5891 ^ n998 ^ 1'b0 ;
  assign n16963 = n6606 | n16962 ;
  assign n16964 = n4488 & ~n16963 ;
  assign n16965 = ( n1416 & n1830 ) | ( n1416 & ~n15394 ) | ( n1830 & ~n15394 ) ;
  assign n16966 = ~n14728 & n16965 ;
  assign n16967 = ~n1093 & n16966 ;
  assign n16968 = n3050 & n4077 ;
  assign n16969 = n16968 ^ n12580 ^ 1'b0 ;
  assign n16970 = n9526 & n14633 ;
  assign n16971 = n8435 & n15630 ;
  assign n16972 = n16971 ^ n16048 ^ 1'b0 ;
  assign n16973 = n9628 & ~n16080 ;
  assign n16974 = n3596 & n16973 ;
  assign n16975 = n1890 & ~n2186 ;
  assign n16976 = n16975 ^ n13364 ^ 1'b0 ;
  assign n16980 = n3597 ^ n2331 ^ 1'b0 ;
  assign n16977 = n3651 & n9524 ;
  assign n16978 = n16977 ^ n1972 ^ 1'b0 ;
  assign n16979 = n3952 | n16978 ;
  assign n16981 = n16980 ^ n16979 ^ 1'b0 ;
  assign n16982 = n1963 ^ n638 ^ 1'b0 ;
  assign n16983 = n15132 & ~n16982 ;
  assign n16984 = n11118 | n16983 ;
  assign n16985 = n131 & ~n1895 ;
  assign n16986 = n16985 ^ n6195 ^ 1'b0 ;
  assign n16987 = n1173 | n16986 ;
  assign n16988 = n15086 ^ n13767 ^ 1'b0 ;
  assign n16989 = n16987 & ~n16988 ;
  assign n16990 = n4621 | n6526 ;
  assign n16991 = n8693 | n16990 ;
  assign n16992 = ( n1470 & n8253 ) | ( n1470 & n16991 ) | ( n8253 & n16991 ) ;
  assign n16993 = n14994 ^ n9174 ^ 1'b0 ;
  assign n16994 = n16992 & ~n16993 ;
  assign n16995 = ~n2730 & n5405 ;
  assign n16996 = ~n3255 & n16995 ;
  assign n16997 = n15854 & ~n16996 ;
  assign n16998 = n16997 ^ n4029 ^ 1'b0 ;
  assign n16999 = n16994 & ~n16998 ;
  assign n17000 = n1178 | n1796 ;
  assign n17001 = n2864 | n6335 ;
  assign n17002 = n17001 ^ n1800 ^ 1'b0 ;
  assign n17003 = x16 & ~n868 ;
  assign n17004 = n3201 & n17003 ;
  assign n17005 = ( n16440 & ~n17002 ) | ( n16440 & n17004 ) | ( ~n17002 & n17004 ) ;
  assign n17006 = ~n8749 & n12196 ;
  assign n17007 = ~n5632 & n17006 ;
  assign n17008 = n10085 ^ n4366 ^ 1'b0 ;
  assign n17009 = ~n1945 & n17008 ;
  assign n17010 = n17009 ^ n2767 ^ 1'b0 ;
  assign n17011 = n10686 | n17010 ;
  assign n17012 = n8205 ^ n6731 ^ 1'b0 ;
  assign n17013 = ~n4384 & n6401 ;
  assign n17014 = n17013 ^ n16266 ^ n3833 ;
  assign n17017 = n7244 & ~n9954 ;
  assign n17018 = n17017 ^ n950 ^ 1'b0 ;
  assign n17015 = n613 & n14279 ;
  assign n17016 = n4729 & n17015 ;
  assign n17019 = n17018 ^ n17016 ^ 1'b0 ;
  assign n17020 = n17014 & ~n17019 ;
  assign n17021 = ~n7292 & n9227 ;
  assign n17022 = n17021 ^ n14440 ^ 1'b0 ;
  assign n17025 = n7732 | n8080 ;
  assign n17023 = x22 & ~n6406 ;
  assign n17024 = n17023 ^ n6789 ^ 1'b0 ;
  assign n17026 = n17025 ^ n17024 ^ 1'b0 ;
  assign n17027 = n6562 ^ n1997 ^ 1'b0 ;
  assign n17028 = n7678 | n17027 ;
  assign n17029 = n5129 & ~n17028 ;
  assign n17030 = n5383 & n9734 ;
  assign n17031 = n5984 | n6537 ;
  assign n17032 = n2854 & ~n10896 ;
  assign n17033 = ~x42 & n17032 ;
  assign n17034 = ( n3401 & ~n17031 ) | ( n3401 & n17033 ) | ( ~n17031 & n17033 ) ;
  assign n17036 = n3512 & n6942 ;
  assign n17037 = n1558 & n17036 ;
  assign n17035 = n2621 & ~n5159 ;
  assign n17038 = n17037 ^ n17035 ^ 1'b0 ;
  assign n17045 = ~n632 & n3443 ;
  assign n17041 = n5381 & ~n5603 ;
  assign n17042 = n17041 ^ n4303 ^ 1'b0 ;
  assign n17039 = n9289 ^ n2446 ^ 1'b0 ;
  assign n17040 = n701 & n17039 ;
  assign n17043 = n17042 ^ n17040 ^ 1'b0 ;
  assign n17044 = n10588 | n17043 ;
  assign n17046 = n17045 ^ n17044 ^ 1'b0 ;
  assign n17047 = ( ~x3 & n7060 ) | ( ~x3 & n9454 ) | ( n7060 & n9454 ) ;
  assign n17048 = n14026 & n17047 ;
  assign n17049 = n6028 & n17048 ;
  assign n17050 = n11238 ^ n5364 ^ 1'b0 ;
  assign n17051 = n17050 ^ n12661 ^ 1'b0 ;
  assign n17054 = ~n5555 & n7673 ;
  assign n17055 = ~n13633 & n17054 ;
  assign n17052 = ~n1406 & n13418 ;
  assign n17053 = ~n190 & n17052 ;
  assign n17056 = n17055 ^ n17053 ^ n10987 ;
  assign n17057 = n15225 ^ n13169 ^ n3482 ;
  assign n17058 = n5652 ^ n250 ^ 1'b0 ;
  assign n17059 = n15314 & n17058 ;
  assign n17060 = n8296 ^ n6428 ^ 1'b0 ;
  assign n17061 = n6760 | n17060 ;
  assign n17062 = ~n2885 & n5876 ;
  assign n17063 = n614 | n3302 ;
  assign n17064 = n17063 ^ n6522 ^ 1'b0 ;
  assign n17065 = ~n3991 & n15405 ;
  assign n17066 = n17065 ^ n2769 ^ 1'b0 ;
  assign n17067 = n8030 & n17066 ;
  assign n17068 = n11468 ^ n5243 ^ 1'b0 ;
  assign n17069 = ~n8101 & n17068 ;
  assign n17070 = n17069 ^ n920 ^ 1'b0 ;
  assign n17071 = n6690 | n7735 ;
  assign n17072 = ~n6868 & n15476 ;
  assign n17073 = n784 | n9525 ;
  assign n17074 = n17073 ^ n5291 ^ 1'b0 ;
  assign n17075 = n5381 | n17074 ;
  assign n17076 = n6853 ^ n2896 ^ 1'b0 ;
  assign n17077 = ~x86 & n17076 ;
  assign n17078 = n5283 & ~n17077 ;
  assign n17079 = n17078 ^ n12541 ^ 1'b0 ;
  assign n17080 = n808 & n17079 ;
  assign n17081 = n17080 ^ n10037 ^ 1'b0 ;
  assign n17082 = n3030 & ~n15728 ;
  assign n17083 = n7722 ^ n456 ^ 1'b0 ;
  assign n17084 = n3038 & n17083 ;
  assign n17085 = ~n2159 & n17084 ;
  assign n17086 = n17085 ^ n825 ^ 1'b0 ;
  assign n17090 = n12569 ^ n6824 ^ 1'b0 ;
  assign n17087 = n1629 & n11157 ;
  assign n17088 = n4334 & n17087 ;
  assign n17089 = ~n5238 & n17088 ;
  assign n17091 = n17090 ^ n17089 ^ n7383 ;
  assign n17092 = n3950 ^ n2848 ^ 1'b0 ;
  assign n17093 = x75 | n17092 ;
  assign n17094 = n15609 ^ n8190 ^ 1'b0 ;
  assign n17096 = n3069 & n15181 ;
  assign n17097 = n17096 ^ n6886 ^ 1'b0 ;
  assign n17095 = ~n1079 & n7506 ;
  assign n17098 = n17097 ^ n17095 ^ 1'b0 ;
  assign n17099 = n6027 & n13421 ;
  assign n17100 = n2843 & n17099 ;
  assign n17101 = n7361 & ~n11004 ;
  assign n17102 = n17101 ^ n12347 ^ 1'b0 ;
  assign n17103 = ~n3350 & n6126 ;
  assign n17104 = n867 | n15193 ;
  assign n17105 = ~n800 & n13132 ;
  assign n17106 = n17105 ^ n10264 ^ 1'b0 ;
  assign n17107 = n17106 ^ n5708 ^ 1'b0 ;
  assign n17108 = n7700 | n17107 ;
  assign n17109 = n11482 & n14674 ;
  assign n17110 = n2490 | n10147 ;
  assign n17111 = n17110 ^ n294 ^ 1'b0 ;
  assign n17112 = n391 | n8259 ;
  assign n17113 = n17112 ^ n6883 ^ 1'b0 ;
  assign n17114 = n2744 | n10170 ;
  assign n17115 = n10557 ^ n10077 ^ n3500 ;
  assign n17116 = ~n8940 & n17115 ;
  assign n17117 = n1632 & n6394 ;
  assign n17118 = n4648 | n7362 ;
  assign n17119 = n12149 & n17118 ;
  assign n17120 = ~n14623 & n17119 ;
  assign n17121 = n8294 | n17120 ;
  assign n17122 = n4224 & n16713 ;
  assign n17123 = ~n17121 & n17122 ;
  assign n17124 = n4933 | n10234 ;
  assign n17125 = n17124 ^ n8958 ^ 1'b0 ;
  assign n17126 = n17125 ^ x50 ^ 1'b0 ;
  assign n17127 = n17126 ^ n7666 ^ 1'b0 ;
  assign n17128 = n17123 | n17127 ;
  assign n17129 = ~n346 & n1548 ;
  assign n17130 = n3764 | n6789 ;
  assign n17131 = n5197 & ~n17130 ;
  assign n17132 = n17131 ^ n484 ^ 1'b0 ;
  assign n17133 = n12763 | n17132 ;
  assign n17134 = n14288 ^ x11 ^ 1'b0 ;
  assign n17135 = n17134 ^ n13742 ^ 1'b0 ;
  assign n17136 = n1753 ^ n660 ^ 1'b0 ;
  assign n17137 = n13548 & n17136 ;
  assign n17138 = n17137 ^ n9295 ^ x49 ;
  assign n17139 = n2539 & n7626 ;
  assign n17140 = ~n847 & n5202 ;
  assign n17141 = n17140 ^ n4438 ^ 1'b0 ;
  assign n17142 = ~n894 & n17141 ;
  assign n17143 = n17142 ^ n5603 ^ 1'b0 ;
  assign n17144 = ~n4858 & n17143 ;
  assign n17145 = ~n17139 & n17144 ;
  assign n17146 = n12504 & ~n12522 ;
  assign n17147 = n17146 ^ n4288 ^ 1'b0 ;
  assign n17148 = n10489 ^ n6044 ^ 1'b0 ;
  assign n17149 = n14118 & ~n17148 ;
  assign n17150 = n14073 ^ n2409 ^ 1'b0 ;
  assign n17151 = ~n2596 & n17150 ;
  assign n17152 = ~n5259 & n17151 ;
  assign n17153 = ~n10280 & n17152 ;
  assign n17154 = n11375 & ~n17153 ;
  assign n17155 = n4478 | n16672 ;
  assign n17156 = n3031 | n5630 ;
  assign n17157 = n5466 | n17156 ;
  assign n17158 = n782 ^ n613 ^ 1'b0 ;
  assign n17159 = ~n4985 & n7997 ;
  assign n17160 = n17159 ^ n694 ^ 1'b0 ;
  assign n17161 = n1601 & ~n16890 ;
  assign n17162 = n17160 | n17161 ;
  assign n17163 = x16 & n2921 ;
  assign n17164 = ~n13792 & n17163 ;
  assign n17190 = ~n1651 & n4025 ;
  assign n17191 = ~n4025 & n17190 ;
  assign n17192 = n3422 & ~n17191 ;
  assign n17165 = n177 & ~n1341 ;
  assign n17166 = ~n177 & n17165 ;
  assign n17167 = x73 & n152 ;
  assign n17168 = ~n152 & n17167 ;
  assign n17169 = n188 & n17168 ;
  assign n17170 = n161 & ~n238 ;
  assign n17171 = n17169 & n17170 ;
  assign n17172 = x78 & n320 ;
  assign n17173 = ~x78 & n17172 ;
  assign n17174 = n625 | n17173 ;
  assign n17175 = n17173 & ~n17174 ;
  assign n17176 = n480 | n17175 ;
  assign n17177 = n17175 & ~n17176 ;
  assign n17178 = n1146 & ~n17177 ;
  assign n17179 = ~n1146 & n17178 ;
  assign n17180 = n373 | n539 ;
  assign n17181 = n539 & ~n17180 ;
  assign n17182 = n496 | n17181 ;
  assign n17183 = n17181 & ~n17182 ;
  assign n17184 = n17183 ^ n2385 ^ 1'b0 ;
  assign n17185 = n17179 | n17184 ;
  assign n17186 = n17179 & ~n17185 ;
  assign n17187 = n17186 ^ n4802 ^ 1'b0 ;
  assign n17188 = n17171 | n17187 ;
  assign n17189 = n17166 | n17188 ;
  assign n17193 = n17192 ^ n17189 ^ 1'b0 ;
  assign n17194 = n3579 | n17193 ;
  assign n17195 = n2292 | n17194 ;
  assign n17196 = n9139 & n17195 ;
  assign n17197 = ~n2942 & n17196 ;
  assign n17198 = n4287 & ~n16351 ;
  assign n17199 = ~x3 & n17198 ;
  assign n17200 = n5213 | n8673 ;
  assign n17201 = n14399 & n17200 ;
  assign n17202 = n595 & ~n6115 ;
  assign n17203 = n2511 | n17202 ;
  assign n17204 = n9901 | n14769 ;
  assign n17205 = n7017 | n12260 ;
  assign n17206 = n4478 & ~n17205 ;
  assign n17207 = n8918 & ~n9602 ;
  assign n17208 = n17207 ^ n11939 ^ 1'b0 ;
  assign n17209 = n9381 ^ n4307 ^ 1'b0 ;
  assign n17210 = n13560 ^ x71 ^ 1'b0 ;
  assign n17211 = n811 & ~n17210 ;
  assign n17212 = n10568 & n16978 ;
  assign n17213 = n17212 ^ n11467 ^ 1'b0 ;
  assign n17214 = n14871 & ~n17213 ;
  assign n17215 = n5764 & n12576 ;
  assign n17216 = n17215 ^ n967 ^ 1'b0 ;
  assign n17217 = n1080 ^ n942 ^ 1'b0 ;
  assign n17218 = n11599 ^ n10633 ^ 1'b0 ;
  assign n17219 = ~n4411 & n4854 ;
  assign n17220 = n17219 ^ n2842 ^ 1'b0 ;
  assign n17221 = x103 & n2555 ;
  assign n17222 = n16109 ^ n15474 ^ x12 ;
  assign n17223 = n17222 ^ n14920 ^ 1'b0 ;
  assign n17224 = n13935 & n16643 ;
  assign n17225 = ( n6156 & n11281 ) | ( n6156 & ~n11870 ) | ( n11281 & ~n11870 ) ;
  assign n17226 = n4693 & ~n17225 ;
  assign n17227 = n8722 & n17226 ;
  assign n17228 = ( x15 & n6181 ) | ( x15 & ~n11597 ) | ( n6181 & ~n11597 ) ;
  assign n17229 = n633 ^ n632 ^ n427 ;
  assign n17230 = n9391 | n17229 ;
  assign n17231 = n17230 ^ n4025 ^ 1'b0 ;
  assign n17232 = n1874 & n6026 ;
  assign n17233 = ~n17231 & n17232 ;
  assign n17234 = n5467 | n10992 ;
  assign n17235 = n9856 ^ n831 ^ 1'b0 ;
  assign n17236 = n876 & n15682 ;
  assign n17237 = ~n857 & n9910 ;
  assign n17238 = n992 | n17237 ;
  assign n17239 = n17238 ^ n2719 ^ 1'b0 ;
  assign n17240 = n17239 ^ n9081 ^ n4091 ;
  assign n17241 = n5103 | n10822 ;
  assign n17242 = n11006 | n17241 ;
  assign n17243 = n10619 ^ n380 ^ 1'b0 ;
  assign n17244 = ( ~n5099 & n6561 ) | ( ~n5099 & n10393 ) | ( n6561 & n10393 ) ;
  assign n17245 = n5904 & n11006 ;
  assign n17246 = ~n7865 & n17245 ;
  assign n17247 = n17246 ^ n5181 ^ 1'b0 ;
  assign n17248 = ~n4359 & n11901 ;
  assign n17249 = n1430 & n7443 ;
  assign n17250 = n17249 ^ n8137 ^ 1'b0 ;
  assign n17251 = n7247 & ~n13987 ;
  assign n17252 = ~n17250 & n17251 ;
  assign n17254 = n7066 ^ n4318 ^ 1'b0 ;
  assign n17255 = n11220 & ~n17254 ;
  assign n17253 = n6887 & ~n14382 ;
  assign n17256 = n17255 ^ n17253 ^ 1'b0 ;
  assign n17257 = n11409 ^ n9611 ^ 1'b0 ;
  assign n17258 = n10152 & n10823 ;
  assign n17259 = n3079 & n17258 ;
  assign n17260 = ~n15615 & n17259 ;
  assign n17261 = n4296 ^ n2091 ^ n2013 ;
  assign n17262 = n1018 | n13000 ;
  assign n17263 = n15414 & ~n17262 ;
  assign n17264 = n5766 & ~n9642 ;
  assign n17265 = n8496 ^ n7360 ^ 1'b0 ;
  assign n17266 = n4731 ^ x108 ^ 1'b0 ;
  assign n17267 = n2125 ^ n757 ^ 1'b0 ;
  assign n17268 = n10941 ^ n328 ^ 1'b0 ;
  assign n17269 = ~n8673 & n17268 ;
  assign n17270 = n1495 ^ n410 ^ 1'b0 ;
  assign n17271 = ~n2470 & n17270 ;
  assign n17272 = n9150 ^ n2099 ^ 1'b0 ;
  assign n17273 = n17271 & ~n17272 ;
  assign n17274 = ~n571 & n17273 ;
  assign n17275 = n17274 ^ x37 ^ 1'b0 ;
  assign n17276 = n17269 & n17275 ;
  assign n17277 = n169 | n6092 ;
  assign n17278 = n8196 ^ n4966 ^ 1'b0 ;
  assign n17279 = n2091 | n17278 ;
  assign n17280 = n2453 | n17279 ;
  assign n17281 = n8828 ^ n4761 ^ 1'b0 ;
  assign n17282 = n3491 | n8249 ;
  assign n17283 = ~n413 & n4912 ;
  assign n17284 = ~n2434 & n17283 ;
  assign n17285 = n1540 & ~n7552 ;
  assign n17286 = n17284 & n17285 ;
  assign n17287 = ~n9903 & n17286 ;
  assign n17288 = n17287 ^ n3189 ^ 1'b0 ;
  assign n17289 = ~n10695 & n17288 ;
  assign n17290 = n4907 | n9305 ;
  assign n17291 = n17290 ^ n5711 ^ 1'b0 ;
  assign n17292 = n17291 ^ n7867 ^ 1'b0 ;
  assign n17293 = n9983 & ~n11568 ;
  assign n17294 = ~n17292 & n17293 ;
  assign n17295 = n1161 & n14755 ;
  assign n17296 = n17295 ^ n2030 ^ 1'b0 ;
  assign n17297 = n922 | n1204 ;
  assign n17298 = n3527 & ~n8400 ;
  assign n17299 = n17298 ^ n2629 ^ 1'b0 ;
  assign n17300 = n17299 ^ n2155 ^ 1'b0 ;
  assign n17301 = n1073 | n17300 ;
  assign n17302 = n1916 & ~n5527 ;
  assign n17303 = ~n17254 & n17302 ;
  assign n17304 = n17303 ^ n5365 ^ 1'b0 ;
  assign n17305 = ~n2367 & n17258 ;
  assign n17306 = ~x123 & n1827 ;
  assign n17307 = n11505 ^ n3466 ^ 1'b0 ;
  assign n17308 = n1923 | n17307 ;
  assign n17309 = n5532 & ~n10264 ;
  assign n17310 = n17309 ^ n1302 ^ 1'b0 ;
  assign n17311 = n17310 ^ n10014 ^ 1'b0 ;
  assign n17312 = n771 & ~n10092 ;
  assign n17313 = n17312 ^ n8643 ^ 1'b0 ;
  assign n17314 = x20 & ~n17313 ;
  assign n17315 = n851 & ~n10010 ;
  assign n17316 = ~n7044 & n17315 ;
  assign n17317 = n7930 & ~n8501 ;
  assign n17318 = n8324 & n17317 ;
  assign n17319 = ~n2901 & n3322 ;
  assign n17320 = n2394 | n10816 ;
  assign n17321 = n17320 ^ n10693 ^ 1'b0 ;
  assign n17322 = n4796 & ~n6043 ;
  assign n17323 = n806 ^ n272 ^ 1'b0 ;
  assign n17324 = ~n11249 & n17323 ;
  assign n17325 = ~n3669 & n17324 ;
  assign n17326 = ~n1950 & n9351 ;
  assign n17327 = n17326 ^ n272 ^ 1'b0 ;
  assign n17328 = n17327 ^ n926 ^ 1'b0 ;
  assign n17329 = n845 & n17328 ;
  assign n17330 = n17329 ^ n13144 ^ n7073 ;
  assign n17331 = ( n5046 & ~n5121 ) | ( n5046 & n17330 ) | ( ~n5121 & n17330 ) ;
  assign n17332 = n6635 ^ n5217 ^ 1'b0 ;
  assign n17333 = n10633 | n17332 ;
  assign n17334 = ~n8276 & n17200 ;
  assign n17335 = n17334 ^ n13143 ^ 1'b0 ;
  assign n17336 = n845 & ~n17335 ;
  assign n17337 = n632 & n15651 ;
  assign n17338 = ~n17336 & n17337 ;
  assign n17339 = n3859 ^ x104 ^ 1'b0 ;
  assign n17340 = n781 | n17339 ;
  assign n17341 = n4131 ^ n1046 ^ 1'b0 ;
  assign n17342 = n1298 | n1663 ;
  assign n17343 = n9264 | n17342 ;
  assign n17344 = ~x17 & n7129 ;
  assign n17347 = n5283 & n14203 ;
  assign n17348 = ~n6737 & n17347 ;
  assign n17345 = ~n3531 & n5692 ;
  assign n17346 = n4502 | n17345 ;
  assign n17349 = n17348 ^ n17346 ^ 1'b0 ;
  assign n17350 = n17349 ^ n11049 ^ n9683 ;
  assign n17351 = n1156 ^ n409 ^ 1'b0 ;
  assign n17352 = n785 | n17351 ;
  assign n17353 = n17352 ^ n1317 ^ 1'b0 ;
  assign n17354 = n17350 | n17353 ;
  assign n17355 = n9898 ^ n444 ^ 1'b0 ;
  assign n17356 = n1026 & n1279 ;
  assign n17357 = n528 & n3108 ;
  assign n17358 = n5155 & ~n9490 ;
  assign n17359 = ~n497 & n6236 ;
  assign n17360 = ~n10324 & n17359 ;
  assign n17361 = n6002 ^ n1830 ^ 1'b0 ;
  assign n17362 = ~n17360 & n17361 ;
  assign n17364 = n7495 ^ n1020 ^ 1'b0 ;
  assign n17363 = n14969 | n15141 ;
  assign n17365 = n17364 ^ n17363 ^ 1'b0 ;
  assign n17366 = n17365 ^ n6596 ^ 1'b0 ;
  assign n17367 = n4098 & n6042 ;
  assign n17368 = n2647 & ~n17367 ;
  assign n17369 = n17368 ^ n2263 ^ 1'b0 ;
  assign n17370 = n8121 | n17369 ;
  assign n17371 = n17370 ^ n5789 ^ 1'b0 ;
  assign n17372 = n9244 ^ n1289 ^ 1'b0 ;
  assign n17373 = ~n315 & n17372 ;
  assign n17374 = n17373 ^ n11614 ^ 1'b0 ;
  assign n17375 = n17371 | n17374 ;
  assign n17376 = ~n4382 & n17070 ;
  assign n17377 = n17376 ^ n4673 ^ 1'b0 ;
  assign n17378 = n4319 ^ n1808 ^ 1'b0 ;
  assign n17379 = n4103 & n17378 ;
  assign n17381 = n5732 ^ n2614 ^ 1'b0 ;
  assign n17382 = n3780 | n17381 ;
  assign n17380 = n9172 & ~n17126 ;
  assign n17383 = n17382 ^ n17380 ^ 1'b0 ;
  assign n17384 = n11253 ^ n3816 ^ 1'b0 ;
  assign n17385 = n4173 & ~n6014 ;
  assign n17386 = ~n16332 & n17385 ;
  assign n17387 = n15277 | n17386 ;
  assign n17388 = n7865 & ~n13756 ;
  assign n17389 = n17388 ^ n13503 ^ 1'b0 ;
  assign n17390 = n4817 & n6092 ;
  assign n17391 = n13173 & n17390 ;
  assign n17392 = n13087 & n17391 ;
  assign n17393 = ~n2634 & n3538 ;
  assign n17394 = n17393 ^ n7128 ^ n4502 ;
  assign n17395 = n13506 ^ x96 ^ 1'b0 ;
  assign n17399 = n2501 & ~n9955 ;
  assign n17396 = n2392 & ~n4037 ;
  assign n17397 = ~n14118 & n17396 ;
  assign n17398 = n9389 | n17397 ;
  assign n17400 = n17399 ^ n17398 ^ 1'b0 ;
  assign n17401 = ~n686 & n8859 ;
  assign n17402 = ~n5485 & n17401 ;
  assign n17404 = ~n3406 & n5653 ;
  assign n17403 = ~n4576 & n10217 ;
  assign n17405 = n17404 ^ n17403 ^ 1'b0 ;
  assign n17406 = n6239 ^ n5528 ^ 1'b0 ;
  assign n17407 = n433 & n17406 ;
  assign n17408 = n956 & ~n1181 ;
  assign n17409 = n17408 ^ n6311 ^ 1'b0 ;
  assign n17410 = n17409 ^ n879 ^ 1'b0 ;
  assign n17411 = n2344 & n10752 ;
  assign n17412 = n3083 | n11946 ;
  assign n17413 = n5691 | n17412 ;
  assign n17414 = n12147 | n12538 ;
  assign n17415 = n17414 ^ n17024 ^ 1'b0 ;
  assign n17416 = ( ~n14200 & n17413 ) | ( ~n14200 & n17415 ) | ( n17413 & n17415 ) ;
  assign n17417 = n8266 ^ n3156 ^ 1'b0 ;
  assign n17418 = n7535 ^ n3700 ^ 1'b0 ;
  assign n17419 = n12149 & n17418 ;
  assign n17420 = n2658 | n8580 ;
  assign n17421 = n1387 & ~n17420 ;
  assign n17422 = n14702 ^ n967 ^ 1'b0 ;
  assign n17423 = n16041 | n17422 ;
  assign n17424 = n5689 ^ n2686 ^ 1'b0 ;
  assign n17425 = n2697 & ~n17424 ;
  assign n17426 = n5522 ^ n2020 ^ 1'b0 ;
  assign n17427 = ~n16619 & n17426 ;
  assign n17428 = n14678 ^ n181 ^ 1'b0 ;
  assign n17429 = n11481 & ~n17428 ;
  assign n17430 = n15951 ^ n12607 ^ 1'b0 ;
  assign n17431 = n230 | n16462 ;
  assign n17432 = ~n3755 & n3765 ;
  assign n17433 = n17432 ^ n6770 ^ 1'b0 ;
  assign n17434 = n12436 & ~n15104 ;
  assign n17435 = ~n1172 & n17434 ;
  assign n17436 = ~n163 & n17435 ;
  assign n17438 = n14768 ^ n1554 ^ 1'b0 ;
  assign n17437 = n2364 & n6233 ;
  assign n17439 = n17438 ^ n17437 ^ 1'b0 ;
  assign n17440 = n3192 ^ n790 ^ 1'b0 ;
  assign n17441 = n17440 ^ n2924 ^ 1'b0 ;
  assign n17442 = n14755 ^ n886 ^ 1'b0 ;
  assign n17443 = x19 & n17442 ;
  assign n17444 = ~n3358 & n17443 ;
  assign n17445 = n17444 ^ n2257 ^ 1'b0 ;
  assign n17446 = n7572 & ~n17445 ;
  assign n17447 = x1 | n7077 ;
  assign n17448 = n5363 ^ n1803 ^ n666 ;
  assign n17449 = n616 & ~n1604 ;
  assign n17450 = x10 & ~x90 ;
  assign n17451 = n17450 ^ n8490 ^ n2035 ;
  assign n17452 = n9868 ^ n169 ^ 1'b0 ;
  assign n17453 = n17452 ^ n6525 ^ 1'b0 ;
  assign n17454 = n1887 | n2632 ;
  assign n17455 = n17454 ^ n2934 ^ 1'b0 ;
  assign n17456 = n11915 ^ n7206 ^ 1'b0 ;
  assign n17457 = ~n17455 & n17456 ;
  assign n17458 = n1637 & ~n4357 ;
  assign n17459 = n10191 ^ n8655 ^ 1'b0 ;
  assign n17460 = n8521 ^ n2433 ^ 1'b0 ;
  assign n17461 = n2775 & n17460 ;
  assign n17462 = n5413 ^ n5257 ^ 1'b0 ;
  assign n17463 = n17075 | n17462 ;
  assign n17464 = n1331 | n17463 ;
  assign n17465 = n5586 & n13230 ;
  assign n17466 = n5492 & n17465 ;
  assign n17467 = ~n700 & n7456 ;
  assign n17468 = n17466 & n17467 ;
  assign n17469 = n16386 ^ n14497 ^ 1'b0 ;
  assign n17470 = ~n6456 & n9792 ;
  assign n17471 = n17470 ^ n2087 ^ 1'b0 ;
  assign n17472 = n14915 ^ n12560 ^ 1'b0 ;
  assign n17473 = n11914 & n17472 ;
  assign n17474 = n17473 ^ n11637 ^ 1'b0 ;
  assign n17475 = n2667 & n17474 ;
  assign n17476 = n1378 & ~n2615 ;
  assign n17478 = n387 & n13278 ;
  assign n17479 = n1786 & n6057 ;
  assign n17480 = n17478 & ~n17479 ;
  assign n17477 = ~n3028 & n4682 ;
  assign n17481 = n17480 ^ n17477 ^ 1'b0 ;
  assign n17482 = n4226 & ~n9590 ;
  assign n17483 = n12054 ^ n7222 ^ 1'b0 ;
  assign n17484 = n613 | n17483 ;
  assign n17485 = n5427 & ~n6714 ;
  assign n17486 = n7702 & n8397 ;
  assign n17487 = n4236 & n17486 ;
  assign n17488 = n750 & n11529 ;
  assign n17489 = n10999 ^ n9557 ^ 1'b0 ;
  assign n17490 = n4521 & n17489 ;
  assign n17491 = n8326 & ~n9067 ;
  assign n17492 = n9692 ^ n2344 ^ 1'b0 ;
  assign n17493 = ~n5043 & n17492 ;
  assign n17494 = n2998 & n17493 ;
  assign n17495 = x7 & n17494 ;
  assign n17496 = n15528 ^ n778 ^ 1'b0 ;
  assign n17497 = n1659 | n10861 ;
  assign n17498 = n17497 ^ n14156 ^ 1'b0 ;
  assign n17499 = n727 & ~n14322 ;
  assign n17500 = n1808 & n17499 ;
  assign n17501 = n17500 ^ n428 ^ 1'b0 ;
  assign n17502 = n6309 & ~n8673 ;
  assign n17503 = n3398 & n17502 ;
  assign n17504 = n12291 ^ n5965 ^ n2146 ;
  assign n17505 = n15799 & n17504 ;
  assign n17506 = n10989 & n16897 ;
  assign n17507 = n17506 ^ n6038 ^ 1'b0 ;
  assign n17508 = n4832 ^ n3165 ^ 1'b0 ;
  assign n17509 = ~n10006 & n17508 ;
  assign n17510 = n8111 | n12025 ;
  assign n17511 = n1880 & n7114 ;
  assign n17512 = n1736 | n11796 ;
  assign n17513 = n12903 & ~n14602 ;
  assign n17514 = n5724 & n11804 ;
  assign n17515 = ~n11676 & n17514 ;
  assign n17516 = n2993 | n6502 ;
  assign n17517 = n12271 & ~n17516 ;
  assign n17518 = ~n10530 & n17517 ;
  assign n17519 = n16529 ^ n11418 ^ 1'b0 ;
  assign n17520 = n7123 & ~n17519 ;
  assign n17521 = n4390 | n16035 ;
  assign n17522 = n13394 ^ n5005 ^ 1'b0 ;
  assign n17523 = n7944 | n17522 ;
  assign n17524 = n17523 ^ n2399 ^ 1'b0 ;
  assign n17525 = n12588 ^ n3356 ^ 1'b0 ;
  assign n17527 = n5968 | n8769 ;
  assign n17528 = n12539 & ~n17527 ;
  assign n17529 = ~n5118 & n17528 ;
  assign n17530 = n17529 ^ n3842 ^ 1'b0 ;
  assign n17526 = n11518 | n14001 ;
  assign n17531 = n17530 ^ n17526 ^ 1'b0 ;
  assign n17533 = n1615 ^ n733 ^ 1'b0 ;
  assign n17532 = ~n430 & n9725 ;
  assign n17534 = n17533 ^ n17532 ^ 1'b0 ;
  assign n17535 = n2608 & ~n4751 ;
  assign n17536 = ~n16251 & n17535 ;
  assign n17537 = n5596 | n16092 ;
  assign n17538 = n181 & ~n8608 ;
  assign n17539 = n15040 ^ n12375 ^ 1'b0 ;
  assign n17540 = n17538 | n17539 ;
  assign n17541 = n2682 & ~n16568 ;
  assign n17542 = n17541 ^ n9449 ^ 1'b0 ;
  assign n17543 = ~n4641 & n17542 ;
  assign n17544 = ~n12830 & n17543 ;
  assign n17545 = ~n5680 & n17544 ;
  assign n17546 = n9271 ^ x14 ^ 1'b0 ;
  assign n17547 = n16872 ^ n6610 ^ 1'b0 ;
  assign n17548 = n17546 | n17547 ;
  assign n17549 = n7133 ^ x11 ^ 1'b0 ;
  assign n17550 = x42 & ~n17549 ;
  assign n17551 = n2248 | n14427 ;
  assign n17552 = n9779 & ~n16397 ;
  assign n17553 = ~n5582 & n17552 ;
  assign n17554 = n1694 & ~n6280 ;
  assign n17555 = n6223 & n9734 ;
  assign n17556 = n17555 ^ n3350 ^ 1'b0 ;
  assign n17557 = n2942 ^ n2198 ^ 1'b0 ;
  assign n17558 = n17557 ^ n14657 ^ 1'b0 ;
  assign n17559 = n9756 ^ n1178 ^ 1'b0 ;
  assign n17560 = n13549 & ~n17559 ;
  assign n17561 = n7137 ^ n6095 ^ n430 ;
  assign n17562 = n1154 & ~n17561 ;
  assign n17563 = n6324 | n17562 ;
  assign n17564 = ~n696 & n7695 ;
  assign n17565 = n5727 & n17564 ;
  assign n17566 = n2264 & n5273 ;
  assign n17567 = n2016 & ~n4506 ;
  assign n17569 = n1351 & ~n13552 ;
  assign n17568 = n11613 ^ n7277 ^ 1'b0 ;
  assign n17570 = n17569 ^ n17568 ^ 1'b0 ;
  assign n17571 = n3607 & ~n4454 ;
  assign n17572 = n17571 ^ n10057 ^ 1'b0 ;
  assign n17573 = n14784 ^ n696 ^ 1'b0 ;
  assign n17574 = n13137 & ~n17573 ;
  assign n17575 = n14878 & n17574 ;
  assign n17576 = n17575 ^ n6018 ^ 1'b0 ;
  assign n17577 = n477 | n3504 ;
  assign n17578 = n2459 | n17577 ;
  assign n17579 = n3986 & ~n17578 ;
  assign n17580 = n1329 & ~n2186 ;
  assign n17581 = n17579 & n17580 ;
  assign n17582 = n4120 & ~n5352 ;
  assign n17584 = n2842 & n3539 ;
  assign n17583 = n9247 & n15797 ;
  assign n17585 = n17584 ^ n17583 ^ 1'b0 ;
  assign n17586 = n17585 ^ n10029 ^ 1'b0 ;
  assign n17587 = ( ~n3367 & n17582 ) | ( ~n3367 & n17586 ) | ( n17582 & n17586 ) ;
  assign n17588 = n5448 ^ n272 ^ 1'b0 ;
  assign n17589 = n6304 & ~n17588 ;
  assign n17590 = ~n216 & n3450 ;
  assign n17591 = ~n17589 & n17590 ;
  assign n17592 = n5183 & ~n17591 ;
  assign n17593 = n17581 & n17592 ;
  assign n17594 = n17350 ^ n8689 ^ 1'b0 ;
  assign n17595 = ~n16266 & n17594 ;
  assign n17596 = n1602 & n17595 ;
  assign n17597 = n17596 ^ n13354 ^ 1'b0 ;
  assign n17598 = n3459 ^ n2441 ^ 1'b0 ;
  assign n17600 = n8518 ^ n4106 ^ 1'b0 ;
  assign n17601 = ( n4991 & n5718 ) | ( n4991 & ~n17600 ) | ( n5718 & ~n17600 ) ;
  assign n17599 = n7283 ^ x88 ^ 1'b0 ;
  assign n17602 = n17601 ^ n17599 ^ 1'b0 ;
  assign n17603 = ~n11040 & n17602 ;
  assign n17604 = n17603 ^ n5381 ^ 1'b0 ;
  assign n17605 = n509 & ~n1284 ;
  assign n17606 = n17605 ^ x65 ^ 1'b0 ;
  assign n17607 = n2977 & ~n4484 ;
  assign n17609 = n3816 & ~n6180 ;
  assign n17608 = n3483 & ~n4288 ;
  assign n17610 = n17609 ^ n17608 ^ 1'b0 ;
  assign n17611 = n13278 ^ n2819 ^ 1'b0 ;
  assign n17612 = n4677 & n17611 ;
  assign n17613 = n14576 ^ n13541 ^ 1'b0 ;
  assign n17614 = n6915 & n17613 ;
  assign n17617 = n2089 | n3700 ;
  assign n17615 = n7560 ^ n7347 ^ n2030 ;
  assign n17616 = ~n13948 & n17615 ;
  assign n17618 = n17617 ^ n17616 ^ 1'b0 ;
  assign n17619 = n6017 & ~n11309 ;
  assign n17620 = n17619 ^ n3096 ^ 1'b0 ;
  assign n17621 = n17618 & ~n17620 ;
  assign n17622 = ~n8387 & n12130 ;
  assign n17626 = n2371 | n5763 ;
  assign n17623 = n4929 & n7518 ;
  assign n17624 = ~n4528 & n17623 ;
  assign n17625 = n16461 | n17624 ;
  assign n17627 = n17626 ^ n17625 ^ 1'b0 ;
  assign n17628 = ~n6557 & n7832 ;
  assign n17629 = n12964 & n17628 ;
  assign n17630 = n17629 ^ n5411 ^ 1'b0 ;
  assign n17631 = n3415 | n14828 ;
  assign n17632 = n17631 ^ n14471 ^ 1'b0 ;
  assign n17635 = n4793 | n14252 ;
  assign n17636 = n3640 | n17635 ;
  assign n17633 = n13644 ^ n6766 ^ n2942 ;
  assign n17634 = n11623 & ~n17633 ;
  assign n17637 = n17636 ^ n17634 ^ 1'b0 ;
  assign n17638 = n3045 ^ n1955 ^ 1'b0 ;
  assign n17639 = n846 | n4120 ;
  assign n17640 = n17639 ^ n9511 ^ 1'b0 ;
  assign n17641 = n17638 & ~n17640 ;
  assign n17642 = n9729 ^ n5842 ^ 1'b0 ;
  assign n17643 = n13714 & n17642 ;
  assign n17644 = n11044 | n17643 ;
  assign n17645 = n201 & ~n3977 ;
  assign n17646 = n2432 & n5130 ;
  assign n17647 = n17646 ^ n14111 ^ 1'b0 ;
  assign n17648 = n6826 & ~n17647 ;
  assign n17649 = n4307 ^ n616 ^ 1'b0 ;
  assign n17650 = n15881 ^ n9719 ^ 1'b0 ;
  assign n17651 = n3196 & n17650 ;
  assign n17652 = n17651 ^ n13857 ^ 1'b0 ;
  assign n17653 = ~n3334 & n9571 ;
  assign n17654 = n11117 ^ n1917 ^ 1'b0 ;
  assign n17655 = x53 & n17654 ;
  assign n17656 = n365 & n950 ;
  assign n17657 = n2861 ^ n1226 ^ 1'b0 ;
  assign n17658 = n1070 | n17657 ;
  assign n17659 = n5437 ^ n1497 ^ 1'b0 ;
  assign n17660 = ~n446 & n17659 ;
  assign n17661 = n17660 ^ n10470 ^ 1'b0 ;
  assign n17662 = ~n10209 & n17661 ;
  assign n17663 = n17662 ^ n3409 ^ 1'b0 ;
  assign n17664 = ~n17658 & n17663 ;
  assign n17665 = n5289 & n7456 ;
  assign n17666 = ~n12417 & n17665 ;
  assign n17667 = n4787 | n5965 ;
  assign n17668 = n17667 ^ n15510 ^ 1'b0 ;
  assign n17669 = n4648 & ~n12423 ;
  assign n17670 = n17669 ^ n2043 ^ 1'b0 ;
  assign n17671 = n5804 & ~n17256 ;
  assign n17672 = n4354 ^ n1668 ^ 1'b0 ;
  assign n17673 = ~n279 & n750 ;
  assign n17674 = ~n17672 & n17673 ;
  assign n17675 = n13395 & n17674 ;
  assign n17676 = n7873 & n10427 ;
  assign n17677 = n17444 ^ n2073 ^ 1'b0 ;
  assign n17678 = n4019 & n8608 ;
  assign n17679 = n3204 & n12518 ;
  assign n17680 = n248 & ~n2836 ;
  assign n17681 = n15321 | n17680 ;
  assign n17682 = n17679 | n17681 ;
  assign n17683 = n323 & n7280 ;
  assign n17684 = n4645 | n13742 ;
  assign n17685 = n17684 ^ n17016 ^ 1'b0 ;
  assign n17686 = n1367 | n3454 ;
  assign n17687 = x105 & n7361 ;
  assign n17688 = n480 & n17687 ;
  assign n17689 = n2615 | n17688 ;
  assign n17690 = n17689 ^ n9864 ^ 1'b0 ;
  assign n17691 = n10305 & n17690 ;
  assign n17692 = n885 | n12045 ;
  assign n17693 = n5016 & ~n9651 ;
  assign n17694 = n7270 & n17693 ;
  assign n17695 = ~n4768 & n17221 ;
  assign n17696 = n4014 ^ n2402 ^ 1'b0 ;
  assign n17697 = ~n2087 & n17696 ;
  assign n17698 = ~n15386 & n17697 ;
  assign n17699 = n17698 ^ n1381 ^ 1'b0 ;
  assign n17700 = n1526 | n3905 ;
  assign n17701 = n17700 ^ n3319 ^ 1'b0 ;
  assign n17702 = n10478 & ~n12832 ;
  assign n17703 = n17702 ^ n8324 ^ 1'b0 ;
  assign n17704 = n15482 ^ n12029 ^ 1'b0 ;
  assign n17705 = n16698 ^ n9047 ^ 1'b0 ;
  assign n17706 = n7167 | n14066 ;
  assign n17707 = n17706 ^ n16103 ^ 1'b0 ;
  assign n17708 = ~n3238 & n17707 ;
  assign n17709 = n230 & n277 ;
  assign n17710 = n552 & n17709 ;
  assign n17711 = n1774 & n17710 ;
  assign n17712 = n17711 ^ n4112 ^ 1'b0 ;
  assign n17713 = n14009 & n17712 ;
  assign n17714 = n13782 ^ n4661 ^ n978 ;
  assign n17715 = n2667 & n13327 ;
  assign n17716 = n17126 & n17715 ;
  assign n17717 = n13099 ^ n9119 ^ 1'b0 ;
  assign n17718 = n17200 & n17717 ;
  assign n17719 = n4919 ^ n2799 ^ 1'b0 ;
  assign n17720 = n4371 & ~n10329 ;
  assign n17721 = n639 ^ n150 ^ 1'b0 ;
  assign n17722 = n17721 ^ n14270 ^ n3289 ;
  assign n17723 = n17722 ^ n12727 ^ 1'b0 ;
  assign n17724 = ~n198 & n10203 ;
  assign n17725 = n5539 | n9853 ;
  assign n17726 = n17725 ^ n8046 ^ 1'b0 ;
  assign n17727 = n1452 & ~n17726 ;
  assign n17728 = n1866 & ~n16501 ;
  assign n17729 = ~n13983 & n17728 ;
  assign n17730 = n6360 ^ n5317 ^ 1'b0 ;
  assign n17731 = n3977 | n17730 ;
  assign n17732 = n6728 & ~n17731 ;
  assign n17733 = ~n2579 & n10425 ;
  assign n17734 = ( n1795 & n1993 ) | ( n1795 & ~n14955 ) | ( n1993 & ~n14955 ) ;
  assign n17735 = n16110 ^ n14914 ^ 1'b0 ;
  assign n17736 = n1542 ^ n800 ^ 1'b0 ;
  assign n17737 = n586 & n17736 ;
  assign n17738 = n15434 & n17737 ;
  assign n17739 = n3823 & ~n7841 ;
  assign n17740 = n17739 ^ n15030 ^ 1'b0 ;
  assign n17741 = n10006 ^ n3392 ^ 1'b0 ;
  assign n17742 = n2409 & ~n17741 ;
  assign n17743 = n7694 ^ n1983 ^ 1'b0 ;
  assign n17744 = x100 | n17743 ;
  assign n17745 = n17744 ^ n8767 ^ 1'b0 ;
  assign n17746 = n12027 ^ n1656 ^ 1'b0 ;
  assign n17747 = n5504 ^ n4767 ^ 1'b0 ;
  assign n17748 = n1751 | n3559 ;
  assign n17749 = n17748 ^ n870 ^ 1'b0 ;
  assign n17750 = ~n16298 & n17749 ;
  assign n17751 = n9856 ^ x85 ^ 1'b0 ;
  assign n17752 = n11586 | n15409 ;
  assign n17753 = n17752 ^ n5862 ^ 1'b0 ;
  assign n17754 = n1663 & ~n7383 ;
  assign n17755 = n7371 ^ n5595 ^ 1'b0 ;
  assign n17756 = n14823 & n17755 ;
  assign n17757 = n3489 & n12776 ;
  assign n17758 = ~n17756 & n17757 ;
  assign n17759 = n2253 ^ n1491 ^ n932 ;
  assign n17760 = x80 & n16529 ;
  assign n17761 = n17760 ^ n1432 ^ 1'b0 ;
  assign n17762 = n14856 | n17761 ;
  assign n17763 = n17762 ^ n8885 ^ 1'b0 ;
  assign n17764 = n5347 ^ n707 ^ 1'b0 ;
  assign n17765 = n7037 & n17764 ;
  assign n17766 = ( n4465 & n11364 ) | ( n4465 & ~n17765 ) | ( n11364 & ~n17765 ) ;
  assign n17767 = n3108 | n11170 ;
  assign n17768 = n535 & n7785 ;
  assign n17769 = n9553 & n17768 ;
  assign n17770 = n5617 ^ n2091 ^ 1'b0 ;
  assign n17771 = n9047 ^ n7222 ^ 1'b0 ;
  assign n17772 = n6190 & n15340 ;
  assign n17773 = n12655 & n17772 ;
  assign n17777 = n3843 ^ n1958 ^ 1'b0 ;
  assign n17774 = n5239 ^ n4204 ^ 1'b0 ;
  assign n17775 = n17774 ^ n1618 ^ 1'b0 ;
  assign n17776 = ~n4070 & n17775 ;
  assign n17778 = n17777 ^ n17776 ^ 1'b0 ;
  assign n17779 = n2381 & n4345 ;
  assign n17780 = n169 | n16071 ;
  assign n17781 = n11624 ^ n1329 ^ 1'b0 ;
  assign n17782 = n8322 ^ x8 ^ 1'b0 ;
  assign n17783 = ~n4908 & n17782 ;
  assign n17784 = n17781 & ~n17783 ;
  assign n17785 = n12958 & ~n16501 ;
  assign n17786 = n17785 ^ n828 ^ 1'b0 ;
  assign n17787 = n1317 | n13604 ;
  assign n17788 = n8193 & ~n17787 ;
  assign n17789 = n2331 | n6086 ;
  assign n17790 = n17789 ^ n1979 ^ 1'b0 ;
  assign n17791 = n12113 ^ n2005 ^ 1'b0 ;
  assign n17792 = n17790 | n17791 ;
  assign n17793 = ~n13945 & n15423 ;
  assign n17794 = n17792 & n17793 ;
  assign n17795 = n7911 ^ n7242 ^ 1'b0 ;
  assign n17796 = n10280 & n17795 ;
  assign n17797 = n17796 ^ n12585 ^ 1'b0 ;
  assign n17798 = n17797 ^ n1116 ^ 1'b0 ;
  assign n17799 = ~n287 & n17798 ;
  assign n17800 = x100 & n8022 ;
  assign n17801 = n9638 ^ n3158 ^ 1'b0 ;
  assign n17802 = n17800 & ~n17801 ;
  assign n17803 = n3976 ^ n1574 ^ 1'b0 ;
  assign n17804 = n17802 & ~n17803 ;
  assign n17805 = n14198 & n17804 ;
  assign n17806 = n9572 ^ n6011 ^ 1'b0 ;
  assign n17807 = n5097 & n8709 ;
  assign n17808 = ~n4621 & n12682 ;
  assign n17809 = n6239 & ~n17808 ;
  assign n17810 = n3611 & ~n13969 ;
  assign n17811 = n9343 ^ n9196 ^ 1'b0 ;
  assign n17812 = n335 & n17811 ;
  assign n17813 = n2023 & n17812 ;
  assign n17814 = ~n2364 & n17813 ;
  assign n17815 = ( n1589 & n6474 ) | ( n1589 & ~n15423 ) | ( n6474 & ~n15423 ) ;
  assign n17816 = n5352 | n17815 ;
  assign n17817 = n2749 | n17816 ;
  assign n17818 = n17817 ^ n8271 ^ 1'b0 ;
  assign n17819 = n16835 & ~n17818 ;
  assign n17820 = ( n6917 & n11505 ) | ( n6917 & n12972 ) | ( n11505 & n12972 ) ;
  assign n17821 = n6926 | n14860 ;
  assign n17822 = n16236 ^ n1830 ^ 1'b0 ;
  assign n17823 = n1395 & n9490 ;
  assign n17824 = n5245 & n6017 ;
  assign n17825 = n17480 & ~n17824 ;
  assign n17826 = n17825 ^ n15615 ^ 1'b0 ;
  assign n17827 = n17582 ^ n13195 ^ 1'b0 ;
  assign n17828 = ~n4354 & n7705 ;
  assign n17829 = n4809 & ~n12270 ;
  assign n17830 = n4492 & ~n10234 ;
  assign n17831 = n17830 ^ n10937 ^ 1'b0 ;
  assign n17832 = n3840 | n9430 ;
  assign n17833 = n7821 & ~n17832 ;
  assign n17834 = n1830 & ~n17833 ;
  assign n17835 = n1990 | n13527 ;
  assign n17836 = n2630 | n17835 ;
  assign n17837 = n1918 & n5705 ;
  assign n17838 = n17837 ^ n5380 ^ 1'b0 ;
  assign n17839 = n967 | n5392 ;
  assign n17840 = n17839 ^ n2073 ^ 1'b0 ;
  assign n17841 = n17840 ^ n14299 ^ 1'b0 ;
  assign n17842 = ~n1683 & n9261 ;
  assign n17843 = n5337 | n17842 ;
  assign n17844 = n1177 & ~n6703 ;
  assign n17845 = n17844 ^ n547 ^ 1'b0 ;
  assign n17846 = n3204 ^ n2655 ^ 1'b0 ;
  assign n17847 = n14893 ^ n5622 ^ 1'b0 ;
  assign n17848 = n5860 & ~n17847 ;
  assign n17849 = n7298 ^ n2436 ^ 1'b0 ;
  assign n17850 = n4467 & ~n17849 ;
  assign n17851 = n2115 & ~n2361 ;
  assign n17852 = n17851 ^ n3567 ^ 1'b0 ;
  assign n17853 = n7622 | n17852 ;
  assign n17854 = n4525 | n17853 ;
  assign n17855 = n17711 ^ n7600 ^ 1'b0 ;
  assign n17856 = n9268 & n17855 ;
  assign n17857 = n17856 ^ n12457 ^ n6398 ;
  assign n17858 = n17857 ^ n2238 ^ 1'b0 ;
  assign n17859 = n3544 ^ n707 ^ 1'b0 ;
  assign n17860 = n10591 | n17859 ;
  assign n17861 = n17860 ^ n7756 ^ x118 ;
  assign n17862 = n16944 ^ n7607 ^ 1'b0 ;
  assign n17863 = n15115 | n17246 ;
  assign n17864 = n2931 & n10619 ;
  assign n17865 = n17863 & n17864 ;
  assign n17866 = ( n1177 & n5615 ) | ( n1177 & ~n8021 ) | ( n5615 & ~n8021 ) ;
  assign n17867 = n5605 ^ n2117 ^ 1'b0 ;
  assign n17868 = ~n17866 & n17867 ;
  assign n17869 = n17868 ^ n12784 ^ 1'b0 ;
  assign n17870 = n17869 ^ n15995 ^ 1'b0 ;
  assign n17871 = n2604 & ~n10595 ;
  assign n17872 = n3840 & ~n16891 ;
  assign n17873 = n9760 ^ n6257 ^ 1'b0 ;
  assign n17874 = n4784 & ~n16713 ;
  assign n17878 = n7436 ^ n409 ^ 1'b0 ;
  assign n17879 = ~n8185 & n17878 ;
  assign n17875 = n788 & ~n3950 ;
  assign n17876 = n17875 ^ n2384 ^ 1'b0 ;
  assign n17877 = n10812 & n17876 ;
  assign n17880 = n17879 ^ n17877 ^ 1'b0 ;
  assign n17881 = n14823 ^ n14478 ^ 1'b0 ;
  assign n17882 = n5898 & ~n13955 ;
  assign n17883 = n8747 ^ n6528 ^ n6355 ;
  assign n17884 = ~n4556 & n12146 ;
  assign n17885 = ~n16897 & n17884 ;
  assign n17886 = n1602 & ~n11014 ;
  assign n17887 = n16576 ^ n7020 ^ 1'b0 ;
  assign n17888 = ~n7573 & n17887 ;
  assign n17889 = n6348 ^ n4747 ^ 1'b0 ;
  assign n17890 = n3063 & ~n17889 ;
  assign n17891 = n5568 ^ n632 ^ n623 ;
  assign n17892 = n3180 | n12015 ;
  assign n17893 = ~n2898 & n5476 ;
  assign n17894 = n17892 & n17893 ;
  assign n17895 = n5886 ^ n3085 ^ 1'b0 ;
  assign n17896 = n3353 & n13938 ;
  assign n17897 = ~n15569 & n17896 ;
  assign n17898 = n11164 ^ n1913 ^ 1'b0 ;
  assign n17899 = ~n3454 & n8892 ;
  assign n17900 = n17899 ^ n4602 ^ 1'b0 ;
  assign n17901 = n3041 | n17900 ;
  assign n17902 = n3484 ^ n1260 ^ 1'b0 ;
  assign n17903 = n5239 & n17902 ;
  assign n17904 = n15467 ^ n721 ^ 1'b0 ;
  assign n17905 = n17903 | n17904 ;
  assign n17906 = n17901 & ~n17905 ;
  assign n17907 = ~n15066 & n17906 ;
  assign n17908 = n4459 ^ n520 ^ 1'b0 ;
  assign n17911 = n5562 | n6221 ;
  assign n17909 = ~n2349 & n6688 ;
  assign n17910 = ( n11155 & n14327 ) | ( n11155 & ~n17909 ) | ( n14327 & ~n17909 ) ;
  assign n17912 = n17911 ^ n17910 ^ 1'b0 ;
  assign n17913 = ~n12063 & n17912 ;
  assign n17914 = n17913 ^ x41 ^ 1'b0 ;
  assign n17915 = ~n660 & n6094 ;
  assign n17916 = n17915 ^ n6565 ^ 1'b0 ;
  assign n17917 = n6813 | n10470 ;
  assign n17919 = ~n5771 & n15569 ;
  assign n17918 = n3217 & n14878 ;
  assign n17920 = n17919 ^ n17918 ^ 1'b0 ;
  assign n17921 = n4589 ^ n1808 ^ 1'b0 ;
  assign n17922 = n14842 & n17921 ;
  assign n17923 = ~n13330 & n17922 ;
  assign n17924 = ~n3526 & n3804 ;
  assign n17925 = n17924 ^ n8531 ^ 1'b0 ;
  assign n17926 = n9205 & n17925 ;
  assign n17928 = ~n978 & n2203 ;
  assign n17929 = ~n2203 & n17928 ;
  assign n17930 = ~n1089 & n17929 ;
  assign n17931 = n6158 ^ n2564 ^ 1'b0 ;
  assign n17932 = n17930 & n17931 ;
  assign n17933 = ~n6698 & n17932 ;
  assign n17934 = n1344 & ~n3651 ;
  assign n17935 = n3651 & n17934 ;
  assign n17936 = n571 | n17935 ;
  assign n17937 = n571 & ~n17936 ;
  assign n17938 = n17933 | n17937 ;
  assign n17939 = n17933 & ~n17938 ;
  assign n17940 = n1199 & ~n4555 ;
  assign n17941 = n4555 & n17940 ;
  assign n17942 = n17941 ^ n14828 ^ 1'b0 ;
  assign n17943 = n9636 & ~n17942 ;
  assign n17944 = n17939 & n17943 ;
  assign n17927 = n4974 & ~n9736 ;
  assign n17945 = n17944 ^ n17927 ^ 1'b0 ;
  assign n17946 = n4289 & ~n4615 ;
  assign n17947 = ~n4289 & n17946 ;
  assign n17948 = n373 & ~n13811 ;
  assign n17949 = n17947 & n17948 ;
  assign n17950 = n17945 & ~n17949 ;
  assign n17951 = ~n17945 & n17950 ;
  assign n17952 = n6430 | n11496 ;
  assign n17953 = n6289 & ~n17952 ;
  assign n17954 = ~n3637 & n12201 ;
  assign n17955 = n17954 ^ n6278 ^ 1'b0 ;
  assign n17956 = n17953 | n17955 ;
  assign n17957 = n3169 & ~n17956 ;
  assign n17958 = n9170 ^ n983 ^ 1'b0 ;
  assign n17959 = n1773 | n3045 ;
  assign n17960 = n4445 & ~n10182 ;
  assign n17961 = ~n5369 & n17960 ;
  assign n17962 = ~n1133 & n8599 ;
  assign n17963 = n967 & n17962 ;
  assign n17964 = n12721 ^ n5723 ^ 1'b0 ;
  assign n17965 = n6026 & ~n7965 ;
  assign n17966 = ~n1560 & n17965 ;
  assign n17967 = n5283 & n7203 ;
  assign n17968 = n13251 & ~n17538 ;
  assign n17969 = n1298 & n10937 ;
  assign n17970 = n1788 & ~n17969 ;
  assign n17971 = n13153 ^ n6575 ^ 1'b0 ;
  assign n17972 = n5550 & n17413 ;
  assign n17973 = ~n4920 & n9521 ;
  assign n17974 = n2518 | n15403 ;
  assign n17975 = n13236 ^ n8183 ^ 1'b0 ;
  assign n17976 = n3149 & n4391 ;
  assign n17977 = n17976 ^ n4408 ^ 1'b0 ;
  assign n17978 = n3979 ^ n3829 ^ 1'b0 ;
  assign n17979 = ~n8522 & n8902 ;
  assign n17980 = n3941 & ~n10526 ;
  assign n17981 = n9308 ^ n632 ^ 1'b0 ;
  assign n17982 = n17981 ^ n522 ^ 1'b0 ;
  assign n17983 = ~n4923 & n17982 ;
  assign n17984 = ~n2634 & n3499 ;
  assign n17985 = n6423 & n17984 ;
  assign n17986 = n17985 ^ n1773 ^ 1'b0 ;
  assign n17987 = n7658 | n11527 ;
  assign n17988 = n17987 ^ n4443 ^ 1'b0 ;
  assign n17989 = n4343 & ~n17988 ;
  assign n17990 = ~n828 & n15969 ;
  assign n17991 = n17990 ^ n11696 ^ 1'b0 ;
  assign n17992 = n8278 ^ n5618 ^ 1'b0 ;
  assign n17993 = n5102 | n17617 ;
  assign n17994 = n7796 | n17993 ;
  assign n17995 = n14711 & ~n17907 ;
  assign n17996 = n17995 ^ n8058 ^ 1'b0 ;
  assign n17997 = n10006 ^ n7347 ^ 1'b0 ;
  assign n17998 = ~n15650 & n17997 ;
  assign n17999 = n5268 & ~n5425 ;
  assign n18000 = n17999 ^ n16146 ^ 1'b0 ;
  assign n18001 = n3430 & ~n18000 ;
  assign n18002 = n7236 ^ n6607 ^ 1'b0 ;
  assign n18003 = n7899 & n15299 ;
  assign n18004 = n5907 ^ x9 ^ 1'b0 ;
  assign n18005 = n6947 & ~n18004 ;
  assign n18006 = n4507 & ~n8501 ;
  assign n18007 = n18006 ^ n1262 ^ 1'b0 ;
  assign n18008 = ~n7809 & n9815 ;
  assign n18010 = n3077 ^ x96 ^ 1'b0 ;
  assign n18009 = n12916 | n13149 ;
  assign n18011 = n18010 ^ n18009 ^ 1'b0 ;
  assign n18012 = n2718 & n3462 ;
  assign n18013 = n18012 ^ n1335 ^ 1'b0 ;
  assign n18014 = ~n3890 & n18013 ;
  assign n18015 = n693 | n2127 ;
  assign n18016 = n9836 & n18015 ;
  assign n18017 = ~n18014 & n18016 ;
  assign n18018 = n3812 ^ n2659 ^ 1'b0 ;
  assign n18019 = n8980 & ~n13185 ;
  assign n18020 = n2969 ^ n2215 ^ 1'b0 ;
  assign n18021 = n9940 & n12215 ;
  assign n18022 = n18020 & n18021 ;
  assign n18023 = ~n3269 & n10142 ;
  assign n18024 = n18023 ^ n5181 ^ 1'b0 ;
  assign n18025 = n5451 ^ n2782 ^ 1'b0 ;
  assign n18026 = n18025 ^ n2002 ^ 1'b0 ;
  assign n18027 = n9105 ^ n6665 ^ n6421 ;
  assign n18028 = n8142 ^ n1270 ^ 1'b0 ;
  assign n18029 = n6333 & n18028 ;
  assign n18030 = ~n2470 & n10878 ;
  assign n18031 = n13103 ^ n6084 ^ 1'b0 ;
  assign n18032 = n10876 | n18031 ;
  assign n18033 = n6902 & ~n18032 ;
  assign n18034 = n3592 & n9161 ;
  assign n18035 = n907 | n9874 ;
  assign n18036 = n18035 ^ n3677 ^ 1'b0 ;
  assign n18037 = n3635 & ~n5981 ;
  assign n18038 = n9648 ^ n8655 ^ 1'b0 ;
  assign n18039 = ~n6260 & n18038 ;
  assign n18040 = n259 & n3697 ;
  assign n18041 = n2386 | n11582 ;
  assign n18042 = n782 & ~n9069 ;
  assign n18043 = n18042 ^ n9031 ^ 1'b0 ;
  assign n18044 = n18043 ^ n7138 ^ 1'b0 ;
  assign n18045 = n1597 | n11482 ;
  assign n18046 = n1714 | n18045 ;
  assign n18047 = n8047 ^ n504 ^ 1'b0 ;
  assign n18048 = n7690 & n17509 ;
  assign n18049 = ~n677 & n4267 ;
  assign n18050 = n11515 & n18049 ;
  assign n18051 = n17632 & ~n18050 ;
  assign n18052 = n3270 & n18051 ;
  assign n18053 = n11573 ^ n8107 ^ 1'b0 ;
  assign n18056 = n394 & ~n11901 ;
  assign n18057 = n18056 ^ n16242 ^ 1'b0 ;
  assign n18054 = n5929 | n7383 ;
  assign n18055 = n3210 & ~n18054 ;
  assign n18058 = n18057 ^ n18055 ^ 1'b0 ;
  assign n18059 = n3572 | n9417 ;
  assign n18060 = n18059 ^ n629 ^ 1'b0 ;
  assign n18061 = n2248 & n13828 ;
  assign n18062 = ~n15821 & n18061 ;
  assign n18063 = n18062 ^ n10980 ^ 1'b0 ;
  assign n18064 = n3846 ^ n1280 ^ 1'b0 ;
  assign n18065 = ~n171 & n6474 ;
  assign n18066 = ~n18064 & n18065 ;
  assign n18067 = n8958 & ~n14061 ;
  assign n18068 = ~n13715 & n18067 ;
  assign n18069 = n16438 ^ n15890 ^ n12136 ;
  assign n18070 = n13418 | n16100 ;
  assign n18071 = n6147 & ~n7647 ;
  assign n18072 = n1816 & ~n12585 ;
  assign n18073 = n18072 ^ n12101 ^ 1'b0 ;
  assign n18074 = ~n4696 & n18073 ;
  assign n18075 = n1913 & n3147 ;
  assign n18076 = n18075 ^ n4880 ^ 1'b0 ;
  assign n18077 = n12474 & ~n18076 ;
  assign n18078 = ~n6958 & n18077 ;
  assign n18082 = ~n2936 & n6167 ;
  assign n18079 = ~n5711 & n10725 ;
  assign n18080 = n5213 & ~n9256 ;
  assign n18081 = ~n18079 & n18080 ;
  assign n18083 = n18082 ^ n18081 ^ n8772 ;
  assign n18084 = n4114 ^ n965 ^ 1'b0 ;
  assign n18085 = n16174 & ~n18084 ;
  assign n18086 = ~n3021 & n12344 ;
  assign n18087 = n18086 ^ n704 ^ 1'b0 ;
  assign n18088 = n3034 & ~n18087 ;
  assign n18089 = n6056 & ~n9474 ;
  assign n18090 = ~n10163 & n18089 ;
  assign n18091 = n4450 & ~n11469 ;
  assign n18092 = n17639 ^ n1199 ^ 1'b0 ;
  assign n18093 = n4431 | n9816 ;
  assign n18094 = n18093 ^ n2525 ^ 1'b0 ;
  assign n18095 = n18094 ^ n13880 ^ 1'b0 ;
  assign n18096 = n18095 ^ n514 ^ 1'b0 ;
  assign n18097 = n583 & ~n18096 ;
  assign n18098 = n806 & ~n4846 ;
  assign n18099 = ~n6729 & n18098 ;
  assign n18100 = n12687 ^ n3819 ^ 1'b0 ;
  assign n18101 = n18099 & ~n18100 ;
  assign n18102 = n16959 ^ n9641 ^ 1'b0 ;
  assign n18103 = n1470 & n3843 ;
  assign n18104 = ~n3215 & n18103 ;
  assign n18105 = n8021 & ~n18104 ;
  assign n18107 = n1579 ^ n439 ^ 1'b0 ;
  assign n18106 = ~n15147 & n15682 ;
  assign n18108 = n18107 ^ n18106 ^ 1'b0 ;
  assign n18109 = ~n704 & n10017 ;
  assign n18110 = n3066 | n4301 ;
  assign n18111 = n6563 & ~n18110 ;
  assign n18112 = n1950 | n18111 ;
  assign n18113 = n11597 ^ n1685 ^ 1'b0 ;
  assign n18114 = ~n2872 & n3581 ;
  assign n18115 = n18114 ^ n9347 ^ 1'b0 ;
  assign n18116 = n18115 ^ n14650 ^ 1'b0 ;
  assign n18117 = n8529 | n18116 ;
  assign n18118 = ~x37 & n1046 ;
  assign n18119 = ~n14556 & n18118 ;
  assign n18120 = n666 & n1566 ;
  assign n18121 = n18120 ^ n330 ^ 1'b0 ;
  assign n18122 = n624 & n18121 ;
  assign n18123 = n6212 ^ n3482 ^ 1'b0 ;
  assign n18124 = n4363 ^ n1452 ^ 1'b0 ;
  assign n18125 = n1571 | n18124 ;
  assign n18126 = n18125 ^ n9459 ^ 1'b0 ;
  assign n18127 = n11151 ^ n9047 ^ 1'b0 ;
  assign n18128 = n4100 | n18127 ;
  assign n18130 = n1972 | n13039 ;
  assign n18129 = ~n2448 & n3529 ;
  assign n18131 = n18130 ^ n18129 ^ 1'b0 ;
  assign n18132 = ~n1290 & n18131 ;
  assign n18133 = n7266 & n17589 ;
  assign n18134 = ~n18132 & n18133 ;
  assign n18135 = n7829 ^ n192 ^ 1'b0 ;
  assign n18136 = ~n1165 & n5589 ;
  assign n18137 = n18136 ^ n17358 ^ n14242 ;
  assign n18138 = n1205 & ~n5276 ;
  assign n18139 = n17907 & n18138 ;
  assign n18140 = x33 & n8425 ;
  assign n18141 = n4919 & n18140 ;
  assign n18142 = n14200 ^ n6495 ^ 1'b0 ;
  assign n18143 = ( n1260 & n18141 ) | ( n1260 & ~n18142 ) | ( n18141 & ~n18142 ) ;
  assign n18144 = n984 & ~n17630 ;
  assign n18145 = n18144 ^ n1344 ^ 1'b0 ;
  assign n18146 = n6788 | n16266 ;
  assign n18147 = n17643 ^ n198 ^ 1'b0 ;
  assign n18148 = n3595 | n18147 ;
  assign n18149 = n2518 & ~n18148 ;
  assign n18150 = n4816 ^ n806 ^ 1'b0 ;
  assign n18151 = n5522 ^ n4579 ^ 1'b0 ;
  assign n18152 = n18151 ^ n17120 ^ 1'b0 ;
  assign n18153 = n18150 & n18152 ;
  assign n18154 = n13713 ^ n9456 ^ 1'b0 ;
  assign n18155 = n12486 | n12830 ;
  assign n18156 = n5235 & ~n18155 ;
  assign n18157 = n13972 ^ n340 ^ 1'b0 ;
  assign n18158 = n4811 & n18157 ;
  assign n18159 = n2484 | n2759 ;
  assign n18160 = n18159 ^ n3826 ^ 1'b0 ;
  assign n18161 = n2711 & n8795 ;
  assign n18162 = ~n18160 & n18161 ;
  assign n18163 = n5337 ^ n4144 ^ 1'b0 ;
  assign n18164 = n7563 & n18163 ;
  assign n18165 = n6962 & n8725 ;
  assign n18166 = ~n1491 & n11961 ;
  assign n18167 = n18165 & n18166 ;
  assign n18168 = n4643 & ~n10629 ;
  assign n18169 = n4970 & n6549 ;
  assign n18170 = ~n18168 & n18169 ;
  assign n18171 = n18170 ^ n16612 ^ 1'b0 ;
  assign n18172 = n9292 & n18171 ;
  assign n18173 = n18172 ^ n3030 ^ 1'b0 ;
  assign n18174 = n11927 | n13096 ;
  assign n18175 = n4032 ^ n1632 ^ 1'b0 ;
  assign n18176 = ~n6482 & n8059 ;
  assign n18177 = ~n18175 & n18176 ;
  assign n18178 = n18177 ^ n17077 ^ n6541 ;
  assign n18179 = n5634 & ~n7271 ;
  assign n18180 = n18179 ^ n4555 ^ 1'b0 ;
  assign n18181 = n731 | n9220 ;
  assign n18182 = n8407 & ~n18181 ;
  assign n18183 = n10696 | n18182 ;
  assign n18184 = n2385 | n18183 ;
  assign n18185 = n358 ^ x109 ^ 1'b0 ;
  assign n18186 = ~n8087 & n18185 ;
  assign n18187 = n18186 ^ n4013 ^ 1'b0 ;
  assign n18188 = n574 & n2068 ;
  assign n18189 = n4589 & n18188 ;
  assign n18190 = n18189 ^ n4720 ^ 1'b0 ;
  assign n18191 = ~n16324 & n18190 ;
  assign n18192 = n185 & n3938 ;
  assign n18193 = n12304 & n14186 ;
  assign n18194 = n13063 ^ n11648 ^ 1'b0 ;
  assign n18195 = n4213 | n14157 ;
  assign n18196 = n18195 ^ n4232 ^ 1'b0 ;
  assign n18197 = ( ~n2440 & n4434 ) | ( ~n2440 & n17089 ) | ( n4434 & n17089 ) ;
  assign n18198 = n8918 ^ n5622 ^ 1'b0 ;
  assign n18199 = n3805 | n18198 ;
  assign n18200 = n18199 ^ n8136 ^ 1'b0 ;
  assign n18201 = n8958 & n18200 ;
  assign n18202 = n18201 ^ n1401 ^ 1'b0 ;
  assign n18203 = ~n15353 & n18202 ;
  assign n18204 = n11601 ^ n11111 ^ 1'b0 ;
  assign n18205 = n2355 & n6256 ;
  assign n18206 = ~n446 & n13092 ;
  assign n18207 = ~n16369 & n18206 ;
  assign n18208 = n18207 ^ n1037 ^ 1'b0 ;
  assign n18209 = ~n9480 & n12001 ;
  assign n18210 = n3271 | n8095 ;
  assign n18211 = ~n13444 & n18168 ;
  assign n18212 = n724 & n18211 ;
  assign n18213 = n6266 ^ n2085 ^ 1'b0 ;
  assign n18214 = ~n6423 & n18213 ;
  assign n18215 = n18214 ^ n6027 ^ 1'b0 ;
  assign n18216 = ~n1064 & n2404 ;
  assign n18217 = ~n14355 & n18216 ;
  assign n18218 = x101 & n18217 ;
  assign n18219 = n18215 & n18218 ;
  assign n18220 = ~n8170 & n8316 ;
  assign n18221 = ~n7617 & n18220 ;
  assign n18222 = ~n10526 & n15303 ;
  assign n18223 = n408 & ~n3130 ;
  assign n18224 = n17010 & ~n18223 ;
  assign n18226 = n13503 ^ n1477 ^ 1'b0 ;
  assign n18227 = n13676 & n18226 ;
  assign n18225 = n4005 & n6575 ;
  assign n18228 = n18227 ^ n18225 ^ n16177 ;
  assign n18229 = n17255 ^ n16295 ^ 1'b0 ;
  assign n18230 = ~n2988 & n18229 ;
  assign n18231 = n11062 ^ n830 ^ 1'b0 ;
  assign n18232 = n3853 ^ n2675 ^ 1'b0 ;
  assign n18233 = n12062 ^ n6051 ^ 1'b0 ;
  assign n18234 = n15652 ^ n6862 ^ n277 ;
  assign n18235 = n18233 & n18234 ;
  assign n18236 = ~n5895 & n18235 ;
  assign n18237 = n387 & n9843 ;
  assign n18238 = n8717 & n18237 ;
  assign n18239 = n14497 ^ n1069 ^ 1'b0 ;
  assign n18240 = n7203 & ~n18239 ;
  assign n18241 = n5464 | n18240 ;
  assign n18243 = n3818 & ~n10498 ;
  assign n18242 = n6167 ^ n2385 ^ n652 ;
  assign n18244 = n18243 ^ n18242 ^ n8803 ;
  assign n18245 = n9779 ^ x125 ^ 1'b0 ;
  assign n18246 = n7664 & ~n10818 ;
  assign n18247 = n1784 & ~n4061 ;
  assign n18248 = n18247 ^ n3312 ^ 1'b0 ;
  assign n18249 = n14950 & n18248 ;
  assign n18250 = n3620 ^ n3271 ^ 1'b0 ;
  assign n18251 = n1821 & ~n18250 ;
  assign n18252 = n18249 & ~n18251 ;
  assign n18253 = n4991 & ~n14370 ;
  assign n18254 = ~x101 & n18253 ;
  assign n18255 = n6918 | n18254 ;
  assign n18256 = n6311 | n18255 ;
  assign n18257 = x18 & n928 ;
  assign n18258 = ~n18256 & n18257 ;
  assign n18259 = ~n3057 & n16203 ;
  assign n18260 = n7617 & ~n15244 ;
  assign n18261 = n1618 & ~n12417 ;
  assign n18262 = n784 | n8210 ;
  assign n18263 = n18262 ^ n926 ^ 1'b0 ;
  assign n18264 = n18263 ^ n5432 ^ 1'b0 ;
  assign n18265 = ~n14804 & n18264 ;
  assign n18266 = n8767 & ~n11882 ;
  assign n18267 = n9310 & ~n18266 ;
  assign n18268 = ~n332 & n18267 ;
  assign n18269 = ( n2392 & n9712 ) | ( n2392 & n11039 ) | ( n9712 & n11039 ) ;
  assign n18270 = n10551 | n18269 ;
  assign n18271 = n870 | n1020 ;
  assign n18272 = n18271 ^ n13466 ^ 1'b0 ;
  assign n18274 = n3242 & ~n12892 ;
  assign n18275 = n1632 & ~n3602 ;
  assign n18276 = ~n18274 & n18275 ;
  assign n18273 = n8314 & ~n11426 ;
  assign n18277 = n18276 ^ n18273 ^ 1'b0 ;
  assign n18278 = n7744 ^ n2821 ^ 1'b0 ;
  assign n18279 = ~n5259 & n18278 ;
  assign n18280 = n18279 ^ n9213 ^ 1'b0 ;
  assign n18281 = n4664 | n4749 ;
  assign n18282 = ( n2650 & ~n7009 ) | ( n2650 & n18281 ) | ( ~n7009 & n18281 ) ;
  assign n18283 = n13429 ^ n6457 ^ 1'b0 ;
  assign n18284 = ~n3453 & n18283 ;
  assign n18285 = n3212 & n18284 ;
  assign n18286 = n15596 ^ n7724 ^ 1'b0 ;
  assign n18287 = n999 ^ x73 ^ 1'b0 ;
  assign n18288 = ~n2809 & n18287 ;
  assign n18289 = n16761 ^ n4671 ^ 1'b0 ;
  assign n18290 = n18288 & ~n18289 ;
  assign n18291 = n5258 & ~n7085 ;
  assign n18292 = n3302 & n18291 ;
  assign n18293 = n6957 | n18292 ;
  assign n18294 = n1422 | n18293 ;
  assign n18295 = n4376 | n14761 ;
  assign n18296 = n2144 & n3591 ;
  assign n18297 = n2994 ^ n1530 ^ 1'b0 ;
  assign n18298 = n942 & ~n18297 ;
  assign n18299 = n18298 ^ n4233 ^ 1'b0 ;
  assign n18300 = n10264 ^ n4523 ^ 1'b0 ;
  assign n18301 = n4819 & ~n18300 ;
  assign n18302 = n6215 | n14618 ;
  assign n18303 = n4878 & ~n18302 ;
  assign n18304 = n18303 ^ n11768 ^ 1'b0 ;
  assign n18305 = ~n784 & n9088 ;
  assign n18306 = ~n6841 & n18305 ;
  assign n18307 = ~n10696 & n13321 ;
  assign n18308 = n18307 ^ n2371 ^ 1'b0 ;
  assign n18309 = n4375 & n18308 ;
  assign n18310 = ~n4093 & n18309 ;
  assign n18312 = n2523 | n16292 ;
  assign n18311 = n2943 | n5165 ;
  assign n18313 = n18312 ^ n18311 ^ 1'b0 ;
  assign n18314 = n7134 | n11228 ;
  assign n18315 = ~n3950 & n6474 ;
  assign n18316 = n18315 ^ n8095 ^ 1'b0 ;
  assign n18317 = n18316 ^ n6723 ^ n650 ;
  assign n18318 = n2873 & ~n9239 ;
  assign n18319 = n5984 & n18318 ;
  assign n18320 = n8987 & n18319 ;
  assign n18321 = n5904 ^ n3307 ^ 1'b0 ;
  assign n18322 = ~n9192 & n18321 ;
  assign n18323 = n18322 ^ n14618 ^ 1'b0 ;
  assign n18324 = n3246 & ~n18323 ;
  assign n18325 = n18324 ^ n5007 ^ 1'b0 ;
  assign n18326 = n13290 ^ n8506 ^ 1'b0 ;
  assign n18327 = n18325 & ~n18326 ;
  assign n18328 = n2944 | n9075 ;
  assign n18329 = n3462 & ~n6638 ;
  assign n18330 = n1744 & ~n9253 ;
  assign n18331 = n1181 | n18330 ;
  assign n18332 = ( n1905 & n6221 ) | ( n1905 & ~n18331 ) | ( n6221 & ~n18331 ) ;
  assign n18333 = n11309 ^ n974 ^ 1'b0 ;
  assign n18334 = n14872 ^ n1854 ^ 1'b0 ;
  assign n18335 = n14124 ^ n911 ^ 1'b0 ;
  assign n18336 = n7829 & ~n18335 ;
  assign n18337 = n8161 ^ n5120 ^ 1'b0 ;
  assign n18338 = ~n17889 & n18337 ;
  assign n18339 = ~n1060 & n18338 ;
  assign n18340 = n2818 | n9399 ;
  assign n18341 = n1329 & n5038 ;
  assign n18342 = n18341 ^ n9293 ^ 1'b0 ;
  assign n18343 = ~n2948 & n14902 ;
  assign n18344 = ~n1536 & n18343 ;
  assign n18345 = ~n12357 & n18344 ;
  assign n18346 = ~n11148 & n13632 ;
  assign n18347 = n18346 ^ n2591 ^ 1'b0 ;
  assign n18348 = n3415 | n18347 ;
  assign n18349 = n5195 & ~n7654 ;
  assign n18350 = ~n4791 & n5273 ;
  assign n18351 = ~n5273 & n18350 ;
  assign n18352 = n13331 | n18351 ;
  assign n18353 = n18351 & ~n18352 ;
  assign n18354 = n2193 ^ n974 ^ 1'b0 ;
  assign n18355 = n4346 & n18354 ;
  assign n18356 = n4998 & n18355 ;
  assign n18357 = ~n2179 & n18356 ;
  assign n18358 = n8930 ^ n4496 ^ 1'b0 ;
  assign n18359 = n2701 ^ n669 ^ 1'b0 ;
  assign n18360 = n18359 ^ n5115 ^ x23 ;
  assign n18361 = n9832 & n12011 ;
  assign n18362 = n3320 & n9258 ;
  assign n18363 = n330 & ~n18362 ;
  assign n18364 = n18363 ^ n1491 ^ 1'b0 ;
  assign n18366 = n3400 & ~n3848 ;
  assign n18367 = n18366 ^ n7595 ^ 1'b0 ;
  assign n18365 = n5749 & n6313 ;
  assign n18368 = n18367 ^ n18365 ^ 1'b0 ;
  assign n18369 = n3953 | n15232 ;
  assign n18372 = n2478 | n6864 ;
  assign n18373 = n2478 & ~n18372 ;
  assign n18374 = n3751 | n18373 ;
  assign n18375 = n3751 & ~n18374 ;
  assign n18370 = n15894 ^ n5903 ^ 1'b0 ;
  assign n18371 = n5046 | n18370 ;
  assign n18376 = n18375 ^ n18371 ^ n6921 ;
  assign n18377 = n3446 | n7232 ;
  assign n18378 = n18377 ^ n13649 ^ 1'b0 ;
  assign n18379 = n8945 | n10476 ;
  assign n18380 = n18379 ^ n444 ^ 1'b0 ;
  assign n18381 = ~n1762 & n2330 ;
  assign n18382 = ~n9174 & n18381 ;
  assign n18383 = n8713 ^ n8107 ^ 1'b0 ;
  assign n18384 = n3833 & ~n4976 ;
  assign n18385 = n18384 ^ n14074 ^ 1'b0 ;
  assign n18386 = n1665 & n18385 ;
  assign n18387 = n10010 | n14913 ;
  assign n18388 = n3527 | n18387 ;
  assign n18389 = n11128 & n18388 ;
  assign n18390 = ~n7569 & n18389 ;
  assign n18391 = n13921 ^ n7760 ^ 1'b0 ;
  assign n18392 = n9981 | n18391 ;
  assign n18393 = n4573 & ~n18392 ;
  assign n18394 = n12769 & ~n18393 ;
  assign n18395 = n18394 ^ n4457 ^ 1'b0 ;
  assign n18396 = ( x39 & n2539 ) | ( x39 & ~n4306 ) | ( n2539 & ~n4306 ) ;
  assign n18397 = n13554 & ~n18396 ;
  assign n18398 = n7467 ^ n7245 ^ n1651 ;
  assign n18399 = ~x68 & n2062 ;
  assign n18400 = n18399 ^ n2469 ^ 1'b0 ;
  assign n18401 = n18400 ^ n3422 ^ 1'b0 ;
  assign n18402 = n894 ^ n430 ^ 1'b0 ;
  assign n18403 = n17039 & n18402 ;
  assign n18404 = n15986 & ~n18403 ;
  assign n18405 = n4047 ^ n1064 ^ 1'b0 ;
  assign n18406 = n5759 & n18405 ;
  assign n18407 = n9500 ^ n6735 ^ 1'b0 ;
  assign n18408 = n2087 | n18407 ;
  assign n18409 = n2428 | n6393 ;
  assign n18410 = n18409 ^ n8699 ^ 1'b0 ;
  assign n18411 = n14391 ^ n8722 ^ 1'b0 ;
  assign n18412 = n12272 | n18411 ;
  assign n18413 = n8617 ^ n3454 ^ 1'b0 ;
  assign n18414 = ~n4480 & n9489 ;
  assign n18415 = n16509 & n18414 ;
  assign n18416 = n1264 & ~n11995 ;
  assign n18417 = n18416 ^ n1010 ^ 1'b0 ;
  assign n18418 = n1401 ^ n335 ^ 1'b0 ;
  assign n18419 = ~n18417 & n18418 ;
  assign n18420 = n13656 & n18419 ;
  assign n18421 = ~n13831 & n18420 ;
  assign n18424 = n150 | n911 ;
  assign n18422 = n6325 ^ n6241 ^ 1'b0 ;
  assign n18423 = n414 & n18422 ;
  assign n18425 = n18424 ^ n18423 ^ n8047 ;
  assign n18426 = n629 & ~n3772 ;
  assign n18427 = n5898 ^ n3591 ^ 1'b0 ;
  assign n18428 = n18426 & n18427 ;
  assign n18429 = n10780 ^ n9235 ^ 1'b0 ;
  assign n18430 = n5469 & ~n8694 ;
  assign n18431 = ~n13168 & n16411 ;
  assign n18432 = n18430 & ~n18431 ;
  assign n18433 = n18432 ^ n238 ^ 1'b0 ;
  assign n18436 = n13716 ^ n13356 ^ 1'b0 ;
  assign n18434 = ~n11880 & n12324 ;
  assign n18435 = n18434 ^ n5953 ^ 1'b0 ;
  assign n18437 = n18436 ^ n18435 ^ n6934 ;
  assign n18438 = ~n11072 & n15898 ;
  assign n18439 = n4047 | n9662 ;
  assign n18440 = n6064 | n18439 ;
  assign n18441 = n18440 ^ n17050 ^ 1'b0 ;
  assign n18442 = n2570 | n17907 ;
  assign n18443 = n3445 & n14179 ;
  assign n18444 = n5902 ^ x108 ^ 1'b0 ;
  assign n18445 = ~n18417 & n18444 ;
  assign n18446 = n7484 & ~n16890 ;
  assign n18447 = n6325 ^ n1395 ^ 1'b0 ;
  assign n18448 = n11915 | n18447 ;
  assign n18449 = n1224 & ~n15581 ;
  assign n18450 = ~n1754 & n7133 ;
  assign n18451 = n18450 ^ n8823 ^ 1'b0 ;
  assign n18452 = n18451 ^ n7211 ^ 1'b0 ;
  assign n18453 = ( n1829 & n4143 ) | ( n1829 & n9351 ) | ( n4143 & n9351 ) ;
  assign n18454 = ( n1510 & ~n15611 ) | ( n1510 & n18453 ) | ( ~n15611 & n18453 ) ;
  assign n18455 = ( n5137 & n14211 ) | ( n5137 & ~n18454 ) | ( n14211 & ~n18454 ) ;
  assign n18456 = n2263 ^ n890 ^ 1'b0 ;
  assign n18457 = n11516 | n18456 ;
  assign n18458 = ~n8994 & n10493 ;
  assign n18459 = n1161 | n7624 ;
  assign n18460 = n18459 ^ n8476 ^ 1'b0 ;
  assign n18461 = n17140 ^ n8270 ^ 1'b0 ;
  assign n18462 = n14868 ^ n2977 ^ 1'b0 ;
  assign n18463 = n1274 | n18462 ;
  assign n18464 = n2707 ^ n1839 ^ 1'b0 ;
  assign n18465 = ~n1349 & n18464 ;
  assign n18466 = n18465 ^ n6817 ^ 1'b0 ;
  assign n18467 = n12553 & n18466 ;
  assign n18468 = n3622 ^ n984 ^ 1'b0 ;
  assign n18469 = n1825 | n18468 ;
  assign n18470 = n3034 & n4215 ;
  assign n18471 = n9675 ^ n1529 ^ 1'b0 ;
  assign n18472 = n9660 & ~n18471 ;
  assign n18473 = n18470 & n18472 ;
  assign n18474 = n15650 ^ n4935 ^ 1'b0 ;
  assign n18475 = n18474 ^ n547 ^ 1'b0 ;
  assign n18476 = n9175 ^ n1436 ^ 1'b0 ;
  assign n18477 = x121 & n18476 ;
  assign n18478 = n756 & n3382 ;
  assign n18479 = n15737 | n16276 ;
  assign n18480 = n18478 & ~n18479 ;
  assign n18481 = n4098 & ~n10334 ;
  assign n18482 = n5440 & ~n6244 ;
  assign n18483 = n18482 ^ n5426 ^ 1'b0 ;
  assign n18484 = n11344 ^ n10126 ^ 1'b0 ;
  assign n18485 = ~n3838 & n5036 ;
  assign n18486 = n3300 | n7715 ;
  assign n18487 = n18486 ^ n3253 ^ 1'b0 ;
  assign n18488 = ~n5766 & n7275 ;
  assign n18489 = n2091 & n18488 ;
  assign n18490 = n11705 ^ n5123 ^ 1'b0 ;
  assign n18491 = n378 & ~n4014 ;
  assign n18492 = n18491 ^ n2839 ^ 1'b0 ;
  assign n18493 = n696 | n1052 ;
  assign n18494 = ~n11959 & n12525 ;
  assign n18495 = n7130 & ~n15522 ;
  assign n18496 = n18495 ^ n9483 ^ 1'b0 ;
  assign n18497 = n15802 ^ n6576 ^ 1'b0 ;
  assign n18498 = n8093 & ~n16192 ;
  assign n18499 = ~n757 & n2750 ;
  assign n18500 = n14578 ^ n7364 ^ 1'b0 ;
  assign n18501 = n18499 & ~n18500 ;
  assign n18502 = n18501 ^ n4753 ^ 1'b0 ;
  assign n18503 = n18502 ^ n8947 ^ 1'b0 ;
  assign n18504 = n17525 & ~n18503 ;
  assign n18505 = n7545 & ~n13559 ;
  assign n18506 = n8170 & n15795 ;
  assign n18507 = n1443 & n7433 ;
  assign n18508 = ~n11875 & n18507 ;
  assign n18509 = n5929 | n6391 ;
  assign n18510 = n18509 ^ n16865 ^ 1'b0 ;
  assign n18511 = n18508 | n18510 ;
  assign n18512 = n3730 & ~n11022 ;
  assign n18513 = n15951 & ~n18512 ;
  assign n18514 = n18513 ^ n16077 ^ 1'b0 ;
  assign n18515 = n11044 & n13636 ;
  assign n18516 = n18515 ^ n1786 ^ 1'b0 ;
  assign n18517 = n502 & ~n18516 ;
  assign n18518 = n3899 & ~n7597 ;
  assign n18519 = ~n5388 & n16038 ;
  assign n18520 = n4086 & ~n12825 ;
  assign n18521 = n9904 & n17747 ;
  assign n18522 = ~n6722 & n18521 ;
  assign n18523 = n1539 & n3629 ;
  assign n18524 = n18523 ^ n17055 ^ 1'b0 ;
  assign n18525 = n1788 ^ x104 ^ 1'b0 ;
  assign n18526 = n10607 ^ n6575 ^ 1'b0 ;
  assign n18527 = x23 & n18526 ;
  assign n18528 = ~n2658 & n7810 ;
  assign n18529 = n8945 ^ n2738 ^ 1'b0 ;
  assign n18530 = n12768 & ~n18529 ;
  assign n18531 = n2323 & ~n2664 ;
  assign n18532 = n10856 | n18531 ;
  assign n18533 = n4832 | n18532 ;
  assign n18534 = n9326 | n16947 ;
  assign n18535 = n18534 ^ n11405 ^ 1'b0 ;
  assign n18536 = n3031 ^ n2675 ^ 1'b0 ;
  assign n18537 = n1768 | n18536 ;
  assign n18538 = n1387 & n6575 ;
  assign n18539 = n571 & ~n5749 ;
  assign n18540 = n18539 ^ n11827 ^ 1'b0 ;
  assign n18541 = n5273 & n17651 ;
  assign n18542 = ~n11295 & n18541 ;
  assign n18543 = n1329 | n1344 ;
  assign n18544 = n18543 ^ x87 ^ 1'b0 ;
  assign n18545 = n18544 ^ n4388 ^ 1'b0 ;
  assign n18546 = n5358 ^ n3558 ^ 1'b0 ;
  assign n18547 = n18545 & n18546 ;
  assign n18548 = n9551 | n18547 ;
  assign n18549 = n5962 & n18284 ;
  assign n18550 = ~n5340 & n18549 ;
  assign n18551 = n18550 ^ n7381 ^ 1'b0 ;
  assign n18552 = n5151 ^ n528 ^ 1'b0 ;
  assign n18553 = x95 & n998 ;
  assign n18554 = n18553 ^ n8662 ^ 1'b0 ;
  assign n18555 = n17831 ^ n3714 ^ n3615 ;
  assign n18556 = n9934 ^ n3281 ^ 1'b0 ;
  assign n18557 = ~n7222 & n18556 ;
  assign n18558 = n14228 & n18557 ;
  assign n18559 = n15899 ^ n4371 ^ 1'b0 ;
  assign n18560 = ~n198 & n8889 ;
  assign n18561 = n15854 ^ n5099 ^ 1'b0 ;
  assign n18562 = ~n2086 & n6284 ;
  assign n18563 = n9176 | n16217 ;
  assign n18564 = n10535 ^ n841 ^ 1'b0 ;
  assign n18565 = n13198 ^ n5632 ^ 1'b0 ;
  assign n18566 = n6916 & n18565 ;
  assign n18567 = n15889 ^ n9091 ^ 1'b0 ;
  assign n18568 = n1447 & ~n18567 ;
  assign n18569 = n18568 ^ n7626 ^ 1'b0 ;
  assign n18574 = n7466 & ~n14517 ;
  assign n18570 = n2775 & n7572 ;
  assign n18571 = n18570 ^ n18416 ^ 1'b0 ;
  assign n18572 = n18571 ^ n15543 ^ 1'b0 ;
  assign n18573 = ~n7100 & n18572 ;
  assign n18575 = n18574 ^ n18573 ^ 1'b0 ;
  assign n18576 = n1788 & n18575 ;
  assign n18577 = n16459 ^ n6267 ^ 1'b0 ;
  assign n18578 = n10864 & ~n18577 ;
  assign n18579 = ~n4819 & n18578 ;
  assign n18580 = n8057 ^ n3338 ^ 1'b0 ;
  assign n18581 = n7486 & ~n18580 ;
  assign n18582 = n11820 ^ n11474 ^ 1'b0 ;
  assign n18587 = n3142 & n7174 ;
  assign n18586 = n3712 & n4040 ;
  assign n18588 = n18587 ^ n18586 ^ 1'b0 ;
  assign n18583 = n10903 ^ n6228 ^ 1'b0 ;
  assign n18584 = n256 & ~n18583 ;
  assign n18585 = n11635 & n18584 ;
  assign n18589 = n18588 ^ n18585 ^ 1'b0 ;
  assign n18590 = n7601 & ~n10633 ;
  assign n18591 = n14610 ^ n8738 ^ 1'b0 ;
  assign n18592 = n1230 & n18591 ;
  assign n18593 = n16251 ^ n7421 ^ 1'b0 ;
  assign n18594 = ~n1979 & n18593 ;
  assign n18595 = n8016 ^ n4067 ^ 1'b0 ;
  assign n18596 = n1079 ^ n387 ^ 1'b0 ;
  assign n18597 = n1015 & ~n15948 ;
  assign n18598 = n18597 ^ n15625 ^ 1'b0 ;
  assign n18599 = n2958 & n18598 ;
  assign n18600 = n3364 & ~n18599 ;
  assign n18601 = n450 & ~n3196 ;
  assign n18602 = n18601 ^ n3662 ^ 1'b0 ;
  assign n18603 = x119 | n14517 ;
  assign n18604 = n18603 ^ n8015 ^ 1'b0 ;
  assign n18605 = ~n18602 & n18604 ;
  assign n18606 = n6501 ^ n813 ^ 1'b0 ;
  assign n18607 = n5613 | n18606 ;
  assign n18608 = n8273 ^ n5253 ^ 1'b0 ;
  assign n18609 = n1245 & ~n18608 ;
  assign n18610 = n6369 ^ n1519 ^ 1'b0 ;
  assign n18611 = n14383 & n18610 ;
  assign n18612 = n9145 & ~n18611 ;
  assign n18613 = n14427 & ~n16690 ;
  assign n18614 = n1147 & ~n10352 ;
  assign n18615 = n5546 ^ n1420 ^ 1'b0 ;
  assign n18616 = n1552 & n18615 ;
  assign n18617 = n18616 ^ n13636 ^ n4172 ;
  assign n18618 = n4141 | n10086 ;
  assign n18619 = n10184 & n18618 ;
  assign n18620 = n7100 ^ n717 ^ 1'b0 ;
  assign n18621 = ~n8302 & n18620 ;
  assign n18622 = ~n2394 & n4835 ;
  assign n18623 = n18622 ^ n10143 ^ 1'b0 ;
  assign n18624 = n13285 ^ n1304 ^ 1'b0 ;
  assign n18625 = n1736 & ~n2739 ;
  assign n18626 = n16822 ^ n5976 ^ 1'b0 ;
  assign n18627 = ~n502 & n3575 ;
  assign n18628 = n18627 ^ n2858 ^ 1'b0 ;
  assign n18629 = n18628 ^ n3401 ^ 1'b0 ;
  assign n18630 = n18629 ^ n15032 ^ 1'b0 ;
  assign n18631 = ~n12164 & n13835 ;
  assign n18632 = n18631 ^ n1133 ^ 1'b0 ;
  assign n18633 = n18632 ^ n9305 ^ 1'b0 ;
  assign n18634 = n4551 & ~n11834 ;
  assign n18635 = n18634 ^ n882 ^ 1'b0 ;
  assign n18636 = n3651 & ~n18635 ;
  assign n18639 = n2037 & ~n13670 ;
  assign n18637 = n4296 ^ n1805 ^ 1'b0 ;
  assign n18638 = ~x123 & n18637 ;
  assign n18640 = n18639 ^ n18638 ^ 1'b0 ;
  assign n18641 = n1724 | n18640 ;
  assign n18642 = n18636 & ~n18641 ;
  assign n18643 = n13902 ^ n6956 ^ 1'b0 ;
  assign n18645 = n499 & n7037 ;
  assign n18644 = ~n5876 & n9107 ;
  assign n18646 = n18645 ^ n18644 ^ 1'b0 ;
  assign n18647 = n6011 ^ n4521 ^ 1'b0 ;
  assign n18648 = n2264 & n18647 ;
  assign n18649 = ~n3751 & n12322 ;
  assign n18650 = n18649 ^ n12908 ^ n12734 ;
  assign n18651 = n8398 | n18650 ;
  assign n18652 = x105 | n9848 ;
  assign n18653 = ( n8095 & n18651 ) | ( n8095 & n18652 ) | ( n18651 & n18652 ) ;
  assign n18654 = n18653 ^ n15621 ^ 1'b0 ;
  assign n18655 = x7 & n18654 ;
  assign n18656 = n16194 ^ n8392 ^ 1'b0 ;
  assign n18657 = n2594 & n18247 ;
  assign n18658 = n10932 ^ n5987 ^ 1'b0 ;
  assign n18659 = n5347 ^ n305 ^ 1'b0 ;
  assign n18660 = ~n8442 & n18659 ;
  assign n18661 = ( n4241 & ~n5148 ) | ( n4241 & n15316 ) | ( ~n5148 & n15316 ) ;
  assign n18662 = n17674 & n18661 ;
  assign n18663 = n4746 & n12604 ;
  assign n18664 = n7272 & n13275 ;
  assign n18665 = n18664 ^ n11241 ^ 1'b0 ;
  assign n18666 = n18663 | n18665 ;
  assign n18667 = n9899 ^ n8050 ^ 1'b0 ;
  assign n18668 = ~n3195 & n4572 ;
  assign n18669 = n4828 | n18668 ;
  assign n18670 = n2880 & n5268 ;
  assign n18671 = n2335 & n18670 ;
  assign n18672 = n10292 & n14760 ;
  assign n18673 = n3286 & n10985 ;
  assign n18674 = n18673 ^ n13948 ^ 1'b0 ;
  assign n18675 = n3925 & n4578 ;
  assign n18676 = n18675 ^ x10 ^ 1'b0 ;
  assign n18677 = n3949 ^ n735 ^ 1'b0 ;
  assign n18678 = n16778 & n18677 ;
  assign n18679 = n8724 & n18678 ;
  assign n18682 = n6473 & ~n16673 ;
  assign n18683 = n18682 ^ n11387 ^ 1'b0 ;
  assign n18684 = n6268 | n18683 ;
  assign n18685 = n3272 | n18684 ;
  assign n18686 = ~n7933 & n18247 ;
  assign n18687 = ~n18685 & n18686 ;
  assign n18680 = n3608 ^ n3087 ^ 1'b0 ;
  assign n18681 = ~n10869 & n18680 ;
  assign n18688 = n18687 ^ n18681 ^ 1'b0 ;
  assign n18689 = n576 | n15697 ;
  assign n18690 = n11344 & ~n18689 ;
  assign n18691 = n10151 & ~n18690 ;
  assign n18692 = n18691 ^ n5683 ^ 1'b0 ;
  assign n18693 = n6607 ^ n2233 ^ 1'b0 ;
  assign n18694 = n7997 & n11218 ;
  assign n18695 = n18694 ^ n11108 ^ 1'b0 ;
  assign n18696 = n18695 ^ n562 ^ 1'b0 ;
  assign n18697 = n2043 & n3362 ;
  assign n18698 = n2529 & n18697 ;
  assign n18699 = n9725 & ~n17954 ;
  assign n18700 = n15937 ^ n4212 ^ 1'b0 ;
  assign n18701 = n17513 ^ n11030 ^ 1'b0 ;
  assign n18702 = n15795 ^ n5039 ^ 1'b0 ;
  assign n18703 = ~n3831 & n16075 ;
  assign n18704 = n12047 & n18703 ;
  assign n18705 = n4300 | n15873 ;
  assign n18706 = n5669 | n18705 ;
  assign n18707 = n5532 | n14599 ;
  assign n18708 = n18707 ^ n11032 ^ 1'b0 ;
  assign n18709 = n15419 & ~n16274 ;
  assign n18710 = n8709 & n10562 ;
  assign n18711 = n8280 & n18710 ;
  assign n18712 = n18711 ^ n3038 ^ 1'b0 ;
  assign n18713 = n7513 | n18712 ;
  assign n18714 = n15113 | n15322 ;
  assign n18715 = n3138 ^ n420 ^ 1'b0 ;
  assign n18716 = n12736 ^ n5720 ^ 1'b0 ;
  assign n18717 = ~n2732 & n18716 ;
  assign n18718 = n2398 ^ n984 ^ 1'b0 ;
  assign n18719 = n18717 & ~n18718 ;
  assign n18720 = ~n201 & n16655 ;
  assign n18721 = ~n1604 & n12769 ;
  assign n18722 = n18721 ^ n11445 ^ 1'b0 ;
  assign n18723 = n13996 ^ n7770 ^ 1'b0 ;
  assign n18724 = ~n5741 & n6064 ;
  assign n18725 = ( n9689 & n10145 ) | ( n9689 & ~n18724 ) | ( n10145 & ~n18724 ) ;
  assign n18726 = x22 & n7465 ;
  assign n18727 = n11563 & ~n18726 ;
  assign n18728 = ~n2472 & n5108 ;
  assign n18729 = n13655 ^ n8343 ^ 1'b0 ;
  assign n18730 = n18729 ^ n11052 ^ 1'b0 ;
  assign n18731 = n18728 | n18730 ;
  assign n18732 = n4224 | n10438 ;
  assign n18733 = n503 & ~n8723 ;
  assign n18734 = n18733 ^ n14031 ^ 1'b0 ;
  assign n18735 = n18734 ^ n5039 ^ 1'b0 ;
  assign n18736 = n3458 & n18735 ;
  assign n18738 = n3804 ^ n2222 ^ 1'b0 ;
  assign n18739 = n3748 & n18738 ;
  assign n18737 = n8940 | n13033 ;
  assign n18740 = n18739 ^ n18737 ^ 1'b0 ;
  assign n18741 = ~n18599 & n18740 ;
  assign n18742 = n6590 ^ n930 ^ 1'b0 ;
  assign n18743 = n1423 | n7004 ;
  assign n18744 = n2219 & ~n18743 ;
  assign n18745 = n11399 & n13333 ;
  assign n18746 = ~n8359 & n18745 ;
  assign n18747 = n512 & ~n14755 ;
  assign n18748 = n2323 & n8655 ;
  assign n18749 = n8691 & n18748 ;
  assign n18750 = ~n3917 & n18749 ;
  assign n18751 = n10868 & ~n14129 ;
  assign n18752 = n18751 ^ n570 ^ 1'b0 ;
  assign n18753 = n1984 & n10597 ;
  assign n18754 = ~n10338 & n18753 ;
  assign n18755 = n18754 ^ n1124 ^ 1'b0 ;
  assign n18756 = n16438 ^ n277 ^ 1'b0 ;
  assign n18757 = n1945 | n18756 ;
  assign n18758 = n18757 ^ n14861 ^ 1'b0 ;
  assign n18759 = n1170 & n5924 ;
  assign n18760 = n9103 & n13279 ;
  assign n18761 = n18760 ^ n16314 ^ 1'b0 ;
  assign n18762 = n252 & n18761 ;
  assign n18763 = n1114 | n15697 ;
  assign n18764 = n8537 & ~n18763 ;
  assign n18765 = n13731 ^ n5641 ^ 1'b0 ;
  assign n18766 = ~n14229 & n18765 ;
  assign n18767 = n2641 | n8113 ;
  assign n18768 = n18767 ^ n11992 ^ 1'b0 ;
  assign n18769 = ~n9232 & n18768 ;
  assign n18770 = n12473 ^ n11594 ^ 1'b0 ;
  assign n18771 = n1941 | n3292 ;
  assign n18772 = n18770 | n18771 ;
  assign n18773 = n7242 & n12073 ;
  assign n18774 = n7736 & n18773 ;
  assign n18775 = n13936 ^ n482 ^ 1'b0 ;
  assign n18776 = ~x4 & n11057 ;
  assign n18777 = n8005 ^ n1663 ^ 1'b0 ;
  assign n18778 = n10240 | n18777 ;
  assign n18779 = n17161 ^ n15790 ^ n12509 ;
  assign n18780 = ~n1779 & n5525 ;
  assign n18781 = n18780 ^ n13765 ^ 1'b0 ;
  assign n18782 = n18781 ^ n18251 ^ 1'b0 ;
  assign n18783 = n15602 ^ n14755 ^ 1'b0 ;
  assign n18784 = n217 & n1016 ;
  assign n18785 = n18784 ^ n15898 ^ 1'b0 ;
  assign n18786 = n6887 ^ n5606 ^ 1'b0 ;
  assign n18787 = n5050 & n18786 ;
  assign n18788 = n14617 & n18787 ;
  assign n18789 = n3193 | n5243 ;
  assign n18790 = n1051 | n8121 ;
  assign n18791 = n1361 | n3721 ;
  assign n18792 = n5313 ^ n330 ^ 1'b0 ;
  assign n18793 = n1601 & ~n18792 ;
  assign n18794 = n18793 ^ n5885 ^ 1'b0 ;
  assign n18795 = n5708 | n18794 ;
  assign n18796 = n17710 ^ n15488 ^ 1'b0 ;
  assign n18797 = n15720 ^ n2928 ^ 1'b0 ;
  assign n18798 = n12756 ^ n4472 ^ 1'b0 ;
  assign n18799 = n5453 ^ n2037 ^ n984 ;
  assign n18800 = n18799 ^ n16162 ^ 1'b0 ;
  assign n18801 = ~n9130 & n18800 ;
  assign n18802 = n5613 & n7223 ;
  assign n18803 = n18802 ^ n4440 ^ 1'b0 ;
  assign n18804 = ~n1630 & n3422 ;
  assign n18805 = ~n2818 & n18804 ;
  assign n18806 = n2496 ^ n2426 ^ 1'b0 ;
  assign n18807 = n14198 | n15279 ;
  assign n18808 = n18806 | n18807 ;
  assign n18809 = n8917 ^ n4798 ^ 1'b0 ;
  assign n18810 = ~n7905 & n18809 ;
  assign n18811 = ~n8007 & n14852 ;
  assign n18812 = n18811 ^ n1860 ^ 1'b0 ;
  assign n18813 = n4287 & ~n6935 ;
  assign n18814 = n18813 ^ n934 ^ 1'b0 ;
  assign n18815 = n5817 & ~n10383 ;
  assign n18816 = ~n18814 & n18815 ;
  assign n18817 = n3012 & n14831 ;
  assign n18818 = n18817 ^ n13057 ^ 1'b0 ;
  assign n18819 = n11474 & n18818 ;
  assign n18820 = n10498 ^ n8829 ^ 1'b0 ;
  assign n18821 = n7146 ^ n4636 ^ 1'b0 ;
  assign n18822 = n831 | n4185 ;
  assign n18823 = ~n696 & n1170 ;
  assign n18824 = n5023 & n18823 ;
  assign n18825 = n13803 | n18824 ;
  assign n18826 = n18825 ^ n8235 ^ 1'b0 ;
  assign n18827 = n9764 ^ n6070 ^ 1'b0 ;
  assign n18828 = n1816 & ~n13024 ;
  assign n18829 = n1491 & n18828 ;
  assign n18830 = n1784 ^ n1467 ^ 1'b0 ;
  assign n18831 = n10553 | n18830 ;
  assign n18832 = n18831 ^ n5927 ^ 1'b0 ;
  assign n18833 = n5096 ^ n2024 ^ 1'b0 ;
  assign n18834 = n17559 | n18833 ;
  assign n18835 = ( ~n886 & n2107 ) | ( ~n886 & n9876 ) | ( n2107 & n9876 ) ;
  assign n18836 = n8948 ^ n7126 ^ 1'b0 ;
  assign n18837 = n950 & n16629 ;
  assign n18838 = n18836 & n18837 ;
  assign n18839 = n15858 ^ n4337 ^ 1'b0 ;
  assign n18840 = n5709 & ~n17093 ;
  assign n18841 = n17765 & ~n18840 ;
  assign n18842 = n2323 & ~n14900 ;
  assign n18843 = n146 & n7707 ;
  assign n18844 = n10216 & ~n18843 ;
  assign n18845 = n2291 & ~n18844 ;
  assign n18846 = ~n824 & n3195 ;
  assign n18847 = n18846 ^ n13144 ^ n5950 ;
  assign n18848 = n5891 | n17509 ;
  assign n18849 = n18848 ^ n2851 ^ 1'b0 ;
  assign n18850 = n2232 & n2441 ;
  assign n18851 = n18850 ^ n1604 ^ 1'b0 ;
  assign n18852 = n18851 ^ n256 ^ 1'b0 ;
  assign n18853 = ( n5705 & ~n12799 ) | ( n5705 & n18852 ) | ( ~n12799 & n18852 ) ;
  assign n18854 = ~n696 & n7037 ;
  assign n18855 = ~x16 & n18854 ;
  assign n18856 = n2364 & n2684 ;
  assign n18857 = n16576 & n18856 ;
  assign n18858 = n18855 & ~n18857 ;
  assign n18859 = n9628 & n9899 ;
  assign n18860 = n18859 ^ n3080 ^ 1'b0 ;
  assign n18861 = n8985 & ~n18860 ;
  assign n18862 = n2283 & ~n6212 ;
  assign n18863 = n16913 ^ n3744 ^ 1'b0 ;
  assign n18864 = n13549 & n15917 ;
  assign n18865 = ~n15986 & n18864 ;
  assign n18866 = n2941 | n6880 ;
  assign n18867 = n3271 & n16296 ;
  assign n18868 = n8508 & n9787 ;
  assign n18869 = n2582 & n3651 ;
  assign n18870 = n18869 ^ n7847 ^ 1'b0 ;
  assign n18871 = ~n1033 & n1983 ;
  assign n18872 = n897 & n6732 ;
  assign n18873 = n18872 ^ n1714 ^ 1'b0 ;
  assign n18874 = n3108 ^ n790 ^ 1'b0 ;
  assign n18875 = ~n7683 & n18781 ;
  assign n18876 = ~n1887 & n5018 ;
  assign n18877 = ~n18875 & n18876 ;
  assign n18878 = n2122 & n13268 ;
  assign n18879 = n18878 ^ n5007 ^ 1'b0 ;
  assign n18880 = n8028 | n16344 ;
  assign n18881 = n18880 ^ n17879 ^ 1'b0 ;
  assign n18882 = ~n4190 & n18881 ;
  assign n18883 = n12018 & n18882 ;
  assign n18884 = n12815 ^ n391 ^ 1'b0 ;
  assign n18885 = n13294 ^ n1655 ^ 1'b0 ;
  assign n18887 = ~n2905 & n13924 ;
  assign n18886 = n11925 | n11928 ;
  assign n18888 = n18887 ^ n18886 ^ 1'b0 ;
  assign n18889 = n15002 ^ n9761 ^ 1'b0 ;
  assign n18890 = n17097 & ~n18889 ;
  assign n18891 = n2515 & ~n5647 ;
  assign n18892 = n18804 ^ n16882 ^ n7414 ;
  assign n18893 = ~n6813 & n10131 ;
  assign n18894 = n18893 ^ n980 ^ 1'b0 ;
  assign n18895 = n18894 ^ n4025 ^ 1'b0 ;
  assign n18896 = n2601 & n5336 ;
  assign n18897 = n18896 ^ n924 ^ 1'b0 ;
  assign n18898 = n18897 ^ n6596 ^ 1'b0 ;
  assign n18899 = n15039 ^ n1691 ^ 1'b0 ;
  assign n18900 = n3462 & n18899 ;
  assign n18901 = ~n4602 & n18900 ;
  assign n18902 = n1280 ^ n857 ^ 1'b0 ;
  assign n18903 = n18902 ^ n6149 ^ 1'b0 ;
  assign n18904 = ~n16884 & n18903 ;
  assign n18905 = n7104 & n7199 ;
  assign n18906 = ~n1923 & n18905 ;
  assign n18907 = n1576 ^ n397 ^ 1'b0 ;
  assign n18908 = n18907 ^ n7816 ^ 1'b0 ;
  assign n18909 = n11681 ^ n3500 ^ 1'b0 ;
  assign n18910 = n999 ^ x87 ^ 1'b0 ;
  assign n18911 = n7543 ^ n5000 ^ 1'b0 ;
  assign n18912 = n1958 & n18911 ;
  assign n18913 = ( ~n889 & n2943 ) | ( ~n889 & n7055 ) | ( n2943 & n7055 ) ;
  assign n18914 = n12910 ^ n4253 ^ 1'b0 ;
  assign n18915 = n18913 | n18914 ;
  assign n18916 = n5016 | n8494 ;
  assign n18917 = n552 & n17311 ;
  assign n18918 = n6331 ^ n4222 ^ 1'b0 ;
  assign n18919 = n8887 & ~n18918 ;
  assign n18920 = n16573 ^ n2660 ^ 1'b0 ;
  assign n18921 = n18920 ^ n15211 ^ 1'b0 ;
  assign n18922 = x58 | n1304 ;
  assign n18923 = n1351 | n4306 ;
  assign n18924 = n5469 & ~n18923 ;
  assign n18925 = n3721 & ~n18924 ;
  assign n18926 = n18925 ^ n17641 ^ 1'b0 ;
  assign n18927 = n6064 & n13317 ;
  assign n18928 = ~n2178 & n18927 ;
  assign n18929 = n949 & ~n1918 ;
  assign n18930 = n7523 ^ n2087 ^ 1'b0 ;
  assign n18931 = n18930 ^ n2959 ^ 1'b0 ;
  assign n18933 = n1169 & ~n7742 ;
  assign n18932 = n6034 & ~n15148 ;
  assign n18934 = n18933 ^ n18932 ^ 1'b0 ;
  assign n18935 = n2505 & ~n2757 ;
  assign n18936 = n18935 ^ n12245 ^ 1'b0 ;
  assign n18937 = n5801 & ~n6514 ;
  assign n18938 = ~n11911 & n18937 ;
  assign n18939 = n18938 ^ n5166 ^ n371 ;
  assign n18940 = ~n18936 & n18939 ;
  assign n18941 = ~n10726 & n18940 ;
  assign n18942 = ( n4065 & n6003 ) | ( n4065 & ~n13629 ) | ( n6003 & ~n13629 ) ;
  assign n18943 = n11437 ^ n8188 ^ 1'b0 ;
  assign n18944 = n14784 & n18943 ;
  assign n18945 = n8121 | n11618 ;
  assign n18946 = n18945 ^ n7052 ^ 1'b0 ;
  assign n18947 = n4579 ^ n788 ^ 1'b0 ;
  assign n18948 = x35 & n18947 ;
  assign n18949 = n1521 & ~n18948 ;
  assign n18950 = n18949 ^ n5985 ^ 1'b0 ;
  assign n18951 = n6449 & ~n7807 ;
  assign n18952 = n18951 ^ n10512 ^ 1'b0 ;
  assign n18953 = n15843 ^ n15198 ^ 1'b0 ;
  assign n18954 = n12181 & ~n18953 ;
  assign n18955 = ~x76 & n18954 ;
  assign n18956 = n15448 ^ n7213 ^ n922 ;
  assign n18957 = n1147 | n5321 ;
  assign n18958 = n18957 ^ n5259 ^ 1'b0 ;
  assign n18959 = n4471 & ~n17546 ;
  assign n18960 = n3667 ^ x24 ^ 1'b0 ;
  assign n18961 = n5347 | n18960 ;
  assign n18962 = n17455 & ~n18961 ;
  assign n18963 = n2051 & n3778 ;
  assign n18964 = n16106 ^ n5652 ^ 1'b0 ;
  assign n18965 = n3509 | n18964 ;
  assign n18966 = ~n4011 & n14932 ;
  assign n18967 = n3723 & ~n16021 ;
  assign n18968 = n3300 & ~n18810 ;
  assign n18969 = n3904 ^ n190 ^ 1'b0 ;
  assign n18970 = n18968 & ~n18969 ;
  assign n18971 = n10890 & ~n13314 ;
  assign n18972 = ~n744 & n2697 ;
  assign n18973 = n18972 ^ n1301 ^ 1'b0 ;
  assign n18974 = n2506 & ~n13159 ;
  assign n18975 = n18974 ^ n528 ^ 1'b0 ;
  assign n18976 = n15664 ^ n9458 ^ 1'b0 ;
  assign n18977 = ~n1291 & n13150 ;
  assign n18990 = ~n5494 & n7676 ;
  assign n18984 = n1329 & n1833 ;
  assign n18985 = ~n1329 & n18984 ;
  assign n18986 = ~n4153 & n18985 ;
  assign n18987 = n4153 & n18986 ;
  assign n18983 = n16474 ^ n11645 ^ 1'b0 ;
  assign n18988 = n18987 ^ n18983 ^ 1'b0 ;
  assign n18978 = n1792 & n2513 ;
  assign n18979 = ~n1792 & n18978 ;
  assign n18980 = n1464 | n5492 ;
  assign n18981 = n18979 & ~n18980 ;
  assign n18982 = n12235 | n18981 ;
  assign n18989 = n18988 ^ n18982 ^ 1'b0 ;
  assign n18991 = n18990 ^ n18989 ^ 1'b0 ;
  assign n18992 = n12878 & ~n18991 ;
  assign n18993 = n2620 & n18992 ;
  assign n18994 = ~n14109 & n18993 ;
  assign n18995 = n1625 & n8314 ;
  assign n18996 = n13446 & n18995 ;
  assign n18997 = ~n1786 & n4005 ;
  assign n18998 = n722 & n5589 ;
  assign n18999 = x10 & n6537 ;
  assign n19000 = ( x33 & n5937 ) | ( x33 & ~n18999 ) | ( n5937 & ~n18999 ) ;
  assign n19001 = n1161 & n6688 ;
  assign n19002 = n237 & n246 ;
  assign n19003 = ~n246 & n19002 ;
  assign n19004 = n652 & ~n19003 ;
  assign n19005 = n19003 & n19004 ;
  assign n19014 = n808 & n2067 ;
  assign n19015 = n19005 & n19014 ;
  assign n19006 = n1387 | n19005 ;
  assign n19007 = n19005 & ~n19006 ;
  assign n19008 = n408 & n627 ;
  assign n19009 = ~n627 & n19008 ;
  assign n19010 = n19009 ^ n4072 ^ 1'b0 ;
  assign n19011 = n9432 & n19010 ;
  assign n19012 = n19007 & n19011 ;
  assign n19013 = n15381 | n19012 ;
  assign n19016 = n19015 ^ n19013 ^ 1'b0 ;
  assign n19017 = n2200 | n19016 ;
  assign n19018 = n19017 ^ n1001 ^ 1'b0 ;
  assign n19019 = n18609 & ~n19018 ;
  assign n19020 = n3794 | n4110 ;
  assign n19021 = n3247 | n6558 ;
  assign n19022 = n17397 ^ n8955 ^ n2160 ;
  assign n19023 = n2704 & n16217 ;
  assign n19024 = n18499 ^ n7238 ^ 1'b0 ;
  assign n19025 = n4452 & ~n19024 ;
  assign n19026 = n754 | n1829 ;
  assign n19027 = n19026 ^ n4558 ^ 1'b0 ;
  assign n19028 = n10862 ^ n6716 ^ 1'b0 ;
  assign n19029 = n19027 & ~n19028 ;
  assign n19030 = ~n18760 & n19029 ;
  assign n19031 = ~n19025 & n19030 ;
  assign n19032 = ~n8605 & n16849 ;
  assign n19033 = ~n2660 & n19032 ;
  assign n19034 = n19033 ^ n11980 ^ 1'b0 ;
  assign n19035 = n11710 ^ n7698 ^ n1816 ;
  assign n19036 = ~n397 & n8602 ;
  assign n19037 = ~n1529 & n19036 ;
  assign n19038 = n4318 | n19037 ;
  assign n19039 = n2478 | n19038 ;
  assign n19040 = n19039 ^ n9495 ^ n3878 ;
  assign n19041 = ~n2533 & n19040 ;
  assign n19042 = n693 & ~n10978 ;
  assign n19043 = ~n1063 & n7804 ;
  assign n19044 = n19043 ^ n15346 ^ 1'b0 ;
  assign n19045 = n15355 ^ n3486 ^ 1'b0 ;
  assign n19046 = ~n10939 & n19045 ;
  assign n19047 = ~n5789 & n13432 ;
  assign n19048 = n10957 & n17574 ;
  assign n19049 = n1626 & ~n1734 ;
  assign n19050 = ~n15146 & n19049 ;
  assign n19051 = n19050 ^ n18246 ^ 1'b0 ;
  assign n19052 = n1049 | n19051 ;
  assign n19053 = n595 & ~n10887 ;
  assign n19054 = n19053 ^ n7354 ^ n1049 ;
  assign n19055 = n12905 & n13961 ;
  assign n19056 = n3192 ^ n1439 ^ 1'b0 ;
  assign n19057 = n823 & ~n19056 ;
  assign n19058 = n2806 | n16873 ;
  assign n19059 = n19058 ^ n13670 ^ 1'b0 ;
  assign n19060 = n4919 & n6293 ;
  assign n19061 = n164 | n19060 ;
  assign n19062 = n3509 & ~n19061 ;
  assign n19063 = n19062 ^ n967 ^ 1'b0 ;
  assign n19065 = n221 | n3220 ;
  assign n19066 = n4276 | n19065 ;
  assign n19064 = x47 & x84 ;
  assign n19067 = n19066 ^ n19064 ^ 1'b0 ;
  assign n19069 = n12367 ^ n5889 ^ 1'b0 ;
  assign n19070 = ~n1867 & n19069 ;
  assign n19068 = n8396 | n9349 ;
  assign n19071 = n19070 ^ n19068 ^ 1'b0 ;
  assign n19072 = n6857 ^ n1908 ^ 1'b0 ;
  assign n19073 = n16182 ^ n4668 ^ 1'b0 ;
  assign n19074 = n4573 & n19073 ;
  assign n19075 = ~n5693 & n15137 ;
  assign n19076 = n19075 ^ n9391 ^ 1'b0 ;
  assign n19077 = n11246 | n14819 ;
  assign n19078 = ~n4618 & n19077 ;
  assign n19079 = n855 | n18564 ;
  assign n19080 = n4267 & n5186 ;
  assign n19081 = n19080 ^ n14871 ^ 1'b0 ;
  assign n19082 = n2683 | n8959 ;
  assign n19083 = n14394 & ~n19082 ;
  assign n19084 = n4069 ^ n3409 ^ 1'b0 ;
  assign n19085 = n859 & ~n19084 ;
  assign n19086 = n13724 ^ n6862 ^ 1'b0 ;
  assign n19087 = n10639 & n19086 ;
  assign n19088 = n5954 ^ n1325 ^ 1'b0 ;
  assign n19089 = ~n10212 & n10528 ;
  assign n19090 = n19088 & n19089 ;
  assign n19091 = n12910 | n19090 ;
  assign n19092 = n9774 | n19091 ;
  assign n19093 = n15177 | n17415 ;
  assign n19094 = ~n6213 & n8235 ;
  assign n19095 = n19094 ^ n410 ^ 1'b0 ;
  assign n19096 = n10528 ^ n707 ^ 1'b0 ;
  assign n19097 = n13234 & n19096 ;
  assign n19098 = n12195 & n19094 ;
  assign n19099 = n1042 & n19098 ;
  assign n19100 = n7361 & n19099 ;
  assign n19101 = n722 & ~n5474 ;
  assign n19102 = n19101 ^ n7643 ^ 1'b0 ;
  assign n19103 = n11989 & n13365 ;
  assign n19104 = n2273 & ~n8933 ;
  assign n19105 = ( ~n3498 & n9763 ) | ( ~n3498 & n19104 ) | ( n9763 & n19104 ) ;
  assign n19106 = n5118 ^ n1226 ^ 1'b0 ;
  assign n19107 = n833 & ~n19106 ;
  assign n19108 = n1905 & n19107 ;
  assign n19109 = n11269 & n19108 ;
  assign n19110 = n2026 & ~n5534 ;
  assign n19111 = n5970 & n5986 ;
  assign n19112 = n6782 & n19111 ;
  assign n19113 = n4898 ^ n560 ^ 1'b0 ;
  assign n19114 = n19112 | n19113 ;
  assign n19115 = ~n12045 & n19114 ;
  assign n19116 = n8789 ^ n5552 ^ 1'b0 ;
  assign n19117 = n6706 | n19116 ;
  assign n19118 = n19117 ^ n2427 ^ 1'b0 ;
  assign n19119 = n5349 & ~n19118 ;
  assign n19120 = n12081 ^ n11249 ^ 1'b0 ;
  assign n19121 = n5686 & ~n7268 ;
  assign n19122 = n19121 ^ n14196 ^ n2906 ;
  assign n19123 = n5693 | n8056 ;
  assign n19124 = n19123 ^ n6887 ^ 1'b0 ;
  assign n19125 = ~n8608 & n19124 ;
  assign n19127 = n12196 ^ n8028 ^ 1'b0 ;
  assign n19128 = n6525 & n19127 ;
  assign n19126 = n8977 & n11829 ;
  assign n19129 = n19128 ^ n19126 ^ 1'b0 ;
  assign n19130 = n13450 ^ n763 ^ 1'b0 ;
  assign n19131 = ~n12765 & n19130 ;
  assign n19132 = n4415 & n5794 ;
  assign n19133 = n19132 ^ n8811 ^ 1'b0 ;
  assign n19134 = ~n2943 & n4384 ;
  assign n19135 = ( n1221 & n4694 ) | ( n1221 & n19134 ) | ( n4694 & n19134 ) ;
  assign n19136 = n5438 ^ n5196 ^ 1'b0 ;
  assign n19137 = n18188 | n19136 ;
  assign n19138 = n19137 ^ n2174 ^ 1'b0 ;
  assign n19139 = ~n19135 & n19138 ;
  assign n19140 = ~n3030 & n17737 ;
  assign n19141 = n19140 ^ n8337 ^ 1'b0 ;
  assign n19142 = n8387 ^ n7603 ^ 1'b0 ;
  assign n19145 = n9257 | n11825 ;
  assign n19143 = n3354 ^ n2389 ^ 1'b0 ;
  assign n19144 = n8014 & ~n19143 ;
  assign n19146 = n19145 ^ n19144 ^ 1'b0 ;
  assign n19147 = n8284 ^ n4706 ^ 1'b0 ;
  assign n19148 = n1072 | n19147 ;
  assign n19149 = n11397 & ~n19148 ;
  assign n19150 = n6934 & ~n15483 ;
  assign n19151 = n4169 & ~n5276 ;
  assign n19152 = ( n3130 & n5878 ) | ( n3130 & n19151 ) | ( n5878 & n19151 ) ;
  assign n19153 = n19152 ^ n3289 ^ n998 ;
  assign n19154 = n741 & n1344 ;
  assign n19155 = n6496 & ~n7806 ;
  assign n19156 = n19155 ^ n15348 ^ 1'b0 ;
  assign n19157 = n12708 ^ n6718 ^ 1'b0 ;
  assign n19158 = ~n6245 & n19157 ;
  assign n19159 = n15652 ^ n277 ^ 1'b0 ;
  assign n19160 = n19159 ^ n8048 ^ 1'b0 ;
  assign n19161 = n9500 & n19160 ;
  assign n19162 = ~n2438 & n13716 ;
  assign n19163 = n19162 ^ n6184 ^ 1'b0 ;
  assign n19164 = n2667 & n8176 ;
  assign n19165 = n19164 ^ n11281 ^ n7547 ;
  assign n19166 = n15321 ^ n11929 ^ n992 ;
  assign n19167 = n12676 & n13824 ;
  assign n19168 = n16585 ^ n9551 ^ 1'b0 ;
  assign n19169 = ~n11241 & n19168 ;
  assign n19170 = n19169 ^ n18797 ^ 1'b0 ;
  assign n19171 = ~n7465 & n14689 ;
  assign n19172 = n19171 ^ n5583 ^ 1'b0 ;
  assign n19173 = n19172 ^ n11295 ^ 1'b0 ;
  assign n19174 = n3196 ^ n2604 ^ 1'b0 ;
  assign n19175 = n18227 ^ n13841 ^ 1'b0 ;
  assign n19176 = n5940 | n19175 ;
  assign n19177 = n2944 & ~n19176 ;
  assign n19178 = n2178 & n11344 ;
  assign n19179 = n2048 & ~n19178 ;
  assign n19180 = ~n6531 & n19179 ;
  assign n19181 = n5944 & n14643 ;
  assign n19182 = ~n5405 & n9560 ;
  assign n19183 = n2160 ^ n538 ^ 1'b0 ;
  assign n19184 = n135 & ~n19183 ;
  assign n19185 = n19184 ^ n17521 ^ 1'b0 ;
  assign n19186 = n1645 | n12100 ;
  assign n19188 = ~n1774 & n13611 ;
  assign n19187 = n1129 | n4790 ;
  assign n19189 = n19188 ^ n19187 ^ n14468 ;
  assign n19190 = n4065 | n5596 ;
  assign n19191 = n6592 | n19190 ;
  assign n19192 = ~n6644 & n19191 ;
  assign n19193 = n1124 & n2161 ;
  assign n19194 = ~n1416 & n7731 ;
  assign n19195 = ~n7731 & n19194 ;
  assign n19196 = ~n7242 & n19195 ;
  assign n19197 = n18431 & ~n19196 ;
  assign n19198 = n11744 & ~n19197 ;
  assign n19199 = ~n10812 & n19198 ;
  assign n19200 = n2396 ^ n1515 ^ 1'b0 ;
  assign n19201 = ~n7335 & n19200 ;
  assign n19202 = ~n177 & n19201 ;
  assign n19203 = n19202 ^ n954 ^ 1'b0 ;
  assign n19204 = n797 & n12519 ;
  assign n19205 = ~n13308 & n19204 ;
  assign n19206 = n942 & ~n2598 ;
  assign n19207 = ~n830 & n19206 ;
  assign n19208 = n19207 ^ n2349 ^ 1'b0 ;
  assign n19209 = n15306 ^ n8054 ^ n6590 ;
  assign n19210 = n12934 ^ n632 ^ 1'b0 ;
  assign n19211 = n18217 ^ n13832 ^ x54 ;
  assign n19212 = n10811 ^ n667 ^ 1'b0 ;
  assign n19213 = ~n1540 & n19212 ;
  assign n19214 = n5789 & ~n7631 ;
  assign n19215 = ( n7235 & ~n14650 ) | ( n7235 & n19214 ) | ( ~n14650 & n19214 ) ;
  assign n19216 = n15175 ^ n830 ^ 1'b0 ;
  assign n19217 = ~n5141 & n19216 ;
  assign n19218 = n19217 ^ n4261 ^ 1'b0 ;
  assign n19219 = n19215 | n19218 ;
  assign n19220 = n795 & n6234 ;
  assign n19221 = n19220 ^ n12219 ^ 1'b0 ;
  assign n19222 = n19221 ^ n994 ^ 1'b0 ;
  assign n19223 = n2581 & ~n3604 ;
  assign n19224 = n19223 ^ n2542 ^ 1'b0 ;
  assign n19225 = n4710 | n6912 ;
  assign n19226 = n5847 & ~n19225 ;
  assign n19227 = n12286 & n18630 ;
  assign n19228 = n16017 ^ n14301 ^ n11421 ;
  assign n19229 = n11195 ^ n1784 ^ n325 ;
  assign n19230 = n19228 | n19229 ;
  assign n19231 = n1864 | n3584 ;
  assign n19232 = n19231 ^ n17050 ^ 1'b0 ;
  assign n19233 = n12248 | n12785 ;
  assign n19234 = n19232 | n19233 ;
  assign n19235 = n6173 ^ n594 ^ 1'b0 ;
  assign n19236 = n6024 & ~n19235 ;
  assign n19237 = x6 & n19236 ;
  assign n19238 = n19237 ^ n1768 ^ 1'b0 ;
  assign n19239 = n3195 & n4340 ;
  assign n19240 = n6242 & ~n19239 ;
  assign n19241 = n19240 ^ n14310 ^ 1'b0 ;
  assign n19242 = n1635 & n19241 ;
  assign n19243 = n1035 & ~n10094 ;
  assign n19244 = n2159 & n19243 ;
  assign n19245 = n8215 ^ n7454 ^ 1'b0 ;
  assign n19246 = n2981 | n19245 ;
  assign n19247 = ~n1084 & n11081 ;
  assign n19248 = n11082 ^ n4252 ^ 1'b0 ;
  assign n19249 = n6024 & n19248 ;
  assign n19250 = n7364 & n19249 ;
  assign n19251 = n1579 & ~n11337 ;
  assign n19259 = n7900 ^ n270 ^ 1'b0 ;
  assign n19260 = ~n480 & n19259 ;
  assign n19252 = x61 & ~n1301 ;
  assign n19253 = ~n998 & n19252 ;
  assign n19254 = n7698 ^ n1381 ^ 1'b0 ;
  assign n19255 = n7444 | n19254 ;
  assign n19256 = n15232 | n19255 ;
  assign n19257 = n18930 & ~n19256 ;
  assign n19258 = n19253 & n19257 ;
  assign n19261 = n19260 ^ n19258 ^ 1'b0 ;
  assign n19262 = ( n8535 & ~n14983 ) | ( n8535 & n19261 ) | ( ~n14983 & n19261 ) ;
  assign n19263 = n2584 & n6540 ;
  assign n19264 = n5035 & ~n19263 ;
  assign n19265 = n14361 ^ n9698 ^ n6057 ;
  assign n19266 = ~n1315 & n15645 ;
  assign n19267 = n1467 & n19266 ;
  assign n19268 = x16 & n5016 ;
  assign n19269 = n19268 ^ n18652 ^ 1'b0 ;
  assign n19270 = n5356 & ~n15440 ;
  assign n19271 = ~n14537 & n17978 ;
  assign n19272 = n19271 ^ n8015 ^ 1'b0 ;
  assign n19273 = n4555 ^ n2726 ^ 1'b0 ;
  assign n19274 = n5349 & ~n19273 ;
  assign n19275 = ~n15391 & n19274 ;
  assign n19276 = n19275 ^ n16390 ^ 1'b0 ;
  assign n19277 = n3697 ^ n1691 ^ 1'b0 ;
  assign n19278 = n936 ^ n867 ^ 1'b0 ;
  assign n19279 = ~n15873 & n19278 ;
  assign n19280 = ~n512 & n19279 ;
  assign n19281 = n12569 ^ n8724 ^ 1'b0 ;
  assign n19282 = n10923 & n19281 ;
  assign n19283 = n14529 | n17442 ;
  assign n19284 = n9056 ^ n7788 ^ 1'b0 ;
  assign n19285 = n6272 & ~n15620 ;
  assign n19286 = n3718 ^ n3339 ^ 1'b0 ;
  assign n19287 = n5538 & ~n19286 ;
  assign n19288 = ~n502 & n19287 ;
  assign n19289 = n6425 & n19288 ;
  assign n19290 = n11280 | n19289 ;
  assign n19291 = n19290 ^ n962 ^ 1'b0 ;
  assign n19292 = ~n3267 & n19291 ;
  assign n19293 = ~n13944 & n19292 ;
  assign n19294 = n1624 & n6522 ;
  assign n19295 = n19294 ^ n17444 ^ 1'b0 ;
  assign n19297 = n835 & ~n1552 ;
  assign n19296 = n1268 & ~n16250 ;
  assign n19298 = n19297 ^ n19296 ^ 1'b0 ;
  assign n19299 = n12425 ^ n2062 ^ 1'b0 ;
  assign n19300 = ~n4457 & n19299 ;
  assign n19301 = n14549 ^ n325 ^ 1'b0 ;
  assign n19302 = ~n3324 & n19301 ;
  assign n19303 = n693 & ~n1716 ;
  assign n19304 = n9252 ^ n2942 ^ 1'b0 ;
  assign n19305 = ~n1604 & n19304 ;
  assign n19306 = n19305 ^ x87 ^ 1'b0 ;
  assign n19307 = n245 & n11188 ;
  assign n19308 = n238 & ~n19307 ;
  assign n19309 = ~x90 & n5543 ;
  assign n19310 = ~n9435 & n12315 ;
  assign n19311 = n741 & ~n1935 ;
  assign n19312 = n19311 ^ n7595 ^ 1'b0 ;
  assign n19313 = ~n2340 & n12862 ;
  assign n19314 = n14763 & ~n17352 ;
  assign n19315 = n7688 ^ n6562 ^ 1'b0 ;
  assign n19316 = n9945 | n19315 ;
  assign n19317 = n835 ^ x22 ^ 1'b0 ;
  assign n19318 = n15995 ^ n8055 ^ 1'b0 ;
  assign n19319 = ~n7905 & n13333 ;
  assign n19320 = n19319 ^ x69 ^ 1'b0 ;
  assign n19321 = n14731 & n19320 ;
  assign n19322 = n6054 & ~n6370 ;
  assign n19323 = n19322 ^ n1070 ^ 1'b0 ;
  assign n19324 = n19323 ^ n14633 ^ n11331 ;
  assign n19325 = n9544 & ~n10157 ;
  assign n19326 = n4690 & n19325 ;
  assign n19327 = n12629 & n19326 ;
  assign n19328 = ~n4091 & n12696 ;
  assign n19329 = n11517 | n12444 ;
  assign n19330 = ~n11363 & n17478 ;
  assign n19331 = ~n14071 & n19330 ;
  assign n19332 = n12942 | n14649 ;
  assign n19333 = n19332 ^ n4112 ^ 1'b0 ;
  assign n19334 = n4998 & ~n9241 ;
  assign n19335 = n8787 & ~n19334 ;
  assign n19336 = n11503 ^ n2835 ^ 1'b0 ;
  assign n19337 = ~n10983 & n19336 ;
  assign n19338 = ~n7391 & n19337 ;
  assign n19339 = n10987 & n19338 ;
  assign n19340 = n19339 ^ n12551 ^ 1'b0 ;
  assign n19342 = ~n6272 & n16553 ;
  assign n19341 = n1648 | n6931 ;
  assign n19343 = n19342 ^ n19341 ^ 1'b0 ;
  assign n19344 = n5268 & ~n7259 ;
  assign n19345 = n847 | n8589 ;
  assign n19346 = n6540 ^ n6197 ^ 1'b0 ;
  assign n19347 = n19346 ^ n16576 ^ n11265 ;
  assign n19348 = n2765 & ~n10669 ;
  assign n19349 = n14329 & ~n14654 ;
  assign n19350 = n19348 & n19349 ;
  assign n19351 = n246 & ~n6059 ;
  assign n19352 = n14745 | n19351 ;
  assign n19353 = n4430 | n5876 ;
  assign n19354 = n19352 & n19353 ;
  assign n19355 = n8518 & n11186 ;
  assign n19356 = n625 & n19355 ;
  assign n19357 = n19042 ^ n196 ^ 1'b0 ;
  assign n19358 = n9465 & ~n18897 ;
  assign n19359 = ~n6756 & n19358 ;
  assign n19360 = n11879 ^ n342 ^ 1'b0 ;
  assign n19361 = n10791 | n19360 ;
  assign n19362 = n19361 ^ n3256 ^ 1'b0 ;
  assign n19363 = ~n9410 & n19362 ;
  assign n19364 = n1356 & n3269 ;
  assign n19365 = n19364 ^ x80 ^ 1'b0 ;
  assign n19366 = n19365 ^ n1008 ^ 1'b0 ;
  assign n19367 = ~n5613 & n19366 ;
  assign n19368 = n14205 | n14578 ;
  assign n19369 = ~n7259 & n19368 ;
  assign n19370 = n5008 ^ n970 ^ 1'b0 ;
  assign n19371 = n15206 ^ n7564 ^ 1'b0 ;
  assign n19372 = n19370 | n19371 ;
  assign n19373 = n1147 & n19372 ;
  assign n19374 = n2794 & ~n19373 ;
  assign n19379 = n502 & ~n4985 ;
  assign n19375 = ( n1348 & n6439 ) | ( n1348 & n7894 ) | ( n6439 & n7894 ) ;
  assign n19376 = n711 & ~n19375 ;
  assign n19377 = n19376 ^ n11677 ^ 1'b0 ;
  assign n19378 = ~n18212 & n19377 ;
  assign n19380 = n19379 ^ n19378 ^ 1'b0 ;
  assign n19381 = n11461 ^ n7467 ^ 1'b0 ;
  assign n19382 = n7439 ^ n6829 ^ 1'b0 ;
  assign n19383 = n19221 ^ n3291 ^ 1'b0 ;
  assign n19384 = ~n19382 & n19383 ;
  assign n19385 = n6890 & ~n13215 ;
  assign n19386 = n7467 | n10305 ;
  assign n19387 = n19385 | n19386 ;
  assign n19388 = n5804 | n9787 ;
  assign n19389 = n19388 ^ n6511 ^ 1'b0 ;
  assign n19390 = ( n2897 & n2986 ) | ( n2897 & ~n3347 ) | ( n2986 & ~n3347 ) ;
  assign n19391 = n19390 ^ n1957 ^ 1'b0 ;
  assign n19392 = n13138 & ~n18663 ;
  assign n19393 = n2669 & ~n5572 ;
  assign n19394 = ~n3353 & n19393 ;
  assign n19395 = n14614 ^ n9441 ^ n4027 ;
  assign n19397 = n8126 & ~n19117 ;
  assign n19396 = n11293 ^ n9145 ^ n972 ;
  assign n19398 = n19397 ^ n19396 ^ 1'b0 ;
  assign n19399 = n14456 ^ n788 ^ 1'b0 ;
  assign n19400 = n5716 & n19399 ;
  assign n19401 = ~n788 & n19400 ;
  assign n19402 = n10313 & n19401 ;
  assign n19403 = n1208 | n6190 ;
  assign n19404 = ~n3708 & n6211 ;
  assign n19405 = n12308 & n19404 ;
  assign n19406 = n1102 & n19131 ;
  assign n19407 = n14760 ^ n1185 ^ 1'b0 ;
  assign n19408 = n307 & ~n15948 ;
  assign n19409 = n16855 & ~n19408 ;
  assign n19410 = ~n5360 & n11838 ;
  assign n19411 = n9791 ^ n2800 ^ 1'b0 ;
  assign n19412 = n3999 ^ n2171 ^ 1'b0 ;
  assign n19413 = n5005 & ~n19412 ;
  assign n19414 = ~n10006 & n19413 ;
  assign n19415 = ~n19411 & n19414 ;
  assign n19416 = n2752 | n19129 ;
  assign n19417 = n19416 ^ n8044 ^ 1'b0 ;
  assign n19418 = n12803 & ~n18204 ;
  assign n19419 = n5455 & ~n6514 ;
  assign n19420 = n326 & n19419 ;
  assign n19421 = n19420 ^ n4819 ^ 1'b0 ;
  assign n19422 = n17027 ^ n10320 ^ n4682 ;
  assign n19423 = n5031 ^ n2795 ^ 1'b0 ;
  assign n19424 = n13127 ^ n2347 ^ n1188 ;
  assign n19425 = n19423 & n19424 ;
  assign n19426 = n6902 ^ n307 ^ 1'b0 ;
  assign n19427 = n18607 | n19426 ;
  assign n19428 = n2136 | n4197 ;
  assign n19429 = n12207 & ~n16065 ;
  assign n19430 = n19429 ^ n5605 ^ 1'b0 ;
  assign n19431 = ~n5596 & n19430 ;
  assign n19432 = n6607 & n6667 ;
  assign n19433 = ~n11822 & n19432 ;
  assign n19434 = n3874 | n19433 ;
  assign n19435 = n6871 ^ n5836 ^ n4635 ;
  assign n19436 = n7231 & n19435 ;
  assign n19437 = n5735 | n18936 ;
  assign n19438 = n19437 ^ n6239 ^ 1'b0 ;
  assign n19439 = n19438 ^ n17737 ^ 1'b0 ;
  assign n19440 = n19439 ^ n15650 ^ 1'b0 ;
  assign n19441 = n19436 & n19440 ;
  assign n19442 = n16244 ^ n3981 ^ n289 ;
  assign n19443 = n4328 & ~n12308 ;
  assign n19444 = n13864 & n19443 ;
  assign n19445 = n19444 ^ n831 ^ 1'b0 ;
  assign n19446 = n12698 ^ n6816 ^ 1'b0 ;
  assign n19447 = n6934 | n19446 ;
  assign n19449 = n8171 & n12685 ;
  assign n19450 = n1837 & n19449 ;
  assign n19448 = ( n9784 & n11348 ) | ( n9784 & n11881 ) | ( n11348 & n11881 ) ;
  assign n19451 = n19450 ^ n19448 ^ 1'b0 ;
  assign n19452 = n3136 & n8145 ;
  assign n19453 = n19452 ^ n10152 ^ 1'b0 ;
  assign n19454 = n6987 & n17478 ;
  assign n19455 = n8615 & n19454 ;
  assign n19456 = n13382 ^ n8005 ^ 1'b0 ;
  assign n19457 = x73 & ~n211 ;
  assign n19458 = n360 & ~n14865 ;
  assign n19459 = n9709 ^ n6991 ^ 1'b0 ;
  assign n19460 = n11240 & ~n19459 ;
  assign n19461 = n1040 & n11840 ;
  assign n19462 = n19461 ^ n3521 ^ 1'b0 ;
  assign n19463 = n5125 ^ n897 ^ 1'b0 ;
  assign n19464 = n5426 | n13851 ;
  assign n19465 = n2673 & ~n7736 ;
  assign n19466 = n19465 ^ n5410 ^ 1'b0 ;
  assign n19467 = n9142 & ~n15062 ;
  assign n19468 = n19466 & n19467 ;
  assign n19469 = n2838 ^ x38 ^ 1'b0 ;
  assign n19470 = n2691 ^ n604 ^ 1'b0 ;
  assign n19471 = ~n19469 & n19470 ;
  assign n19472 = n4661 | n11024 ;
  assign n19473 = n7855 & ~n17508 ;
  assign n19474 = n19473 ^ n1714 ^ 1'b0 ;
  assign n19475 = n5414 | n15911 ;
  assign n19476 = n1005 & n10142 ;
  assign n19477 = ~n3238 & n19476 ;
  assign n19478 = n775 | n5214 ;
  assign n19479 = n11715 & ~n19478 ;
  assign n19480 = n19479 ^ n16041 ^ 1'b0 ;
  assign n19481 = n2224 ^ n373 ^ 1'b0 ;
  assign n19482 = n2694 & n7933 ;
  assign n19483 = n12484 ^ n4708 ^ n3499 ;
  assign n19484 = n3975 | n10196 ;
  assign n19485 = n648 ^ n492 ^ 1'b0 ;
  assign n19486 = n19485 ^ n8194 ^ n2893 ;
  assign n19487 = n2898 | n17237 ;
  assign n19488 = n19487 ^ n10352 ^ 1'b0 ;
  assign n19489 = n3613 & n10864 ;
  assign n19490 = n7349 & n19489 ;
  assign n19491 = n1792 & n9265 ;
  assign n19492 = ~n11385 & n19491 ;
  assign n19493 = n12090 & ~n13688 ;
  assign n19494 = n2669 & n19493 ;
  assign n19495 = n19494 ^ n2113 ^ 1'b0 ;
  assign n19496 = n3580 & n8398 ;
  assign n19497 = n19496 ^ n18925 ^ 1'b0 ;
  assign n19498 = n4459 ^ n3764 ^ 1'b0 ;
  assign n19499 = n3082 | n19498 ;
  assign n19502 = n198 | n2044 ;
  assign n19503 = n6421 & ~n19502 ;
  assign n19504 = n7468 & ~n19503 ;
  assign n19500 = n4238 | n8980 ;
  assign n19501 = n19500 ^ n8067 ^ 1'b0 ;
  assign n19505 = n19504 ^ n19501 ^ 1'b0 ;
  assign n19506 = n5087 ^ n4749 ^ 1'b0 ;
  assign n19507 = n10058 | n10263 ;
  assign n19508 = n19507 ^ n10777 ^ 1'b0 ;
  assign n19509 = n19506 | n19508 ;
  assign n19510 = n14166 | n19509 ;
  assign n19511 = n1414 & n2775 ;
  assign n19512 = ~n3047 & n19511 ;
  assign n19513 = ~x100 & n5098 ;
  assign n19514 = n333 & n3859 ;
  assign n19515 = n2713 ^ n893 ^ 1'b0 ;
  assign n19516 = n19514 & ~n19515 ;
  assign n19517 = ~n19513 & n19516 ;
  assign n19518 = n3785 & n9005 ;
  assign n19519 = ~n15645 & n19518 ;
  assign n19520 = n3302 & n7685 ;
  assign n19521 = n2999 & n8022 ;
  assign n19522 = n19521 ^ x17 ^ 1'b0 ;
  assign n19523 = n19522 ^ n5363 ^ 1'b0 ;
  assign n19524 = n1329 & n9602 ;
  assign n19525 = n16585 ^ n3418 ^ n2091 ;
  assign n19526 = n5844 & n19525 ;
  assign n19527 = n3153 & ~n14497 ;
  assign n19528 = ~n16902 & n17473 ;
  assign n19529 = n18756 & n19528 ;
  assign n19530 = n2048 & n12083 ;
  assign n19531 = ~n9217 & n19530 ;
  assign n19532 = n16182 | n19531 ;
  assign n19533 = n19532 ^ n10586 ^ n9791 ;
  assign n19534 = n19533 ^ n16434 ^ 1'b0 ;
  assign n19535 = n3112 & n19534 ;
  assign n19536 = n2328 | n10198 ;
  assign n19537 = ~n19535 & n19536 ;
  assign n19538 = ~n13082 & n16313 ;
  assign n19539 = n11124 ^ n507 ^ 1'b0 ;
  assign n19540 = n2317 | n19539 ;
  assign n19541 = n1467 | n11404 ;
  assign n19542 = n19541 ^ n5488 ^ 1'b0 ;
  assign n19543 = n7942 ^ n198 ^ 1'b0 ;
  assign n19544 = n14118 | n19543 ;
  assign n19545 = n4323 & ~n19544 ;
  assign n19546 = n15697 | n19545 ;
  assign n19547 = n3525 ^ n1984 ^ 1'b0 ;
  assign n19548 = n19546 & ~n19547 ;
  assign n19549 = n19323 ^ n4654 ^ 1'b0 ;
  assign n19550 = n15901 ^ x11 ^ 1'b0 ;
  assign n19551 = n12796 & ~n19550 ;
  assign n19552 = ~n8506 & n14586 ;
  assign n19553 = n19552 ^ n5245 ^ 1'b0 ;
  assign n19554 = n18608 & n19553 ;
  assign n19555 = n3428 & ~n11433 ;
  assign n19556 = ~n6338 & n19555 ;
  assign n19557 = n12984 ^ n1904 ^ 1'b0 ;
  assign n19558 = n14808 ^ n10563 ^ 1'b0 ;
  assign n19563 = n3722 & ~n4863 ;
  assign n19559 = n16203 ^ n9367 ^ 1'b0 ;
  assign n19560 = n2129 & ~n19559 ;
  assign n19561 = x103 & ~n19560 ;
  assign n19562 = n19561 ^ n5705 ^ n3070 ;
  assign n19564 = n19563 ^ n19562 ^ 1'b0 ;
  assign n19565 = n10382 ^ n8083 ^ n6333 ;
  assign n19566 = ~n2043 & n19565 ;
  assign n19567 = n1449 & ~n1662 ;
  assign n19568 = n6018 | n19567 ;
  assign n19569 = n19568 ^ n9801 ^ 1'b0 ;
  assign n19570 = ( n427 & n886 ) | ( n427 & n6617 ) | ( n886 & n6617 ) ;
  assign n19571 = n19570 ^ n6901 ^ 1'b0 ;
  assign n19572 = n3353 ^ n1623 ^ 1'b0 ;
  assign n19573 = n3238 & ~n19572 ;
  assign n19574 = n7573 ^ n6214 ^ 1'b0 ;
  assign n19575 = n2707 & ~n19574 ;
  assign n19576 = ~n865 & n3429 ;
  assign n19577 = ~n18429 & n19576 ;
  assign n19578 = ~n19575 & n19577 ;
  assign n19579 = n15818 | n18729 ;
  assign n19580 = n4240 & ~n19579 ;
  assign n19581 = n7338 ^ n5722 ^ 1'b0 ;
  assign n19582 = n1001 & n19581 ;
  assign n19583 = n19582 ^ n5929 ^ 1'b0 ;
  assign n19584 = n814 | n19365 ;
  assign n19586 = n2329 ^ n399 ^ 1'b0 ;
  assign n19585 = n8244 & n12436 ;
  assign n19587 = n19586 ^ n19585 ^ 1'b0 ;
  assign n19588 = n12271 ^ n10831 ^ n5688 ;
  assign n19589 = n6566 & ~n13701 ;
  assign n19590 = n19589 ^ n6384 ^ 1'b0 ;
  assign n19591 = n8009 ^ n1228 ^ 1'b0 ;
  assign n19592 = n1558 & ~n2309 ;
  assign n19593 = n19592 ^ n4978 ^ 1'b0 ;
  assign n19594 = n5525 & ~n19593 ;
  assign n19598 = n1436 & ~n4621 ;
  assign n19595 = n9218 ^ n6933 ^ 1'b0 ;
  assign n19596 = n11499 & n19595 ;
  assign n19597 = ~n7535 & n19596 ;
  assign n19599 = n19598 ^ n19597 ^ 1'b0 ;
  assign n19600 = n8874 | n18939 ;
  assign n19601 = n156 & n9647 ;
  assign n19602 = n4901 & n7673 ;
  assign n19603 = n19602 ^ n1185 ^ 1'b0 ;
  assign n19604 = ~n8813 & n15251 ;
  assign n19605 = n19604 ^ n14209 ^ 1'b0 ;
  assign n19606 = n11873 ^ n10497 ^ 1'b0 ;
  assign n19607 = ~n8237 & n11047 ;
  assign n19608 = n19607 ^ n14465 ^ 1'b0 ;
  assign n19609 = n19608 ^ n13663 ^ 1'b0 ;
  assign n19610 = ~n18188 & n19609 ;
  assign n19611 = n6336 & ~n9541 ;
  assign n19612 = ~n5121 & n19261 ;
  assign n19613 = ~n5096 & n19612 ;
  assign n19614 = n4933 | n5165 ;
  assign n19616 = n8488 & ~n10887 ;
  assign n19617 = n19616 ^ n3746 ^ 1'b0 ;
  assign n19615 = n9059 & ~n11677 ;
  assign n19618 = n19617 ^ n19615 ^ n9858 ;
  assign n19619 = n9071 ^ n6861 ^ 1'b0 ;
  assign n19620 = n12882 & ~n19619 ;
  assign n19621 = ~n2716 & n2925 ;
  assign n19622 = n709 & n19621 ;
  assign n19623 = n1632 & n19370 ;
  assign n19624 = n19623 ^ n9190 ^ 1'b0 ;
  assign n19625 = n2002 & ~n19624 ;
  assign n19626 = n19625 ^ n7037 ^ 1'b0 ;
  assign n19627 = n7935 ^ n5113 ^ n1548 ;
  assign n19628 = x46 & n4647 ;
  assign n19629 = n10918 & n19628 ;
  assign n19630 = n19185 ^ n15813 ^ 1'b0 ;
  assign n19631 = ~n2669 & n19630 ;
  assign n19632 = n3371 | n14093 ;
  assign n19633 = n19632 ^ n11164 ^ 1'b0 ;
  assign n19634 = n825 & ~n11309 ;
  assign n19635 = n19634 ^ n733 ^ 1'b0 ;
  assign n19636 = n9913 ^ n2155 ^ 1'b0 ;
  assign n19637 = n16822 ^ n11853 ^ 1'b0 ;
  assign n19638 = ~n15652 & n19637 ;
  assign n19639 = n11399 | n14209 ;
  assign n19640 = n3917 & ~n19639 ;
  assign n19641 = n1321 ^ n888 ^ 1'b0 ;
  assign n19642 = n12696 & ~n19641 ;
  assign n19643 = n9780 & ~n14092 ;
  assign n19644 = n1170 | n19490 ;
  assign n19645 = n19644 ^ n17500 ^ 1'b0 ;
  assign n19646 = n4694 | n4816 ;
  assign n19647 = n19646 ^ n10666 ^ 1'b0 ;
  assign n19648 = n7926 ^ n7905 ^ 1'b0 ;
  assign n19649 = n5749 & ~n19648 ;
  assign n19650 = n3144 & ~n6303 ;
  assign n19651 = n14034 & n19650 ;
  assign n19652 = n2598 & ~n19651 ;
  assign n19653 = n2944 | n8356 ;
  assign n19654 = n12172 ^ n3521 ^ 1'b0 ;
  assign n19655 = n1724 & ~n5977 ;
  assign n19656 = n19655 ^ n2641 ^ 1'b0 ;
  assign n19657 = x77 & n8958 ;
  assign n19658 = n2154 & n19657 ;
  assign n19659 = n2987 | n12025 ;
  assign n19660 = ~n19658 & n19659 ;
  assign n19661 = n19660 ^ n2949 ^ 1'b0 ;
  assign n19662 = n18086 ^ n365 ^ 1'b0 ;
  assign n19667 = n8067 ^ n1924 ^ 1'b0 ;
  assign n19666 = n8055 ^ n7232 ^ 1'b0 ;
  assign n19663 = n624 & ~n1545 ;
  assign n19664 = n6934 | n8021 ;
  assign n19665 = n19663 & ~n19664 ;
  assign n19668 = n19667 ^ n19666 ^ n19665 ;
  assign n19669 = n12964 ^ n9475 ^ 1'b0 ;
  assign n19670 = n12984 | n19669 ;
  assign n19671 = n2396 & ~n17013 ;
  assign n19672 = ( ~n3852 & n4114 ) | ( ~n3852 & n14913 ) | ( n4114 & n14913 ) ;
  assign n19673 = n4469 & ~n4900 ;
  assign n19674 = n19672 | n19673 ;
  assign n19675 = ~n1031 & n2873 ;
  assign n19676 = n19675 ^ n8874 ^ 1'b0 ;
  assign n19677 = n2056 & ~n4469 ;
  assign n19678 = n19677 ^ n4556 ^ 1'b0 ;
  assign n19679 = n13802 | n19678 ;
  assign n19680 = n314 & ~n1671 ;
  assign n19681 = n15805 ^ n11698 ^ 1'b0 ;
  assign n19682 = n5115 | n14839 ;
  assign n19683 = n18302 & ~n19682 ;
  assign n19684 = n19683 ^ n512 ^ 1'b0 ;
  assign n19685 = n3910 & n9145 ;
  assign n19686 = ~n7637 & n19685 ;
  assign n19687 = n19686 ^ n19240 ^ 1'b0 ;
  assign n19688 = n19687 ^ n15105 ^ 1'b0 ;
  assign n19689 = ( n1574 & n6851 ) | ( n1574 & n13149 ) | ( n6851 & n13149 ) ;
  assign n19690 = n19689 ^ n17279 ^ 1'b0 ;
  assign n19691 = ~n9623 & n14232 ;
  assign n19692 = n9505 | n12817 ;
  assign n19693 = n9074 | n9749 ;
  assign n19694 = ~n6992 & n13134 ;
  assign n19695 = n143 | n19694 ;
  assign n19696 = n2896 & ~n5630 ;
  assign n19697 = n16934 ^ n15897 ^ 1'b0 ;
  assign n19698 = ~n11654 & n19697 ;
  assign n19699 = n9839 & n17508 ;
  assign n19700 = n1201 | n4022 ;
  assign n19701 = n19699 & ~n19700 ;
  assign n19702 = ~n14685 & n19701 ;
  assign n19703 = n2291 & ~n8055 ;
  assign n19704 = ~n2954 & n19703 ;
  assign n19705 = ~n17256 & n19704 ;
  assign n19706 = n13782 ^ n1493 ^ 1'b0 ;
  assign n19707 = n4716 & n12120 ;
  assign n19708 = n992 & ~n12731 ;
  assign n19709 = n19708 ^ n3236 ^ 1'b0 ;
  assign n19710 = ~n2148 & n5634 ;
  assign n19711 = n19710 ^ n13431 ^ 1'b0 ;
  assign n19712 = n6456 ^ n5819 ^ 1'b0 ;
  assign n19713 = n1351 & ~n8400 ;
  assign n19714 = n19713 ^ n13983 ^ 1'b0 ;
  assign n19715 = n5432 ^ n2940 ^ 1'b0 ;
  assign n19716 = x97 & ~n1898 ;
  assign n19717 = n19715 & n19716 ;
  assign n19718 = n13108 | n19717 ;
  assign n19719 = n19714 & ~n19718 ;
  assign n19720 = n9744 ^ n1002 ^ 1'b0 ;
  assign n19721 = n13077 & n19720 ;
  assign n19722 = n10963 ^ n6320 ^ 1'b0 ;
  assign n19723 = n19721 & n19722 ;
  assign n19724 = n9632 | n12001 ;
  assign n19725 = n7836 & ~n12717 ;
  assign n19728 = n2129 & n5669 ;
  assign n19729 = n19728 ^ n15346 ^ 1'b0 ;
  assign n19730 = n13022 ^ n424 ^ 1'b0 ;
  assign n19731 = n19729 & n19730 ;
  assign n19726 = n15908 ^ n1189 ^ 1'b0 ;
  assign n19727 = ~n11710 & n19726 ;
  assign n19732 = n19731 ^ n19727 ^ n487 ;
  assign n19733 = n436 & ~n948 ;
  assign n19734 = ~n632 & n19733 ;
  assign n19735 = ~x9 & n18122 ;
  assign n19736 = n6271 | n11118 ;
  assign n19737 = n542 & ~n4335 ;
  assign n19738 = ~x9 & n19737 ;
  assign n19739 = n3577 & n19738 ;
  assign n19740 = n19739 ^ n7043 ^ n1718 ;
  assign n19741 = n5404 ^ n4384 ^ 1'b0 ;
  assign n19742 = n14427 ^ n2193 ^ 1'b0 ;
  assign n19743 = n12292 ^ n6945 ^ 1'b0 ;
  assign n19744 = n16454 ^ n3824 ^ 1'b0 ;
  assign n19745 = n16047 | n19744 ;
  assign n19746 = x37 & ~n3071 ;
  assign n19747 = n6091 ^ n992 ^ 1'b0 ;
  assign n19748 = n11469 ^ n9632 ^ 1'b0 ;
  assign n19749 = n19747 & n19748 ;
  assign n19750 = n13594 ^ n7404 ^ 1'b0 ;
  assign n19751 = ( n3952 & ~n6907 ) | ( n3952 & n19750 ) | ( ~n6907 & n19750 ) ;
  assign n19752 = ~n468 & n9848 ;
  assign n19753 = n12203 ^ n8837 ^ 1'b0 ;
  assign n19754 = n6971 & n10211 ;
  assign n19755 = n8286 & n19754 ;
  assign n19756 = n19755 ^ n428 ^ 1'b0 ;
  assign n19757 = n3908 ^ n221 ^ 1'b0 ;
  assign n19758 = n359 | n19757 ;
  assign n19759 = n4337 & ~n10512 ;
  assign n19760 = n9069 ^ n1126 ^ 1'b0 ;
  assign n19761 = n8961 & n19760 ;
  assign n19762 = n19761 ^ n17074 ^ 1'b0 ;
  assign n19763 = n5096 & ~n11735 ;
  assign n19764 = n3672 | n19763 ;
  assign n19765 = n2413 & ~n10688 ;
  assign n19766 = n4289 ^ n4033 ^ 1'b0 ;
  assign n19767 = n5014 & n19766 ;
  assign n19768 = n19767 ^ n9433 ^ 1'b0 ;
  assign n19769 = n13839 | n14886 ;
  assign n19770 = n19769 ^ n7973 ^ 1'b0 ;
  assign n19771 = n4106 & n16901 ;
  assign n19772 = n6948 & ~n9349 ;
  assign n19773 = n19772 ^ n2958 ^ 1'b0 ;
  assign n19774 = n19773 ^ n13715 ^ n7206 ;
  assign n19776 = ~n10695 & n11116 ;
  assign n19777 = n4167 | n19776 ;
  assign n19775 = ~n3035 & n17912 ;
  assign n19778 = n19777 ^ n19775 ^ 1'b0 ;
  assign n19779 = n9383 ^ n5611 ^ 1'b0 ;
  assign n19780 = n4643 & ~n10078 ;
  assign n19781 = n739 & n6361 ;
  assign n19782 = n9364 & n9410 ;
  assign n19783 = n19782 ^ n1833 ^ 1'b0 ;
  assign n19784 = n2811 | n4112 ;
  assign n19785 = n10149 & ~n15083 ;
  assign n19786 = n19785 ^ n18806 ^ 1'b0 ;
  assign n19787 = n6736 | n9784 ;
  assign n19788 = n19787 ^ n7195 ^ 1'b0 ;
  assign n19790 = n1526 ^ n1364 ^ 1'b0 ;
  assign n19791 = n1118 | n19790 ;
  assign n19792 = n18907 ^ x52 ^ 1'b0 ;
  assign n19793 = ~n19791 & n19792 ;
  assign n19789 = ~n1644 & n2574 ;
  assign n19794 = n19793 ^ n19789 ^ 1'b0 ;
  assign n19795 = n2941 ^ n984 ^ 1'b0 ;
  assign n19796 = n18050 | n19795 ;
  assign n19797 = n19796 ^ n1805 ^ 1'b0 ;
  assign n19798 = n2234 | n9600 ;
  assign n19799 = n7188 & ~n19798 ;
  assign n19800 = n19799 ^ n14467 ^ 1'b0 ;
  assign n19801 = n5046 & ~n16081 ;
  assign n19802 = ~n7834 & n19801 ;
  assign n19803 = n19802 ^ n19411 ^ 1'b0 ;
  assign n19804 = n9022 ^ n1986 ^ 1'b0 ;
  assign n19805 = n14441 & n19804 ;
  assign n19806 = n5859 ^ n3813 ^ 1'b0 ;
  assign n19807 = ~n19805 & n19806 ;
  assign n19808 = n19435 ^ n3053 ^ 1'b0 ;
  assign n19809 = n8263 ^ n1702 ^ 1'b0 ;
  assign n19810 = n6907 & ~n18478 ;
  assign n19811 = n4232 & ~n5804 ;
  assign n19812 = n2430 & n19811 ;
  assign n19813 = n19104 ^ n14678 ^ 1'b0 ;
  assign n19814 = n19812 | n19813 ;
  assign n19815 = n10544 ^ n3559 ^ 1'b0 ;
  assign n19816 = ~n11066 & n11801 ;
  assign n19817 = n1807 & n19816 ;
  assign n19818 = n4106 & n19817 ;
  assign n19819 = n2440 ^ n2224 ^ 1'b0 ;
  assign n19820 = n15211 ^ n3160 ^ 1'b0 ;
  assign n19821 = ( n5096 & n11873 ) | ( n5096 & ~n12541 ) | ( n11873 & ~n12541 ) ;
  assign n19822 = n5161 | n8673 ;
  assign n19823 = n3208 & n14937 ;
  assign n19824 = n19823 ^ n8823 ^ 1'b0 ;
  assign n19825 = n696 ^ x22 ^ 1'b0 ;
  assign n19826 = n5007 | n19825 ;
  assign n19827 = ( x17 & n1534 ) | ( x17 & n4746 ) | ( n1534 & n4746 ) ;
  assign n19828 = n19827 ^ n19450 ^ 1'b0 ;
  assign n19829 = x82 | n11245 ;
  assign n19830 = n4274 & ~n19829 ;
  assign n19831 = x55 | n19830 ;
  assign n19832 = n9641 & ~n19831 ;
  assign n19833 = n19832 ^ x83 ^ 1'b0 ;
  assign n19834 = n171 | n11484 ;
  assign n19835 = n14305 ^ n9217 ^ 1'b0 ;
  assign n19837 = n7216 & n9983 ;
  assign n19838 = n10588 & n19837 ;
  assign n19836 = n766 & ~n3179 ;
  assign n19839 = n19838 ^ n19836 ^ 1'b0 ;
  assign n19840 = n4157 | n19839 ;
  assign n19841 = n8176 & n19840 ;
  assign n19842 = ~n1755 & n4224 ;
  assign n19843 = n19842 ^ n11787 ^ n4334 ;
  assign n19844 = n19221 & n19843 ;
  assign n19845 = n5745 & n19844 ;
  assign n19846 = n19845 ^ n9969 ^ 1'b0 ;
  assign n19848 = n4180 & ~n10357 ;
  assign n19847 = n9207 & n11058 ;
  assign n19849 = n19848 ^ n19847 ^ 1'b0 ;
  assign n19850 = n391 | n2934 ;
  assign n19851 = n391 & ~n19850 ;
  assign n19852 = n5898 & ~n19851 ;
  assign n19853 = ( ~n8844 & n19729 ) | ( ~n8844 & n19852 ) | ( n19729 & n19852 ) ;
  assign n19854 = n259 & n19853 ;
  assign n19855 = ( ~n4157 & n6864 ) | ( ~n4157 & n7171 ) | ( n6864 & n7171 ) ;
  assign n19856 = ~n502 & n1887 ;
  assign n19857 = n10278 & n14371 ;
  assign n19858 = n19857 ^ n5089 ^ 1'b0 ;
  assign n19859 = n3449 & ~n17455 ;
  assign n19860 = n19859 ^ n1839 ^ 1'b0 ;
  assign n19861 = n1082 & n19860 ;
  assign n19862 = n7712 & ~n10686 ;
  assign n19863 = n19862 ^ n1235 ^ 1'b0 ;
  assign n19864 = ~n6286 & n14449 ;
  assign n19865 = ~n1229 & n19864 ;
  assign n19866 = n1914 | n18490 ;
  assign n19867 = n1204 | n19866 ;
  assign n19868 = n19867 ^ n13532 ^ n4582 ;
  assign n19869 = n1314 | n11463 ;
  assign n19870 = n11015 | n19869 ;
  assign n19871 = n3585 & n19685 ;
  assign n19872 = n19871 ^ n3510 ^ 1'b0 ;
  assign n19873 = n13918 | n19872 ;
  assign n19874 = n1851 & n5450 ;
  assign n19875 = ~n616 & n19874 ;
  assign n19876 = n9001 ^ n6539 ^ 1'b0 ;
  assign n19877 = n12641 & ~n19876 ;
  assign n19878 = n19152 ^ n10165 ^ 1'b0 ;
  assign n19879 = n4146 & ~n19878 ;
  assign n19883 = n900 ^ n632 ^ 1'b0 ;
  assign n19882 = ~n6829 & n7606 ;
  assign n19884 = n19883 ^ n19882 ^ 1'b0 ;
  assign n19880 = ~n6740 & n15349 ;
  assign n19881 = n2937 | n19880 ;
  assign n19885 = n19884 ^ n19881 ^ 1'b0 ;
  assign n19886 = n18638 ^ n6180 ^ n6096 ;
  assign n19888 = n1080 & ~n2432 ;
  assign n19887 = n1583 & ~n19275 ;
  assign n19889 = n19888 ^ n19887 ^ 1'b0 ;
  assign n19890 = ( n814 & n9774 ) | ( n814 & n14755 ) | ( n9774 & n14755 ) ;
  assign n19891 = n19890 ^ n3725 ^ 1'b0 ;
  assign n19892 = ~n7046 & n17104 ;
  assign n19893 = ~n4150 & n19892 ;
  assign n19894 = n19893 ^ n5519 ^ 1'b0 ;
  assign n19895 = ~n14022 & n16250 ;
  assign n19896 = n877 & n16222 ;
  assign n19897 = n2318 | n19896 ;
  assign n19898 = n19897 ^ n7625 ^ 1'b0 ;
  assign n19899 = n8145 ^ n4415 ^ 1'b0 ;
  assign n19900 = n5993 | n6376 ;
  assign n19901 = n6173 & n11228 ;
  assign n19902 = n3244 & n19901 ;
  assign n19903 = n3615 & n19902 ;
  assign n19904 = x122 & ~n8518 ;
  assign n19905 = n2789 | n3819 ;
  assign n19906 = n16533 & ~n19905 ;
  assign n19907 = n1161 ^ n1055 ^ 1'b0 ;
  assign n19908 = n10748 & n19907 ;
  assign n19909 = n19908 ^ n4875 ^ 1'b0 ;
  assign n19910 = n4947 | n8625 ;
  assign n19911 = n19910 ^ n2642 ^ 1'b0 ;
  assign n19912 = n8335 ^ n7902 ^ 1'b0 ;
  assign n19913 = n9459 | n19912 ;
  assign n19914 = n19913 ^ n17525 ^ 1'b0 ;
  assign n19915 = n19911 & ~n19914 ;
  assign n19916 = ~n6562 & n15430 ;
  assign n19917 = n4744 ^ n1589 ^ 1'b0 ;
  assign n19918 = n10994 | n14240 ;
  assign n19919 = n5431 ^ n5412 ^ 1'b0 ;
  assign n19920 = n18393 ^ n4190 ^ 1'b0 ;
  assign n19921 = n13783 ^ n457 ^ 1'b0 ;
  assign n19922 = n5261 & ~n19921 ;
  assign n19923 = n8765 ^ n5538 ^ 1'b0 ;
  assign n19924 = n1038 & n5661 ;
  assign n19925 = n3498 & n19924 ;
  assign n19926 = n1351 | n19925 ;
  assign n19927 = n11722 ^ n7547 ^ n3110 ;
  assign n19928 = n10777 & ~n19927 ;
  assign n19929 = n15734 ^ n7439 ^ 1'b0 ;
  assign n19930 = n12013 & ~n19929 ;
  assign n19931 = n14531 ^ n8968 ^ 1'b0 ;
  assign n19932 = n4340 | n13440 ;
  assign n19933 = n12423 ^ n1146 ^ 1'b0 ;
  assign n19934 = n8178 | n19933 ;
  assign n19935 = n19932 & ~n19934 ;
  assign n19936 = n14237 ^ n2068 ^ 1'b0 ;
  assign n19937 = x54 & n19936 ;
  assign n19938 = n19937 ^ n18797 ^ 1'b0 ;
  assign n19939 = x120 & n747 ;
  assign n19940 = ~n14424 & n17104 ;
  assign n19941 = n19940 ^ n17974 ^ 1'b0 ;
  assign n19942 = ~n6817 & n19941 ;
  assign n19943 = ~n1723 & n7391 ;
  assign n19944 = x125 & ~n1746 ;
  assign n19945 = ~n7588 & n19944 ;
  assign n19946 = n13317 ^ n2221 ^ 1'b0 ;
  assign n19947 = ~n733 & n19946 ;
  assign n19948 = n19947 ^ n5028 ^ 1'b0 ;
  assign n19949 = n5434 & n15818 ;
  assign n19950 = n7876 & n15828 ;
  assign n19951 = ~n17084 & n19950 ;
  assign n19952 = n16571 ^ n8956 ^ 1'b0 ;
  assign n19953 = n19952 ^ n8168 ^ n4929 ;
  assign n19954 = n19953 ^ n11084 ^ 1'b0 ;
  assign n19955 = n19951 | n19954 ;
  assign n19956 = n9242 ^ n5336 ^ 1'b0 ;
  assign n19957 = n19907 & ~n19956 ;
  assign n19958 = n11209 | n19957 ;
  assign n19959 = n19958 ^ n359 ^ 1'b0 ;
  assign n19960 = n13182 & n14950 ;
  assign n19961 = n19960 ^ n3089 ^ 1'b0 ;
  assign n19962 = ~n4706 & n19961 ;
  assign n19963 = x106 & ~n10581 ;
  assign n19964 = n19963 ^ n4878 ^ 1'b0 ;
  assign n19965 = n3340 & n18130 ;
  assign n19966 = n19965 ^ n18902 ^ 1'b0 ;
  assign n19967 = n8292 ^ n2555 ^ 1'b0 ;
  assign n19968 = n6016 | n19967 ;
  assign n19969 = n782 ^ n655 ^ 1'b0 ;
  assign n19970 = ~n5223 & n19969 ;
  assign n19971 = n17725 ^ n10086 ^ 1'b0 ;
  assign n19972 = n7282 & ~n19971 ;
  assign n19973 = n19972 ^ n1378 ^ 1'b0 ;
  assign n19974 = n19973 ^ n15894 ^ n10830 ;
  assign n19975 = ~n1782 & n14126 ;
  assign n19976 = n10333 & n15581 ;
  assign n19977 = ~n16131 & n19976 ;
  assign n19979 = n16124 ^ n11516 ^ 1'b0 ;
  assign n19980 = n10748 & ~n19979 ;
  assign n19978 = n1835 | n8188 ;
  assign n19981 = n19980 ^ n19978 ^ 1'b0 ;
  assign n19982 = ~n13880 & n19981 ;
  assign n19983 = ~n16778 & n19982 ;
  assign n19984 = n1137 | n1825 ;
  assign n19985 = n11710 & ~n19984 ;
  assign n19986 = n14569 ^ n2099 ^ 1'b0 ;
  assign n19987 = ~n1290 & n11805 ;
  assign n19988 = ~n5976 & n19987 ;
  assign n19989 = n19795 | n19988 ;
  assign n19990 = n9047 | n13220 ;
  assign n19991 = n8362 & n8702 ;
  assign n19992 = ~n12154 & n19991 ;
  assign n19993 = ~n11946 & n12621 ;
  assign n19994 = n2373 ^ n1409 ^ 1'b0 ;
  assign n19995 = n19994 ^ n14144 ^ 1'b0 ;
  assign n19996 = n14232 ^ n5059 ^ 1'b0 ;
  assign n19997 = n11076 & n19996 ;
  assign n19998 = n11864 ^ n3803 ^ 1'b0 ;
  assign n19999 = ~x56 & n19998 ;
  assign n20000 = n19999 ^ n8772 ^ 1'b0 ;
  assign n20001 = n14619 ^ n13598 ^ 1'b0 ;
  assign n20002 = ~n3403 & n20001 ;
  assign n20003 = n1667 ^ x28 ^ 1'b0 ;
  assign n20004 = n9757 & ~n20003 ;
  assign n20005 = x88 & ~n13094 ;
  assign n20006 = n4242 | n9185 ;
  assign n20007 = n2515 & ~n20006 ;
  assign n20008 = ~n3494 & n5126 ;
  assign n20009 = ~n3632 & n20008 ;
  assign n20010 = ~n2185 & n2756 ;
  assign n20011 = n1139 & ~n6667 ;
  assign n20012 = n20011 ^ n6240 ^ 1'b0 ;
  assign n20013 = n173 | n20012 ;
  assign n20014 = n1035 & ~n4505 ;
  assign n20015 = n20013 & n20014 ;
  assign n20016 = n5059 ^ n4397 ^ x118 ;
  assign n20017 = n11245 ^ n4521 ^ 1'b0 ;
  assign n20018 = n3224 & ~n20017 ;
  assign n20019 = n19721 & ~n20018 ;
  assign n20020 = n14567 & n17568 ;
  assign n20021 = ~n12530 & n20020 ;
  assign n20022 = n4784 | n12654 ;
  assign n20023 = n1626 & n20022 ;
  assign n20024 = n20021 & n20023 ;
  assign n20025 = ~n1290 & n5545 ;
  assign n20026 = n4129 & n14046 ;
  assign n20027 = n14508 & n20026 ;
  assign n20028 = n10028 ^ n5264 ^ 1'b0 ;
  assign n20029 = ( n800 & n1726 ) | ( n800 & n20028 ) | ( n1726 & n20028 ) ;
  assign n20030 = n16020 ^ n7722 ^ 1'b0 ;
  assign n20031 = x60 & n680 ;
  assign n20032 = n12169 ^ n503 ^ 1'b0 ;
  assign n20033 = n20031 & n20032 ;
  assign n20034 = n739 & ~n4759 ;
  assign n20035 = n9042 ^ n7668 ^ n5950 ;
  assign n20036 = n835 & n19426 ;
  assign n20037 = n20036 ^ n19178 ^ 1'b0 ;
  assign n20038 = n3347 ^ n155 ^ 1'b0 ;
  assign n20039 = n20031 & ~n20038 ;
  assign n20040 = n8354 ^ n6565 ^ 1'b0 ;
  assign n20041 = n2608 | n13149 ;
  assign n20042 = n7473 | n20041 ;
  assign n20043 = n3336 | n11788 ;
  assign n20044 = n20043 ^ n8762 ^ 1'b0 ;
  assign n20045 = n20044 ^ n4384 ^ 1'b0 ;
  assign n20046 = n4071 | n8389 ;
  assign n20047 = n20046 ^ n4378 ^ 1'b0 ;
  assign n20048 = n20047 ^ n16553 ^ n6893 ;
  assign n20049 = n9154 ^ n2525 ^ 1'b0 ;
  assign n20050 = n3426 & ~n20049 ;
  assign n20051 = x35 & ~n6206 ;
  assign n20052 = n14474 ^ n12393 ^ 1'b0 ;
  assign n20053 = n7435 | n20052 ;
  assign n20055 = n6563 & n10129 ;
  assign n20056 = n20055 ^ n390 ^ 1'b0 ;
  assign n20054 = ~n9230 & n17416 ;
  assign n20057 = n20056 ^ n20054 ^ 1'b0 ;
  assign n20058 = n7236 & ~n10339 ;
  assign n20059 = n7679 & ~n20058 ;
  assign n20060 = n20059 ^ n7556 ^ 1'b0 ;
  assign n20061 = n14895 | n20060 ;
  assign n20062 = n20061 ^ n3625 ^ 1'b0 ;
  assign n20063 = n7865 ^ n2646 ^ 1'b0 ;
  assign n20064 = n18840 ^ n17966 ^ 1'b0 ;
  assign n20065 = n2649 & ~n6708 ;
  assign n20066 = n20065 ^ n11135 ^ 1'b0 ;
  assign n20067 = n9435 & ~n10710 ;
  assign n20068 = n10207 & ~n20067 ;
  assign n20069 = x70 & ~n9431 ;
  assign n20070 = n20069 ^ n11637 ^ 1'b0 ;
  assign n20071 = ~n2074 & n20070 ;
  assign n20072 = n4817 | n9000 ;
  assign n20073 = n20072 ^ n18578 ^ 1'b0 ;
  assign n20074 = n1832 | n20073 ;
  assign n20075 = n20074 ^ n6159 ^ 1'b0 ;
  assign n20076 = n16242 | n20075 ;
  assign n20077 = n7081 ^ n2168 ^ 1'b0 ;
  assign n20078 = ~n3642 & n20077 ;
  assign n20079 = n2769 ^ n1728 ^ 1'b0 ;
  assign n20080 = n2929 & n2996 ;
  assign n20081 = n17145 & n20080 ;
  assign n20082 = n8053 ^ n852 ^ 1'b0 ;
  assign n20083 = n1789 | n20082 ;
  assign n20084 = x63 & ~n20083 ;
  assign n20085 = n13404 & n20084 ;
  assign n20086 = n482 | n14618 ;
  assign n20087 = n2818 | n20086 ;
  assign n20088 = n4126 & ~n20087 ;
  assign n20089 = ~n3856 & n11176 ;
  assign n20090 = n20089 ^ n3786 ^ 1'b0 ;
  assign n20091 = ( ~n1691 & n3707 ) | ( ~n1691 & n10222 ) | ( n3707 & n10222 ) ;
  assign n20092 = n3619 & ~n20091 ;
  assign n20093 = n8127 & n20092 ;
  assign n20094 = n20093 ^ n3840 ^ 1'b0 ;
  assign n20095 = n7484 & ~n10324 ;
  assign n20096 = n13540 ^ n8501 ^ n5291 ;
  assign n20097 = ~n8644 & n15198 ;
  assign n20098 = n14760 ^ n3742 ^ 1'b0 ;
  assign n20099 = n18431 ^ n846 ^ 1'b0 ;
  assign n20101 = n1864 | n2535 ;
  assign n20100 = n5369 & ~n6554 ;
  assign n20102 = n20101 ^ n20100 ^ 1'b0 ;
  assign n20103 = n20102 ^ n9830 ^ 1'b0 ;
  assign n20104 = n13360 ^ n1786 ^ 1'b0 ;
  assign n20105 = n9785 ^ n3725 ^ 1'b0 ;
  assign n20106 = n5118 & ~n20105 ;
  assign n20107 = n2656 ^ n1170 ^ 1'b0 ;
  assign n20108 = ~n3037 & n3500 ;
  assign n20109 = n20108 ^ n17706 ^ 1'b0 ;
  assign n20110 = n15512 ^ n428 ^ 1'b0 ;
  assign n20116 = ~n222 & n14299 ;
  assign n20111 = n1026 & ~n13212 ;
  assign n20112 = n20111 ^ n1983 ^ 1'b0 ;
  assign n20113 = n16254 & n20112 ;
  assign n20114 = ~n8958 & n20113 ;
  assign n20115 = n16253 | n20114 ;
  assign n20117 = n20116 ^ n20115 ^ 1'b0 ;
  assign n20118 = n5350 ^ n3104 ^ 1'b0 ;
  assign n20119 = n18431 ^ n5327 ^ 1'b0 ;
  assign n20120 = n14006 & n20119 ;
  assign n20121 = n8201 ^ n7777 ^ 1'b0 ;
  assign n20122 = n1274 | n9459 ;
  assign n20123 = n20121 & ~n20122 ;
  assign n20124 = n13472 ^ n4310 ^ 1'b0 ;
  assign n20125 = n13670 ^ n245 ^ 1'b0 ;
  assign n20126 = n5634 ^ n3607 ^ 1'b0 ;
  assign n20127 = n12653 ^ n11437 ^ 1'b0 ;
  assign n20128 = n4821 | n15149 ;
  assign n20129 = n8124 ^ n6876 ^ 1'b0 ;
  assign n20130 = n20128 | n20129 ;
  assign n20131 = n20127 & ~n20130 ;
  assign n20132 = n579 & n20131 ;
  assign n20133 = n7786 | n14399 ;
  assign n20134 = n20133 ^ n9713 ^ 1'b0 ;
  assign n20135 = n1644 & ~n6782 ;
  assign n20136 = ~n18597 & n20135 ;
  assign n20137 = n5885 & ~n20136 ;
  assign n20138 = n11873 & ~n18545 ;
  assign n20139 = n20138 ^ n6642 ^ n4837 ;
  assign n20140 = n6992 ^ n477 ^ 1'b0 ;
  assign n20141 = n877 | n20140 ;
  assign n20142 = ( n20137 & n20139 ) | ( n20137 & ~n20141 ) | ( n20139 & ~n20141 ) ;
  assign n20143 = n2246 | n4821 ;
  assign n20144 = n3083 & n9026 ;
  assign n20145 = n19635 ^ n9345 ^ 1'b0 ;
  assign n20146 = n15437 & ~n16713 ;
  assign n20147 = n1772 & n20146 ;
  assign n20148 = n20147 ^ n12848 ^ 1'b0 ;
  assign n20150 = n13033 ^ n1716 ^ 1'b0 ;
  assign n20149 = ~n6902 & n7475 ;
  assign n20151 = n20150 ^ n20149 ^ 1'b0 ;
  assign n20152 = n15265 | n20151 ;
  assign n20153 = n980 & ~n5306 ;
  assign n20154 = ~n12972 & n20153 ;
  assign n20155 = ~n7387 & n20154 ;
  assign n20156 = n4662 ^ n3998 ^ 1'b0 ;
  assign n20157 = n15582 ^ n7782 ^ 1'b0 ;
  assign n20158 = n1766 | n20157 ;
  assign n20159 = ~n20156 & n20158 ;
  assign n20160 = n3500 & ~n14654 ;
  assign n20161 = n6805 & ~n12426 ;
  assign n20162 = n4691 & ~n7155 ;
  assign n20163 = ~n4691 & n20162 ;
  assign n20164 = n1109 & ~n9986 ;
  assign n20165 = ~n1109 & n20164 ;
  assign n20166 = ~n1131 & n20165 ;
  assign n20167 = n20166 ^ n7836 ^ 1'b0 ;
  assign n20168 = n20163 | n20167 ;
  assign n20169 = n20163 & ~n20168 ;
  assign n20170 = n4296 | n16095 ;
  assign n20171 = n6155 ^ n4929 ^ 1'b0 ;
  assign n20172 = n7158 & n20171 ;
  assign n20173 = n1726 & ~n2838 ;
  assign n20174 = n11064 ^ n5541 ^ 1'b0 ;
  assign n20175 = ~n8400 & n20174 ;
  assign n20176 = x60 & n15836 ;
  assign n20177 = n20176 ^ n14227 ^ 1'b0 ;
  assign n20178 = n4326 & ~n8573 ;
  assign n20179 = n3874 & ~n19087 ;
  assign n20180 = n20179 ^ n4177 ^ 1'b0 ;
  assign n20181 = n19963 ^ n967 ^ 1'b0 ;
  assign n20182 = n6525 & n20181 ;
  assign n20183 = n11865 ^ n3253 ^ 1'b0 ;
  assign n20184 = ~n12785 & n12937 ;
  assign n20185 = n14663 ^ n7792 ^ 1'b0 ;
  assign n20186 = n14731 & n20185 ;
  assign n20187 = n20186 ^ n6186 ^ 1'b0 ;
  assign n20188 = n9091 ^ n4050 ^ 1'b0 ;
  assign n20189 = ~n4204 & n4720 ;
  assign n20190 = ~n3733 & n20189 ;
  assign n20191 = ~n20188 & n20190 ;
  assign n20192 = n13832 & ~n20191 ;
  assign n20193 = n19524 ^ n8945 ^ 1'b0 ;
  assign n20194 = ~n7853 & n20193 ;
  assign n20195 = n13062 ^ n7451 ^ 1'b0 ;
  assign n20196 = ( x54 & n5625 ) | ( x54 & n20195 ) | ( n5625 & n20195 ) ;
  assign n20197 = n6837 ^ n5570 ^ 1'b0 ;
  assign n20198 = n9189 ^ n7554 ^ n210 ;
  assign n20199 = ~n16009 & n18402 ;
  assign n20200 = n811 & n7195 ;
  assign n20201 = ~n3120 & n20200 ;
  assign n20202 = n20201 ^ n10818 ^ 1'b0 ;
  assign n20203 = n1436 | n5470 ;
  assign n20204 = n2129 & n19213 ;
  assign n20205 = n14427 ^ n12348 ^ n3295 ;
  assign n20206 = n20205 ^ n7556 ^ 1'b0 ;
  assign n20207 = n4357 & ~n4513 ;
  assign n20208 = n5183 ^ n2376 ^ 1'b0 ;
  assign n20209 = n963 & ~n8329 ;
  assign n20210 = ~n2456 & n3926 ;
  assign n20211 = n20192 ^ n9132 ^ 1'b0 ;
  assign n20212 = ~n4146 & n12556 ;
  assign n20213 = n1209 & n3358 ;
  assign n20214 = n20213 ^ n3563 ^ 1'b0 ;
  assign n20215 = n333 & ~n2074 ;
  assign n20216 = n1419 & n20215 ;
  assign n20217 = n20214 & n20216 ;
  assign n20218 = n502 | n5336 ;
  assign n20219 = n3805 ^ n882 ^ 1'b0 ;
  assign n20220 = n17286 ^ n6730 ^ 1'b0 ;
  assign n20221 = n10782 & n20220 ;
  assign n20222 = n18890 ^ n851 ^ 1'b0 ;
  assign n20223 = n984 & n10228 ;
  assign n20224 = n1808 & n20223 ;
  assign n20225 = n12065 | n20224 ;
  assign n20226 = n19192 & ~n20225 ;
  assign n20227 = n741 & n3970 ;
  assign n20228 = n13864 ^ n11538 ^ 1'b0 ;
  assign n20229 = n9111 | n20228 ;
  assign n20230 = n4247 | n6540 ;
  assign n20231 = n642 ^ n297 ^ 1'b0 ;
  assign n20232 = ~n1046 & n3829 ;
  assign n20233 = n3585 | n20232 ;
  assign n20234 = n17740 & ~n20233 ;
  assign n20235 = ~n20231 & n20234 ;
  assign n20236 = n999 & n7127 ;
  assign n20237 = n577 | n20236 ;
  assign n20238 = n7288 ^ n2083 ^ 1'b0 ;
  assign n20239 = n14114 ^ n2198 ^ 1'b0 ;
  assign n20240 = n20238 | n20239 ;
  assign n20241 = n7969 ^ n717 ^ 1'b0 ;
  assign n20242 = n20241 ^ n19633 ^ 1'b0 ;
  assign n20243 = n15064 | n20242 ;
  assign n20244 = n2859 & n6282 ;
  assign n20245 = n5512 & n20244 ;
  assign n20246 = n5517 & ~n6333 ;
  assign n20247 = n3401 & ~n20246 ;
  assign n20248 = n1462 & ~n2221 ;
  assign n20249 = n10067 & n20248 ;
  assign n20250 = ~n5430 & n15686 ;
  assign n20251 = n20249 & n20250 ;
  assign n20252 = ~n528 & n6017 ;
  assign n20253 = ( ~n10131 & n17615 ) | ( ~n10131 & n20252 ) | ( n17615 & n20252 ) ;
  assign n20254 = ~n608 & n11976 ;
  assign n20255 = n4163 | n15633 ;
  assign n20256 = n5250 | n5590 ;
  assign n20257 = n1077 | n20256 ;
  assign n20258 = n3900 & n20257 ;
  assign n20259 = n2752 & ~n5453 ;
  assign n20260 = n3549 | n16734 ;
  assign n20261 = n4385 | n20260 ;
  assign n20262 = n12818 & ~n20261 ;
  assign n20263 = n20262 ^ n9692 ^ 1'b0 ;
  assign n20264 = n924 | n12062 ;
  assign n20265 = ~n4433 & n20264 ;
  assign n20266 = n20265 ^ n1328 ^ 1'b0 ;
  assign n20267 = n20266 ^ n17923 ^ 1'b0 ;
  assign n20268 = n5354 & ~n20267 ;
  assign n20269 = n4576 ^ n1071 ^ 1'b0 ;
  assign n20270 = n1908 ^ x13 ^ 1'b0 ;
  assign n20271 = n20269 | n20270 ;
  assign n20272 = n9625 | n20271 ;
  assign n20273 = n20272 ^ n10650 ^ 1'b0 ;
  assign n20274 = n16298 ^ n3916 ^ 1'b0 ;
  assign n20275 = n5797 ^ n5649 ^ n2454 ;
  assign n20276 = n20275 ^ n8978 ^ 1'b0 ;
  assign n20277 = n5234 ^ n5002 ^ 1'b0 ;
  assign n20278 = ~n6435 & n20277 ;
  assign n20279 = ( n8529 & n9285 ) | ( n8529 & ~n19450 ) | ( n9285 & ~n19450 ) ;
  assign n20280 = n4341 | n13559 ;
  assign n20281 = n1837 & n10295 ;
  assign n20282 = n4032 ^ n2243 ^ 1'b0 ;
  assign n20283 = n208 | n20282 ;
  assign n20284 = n20283 ^ n2942 ^ 1'b0 ;
  assign n20285 = ~n489 & n8810 ;
  assign n20286 = n5470 & n20285 ;
  assign n20287 = n4093 & n18167 ;
  assign n20288 = n20286 & n20287 ;
  assign n20289 = n1290 | n5739 ;
  assign n20290 = n9454 | n20289 ;
  assign n20292 = n18081 ^ n1623 ^ 1'b0 ;
  assign n20291 = ~n7773 & n10950 ;
  assign n20293 = n20292 ^ n20291 ^ 1'b0 ;
  assign n20294 = n5052 & n8217 ;
  assign n20295 = n574 & ~n5948 ;
  assign n20296 = n5388 ^ n1211 ^ 1'b0 ;
  assign n20297 = ~n1738 & n20296 ;
  assign n20298 = n6394 & n20297 ;
  assign n20299 = n20298 ^ n16506 ^ 1'b0 ;
  assign n20300 = n16086 ^ n8909 ^ 1'b0 ;
  assign n20301 = ~n4746 & n20300 ;
  assign n20302 = n831 & ~n20214 ;
  assign n20303 = n4505 ^ n666 ^ 1'b0 ;
  assign n20304 = ~n7060 & n10215 ;
  assign n20305 = n1738 & n20304 ;
  assign n20306 = n9704 | n20305 ;
  assign n20307 = n20303 | n20306 ;
  assign n20308 = n1782 | n11016 ;
  assign n20309 = n16783 ^ n391 ^ 1'b0 ;
  assign n20310 = ~n2371 & n9270 ;
  assign n20311 = n20310 ^ n2604 ^ 1'b0 ;
  assign n20312 = n1299 & ~n2718 ;
  assign n20313 = n1587 & n20312 ;
  assign n20314 = ~n4726 & n12634 ;
  assign n20315 = n10064 & n20314 ;
  assign n20316 = n908 & ~n7816 ;
  assign n20317 = n20316 ^ n4867 ^ 1'b0 ;
  assign n20318 = n4659 & n9892 ;
  assign n20319 = n5168 | n6118 ;
  assign n20320 = n20319 ^ n9057 ^ 1'b0 ;
  assign n20321 = ~n2166 & n5658 ;
  assign n20322 = n20321 ^ n6756 ^ 1'b0 ;
  assign n20323 = n2276 | n5019 ;
  assign n20324 = n20322 | n20323 ;
  assign n20325 = n11654 & ~n12267 ;
  assign n20326 = n13749 ^ n7643 ^ 1'b0 ;
  assign n20327 = ~n3037 & n20326 ;
  assign n20328 = n20327 ^ n6401 ^ 1'b0 ;
  assign n20329 = n20328 ^ n13362 ^ 1'b0 ;
  assign n20330 = ~n8235 & n20329 ;
  assign n20331 = n16777 ^ n12472 ^ 1'b0 ;
  assign n20332 = n9528 | n20331 ;
  assign n20333 = ~n1602 & n20332 ;
  assign n20334 = n17030 & ~n20333 ;
  assign n20335 = n20334 ^ n12661 ^ 1'b0 ;
  assign n20336 = n8498 ^ n2584 ^ 1'b0 ;
  assign n20337 = n5950 ^ n609 ^ 1'b0 ;
  assign n20338 = ~n3937 & n20337 ;
  assign n20339 = n1214 ^ x119 ^ 1'b0 ;
  assign n20340 = n20339 ^ n17876 ^ n1937 ;
  assign n20341 = n4691 ^ n2422 ^ n1430 ;
  assign n20342 = n19205 | n20341 ;
  assign n20343 = n17509 ^ n15904 ^ 1'b0 ;
  assign n20344 = n3193 | n20343 ;
  assign n20345 = n4654 ^ n3664 ^ 1'b0 ;
  assign n20346 = n9708 & n20345 ;
  assign n20347 = n3797 & n12095 ;
  assign n20348 = n5500 & n20347 ;
  assign n20349 = n20348 ^ n3140 ^ 1'b0 ;
  assign n20350 = n1222 | n8246 ;
  assign n20351 = n1284 | n20350 ;
  assign n20352 = n20351 ^ n5268 ^ 1'b0 ;
  assign n20353 = n3320 | n20352 ;
  assign n20354 = ~n7670 & n19509 ;
  assign n20355 = n4114 | n10329 ;
  assign n20356 = n10519 | n15147 ;
  assign n20357 = n3367 & n10587 ;
  assign n20358 = n7167 ^ n630 ^ 1'b0 ;
  assign n20359 = ~n20357 & n20358 ;
  assign n20360 = n321 & n7692 ;
  assign n20361 = n1080 | n3116 ;
  assign n20362 = n5278 | n20361 ;
  assign n20363 = n20362 ^ n7892 ^ 1'b0 ;
  assign n20364 = n20360 & n20363 ;
  assign n20365 = ~n5429 & n14633 ;
  assign n20366 = n2299 & n20365 ;
  assign n20367 = ~n7376 & n20366 ;
  assign n20368 = ( ~n5809 & n14994 ) | ( ~n5809 & n15781 ) | ( n14994 & n15781 ) ;
  assign n20369 = n9364 & ~n20368 ;
  assign n20370 = n20369 ^ n10958 ^ 1'b0 ;
  assign n20371 = n4272 & n13063 ;
  assign n20372 = ~n17037 & n20371 ;
  assign n20373 = n6188 ^ n1788 ^ 1'b0 ;
  assign n20374 = n3426 & n5514 ;
  assign n20375 = n20373 & n20374 ;
  assign n20376 = n15025 & ~n20375 ;
  assign n20377 = n1197 ^ n1020 ^ 1'b0 ;
  assign n20378 = n20377 ^ n16932 ^ n2896 ;
  assign n20379 = n17981 ^ n5575 ^ 1'b0 ;
  assign n20380 = n19062 | n20379 ;
  assign n20381 = n984 ^ n261 ^ 1'b0 ;
  assign n20382 = n5717 | n20381 ;
  assign n20383 = n10077 ^ n6098 ^ 1'b0 ;
  assign n20384 = n12609 & n20383 ;
  assign n20385 = n5120 ^ n4117 ^ 1'b0 ;
  assign n20386 = ~n3468 & n4590 ;
  assign n20387 = n20386 ^ n293 ^ 1'b0 ;
  assign n20388 = n20030 & n20387 ;
  assign n20389 = n20388 ^ n4434 ^ 1'b0 ;
  assign n20390 = ( ~n7821 & n8385 ) | ( ~n7821 & n10317 ) | ( n8385 & n10317 ) ;
  assign n20391 = n788 & ~n2592 ;
  assign n20392 = x58 & n290 ;
  assign n20393 = ~x58 & n20392 ;
  assign n20394 = n721 | n20393 ;
  assign n20395 = n721 & ~n20394 ;
  assign n20396 = x41 & n213 ;
  assign n20397 = n20395 & n20396 ;
  assign n20398 = n7866 | n20397 ;
  assign n20399 = n1035 & ~n5144 ;
  assign n20400 = ~n1035 & n20399 ;
  assign n20401 = n634 & n20400 ;
  assign n20402 = n266 & ~n20401 ;
  assign n20403 = n20401 & n20402 ;
  assign n20404 = n588 | n20403 ;
  assign n20405 = n588 & ~n20404 ;
  assign n20406 = n9185 | n20405 ;
  assign n20407 = n20405 & ~n20406 ;
  assign n20408 = n2047 | n3165 ;
  assign n20409 = n2047 & ~n20408 ;
  assign n20410 = x54 & n20409 ;
  assign n20411 = n20407 & n20410 ;
  assign n20412 = n20398 & ~n20411 ;
  assign n20413 = n20412 ^ n4318 ^ 1'b0 ;
  assign n20414 = ~n20391 & n20413 ;
  assign n20415 = n7059 & n9102 ;
  assign n20416 = ~n10622 & n20415 ;
  assign n20417 = n8007 & ~n20416 ;
  assign n20418 = n6043 | n16390 ;
  assign n20419 = n696 | n4135 ;
  assign n20422 = ~n12556 & n18136 ;
  assign n20423 = ~n10033 & n20422 ;
  assign n20420 = n6069 | n10891 ;
  assign n20421 = n9483 | n20420 ;
  assign n20424 = n20423 ^ n20421 ^ 1'b0 ;
  assign n20425 = ~n1361 & n4344 ;
  assign n20426 = n1796 & n20425 ;
  assign n20427 = ~n5143 & n20426 ;
  assign n20428 = n3422 & n19228 ;
  assign n20429 = ~n20427 & n20428 ;
  assign n20430 = n788 & ~n6001 ;
  assign n20431 = ~n1161 & n20430 ;
  assign n20432 = n15509 ^ n12653 ^ 1'b0 ;
  assign n20433 = n10367 ^ n5356 ^ 1'b0 ;
  assign n20434 = ~n5097 & n7437 ;
  assign n20435 = n20433 | n20434 ;
  assign n20436 = n1302 & ~n19370 ;
  assign n20437 = n20436 ^ n20357 ^ 1'b0 ;
  assign n20438 = ( ~n879 & n971 ) | ( ~n879 & n7523 ) | ( n971 & n7523 ) ;
  assign n20439 = n7484 | n20438 ;
  assign n20440 = n272 | n7038 ;
  assign n20441 = n20440 ^ n2533 ^ 1'b0 ;
  assign n20442 = n11573 & n11786 ;
  assign n20443 = n20441 & n20442 ;
  assign n20444 = n9051 | n13543 ;
  assign n20445 = n13217 ^ n9047 ^ 1'b0 ;
  assign n20446 = n20444 & n20445 ;
  assign n20447 = n7573 & ~n10799 ;
  assign n20448 = n2535 | n6575 ;
  assign n20449 = n20447 | n20448 ;
  assign n20450 = n8627 ^ n1981 ^ 1'b0 ;
  assign n20451 = n10609 & n19678 ;
  assign n20452 = n20323 ^ n14584 ^ n12971 ;
  assign n20453 = n4298 & n7900 ;
  assign n20454 = n20453 ^ n173 ^ 1'b0 ;
  assign n20455 = n5347 | n20454 ;
  assign n20456 = n20455 ^ n12408 ^ 1'b0 ;
  assign n20457 = ~n9176 & n15904 ;
  assign n20458 = n20457 ^ n5417 ^ 1'b0 ;
  assign n20459 = n9421 ^ n5979 ^ n146 ;
  assign n20460 = n8249 | n20459 ;
  assign n20461 = n2010 ^ n361 ^ 1'b0 ;
  assign n20462 = n4497 & n20461 ;
  assign n20463 = n2550 & ~n17513 ;
  assign n20464 = x74 | n15231 ;
  assign n20465 = n20464 ^ n7062 ^ 1'b0 ;
  assign n20466 = n6954 & ~n20188 ;
  assign n20467 = n20466 ^ n4902 ^ 1'b0 ;
  assign n20468 = ~n20465 & n20467 ;
  assign n20469 = n9148 & n10018 ;
  assign n20470 = n17350 & n20469 ;
  assign n20471 = n4425 | n20470 ;
  assign n20472 = n4393 & ~n20471 ;
  assign n20473 = n11205 ^ n4576 ^ 1'b0 ;
  assign n20474 = n5247 & ~n20473 ;
  assign n20475 = n5010 & n17006 ;
  assign n20476 = n4507 ^ n2732 ^ 1'b0 ;
  assign n20477 = n20476 ^ n10518 ^ 1'b0 ;
  assign n20478 = n9785 & n14232 ;
  assign n20479 = n20478 ^ n7237 ^ 1'b0 ;
  assign n20480 = n20479 ^ n16020 ^ 1'b0 ;
  assign n20481 = n10776 | n20434 ;
  assign n20482 = n305 | n20481 ;
  assign n20483 = n6001 ^ n4966 ^ 1'b0 ;
  assign n20484 = ~n20015 & n20483 ;
  assign n20485 = ~n6817 & n7615 ;
  assign n20486 = n6114 | n7898 ;
  assign n20487 = n20486 ^ n851 ^ 1'b0 ;
  assign n20488 = n20485 | n20487 ;
  assign n20489 = n6739 & ~n11557 ;
  assign n20490 = n1751 & n20489 ;
  assign n20491 = n237 & n6308 ;
  assign n20492 = n20491 ^ n6931 ^ 1'b0 ;
  assign n20493 = n6244 | n19486 ;
  assign n20494 = n10295 ^ n9151 ^ 1'b0 ;
  assign n20495 = n448 & n20494 ;
  assign n20496 = ~n1887 & n8235 ;
  assign n20497 = ~n2509 & n20496 ;
  assign n20498 = n13948 | n20497 ;
  assign n20499 = n14039 | n20498 ;
  assign n20500 = n15414 ^ n13930 ^ 1'b0 ;
  assign n20501 = n7495 & n13633 ;
  assign n20502 = n2610 & ~n9211 ;
  assign n20503 = n20502 ^ n18502 ^ 1'b0 ;
  assign n20504 = n1574 & ~n8941 ;
  assign n20505 = n2323 | n4976 ;
  assign n20506 = n3288 & ~n20505 ;
  assign n20507 = n6965 & ~n20506 ;
  assign n20508 = n4974 | n16367 ;
  assign n20509 = n13761 | n20508 ;
  assign n20510 = ~n1950 & n19191 ;
  assign n20511 = n6536 & n20510 ;
  assign n20512 = n4061 & ~n20511 ;
  assign n20513 = n9446 & ~n11475 ;
  assign n20514 = n20513 ^ n9749 ^ 1'b0 ;
  assign n20515 = n18010 ^ n6552 ^ n2389 ;
  assign n20516 = n729 & n9019 ;
  assign n20517 = n20516 ^ n15640 ^ 1'b0 ;
  assign n20518 = n4701 & n10486 ;
  assign n20519 = n20518 ^ n6011 ^ 1'b0 ;
  assign n20520 = n6536 & ~n7465 ;
  assign n20521 = n1329 & n3785 ;
  assign n20522 = n20521 ^ n7093 ^ n6448 ;
  assign n20523 = n10975 ^ n10801 ^ 1'b0 ;
  assign n20524 = n8496 ^ n1892 ^ 1'b0 ;
  assign n20525 = ~n10920 & n20524 ;
  assign n20527 = n6869 & ~n9046 ;
  assign n20528 = n20527 ^ n728 ^ 1'b0 ;
  assign n20529 = n141 & n20528 ;
  assign n20530 = n1691 & n15569 ;
  assign n20531 = ~n20529 & n20530 ;
  assign n20526 = n2297 & n9904 ;
  assign n20532 = n20531 ^ n20526 ^ 1'b0 ;
  assign n20533 = n5532 | n8433 ;
  assign n20534 = n10268 | n20533 ;
  assign n20535 = n18839 ^ n8276 ^ 1'b0 ;
  assign n20536 = n9175 ^ n2604 ^ 1'b0 ;
  assign n20538 = x91 & ~n4013 ;
  assign n20539 = n20538 ^ n9421 ^ 1'b0 ;
  assign n20540 = n20539 ^ n2893 ^ 1'b0 ;
  assign n20541 = n7242 & n20540 ;
  assign n20537 = ~n3299 & n9683 ;
  assign n20542 = n20541 ^ n20537 ^ 1'b0 ;
  assign n20543 = n4643 & ~n8596 ;
  assign n20544 = n8909 & n20543 ;
  assign n20545 = n12005 ^ n1703 ^ 1'b0 ;
  assign n20546 = n2471 | n20545 ;
  assign n20547 = n4022 ^ x115 ^ 1'b0 ;
  assign n20548 = n14991 & ~n20547 ;
  assign n20549 = ~x12 & n524 ;
  assign n20550 = ~n12080 & n20549 ;
  assign n20551 = n3454 & n20550 ;
  assign n20552 = n12779 | n17633 ;
  assign n20553 = n1346 & ~n10295 ;
  assign n20554 = n18659 ^ n13266 ^ n7224 ;
  assign n20557 = n11791 & ~n18557 ;
  assign n20555 = n315 & n3272 ;
  assign n20556 = n19092 & ~n20555 ;
  assign n20558 = n20557 ^ n20556 ^ 1'b0 ;
  assign n20559 = n9414 ^ n6772 ^ 1'b0 ;
  assign n20560 = n1964 | n20559 ;
  assign n20561 = n1157 & ~n2722 ;
  assign n20562 = n20561 ^ n6969 ^ 1'b0 ;
  assign n20563 = n20560 | n20562 ;
  assign n20564 = n595 & n3999 ;
  assign n20565 = n9341 ^ n8800 ^ 1'b0 ;
  assign n20566 = ~n20564 & n20565 ;
  assign n20567 = n8512 & n11038 ;
  assign n20568 = n4390 & ~n6727 ;
  assign n20569 = n3831 | n20568 ;
  assign n20570 = x33 & ~n8800 ;
  assign n20571 = n3789 & n20570 ;
  assign n20572 = n10166 ^ n4057 ^ 1'b0 ;
  assign n20573 = n20571 | n20572 ;
  assign n20574 = n4657 | n6419 ;
  assign n20575 = ~n20390 & n20574 ;
  assign n20577 = n863 & ~n5070 ;
  assign n20576 = ~n3677 & n17660 ;
  assign n20578 = n20577 ^ n20576 ^ 1'b0 ;
  assign n20579 = ~n17075 & n17140 ;
  assign n20580 = n20579 ^ n9749 ^ 1'b0 ;
  assign n20581 = n5833 ^ n1903 ^ 1'b0 ;
  assign n20582 = n6259 & n20581 ;
  assign n20583 = n8728 | n14430 ;
  assign n20584 = n7715 & n18343 ;
  assign n20585 = n3290 | n12971 ;
  assign n20586 = n20585 ^ n16096 ^ 1'b0 ;
  assign n20587 = ~n1807 & n4136 ;
  assign n20588 = n5592 & n20587 ;
  assign n20589 = n20588 ^ n1329 ^ 1'b0 ;
  assign n20590 = n3585 | n7980 ;
  assign n20591 = n1067 | n20590 ;
  assign n20592 = n20589 | n20591 ;
  assign n20593 = n17686 ^ n4980 ^ 1'b0 ;
  assign n20594 = ~n11072 & n20593 ;
  assign n20595 = n1627 & n20594 ;
  assign n20596 = n588 & n20595 ;
  assign n20597 = n9174 & ~n14032 ;
  assign n20598 = n4167 & n20597 ;
  assign n20599 = n19285 ^ n1867 ^ 1'b0 ;
  assign n20600 = n952 & n7165 ;
  assign n20601 = ~n504 & n20600 ;
  assign n20602 = n12984 & n20601 ;
  assign n20603 = n3794 & n14839 ;
  assign n20604 = n4942 & ~n8512 ;
  assign n20605 = n3077 ^ n1147 ^ n1013 ;
  assign n20606 = n5429 & ~n20605 ;
  assign n20607 = n7841 & ~n20606 ;
  assign n20608 = n20607 ^ n9235 ^ 1'b0 ;
  assign n20609 = n1774 & n13885 ;
  assign n20610 = n14194 ^ n10481 ^ 1'b0 ;
  assign n20611 = n13041 | n17043 ;
  assign n20612 = n10363 ^ n1781 ^ 1'b0 ;
  assign n20613 = n5223 & n20612 ;
  assign n20614 = n5744 ^ n1498 ^ 1'b0 ;
  assign n20615 = n20613 & n20614 ;
  assign n20616 = ~n830 & n20615 ;
  assign n20617 = ~n9370 & n19485 ;
  assign n20618 = n16671 & ~n20617 ;
  assign n20619 = n12668 & ~n20552 ;
  assign n20620 = ~x84 & n20619 ;
  assign n20621 = n2658 ^ n1663 ^ 1'b0 ;
  assign n20622 = n6310 & ~n20621 ;
  assign n20623 = n20622 ^ n8249 ^ 1'b0 ;
  assign n20624 = n9514 & n20623 ;
  assign n20625 = ~n5023 & n11858 ;
  assign n20626 = n20625 ^ n17530 ^ 1'b0 ;
  assign n20627 = n3966 & ~n19334 ;
  assign n20628 = n20626 & n20627 ;
  assign n20629 = n14134 ^ n9064 ^ 1'b0 ;
  assign n20630 = n14531 ^ n1323 ^ 1'b0 ;
  assign n20631 = n7879 & n14947 ;
  assign n20632 = ~n6034 & n20631 ;
  assign n20633 = n18523 | n20632 ;
  assign n20634 = n7102 & ~n20633 ;
  assign n20635 = ~n18345 & n20634 ;
  assign n20636 = n5878 & ~n18632 ;
  assign n20637 = ~n2932 & n20636 ;
  assign n20640 = n8174 & n13066 ;
  assign n20638 = n526 | n17284 ;
  assign n20639 = n5553 & ~n20638 ;
  assign n20641 = n20640 ^ n20639 ^ n3395 ;
  assign n20642 = n5243 & n5313 ;
  assign n20643 = n20642 ^ n20594 ^ 1'b0 ;
  assign n20644 = n3322 & ~n3468 ;
  assign n20645 = n11076 & n20644 ;
  assign n20646 = n19210 ^ n10096 ^ n3489 ;
  assign n20647 = n835 & n20646 ;
  assign n20648 = n7503 & ~n8445 ;
  assign n20649 = ~n4298 & n12102 ;
  assign n20650 = ~n20648 & n20649 ;
  assign n20651 = n2229 & n3230 ;
  assign n20652 = ~n12147 & n20651 ;
  assign n20653 = x49 & ~n268 ;
  assign n20654 = n20653 ^ n1201 ^ 1'b0 ;
  assign n20655 = n971 ^ n862 ^ 1'b0 ;
  assign n20656 = n7288 ^ n3503 ^ 1'b0 ;
  assign n20657 = n810 & n20656 ;
  assign n20658 = n3651 & n20657 ;
  assign n20659 = n20658 ^ n11255 ^ 1'b0 ;
  assign n20660 = n20659 ^ n14731 ^ 1'b0 ;
  assign n20661 = n16801 ^ n10932 ^ 1'b0 ;
  assign n20662 = n4988 ^ n2809 ^ 1'b0 ;
  assign n20663 = ~n20661 & n20662 ;
  assign n20664 = n9205 & n20663 ;
  assign n20665 = x119 & ~n2636 ;
  assign n20666 = n15357 ^ n5373 ^ 1'b0 ;
  assign n20667 = n221 & ~n20666 ;
  assign n20668 = n4395 & n5667 ;
  assign n20669 = ~n5985 & n20044 ;
  assign n20670 = n889 & n1913 ;
  assign n20671 = n15191 ^ n1706 ^ 1'b0 ;
  assign n20672 = n20670 & ~n20671 ;
  assign n20673 = ~n5048 & n6818 ;
  assign n20674 = n444 & ~n6091 ;
  assign n20675 = n8775 ^ n4236 ^ n643 ;
  assign n20676 = n14807 ^ n13954 ^ 1'b0 ;
  assign n20677 = ~n6069 & n20676 ;
  assign n20678 = n20465 ^ n6579 ^ 1'b0 ;
  assign n20679 = ~n18362 & n20678 ;
  assign n20680 = n3230 & n20679 ;
  assign n20681 = ~n11624 & n20680 ;
  assign n20682 = ~n3473 & n9490 ;
  assign n20683 = n11231 ^ n1060 ^ 1'b0 ;
  assign n20684 = n12793 ^ n3286 ^ 1'b0 ;
  assign n20685 = n9075 & ~n20684 ;
  assign n20686 = n9102 ^ n4638 ^ 1'b0 ;
  assign n20687 = ~n2771 & n20686 ;
  assign n20688 = n1779 & n4429 ;
  assign n20689 = n20688 ^ n6089 ^ 1'b0 ;
  assign n20690 = n20687 & ~n20689 ;
  assign n20691 = n11128 ^ n3286 ^ 1'b0 ;
  assign n20692 = n593 | n20691 ;
  assign n20693 = n8596 | n20692 ;
  assign n20694 = n13972 ^ n8762 ^ n383 ;
  assign n20695 = n5096 & n11843 ;
  assign n20696 = n20694 & n20695 ;
  assign n20698 = x122 & n1035 ;
  assign n20699 = n20698 ^ n4267 ^ 1'b0 ;
  assign n20697 = n392 | n15751 ;
  assign n20700 = n20699 ^ n20697 ^ 1'b0 ;
  assign n20701 = n167 & ~n4731 ;
  assign n20704 = n3037 ^ n1402 ^ 1'b0 ;
  assign n20702 = n5273 & ~n6801 ;
  assign n20703 = n7655 & ~n20702 ;
  assign n20705 = n20704 ^ n20703 ^ n2471 ;
  assign n20706 = n13198 ^ n892 ^ 1'b0 ;
  assign n20707 = n9916 | n11662 ;
  assign n20710 = ~n3422 & n10987 ;
  assign n20711 = n7689 & n20710 ;
  assign n20709 = n410 & n5014 ;
  assign n20712 = n20711 ^ n20709 ^ 1'b0 ;
  assign n20708 = n942 & n12287 ;
  assign n20713 = n20712 ^ n20708 ^ 1'b0 ;
  assign n20714 = n11613 ^ n788 ^ 1'b0 ;
  assign n20715 = n1554 & ~n2165 ;
  assign n20716 = n18474 & n20715 ;
  assign n20717 = n15863 & ~n16711 ;
  assign n20718 = ~n8055 & n9281 ;
  assign n20719 = ~n7996 & n20718 ;
  assign n20720 = ~n10811 & n17854 ;
  assign n20721 = n7374 & n20720 ;
  assign n20722 = n2809 | n10760 ;
  assign n20723 = ~n13428 & n20722 ;
  assign n20724 = ~n11057 & n20723 ;
  assign n20725 = n13049 ^ n428 ^ n283 ;
  assign n20726 = n1026 & n5751 ;
  assign n20727 = n10548 ^ n828 ^ 1'b0 ;
  assign n20728 = ~n20726 & n20727 ;
  assign n20729 = n1479 & ~n4023 ;
  assign n20730 = n3600 & ~n4846 ;
  assign n20731 = n3029 & n20730 ;
  assign n20732 = n20731 ^ n8362 ^ 1'b0 ;
  assign n20733 = n4524 & ~n20732 ;
  assign n20734 = n371 & n3500 ;
  assign n20735 = n1035 & n1228 ;
  assign n20736 = n18178 ^ n2344 ^ 1'b0 ;
  assign n20737 = n20735 & n20736 ;
  assign n20738 = n3648 | n3782 ;
  assign n20739 = n6126 | n20738 ;
  assign n20740 = ~n7935 & n20739 ;
  assign n20741 = n20740 ^ n19582 ^ 1'b0 ;
  assign n20742 = n20741 ^ n10162 ^ n508 ;
  assign n20743 = n6694 & n12771 ;
  assign n20744 = n3611 ^ n1789 ^ 1'b0 ;
  assign n20745 = n14497 & n20744 ;
  assign n20746 = n9787 & n20745 ;
  assign n20747 = n17151 ^ n4500 ^ 1'b0 ;
  assign n20748 = n7986 & ~n17065 ;
  assign n20749 = n3527 ^ n1867 ^ 1'b0 ;
  assign n20750 = n5568 | n20749 ;
  assign n20751 = n19734 ^ n16741 ^ 1'b0 ;
  assign n20752 = ~n19241 & n20751 ;
  assign n20753 = n7462 ^ n4416 ^ 1'b0 ;
  assign n20754 = n4126 & ~n15763 ;
  assign n20755 = n20754 ^ n1908 ^ 1'b0 ;
  assign n20756 = n20755 ^ n13036 ^ n8707 ;
  assign n20757 = n17891 ^ n16759 ^ 1'b0 ;
  assign n20758 = n7237 & n20757 ;
  assign n20759 = n3902 & n20422 ;
  assign n20760 = n1325 | n1552 ;
  assign n20761 = ~n5727 & n8869 ;
  assign n20762 = ~n5685 & n16835 ;
  assign n20763 = ~n20761 & n20762 ;
  assign n20764 = n7134 ^ n6787 ^ 1'b0 ;
  assign n20765 = n11652 & ~n20764 ;
  assign n20766 = ~n1146 & n15749 ;
  assign n20767 = n19562 ^ n6069 ^ 1'b0 ;
  assign n20768 = ~n512 & n4611 ;
  assign n20769 = n10619 & ~n14618 ;
  assign n20770 = n9784 & n20769 ;
  assign n20771 = n1289 & n4832 ;
  assign n20772 = ~n6116 & n20771 ;
  assign n20773 = n11497 ^ n196 ^ 1'b0 ;
  assign n20774 = n5105 ^ n2718 ^ 1'b0 ;
  assign n20775 = n6647 & n20774 ;
  assign n20776 = n12414 & n15737 ;
  assign n20777 = n14319 ^ n1035 ^ 1'b0 ;
  assign n20778 = n20777 ^ n6654 ^ 1'b0 ;
  assign n20779 = n6625 | n20778 ;
  assign n20780 = n5336 & ~n8917 ;
  assign n20781 = n450 & n20780 ;
  assign n20782 = n11533 & ~n20781 ;
  assign n20783 = ~n8581 & n18150 ;
  assign n20784 = ( n409 & n6523 ) | ( n409 & ~n16081 ) | ( n6523 & ~n16081 ) ;
  assign n20785 = n13658 & ~n20784 ;
  assign n20786 = n2312 ^ n1052 ^ 1'b0 ;
  assign n20787 = n3659 ^ n2967 ^ 1'b0 ;
  assign n20788 = ~n20786 & n20787 ;
  assign n20789 = ~n4042 & n19638 ;
  assign n20790 = n1547 & ~n18810 ;
  assign n20791 = n20790 ^ n7590 ^ 1'b0 ;
  assign n20792 = n1726 & ~n7773 ;
  assign n20793 = n1163 | n3419 ;
  assign n20794 = n13360 | n20793 ;
  assign n20795 = n17533 ^ n16671 ^ 1'b0 ;
  assign n20796 = n12672 | n15032 ;
  assign n20797 = n1953 & ~n20796 ;
  assign n20798 = n5139 ^ n353 ^ 1'b0 ;
  assign n20799 = n9898 ^ n8737 ^ 1'b0 ;
  assign n20800 = ~n20798 & n20799 ;
  assign n20801 = n8496 & ~n19531 ;
  assign n20802 = n5186 & ~n20801 ;
  assign n20803 = n20802 ^ n14371 ^ 1'b0 ;
  assign n20804 = n12160 | n15002 ;
  assign n20805 = ~n259 & n1444 ;
  assign n20806 = n16576 & n20805 ;
  assign n20807 = n11288 | n18906 ;
  assign n20808 = n20806 & ~n20807 ;
  assign n20809 = n7001 ^ n922 ^ 1'b0 ;
  assign n20810 = n1996 | n20809 ;
  assign n20811 = n17473 ^ n17145 ^ 1'b0 ;
  assign n20812 = n20810 | n20811 ;
  assign n20813 = n7069 | n7789 ;
  assign n20814 = n307 & ~n3542 ;
  assign n20815 = n3542 & n20814 ;
  assign n20816 = ~n680 & n3286 ;
  assign n20817 = n680 & n20816 ;
  assign n20818 = n5595 & ~n20817 ;
  assign n20819 = n20815 & n20818 ;
  assign n20820 = n20819 ^ n13237 ^ 1'b0 ;
  assign n20821 = ( n7423 & ~n18084 ) | ( n7423 & n20820 ) | ( ~n18084 & n20820 ) ;
  assign n20822 = n9782 & ~n20821 ;
  assign n20823 = n2295 | n2716 ;
  assign n20824 = n20823 ^ n6579 ^ 1'b0 ;
  assign n20825 = ~n707 & n20824 ;
  assign n20826 = n13831 ^ n7683 ^ 1'b0 ;
  assign n20827 = n20825 | n20826 ;
  assign n20828 = n2390 ^ n1095 ^ 1'b0 ;
  assign n20829 = n17157 & n20828 ;
  assign n20830 = n16924 ^ n9895 ^ 1'b0 ;
  assign n20831 = n1548 & ~n20830 ;
  assign n20832 = n20831 ^ n13392 ^ 1'b0 ;
  assign n20833 = ( n2119 & ~n5235 ) | ( n2119 & n19382 ) | ( ~n5235 & n19382 ) ;
  assign n20834 = n17866 ^ n5191 ^ 1'b0 ;
  assign n20835 = n15561 ^ n1281 ^ 1'b0 ;
  assign n20836 = n20834 | n20835 ;
  assign n20837 = n1864 & n5522 ;
  assign n20838 = n18613 ^ n7191 ^ 1'b0 ;
  assign n20839 = n4860 | n5097 ;
  assign n20840 = x62 | n10726 ;
  assign n20841 = n10228 ^ n7364 ^ 1'b0 ;
  assign n20842 = n2091 & ~n20841 ;
  assign n20843 = n3094 & n20842 ;
  assign n20844 = ~n19598 & n20843 ;
  assign n20845 = n7644 ^ n2543 ^ 1'b0 ;
  assign n20846 = n20845 ^ n7171 ^ 1'b0 ;
  assign n20847 = n8573 & n8705 ;
  assign n20848 = n972 & n18295 ;
  assign n20849 = n20847 & n20848 ;
  assign n20850 = ( ~n4430 & n8720 ) | ( ~n4430 & n10329 ) | ( n8720 & n10329 ) ;
  assign n20851 = n14931 ^ n2291 ^ 1'b0 ;
  assign n20852 = n4051 & ~n20851 ;
  assign n20853 = n3278 & n18839 ;
  assign n20854 = n20853 ^ n16877 ^ 1'b0 ;
  assign n20855 = n11688 ^ n1432 ^ 1'b0 ;
  assign n20856 = n5255 & n20855 ;
  assign n20858 = n17462 ^ n11792 ^ 1'b0 ;
  assign n20857 = n7603 & ~n10297 ;
  assign n20859 = n20858 ^ n20857 ^ 1'b0 ;
  assign n20860 = ~n12643 & n20859 ;
  assign n20861 = ~n3548 & n16904 ;
  assign n20862 = n20861 ^ n5258 ^ 1'b0 ;
  assign n20866 = n16788 ^ n9111 ^ 1'b0 ;
  assign n20863 = n2942 & ~n15108 ;
  assign n20864 = n20863 ^ n10630 ^ 1'b0 ;
  assign n20865 = n7803 & n20864 ;
  assign n20867 = n20866 ^ n20865 ^ 1'b0 ;
  assign n20868 = n10850 ^ n1597 ^ 1'b0 ;
  assign n20869 = n7028 & ~n20868 ;
  assign n20870 = ~n17879 & n20869 ;
  assign n20871 = ~n967 & n20870 ;
  assign n20872 = ~n15456 & n20871 ;
  assign n20873 = ~n10214 & n19617 ;
  assign n20874 = ~n988 & n8140 ;
  assign n20875 = n20874 ^ n8217 ^ 1'b0 ;
  assign n20876 = n1281 & n20875 ;
  assign n20877 = n20876 ^ n13878 ^ 1'b0 ;
  assign n20878 = n20877 ^ n7814 ^ 1'b0 ;
  assign n20879 = ~n1329 & n11714 ;
  assign n20880 = n15195 ^ n8961 ^ 1'b0 ;
  assign n20881 = n18650 ^ n5863 ^ 1'b0 ;
  assign n20882 = n2581 | n4095 ;
  assign n20883 = n20882 ^ n10058 ^ 1'b0 ;
  assign n20884 = n20881 & n20883 ;
  assign n20885 = n2787 ^ n2604 ^ 1'b0 ;
  assign n20886 = n20885 ^ n8902 ^ 1'b0 ;
  assign n20887 = ~n13802 & n20886 ;
  assign n20888 = n6975 ^ n4191 ^ 1'b0 ;
  assign n20889 = n20480 ^ n1882 ^ 1'b0 ;
  assign n20890 = n20888 | n20889 ;
  assign n20891 = n768 & n2010 ;
  assign n20892 = n6239 & n11173 ;
  assign n20893 = n17691 & ~n20485 ;
  assign n20894 = ~n20892 & n20893 ;
  assign n20895 = n17315 ^ n10586 ^ 1'b0 ;
  assign n20896 = ~n3908 & n5229 ;
  assign n20897 = ~n6714 & n20896 ;
  assign n20898 = n1825 | n14355 ;
  assign n20899 = n3191 & n4988 ;
  assign n20900 = n12473 | n20323 ;
  assign n20901 = n2530 ^ n2402 ^ 1'b0 ;
  assign n20902 = n4715 & ~n20901 ;
  assign n20903 = n20902 ^ n3302 ^ 1'b0 ;
  assign n20904 = n19287 & ~n20903 ;
  assign n20905 = n7298 & ~n11038 ;
  assign n20906 = n20905 ^ n3969 ^ 1'b0 ;
  assign n20907 = ~n9253 & n14422 ;
  assign n20908 = ~n4621 & n20907 ;
  assign n20909 = ~n6780 & n17581 ;
  assign n20910 = n11568 ^ n5268 ^ 1'b0 ;
  assign n20911 = ~n6851 & n20910 ;
  assign n20912 = ~n9295 & n20777 ;
  assign n20913 = ~n20911 & n20912 ;
  assign n20914 = n18492 & ~n20913 ;
  assign n20915 = n20914 ^ n3998 ^ 1'b0 ;
  assign n20916 = n2641 & n14329 ;
  assign n20917 = ~n5013 & n20916 ;
  assign n20918 = n13826 ^ n5991 ^ 1'b0 ;
  assign n20919 = ~n15070 & n20918 ;
  assign n20920 = n20919 ^ n17392 ^ 1'b0 ;
  assign n20921 = ~n2687 & n5545 ;
  assign n20922 = n20921 ^ n7509 ^ 1'b0 ;
  assign n20923 = n3071 ^ n1982 ^ 1'b0 ;
  assign n20924 = n7683 | n20923 ;
  assign n20925 = n870 & ~n8339 ;
  assign n20926 = n20780 & ~n20925 ;
  assign n20927 = n5023 & ~n13066 ;
  assign n20928 = n2245 | n7655 ;
  assign n20929 = n7832 & ~n20928 ;
  assign n20930 = n17718 & ~n20929 ;
  assign n20931 = n20930 ^ n12626 ^ 1'b0 ;
  assign n20932 = n15932 ^ n12323 ^ n7190 ;
  assign n20933 = n473 | n20932 ;
  assign n20934 = ~n4128 & n18189 ;
  assign n20935 = n19532 & n20934 ;
  assign n20936 = ~n10067 & n20935 ;
  assign n20937 = n19110 | n20936 ;
  assign n20938 = n20937 ^ n18136 ^ 1'b0 ;
  assign n20939 = n1267 | n7708 ;
  assign n20940 = n3658 & n18680 ;
  assign n20941 = ~n20939 & n20940 ;
  assign n20942 = n9042 | n20941 ;
  assign n20943 = n20942 ^ n588 ^ 1'b0 ;
  assign n20944 = n1718 & n20943 ;
  assign n20945 = n2713 | n16162 ;
  assign n20946 = n9459 & ~n20945 ;
  assign n20947 = n704 & n3230 ;
  assign n20948 = n806 & n20947 ;
  assign n20949 = n20948 ^ n496 ^ 1'b0 ;
  assign n20950 = ~n20946 & n20949 ;
  assign n20951 = n3123 & n3824 ;
  assign n20952 = ~n2951 & n20951 ;
  assign n20953 = n700 & ~n8813 ;
  assign n20954 = n5046 & n12504 ;
  assign n20955 = ~n19315 & n20954 ;
  assign n20956 = n632 | n9000 ;
  assign n20957 = ~n20354 & n20956 ;
  assign n20958 = n20955 & n20957 ;
  assign n20959 = n11885 ^ n7798 ^ 1'b0 ;
  assign n20960 = n8205 ^ n4809 ^ 1'b0 ;
  assign n20961 = n7297 & n17625 ;
  assign n20962 = ~n20960 & n20961 ;
  assign n20963 = n9712 | n17614 ;
  assign n20964 = n3483 & ~n12096 ;
  assign n20965 = ~n20963 & n20964 ;
  assign n20966 = n2505 ^ n1724 ^ 1'b0 ;
  assign n20967 = n18573 ^ n1909 ^ 1'b0 ;
  assign n20968 = n8681 ^ n3999 ^ 1'b0 ;
  assign n20969 = n526 & ~n20968 ;
  assign n20970 = n7690 & n20969 ;
  assign n20971 = ~n4507 & n20970 ;
  assign n20972 = n1808 | n5321 ;
  assign n20973 = n20971 & ~n20972 ;
  assign n20974 = n9596 | n20973 ;
  assign n20975 = n20974 ^ n1035 ^ 1'b0 ;
  assign n20976 = n4924 ^ n1543 ^ 1'b0 ;
  assign n20977 = n2859 ^ n1356 ^ 1'b0 ;
  assign n20978 = n4832 & ~n20977 ;
  assign n20979 = n20978 ^ n5613 ^ 1'b0 ;
  assign n20980 = n1484 & n18054 ;
  assign n20981 = n4086 & n13978 ;
  assign n20982 = ~n9034 & n20981 ;
  assign n20983 = n11183 ^ n1502 ^ 1'b0 ;
  assign n20984 = ~n2730 & n20983 ;
  assign n20985 = n20984 ^ n3184 ^ n1344 ;
  assign n20986 = ~n4876 & n10470 ;
  assign n20987 = n3343 & n20986 ;
  assign n20988 = ~n7283 & n17092 ;
  assign n20989 = n15801 & n20988 ;
  assign n20990 = n20989 ^ n6705 ^ 1'b0 ;
  assign n20991 = n3002 & n13217 ;
  assign n20992 = n20991 ^ n5102 ^ 1'b0 ;
  assign n20993 = n3236 ^ n473 ^ 1'b0 ;
  assign n20994 = n5400 | n20993 ;
  assign n20995 = ~n4465 & n16811 ;
  assign n20996 = n13073 ^ n800 ^ 1'b0 ;
  assign n20997 = n9192 ^ n1158 ^ 1'b0 ;
  assign n20998 = ~n9486 & n20997 ;
  assign n20999 = n17541 ^ n7644 ^ 1'b0 ;
  assign n21000 = ~n14508 & n20999 ;
  assign n21001 = n1409 | n2661 ;
  assign n21002 = n9764 & ~n21001 ;
  assign n21003 = n14127 ^ n2929 ^ 1'b0 ;
  assign n21004 = n9082 ^ n6144 ^ 1'b0 ;
  assign n21005 = ~n1201 & n16644 ;
  assign n21006 = n1485 | n1625 ;
  assign n21007 = n21006 ^ n7437 ^ n2393 ;
  assign n21008 = n5652 | n21007 ;
  assign n21009 = n21008 ^ n13726 ^ n4457 ;
  assign n21010 = ~n409 & n21009 ;
  assign n21011 = n5397 ^ n1571 ^ 1'b0 ;
  assign n21012 = n10563 | n21011 ;
  assign n21013 = n15602 ^ n2416 ^ 1'b0 ;
  assign n21015 = n4600 ^ n2439 ^ 1'b0 ;
  assign n21014 = n2710 & ~n6092 ;
  assign n21016 = n21015 ^ n21014 ^ n15743 ;
  assign n21017 = n13955 ^ n7855 ^ 1'b0 ;
  assign n21018 = n19227 ^ n1872 ^ 1'b0 ;
  assign n21019 = ~n14056 & n21018 ;
  assign n21020 = n12924 & ~n17377 ;
  assign n21021 = n21020 ^ n504 ^ 1'b0 ;
  assign n21022 = n16965 ^ n13094 ^ 1'b0 ;
  assign n21023 = ~n12369 & n21022 ;
  assign n21024 = n6880 | n9229 ;
  assign n21025 = n13302 ^ n1993 ^ 1'b0 ;
  assign n21026 = ~n3569 & n21025 ;
  assign n21027 = n21026 ^ n16454 ^ 1'b0 ;
  assign n21028 = n2948 | n7821 ;
  assign n21029 = n6616 & n15939 ;
  assign n21030 = n21029 ^ n9848 ^ 1'b0 ;
  assign n21031 = n6478 & ~n6831 ;
  assign n21032 = n9987 ^ n7374 ^ n6506 ;
  assign n21033 = n12761 ^ n5234 ^ 1'b0 ;
  assign n21034 = n2608 & ~n15386 ;
  assign n21035 = n5545 ^ n2231 ^ 1'b0 ;
  assign n21036 = n806 | n2528 ;
  assign n21037 = n16628 & ~n21036 ;
  assign n21038 = ~n3291 & n5859 ;
  assign n21039 = ~n13976 & n21038 ;
  assign n21040 = n20529 ^ n2584 ^ 1'b0 ;
  assign n21041 = n11111 & ~n21040 ;
  assign n21042 = n21041 ^ x107 ^ 1'b0 ;
  assign n21043 = n11190 & ~n21042 ;
  assign n21044 = x125 & n21043 ;
  assign n21045 = n9600 ^ x5 ^ 1'b0 ;
  assign n21046 = n5033 ^ n2573 ^ 1'b0 ;
  assign n21047 = n17354 ^ n1722 ^ 1'b0 ;
  assign n21048 = n5951 & n21047 ;
  assign n21049 = n8941 & ~n16065 ;
  assign n21050 = n6950 & n21049 ;
  assign n21051 = ~n8533 & n9415 ;
  assign n21052 = n14015 & ~n18933 ;
  assign n21053 = n17796 ^ n16567 ^ n12585 ;
  assign n21054 = n3859 & ~n21053 ;
  assign n21055 = n2432 | n6190 ;
  assign n21056 = n11222 & n21055 ;
  assign n21057 = n21056 ^ n3733 ^ 1'b0 ;
  assign n21058 = n1691 & ~n18936 ;
  assign n21059 = ~n2964 & n21058 ;
  assign n21060 = n1351 ^ n1069 ^ 1'b0 ;
  assign n21061 = n21059 | n21060 ;
  assign n21062 = n5308 & n18188 ;
  assign n21063 = ~n14822 & n21062 ;
  assign n21065 = n4061 | n8773 ;
  assign n21064 = n15289 ^ n2122 ^ 1'b0 ;
  assign n21066 = n21065 ^ n21064 ^ n15070 ;
  assign n21067 = n3030 | n3403 ;
  assign n21068 = n9913 ^ n3869 ^ 1'b0 ;
  assign n21069 = ~n6004 & n21068 ;
  assign n21070 = n1636 ^ n1419 ^ 1'b0 ;
  assign n21071 = n3989 & n21070 ;
  assign n21072 = n7601 ^ n4853 ^ 1'b0 ;
  assign n21073 = ~n7137 & n21072 ;
  assign n21074 = n4840 & n7658 ;
  assign n21075 = ~n3512 & n21074 ;
  assign n21076 = n7134 ^ n6644 ^ 1'b0 ;
  assign n21077 = n2034 & n3819 ;
  assign n21078 = n21077 ^ n11254 ^ 1'b0 ;
  assign n21079 = n4858 | n21078 ;
  assign n21080 = n21079 ^ n2265 ^ 1'b0 ;
  assign n21081 = ~n1226 & n8494 ;
  assign n21082 = ~n4359 & n7625 ;
  assign n21083 = ~n245 & n7798 ;
  assign n21084 = n4964 | n16258 ;
  assign n21085 = n21083 | n21084 ;
  assign n21086 = ~n2803 & n2860 ;
  assign n21087 = n6975 | n19651 ;
  assign n21088 = n21087 ^ n6984 ^ 1'b0 ;
  assign n21089 = n21088 ^ n15828 ^ n2376 ;
  assign n21090 = n15129 & ~n20810 ;
  assign n21091 = n4404 & n21090 ;
  assign n21092 = n5698 & n17586 ;
  assign n21093 = n2344 ^ n216 ^ 1'b0 ;
  assign n21094 = n4323 ^ x122 ^ 1'b0 ;
  assign n21095 = n21093 & ~n21094 ;
  assign n21096 = n7283 & n21095 ;
  assign n21097 = n8608 | n18888 ;
  assign n21098 = n9349 | n10440 ;
  assign n21099 = n8359 | n21098 ;
  assign n21100 = n21099 ^ n8883 ^ 1'b0 ;
  assign n21101 = ~n5472 & n21100 ;
  assign n21102 = n436 & n21101 ;
  assign n21103 = n7633 & ~n19137 ;
  assign n21104 = n21103 ^ n8454 ^ 1'b0 ;
  assign n21105 = n1669 & n21104 ;
  assign n21106 = n15802 ^ n2267 ^ 1'b0 ;
  assign n21107 = n3972 & ~n13120 ;
  assign n21108 = ~x46 & n16084 ;
  assign n21109 = ( ~n2566 & n7093 ) | ( ~n2566 & n11496 ) | ( n7093 & n11496 ) ;
  assign n21110 = x94 & n4983 ;
  assign n21112 = n9429 & ~n10983 ;
  assign n21111 = ~n294 & n6361 ;
  assign n21113 = n21112 ^ n21111 ^ 1'b0 ;
  assign n21114 = n9832 & ~n18488 ;
  assign n21115 = n1658 & ~n2305 ;
  assign n21116 = n5464 | n6716 ;
  assign n21117 = n21115 | n21116 ;
  assign n21118 = n6073 & ~n6268 ;
  assign n21119 = n8986 | n10052 ;
  assign n21120 = n21119 ^ n2266 ^ 1'b0 ;
  assign n21121 = n21120 ^ n2458 ^ 1'b0 ;
  assign n21122 = n4497 & n18084 ;
  assign n21123 = n21122 ^ n1181 ^ 1'b0 ;
  assign n21124 = n21123 ^ n7223 ^ 1'b0 ;
  assign n21125 = n7733 & ~n19415 ;
  assign n21126 = n21125 ^ n10082 ^ 1'b0 ;
  assign n21127 = n21126 ^ n5300 ^ 1'b0 ;
  assign n21128 = ~n8966 & n21127 ;
  assign n21129 = n9749 & ~n17295 ;
  assign n21130 = n3607 & n21129 ;
  assign n21131 = n4897 | n6249 ;
  assign n21132 = n1808 | n13878 ;
  assign n21133 = n21132 ^ n8835 ^ 1'b0 ;
  assign n21134 = n9854 ^ n1232 ^ 1'b0 ;
  assign n21135 = n6383 | n21134 ;
  assign n21136 = n702 & n16046 ;
  assign n21137 = n4106 & n21136 ;
  assign n21138 = n21135 | n21137 ;
  assign n21139 = ~n1944 & n3439 ;
  assign n21140 = n9378 & n12615 ;
  assign n21141 = n5451 & ~n17299 ;
  assign n21142 = ~n579 & n17840 ;
  assign n21143 = n7028 & ~n10630 ;
  assign n21144 = n21143 ^ n10810 ^ 1'b0 ;
  assign n21145 = n10358 & n21144 ;
  assign n21146 = n14664 & ~n19494 ;
  assign n21147 = ~n2253 & n21146 ;
  assign n21148 = n1737 | n4527 ;
  assign n21149 = n810 & ~n15955 ;
  assign n21150 = n1293 | n11517 ;
  assign n21151 = n6022 & ~n21150 ;
  assign n21152 = n11047 ^ n7898 ^ 1'b0 ;
  assign n21153 = n21152 ^ n5613 ^ 1'b0 ;
  assign n21154 = n21151 | n21153 ;
  assign n21155 = n5093 ^ n2532 ^ 1'b0 ;
  assign n21156 = n5315 ^ n4020 ^ 1'b0 ;
  assign n21157 = ~n21155 & n21156 ;
  assign n21158 = n13269 ^ x88 ^ 1'b0 ;
  assign n21159 = n1149 | n13690 ;
  assign n21160 = n10385 & ~n17389 ;
  assign n21161 = n21159 & n21160 ;
  assign n21162 = n5152 & n6439 ;
  assign n21163 = n21162 ^ n3842 ^ 1'b0 ;
  assign n21166 = n442 & n1652 ;
  assign n21167 = ~n1652 & n21166 ;
  assign n21168 = n3702 & n21167 ;
  assign n21164 = n3998 ^ n3479 ^ 1'b0 ;
  assign n21165 = n9316 & ~n21164 ;
  assign n21169 = n21168 ^ n21165 ^ 1'b0 ;
  assign n21170 = ~n4595 & n11281 ;
  assign n21171 = ~n5820 & n21170 ;
  assign n21172 = ~n299 & n21171 ;
  assign n21173 = n363 | n961 ;
  assign n21174 = n21173 ^ n2819 ^ 1'b0 ;
  assign n21175 = ~x52 & n6811 ;
  assign n21176 = n946 | n7719 ;
  assign n21177 = n4908 | n8356 ;
  assign n21178 = n4449 | n21177 ;
  assign n21179 = n5356 | n20232 ;
  assign n21180 = n21179 ^ n6059 ^ 1'b0 ;
  assign n21182 = ~n8182 & n10515 ;
  assign n21183 = n21182 ^ n3902 ^ 1'b0 ;
  assign n21184 = n3726 & ~n21183 ;
  assign n21185 = n21184 ^ n12794 ^ 1'b0 ;
  assign n21181 = n672 & ~n10500 ;
  assign n21186 = n21185 ^ n21181 ^ 1'b0 ;
  assign n21188 = x75 | n496 ;
  assign n21189 = n21188 ^ n1823 ^ 1'b0 ;
  assign n21190 = n21189 ^ n7772 ^ 1'b0 ;
  assign n21187 = n2295 | n8800 ;
  assign n21191 = n21190 ^ n21187 ^ 1'b0 ;
  assign n21192 = ~n8787 & n9413 ;
  assign n21193 = n1244 | n11925 ;
  assign n21194 = n21193 ^ n4307 ^ 1'b0 ;
  assign n21195 = n1439 & n8606 ;
  assign n21196 = ~n3491 & n11580 ;
  assign n21197 = n21195 & ~n21196 ;
  assign n21198 = n3624 & n15904 ;
  assign n21199 = n4618 & ~n14909 ;
  assign n21200 = n19188 & n21199 ;
  assign n21201 = ~n446 & n949 ;
  assign n21202 = n21201 ^ n2051 ^ 1'b0 ;
  assign n21203 = n4880 ^ n3563 ^ n1808 ;
  assign n21204 = ( n9270 & ~n16573 ) | ( n9270 & n21203 ) | ( ~n16573 & n21203 ) ;
  assign n21205 = n8021 & ~n15621 ;
  assign n21206 = n1856 & ~n2085 ;
  assign n21207 = n9214 & n21206 ;
  assign n21208 = n21207 ^ n567 ^ 1'b0 ;
  assign n21209 = n2148 & ~n10717 ;
  assign n21210 = n21209 ^ n8581 ^ 1'b0 ;
  assign n21211 = n4821 & n5050 ;
  assign n21212 = ~n5050 & n21211 ;
  assign n21213 = n5027 & n19176 ;
  assign n21214 = ( ~n8058 & n21212 ) | ( ~n8058 & n21213 ) | ( n21212 & n21213 ) ;
  assign n21215 = n14801 ^ n13290 ^ 1'b0 ;
  assign n21216 = ~n10958 & n21215 ;
  assign n21217 = n13076 ^ n1224 ^ 1'b0 ;
  assign n21218 = n20104 | n21217 ;
  assign n21219 = n9394 & ~n19151 ;
  assign n21220 = ~n16345 & n21219 ;
  assign n21221 = n17954 & ~n20341 ;
  assign n21222 = n21221 ^ n5771 ^ 1'b0 ;
  assign n21223 = n21222 ^ n8459 ^ 1'b0 ;
  assign n21224 = n16801 ^ n6579 ^ n610 ;
  assign n21225 = n21224 ^ n5395 ^ 1'b0 ;
  assign n21226 = n10312 ^ n3831 ^ 1'b0 ;
  assign n21227 = n8699 & ~n21226 ;
  assign n21228 = n2091 & n6782 ;
  assign n21229 = n16882 ^ n9257 ^ 1'b0 ;
  assign n21230 = n967 | n3266 ;
  assign n21231 = ( n528 & ~n1365 ) | ( n528 & n4105 ) | ( ~n1365 & n4105 ) ;
  assign n21232 = n21231 ^ n5329 ^ 1'b0 ;
  assign n21233 = n20231 | n21232 ;
  assign n21234 = n10478 & ~n14124 ;
  assign n21235 = ~n10677 & n16387 ;
  assign n21236 = n6393 ^ n766 ^ 1'b0 ;
  assign n21237 = n1504 & ~n21236 ;
  assign n21238 = n6716 & n14006 ;
  assign n21239 = ~n4167 & n5043 ;
  assign n21240 = n18839 ^ n18464 ^ 1'b0 ;
  assign n21241 = n14991 ^ n1932 ^ 1'b0 ;
  assign n21243 = n2330 | n5530 ;
  assign n21242 = n5144 | n12661 ;
  assign n21244 = n21243 ^ n21242 ^ 1'b0 ;
  assign n21245 = n21244 ^ n7445 ^ 1'b0 ;
  assign n21246 = n5321 | n21245 ;
  assign n21247 = n20549 ^ n8737 ^ n707 ;
  assign n21248 = n4462 & ~n6703 ;
  assign n21249 = n21248 ^ n16810 ^ 1'b0 ;
  assign n21250 = n15124 & ~n21249 ;
  assign n21251 = n21250 ^ n10220 ^ 1'b0 ;
  assign n21252 = n3972 & n12645 ;
  assign n21253 = ~n3552 & n21252 ;
  assign n21254 = n18936 ^ n4668 ^ 1'b0 ;
  assign n21255 = n6330 ^ n5097 ^ 1'b0 ;
  assign n21256 = ~n1226 & n21255 ;
  assign n21257 = n18920 ^ n1204 ^ 1'b0 ;
  assign n21258 = n17120 ^ n1539 ^ 1'b0 ;
  assign n21259 = n8021 & ~n21258 ;
  assign n21260 = x52 & n10512 ;
  assign n21261 = n5791 & ~n16332 ;
  assign n21264 = n4573 ^ n2255 ^ 1'b0 ;
  assign n21262 = ~n677 & n2704 ;
  assign n21263 = n16265 & ~n21262 ;
  assign n21265 = n21264 ^ n21263 ^ 1'b0 ;
  assign n21266 = ~n6554 & n6982 ;
  assign n21267 = ~n6331 & n21266 ;
  assign n21268 = n10840 ^ n8576 ^ 1'b0 ;
  assign n21269 = ( ~n8927 & n13360 ) | ( ~n8927 & n15863 ) | ( n13360 & n15863 ) ;
  assign n21270 = n7548 ^ n806 ^ 1'b0 ;
  assign n21271 = n15388 | n21270 ;
  assign n21272 = n6166 & ~n21271 ;
  assign n21273 = n13993 ^ n7350 ^ 1'b0 ;
  assign n21274 = n7569 & ~n21273 ;
  assign n21275 = n4205 | n9086 ;
  assign n21276 = n8757 ^ n5648 ^ 1'b0 ;
  assign n21277 = n21275 | n21276 ;
  assign n21278 = ~n8636 & n8958 ;
  assign n21279 = n21278 ^ n12090 ^ 1'b0 ;
  assign n21280 = n4563 | n10318 ;
  assign n21281 = n16867 ^ n10385 ^ x15 ;
  assign n21282 = n21280 & n21281 ;
  assign n21283 = n1919 & n19411 ;
  assign n21284 = n988 & ~n7747 ;
  assign n21285 = ~n2985 & n14424 ;
  assign n21286 = ~n21284 & n21285 ;
  assign n21287 = n8340 ^ n3507 ^ 1'b0 ;
  assign n21288 = n21287 ^ n15751 ^ 1'b0 ;
  assign n21289 = n6822 | n10057 ;
  assign n21290 = ~n13737 & n19081 ;
  assign n21291 = n2310 | n14964 ;
  assign n21292 = n9376 | n12212 ;
  assign n21293 = n991 & n13400 ;
  assign n21294 = n15147 & n21293 ;
  assign n21295 = n21294 ^ n3067 ^ 1'b0 ;
  assign n21296 = n3496 ^ n2689 ^ 1'b0 ;
  assign n21297 = n1334 & n17910 ;
  assign n21298 = n6436 | n11955 ;
  assign n21299 = n21298 ^ n20842 ^ 1'b0 ;
  assign n21300 = n12293 ^ n6404 ^ 1'b0 ;
  assign n21301 = ~n21299 & n21300 ;
  assign n21302 = n14368 ^ n4397 ^ 1'b0 ;
  assign n21303 = n14955 ^ n1258 ^ 1'b0 ;
  assign n21304 = n1240 & ~n7440 ;
  assign n21305 = n15458 | n18866 ;
  assign n21306 = n21304 & ~n21305 ;
  assign n21307 = n2780 & ~n5336 ;
  assign n21308 = n21306 & n21307 ;
  assign n21309 = n20255 ^ n17824 ^ 1'b0 ;
  assign n21310 = n5293 | n21309 ;
  assign n21311 = n7172 ^ n5962 ^ 1'b0 ;
  assign n21312 = n5406 | n21311 ;
  assign n21313 = n1443 | n4002 ;
  assign n21314 = ( n8709 & n9293 ) | ( n8709 & n21313 ) | ( n9293 & n21313 ) ;
  assign n21316 = n2584 ^ n614 ^ 1'b0 ;
  assign n21315 = n1020 & ~n2442 ;
  assign n21317 = n21316 ^ n21315 ^ 1'b0 ;
  assign n21318 = n14147 & ~n21317 ;
  assign n21319 = x9 & ~n21318 ;
  assign n21320 = n4019 ^ n3748 ^ 1'b0 ;
  assign n21321 = n12878 & n21320 ;
  assign n21322 = n539 | n5757 ;
  assign n21323 = n21322 ^ n5737 ^ 1'b0 ;
  assign n21324 = n13567 ^ n6499 ^ 1'b0 ;
  assign n21325 = ~n1053 & n11705 ;
  assign n21326 = n21325 ^ n2224 ^ 1'b0 ;
  assign n21327 = n21142 ^ n7297 ^ 1'b0 ;
  assign n21328 = n666 & n11405 ;
  assign n21329 = n21328 ^ n10884 ^ 1'b0 ;
  assign n21330 = n16997 & ~n21329 ;
  assign n21331 = ~n10173 & n20529 ;
  assign n21332 = n7562 & n9413 ;
  assign n21333 = n1624 & n5526 ;
  assign n21334 = ~n12514 & n21333 ;
  assign n21335 = ~n10613 & n11817 ;
  assign n21336 = n1900 & ~n2757 ;
  assign n21337 = n922 & ~n21336 ;
  assign n21338 = n1993 & n16231 ;
  assign n21342 = n1990 | n7140 ;
  assign n21343 = n2041 | n21342 ;
  assign n21339 = ~n2081 & n3376 ;
  assign n21340 = n4817 & n21339 ;
  assign n21341 = n3873 & ~n21340 ;
  assign n21344 = n21343 ^ n21341 ^ 1'b0 ;
  assign n21345 = ~n5090 & n11254 ;
  assign n21346 = n3917 | n21345 ;
  assign n21347 = n1275 | n21346 ;
  assign n21348 = n1642 | n14974 ;
  assign n21349 = n7926 | n13617 ;
  assign n21350 = n4340 ^ n4267 ^ 1'b0 ;
  assign n21351 = n3813 & ~n21350 ;
  assign n21352 = n21351 ^ n10392 ^ 1'b0 ;
  assign n21353 = n782 & n15899 ;
  assign n21354 = n10609 | n20298 ;
  assign n21355 = n8059 & n21354 ;
  assign n21356 = n20754 ^ n221 ^ 1'b0 ;
  assign n21357 = n4918 & ~n21356 ;
  assign n21358 = n7360 & ~n11703 ;
  assign n21359 = ~n2151 & n21358 ;
  assign n21360 = n1558 ^ n323 ^ 1'b0 ;
  assign n21361 = n16762 ^ n9876 ^ 1'b0 ;
  assign n21362 = n3189 & ~n21361 ;
  assign n21363 = n8414 | n12793 ;
  assign n21364 = ~n2792 & n6457 ;
  assign n21365 = n21363 & n21364 ;
  assign n21366 = n9761 | n21365 ;
  assign n21367 = n1786 & ~n21366 ;
  assign n21368 = ~n1158 & n9394 ;
  assign n21369 = n6603 & ~n21368 ;
  assign n21370 = n3041 ^ n1329 ^ 1'b0 ;
  assign n21371 = n1493 | n9910 ;
  assign n21372 = n21371 ^ n3815 ^ 1'b0 ;
  assign n21375 = n2673 ^ n1103 ^ 1'b0 ;
  assign n21376 = ~n2430 & n21375 ;
  assign n21373 = n3925 & n5426 ;
  assign n21374 = n21373 ^ n2555 ^ 1'b0 ;
  assign n21377 = n21376 ^ n21374 ^ 1'b0 ;
  assign n21378 = n21377 ^ n16944 ^ 1'b0 ;
  assign n21379 = n463 & ~n2512 ;
  assign n21380 = ~n545 & n21379 ;
  assign n21381 = n5194 | n21380 ;
  assign n21382 = n2234 | n21381 ;
  assign n21383 = n13686 | n21382 ;
  assign n21384 = ~n8433 & n14196 ;
  assign n21385 = n21384 ^ n11022 ^ 1'b0 ;
  assign n21386 = n14310 ^ n463 ^ 1'b0 ;
  assign n21387 = ~n4416 & n7777 ;
  assign n21390 = ~n297 & n2511 ;
  assign n21388 = n12682 ^ n3589 ^ 1'b0 ;
  assign n21389 = ~n9452 & n21388 ;
  assign n21391 = n21390 ^ n21389 ^ 1'b0 ;
  assign n21392 = ~n4959 & n20458 ;
  assign n21393 = n1779 ^ n1301 ^ 1'b0 ;
  assign n21394 = ~n6537 & n21393 ;
  assign n21395 = n1885 | n15392 ;
  assign n21396 = n4812 & ~n21395 ;
  assign n21397 = n11423 | n12065 ;
  assign n21398 = n21396 & ~n21397 ;
  assign n21399 = n21398 ^ n2418 ^ 1'b0 ;
  assign n21400 = n2385 ^ n2371 ^ 1'b0 ;
  assign n21401 = n4716 & n21400 ;
  assign n21402 = n21401 ^ n8590 ^ 1'b0 ;
  assign n21403 = n19450 ^ n3230 ^ 1'b0 ;
  assign n21404 = n945 | n12357 ;
  assign n21405 = n9566 | n21404 ;
  assign n21406 = n21405 ^ n6448 ^ 1'b0 ;
  assign n21407 = n4310 | n5682 ;
  assign n21408 = n12272 & ~n18607 ;
  assign n21409 = n21408 ^ n3369 ^ 1'b0 ;
  assign n21410 = n20117 & n21409 ;
  assign n21411 = n9782 ^ n2929 ^ 1'b0 ;
  assign n21412 = n4344 ^ n3764 ^ 1'b0 ;
  assign n21413 = n18739 & ~n21412 ;
  assign n21414 = n21413 ^ n9511 ^ 1'b0 ;
  assign n21415 = n2578 & ~n7202 ;
  assign n21416 = n21415 ^ n5647 ^ 1'b0 ;
  assign n21417 = n5404 & ~n18645 ;
  assign n21418 = n156 & n21417 ;
  assign n21419 = ~n16582 & n21418 ;
  assign n21420 = ~n1781 & n11773 ;
  assign n21421 = ~n5683 & n21420 ;
  assign n21422 = n21421 ^ n18385 ^ 1'b0 ;
  assign n21423 = ~n6471 & n15320 ;
  assign n21424 = ~n1133 & n21423 ;
  assign n21425 = n12261 ^ n11350 ^ 1'b0 ;
  assign n21426 = n1798 ^ n192 ^ 1'b0 ;
  assign n21427 = n7927 | n9763 ;
  assign n21428 = n11380 ^ n466 ^ 1'b0 ;
  assign n21429 = n10884 & ~n21428 ;
  assign n21430 = n21429 ^ n1772 ^ 1'b0 ;
  assign n21431 = n16180 ^ n2174 ^ 1'b0 ;
  assign n21432 = n8450 & n21431 ;
  assign n21433 = n20802 ^ n9507 ^ 1'b0 ;
  assign n21434 = n7081 | n12214 ;
  assign n21435 = n7822 ^ n3242 ^ 1'b0 ;
  assign n21436 = n14552 | n21435 ;
  assign y0 = x1 ;
  assign y1 = x2 ;
  assign y2 = x4 ;
  assign y3 = x6 ;
  assign y4 = x8 ;
  assign y5 = x11 ;
  assign y6 = x15 ;
  assign y7 = x18 ;
  assign y8 = x19 ;
  assign y9 = x20 ;
  assign y10 = x24 ;
  assign y11 = x31 ;
  assign y12 = x33 ;
  assign y13 = x37 ;
  assign y14 = x39 ;
  assign y15 = x42 ;
  assign y16 = x43 ;
  assign y17 = x45 ;
  assign y18 = x50 ;
  assign y19 = x57 ;
  assign y20 = x63 ;
  assign y21 = x65 ;
  assign y22 = x66 ;
  assign y23 = x71 ;
  assign y24 = x74 ;
  assign y25 = x76 ;
  assign y26 = x81 ;
  assign y27 = x82 ;
  assign y28 = x85 ;
  assign y29 = x87 ;
  assign y30 = x92 ;
  assign y31 = x96 ;
  assign y32 = x98 ;
  assign y33 = x100 ;
  assign y34 = x102 ;
  assign y35 = x114 ;
  assign y36 = x116 ;
  assign y37 = x117 ;
  assign y38 = x127 ;
  assign y39 = ~n129 ;
  assign y40 = ~1'b0 ;
  assign y41 = ~n131 ;
  assign y42 = ~n132 ;
  assign y43 = ~n134 ;
  assign y44 = n135 ;
  assign y45 = ~1'b0 ;
  assign y46 = n137 ;
  assign y47 = ~1'b0 ;
  assign y48 = n143 ;
  assign y49 = ~1'b0 ;
  assign y50 = ~n144 ;
  assign y51 = ~n148 ;
  assign y52 = n150 ;
  assign y53 = n152 ;
  assign y54 = ~1'b0 ;
  assign y55 = ~n155 ;
  assign y56 = ~1'b0 ;
  assign y57 = n156 ;
  assign y58 = n158 ;
  assign y59 = n159 ;
  assign y60 = ~n164 ;
  assign y61 = ~n171 ;
  assign y62 = ~n177 ;
  assign y63 = n181 ;
  assign y64 = ~n183 ;
  assign y65 = ~n185 ;
  assign y66 = ~1'b0 ;
  assign y67 = ~n189 ;
  assign y68 = n190 ;
  assign y69 = 1'b0 ;
  assign y70 = ~n192 ;
  assign y71 = ~n196 ;
  assign y72 = n205 ;
  assign y73 = ~n208 ;
  assign y74 = ~n211 ;
  assign y75 = ~x106 ;
  assign y76 = ~n216 ;
  assign y77 = n217 ;
  assign y78 = n220 ;
  assign y79 = ~1'b0 ;
  assign y80 = ~1'b0 ;
  assign y81 = n221 ;
  assign y82 = ~n225 ;
  assign y83 = n235 ;
  assign y84 = n237 ;
  assign y85 = ~1'b0 ;
  assign y86 = ~n238 ;
  assign y87 = ~n243 ;
  assign y88 = n248 ;
  assign y89 = ~n251 ;
  assign y90 = ~1'b0 ;
  assign y91 = ~n258 ;
  assign y92 = ~n259 ;
  assign y93 = ~1'b0 ;
  assign y94 = n270 ;
  assign y95 = ~n273 ;
  assign y96 = ~n287 ;
  assign y97 = ~n288 ;
  assign y98 = ~1'b0 ;
  assign y99 = n289 ;
  assign y100 = ~1'b0 ;
  assign y101 = ~1'b0 ;
  assign y102 = ~1'b0 ;
  assign y103 = ~1'b0 ;
  assign y104 = ~1'b0 ;
  assign y105 = ~n292 ;
  assign y106 = ~1'b0 ;
  assign y107 = n293 ;
  assign y108 = ~n294 ;
  assign y109 = ~1'b0 ;
  assign y110 = ~n216 ;
  assign y111 = ~1'b0 ;
  assign y112 = ~n297 ;
  assign y113 = ~n302 ;
  assign y114 = n304 ;
  assign y115 = ~1'b0 ;
  assign y116 = n308 ;
  assign y117 = ~n310 ;
  assign y118 = n311 ;
  assign y119 = ~n315 ;
  assign y120 = ~n318 ;
  assign y121 = ~n320 ;
  assign y122 = ~n324 ;
  assign y123 = n325 ;
  assign y124 = n326 ;
  assign y125 = ~n328 ;
  assign y126 = n333 ;
  assign y127 = ~1'b0 ;
  assign y128 = n335 ;
  assign y129 = n336 ;
  assign y130 = ~n339 ;
  assign y131 = ~n340 ;
  assign y132 = ~1'b0 ;
  assign y133 = ~x66 ;
  assign y134 = n342 ;
  assign y135 = ~1'b0 ;
  assign y136 = ~1'b0 ;
  assign y137 = ~1'b0 ;
  assign y138 = ~n343 ;
  assign y139 = ~1'b0 ;
  assign y140 = ~1'b0 ;
  assign y141 = ~1'b0 ;
  assign y142 = ~n344 ;
  assign y143 = ~n346 ;
  assign y144 = ~1'b0 ;
  assign y145 = n361 ;
  assign y146 = n365 ;
  assign y147 = ~n369 ;
  assign y148 = ~n375 ;
  assign y149 = ~1'b0 ;
  assign y150 = ~n385 ;
  assign y151 = ~1'b0 ;
  assign y152 = n387 ;
  assign y153 = ~n389 ;
  assign y154 = n336 ;
  assign y155 = ~n390 ;
  assign y156 = 1'b0 ;
  assign y157 = ~n391 ;
  assign y158 = n394 ;
  assign y159 = ~1'b0 ;
  assign y160 = ~n399 ;
  assign y161 = ~1'b0 ;
  assign y162 = n400 ;
  assign y163 = ~n406 ;
  assign y164 = n407 ;
  assign y165 = ~1'b0 ;
  assign y166 = n409 ;
  assign y167 = n410 ;
  assign y168 = ~n412 ;
  assign y169 = ~1'b0 ;
  assign y170 = ~1'b0 ;
  assign y171 = ~n413 ;
  assign y172 = ~1'b0 ;
  assign y173 = ~n417 ;
  assign y174 = ~n173 ;
  assign y175 = n418 ;
  assign y176 = n422 ;
  assign y177 = n424 ;
  assign y178 = ~n427 ;
  assign y179 = ~1'b0 ;
  assign y180 = ~1'b0 ;
  assign y181 = ~n430 ;
  assign y182 = ~n435 ;
  assign y183 = n436 ;
  assign y184 = ~n439 ;
  assign y185 = ~n441 ;
  assign y186 = ~n442 ;
  assign y187 = ~n444 ;
  assign y188 = ~n453 ;
  assign y189 = ~1'b0 ;
  assign y190 = ~1'b0 ;
  assign y191 = n456 ;
  assign y192 = n461 ;
  assign y193 = ~n464 ;
  assign y194 = n467 ;
  assign y195 = ~1'b0 ;
  assign y196 = ~n468 ;
  assign y197 = ~n471 ;
  assign y198 = ~n474 ;
  assign y199 = 1'b0 ;
  assign y200 = ~n373 ;
  assign y201 = ~n478 ;
  assign y202 = ~1'b0 ;
  assign y203 = ~n482 ;
  assign y204 = ~1'b0 ;
  assign y205 = ~1'b0 ;
  assign y206 = ~n484 ;
  assign y207 = n487 ;
  assign y208 = ~n491 ;
  assign y209 = n492 ;
  assign y210 = ~n494 ;
  assign y211 = ~n496 ;
  assign y212 = n503 ;
  assign y213 = ~1'b0 ;
  assign y214 = ~1'b0 ;
  assign y215 = ~n506 ;
  assign y216 = ~1'b0 ;
  assign y217 = ~n508 ;
  assign y218 = ~1'b0 ;
  assign y219 = ~1'b0 ;
  assign y220 = ~1'b0 ;
  assign y221 = ~1'b0 ;
  assign y222 = ~n512 ;
  assign y223 = ~n518 ;
  assign y224 = ~1'b0 ;
  assign y225 = ~1'b0 ;
  assign y226 = n520 ;
  assign y227 = ~n522 ;
  assign y228 = n524 ;
  assign y229 = n530 ;
  assign y230 = n531 ;
  assign y231 = ~1'b0 ;
  assign y232 = ~1'b0 ;
  assign y233 = n533 ;
  assign y234 = ~1'b0 ;
  assign y235 = n540 ;
  assign y236 = n547 ;
  assign y237 = ~n548 ;
  assign y238 = ~n549 ;
  assign y239 = ~1'b0 ;
  assign y240 = ~1'b0 ;
  assign y241 = n550 ;
  assign y242 = ~n558 ;
  assign y243 = n562 ;
  assign y244 = n564 ;
  assign y245 = ~n566 ;
  assign y246 = ~n568 ;
  assign y247 = ~1'b0 ;
  assign y248 = ~n571 ;
  assign y249 = ~n574 ;
  assign y250 = ~1'b0 ;
  assign y251 = ~1'b0 ;
  assign y252 = ~1'b0 ;
  assign y253 = ~n575 ;
  assign y254 = 1'b0 ;
  assign y255 = n576 ;
  assign y256 = ~1'b0 ;
  assign y257 = 1'b0 ;
  assign y258 = ~1'b0 ;
  assign y259 = ~n577 ;
  assign y260 = ~1'b0 ;
  assign y261 = ~n579 ;
  assign y262 = ~n487 ;
  assign y263 = ~1'b0 ;
  assign y264 = ~1'b0 ;
  assign y265 = ~1'b0 ;
  assign y266 = ~n360 ;
  assign y267 = ~1'b0 ;
  assign y268 = ~1'b0 ;
  assign y269 = ~n581 ;
  assign y270 = ~n584 ;
  assign y271 = ~n590 ;
  assign y272 = ~1'b0 ;
  assign y273 = ~1'b0 ;
  assign y274 = ~1'b0 ;
  assign y275 = n594 ;
  assign y276 = ~n245 ;
  assign y277 = n597 ;
  assign y278 = ~1'b0 ;
  assign y279 = n608 ;
  assign y280 = n610 ;
  assign y281 = n612 ;
  assign y282 = n613 ;
  assign y283 = ~1'b0 ;
  assign y284 = ~n624 ;
  assign y285 = n629 ;
  assign y286 = ~n497 ;
  assign y287 = ~1'b0 ;
  assign y288 = ~1'b0 ;
  assign y289 = ~n245 ;
  assign y290 = ~n630 ;
  assign y291 = n633 ;
  assign y292 = n634 ;
  assign y293 = ~1'b0 ;
  assign y294 = ~1'b0 ;
  assign y295 = ~1'b0 ;
  assign y296 = ~1'b0 ;
  assign y297 = ~n636 ;
  assign y298 = ~n640 ;
  assign y299 = n647 ;
  assign y300 = ~1'b0 ;
  assign y301 = ~n656 ;
  assign y302 = ~n663 ;
  assign y303 = n665 ;
  assign y304 = ~1'b0 ;
  assign y305 = n666 ;
  assign y306 = n667 ;
  assign y307 = n671 ;
  assign y308 = ~1'b0 ;
  assign y309 = ~1'b0 ;
  assign y310 = ~n675 ;
  assign y311 = n681 ;
  assign y312 = ~n686 ;
  assign y313 = n690 ;
  assign y314 = ~n692 ;
  assign y315 = ~1'b0 ;
  assign y316 = ~n613 ;
  assign y317 = ~n693 ;
  assign y318 = ~n694 ;
  assign y319 = ~1'b0 ;
  assign y320 = ~1'b0 ;
  assign y321 = ~n695 ;
  assign y322 = ~1'b0 ;
  assign y323 = n696 ;
  assign y324 = n698 ;
  assign y325 = n701 ;
  assign y326 = n702 ;
  assign y327 = n703 ;
  assign y328 = ~1'b0 ;
  assign y329 = ~n704 ;
  assign y330 = ~1'b0 ;
  assign y331 = ~1'b0 ;
  assign y332 = ~1'b0 ;
  assign y333 = n705 ;
  assign y334 = ~n713 ;
  assign y335 = ~1'b0 ;
  assign y336 = n716 ;
  assign y337 = ~n720 ;
  assign y338 = n722 ;
  assign y339 = n727 ;
  assign y340 = n728 ;
  assign y341 = ~n571 ;
  assign y342 = n729 ;
  assign y343 = n731 ;
  assign y344 = ~n735 ;
  assign y345 = ~n742 ;
  assign y346 = ~n744 ;
  assign y347 = ~1'b0 ;
  assign y348 = 1'b0 ;
  assign y349 = ~1'b0 ;
  assign y350 = n745 ;
  assign y351 = ~n749 ;
  assign y352 = n750 ;
  assign y353 = ~1'b0 ;
  assign y354 = ~n757 ;
  assign y355 = ~1'b0 ;
  assign y356 = ~1'b0 ;
  assign y357 = ~n761 ;
  assign y358 = n763 ;
  assign y359 = ~n764 ;
  assign y360 = ~n770 ;
  assign y361 = ~1'b0 ;
  assign y362 = n775 ;
  assign y363 = ~n778 ;
  assign y364 = ~1'b0 ;
  assign y365 = n782 ;
  assign y366 = ~1'b0 ;
  assign y367 = ~n785 ;
  assign y368 = ~n788 ;
  assign y369 = ~n793 ;
  assign y370 = n794 ;
  assign y371 = ~n801 ;
  assign y372 = ~1'b0 ;
  assign y373 = n245 ;
  assign y374 = n802 ;
  assign y375 = ~1'b0 ;
  assign y376 = ~n805 ;
  assign y377 = ~1'b0 ;
  assign y378 = ~n806 ;
  assign y379 = n808 ;
  assign y380 = ~1'b0 ;
  assign y381 = ~1'b0 ;
  assign y382 = ~1'b0 ;
  assign y383 = ~n809 ;
  assign y384 = ~1'b0 ;
  assign y385 = ~1'b0 ;
  assign y386 = n810 ;
  assign y387 = x104 ;
  assign y388 = n237 ;
  assign y389 = n813 ;
  assign y390 = ~1'b0 ;
  assign y391 = n814 ;
  assign y392 = ~n824 ;
  assign y393 = ~1'b0 ;
  assign y394 = n825 ;
  assign y395 = ~1'b0 ;
  assign y396 = n826 ;
  assign y397 = n833 ;
  assign y398 = ~1'b0 ;
  assign y399 = ~n836 ;
  assign y400 = n788 ;
  assign y401 = ~n837 ;
  assign y402 = ~1'b0 ;
  assign y403 = n841 ;
  assign y404 = ~n842 ;
  assign y405 = n844 ;
  assign y406 = n845 ;
  assign y407 = n846 ;
  assign y408 = ~1'b0 ;
  assign y409 = ~1'b0 ;
  assign y410 = ~n853 ;
  assign y411 = ~n510 ;
  assign y412 = ~n854 ;
  assign y413 = n855 ;
  assign y414 = x54 ;
  assign y415 = n858 ;
  assign y416 = ~1'b0 ;
  assign y417 = n861 ;
  assign y418 = ~n866 ;
  assign y419 = ~n867 ;
  assign y420 = ~n868 ;
  assign y421 = n869 ;
  assign y422 = n870 ;
  assign y423 = n876 ;
  assign y424 = n877 ;
  assign y425 = ~1'b0 ;
  assign y426 = ~n879 ;
  assign y427 = n880 ;
  assign y428 = ~n428 ;
  assign y429 = ~n885 ;
  assign y430 = ~1'b0 ;
  assign y431 = n888 ;
  assign y432 = ~n889 ;
  assign y433 = ~n890 ;
  assign y434 = 1'b0 ;
  assign y435 = ~1'b0 ;
  assign y436 = n891 ;
  assign y437 = ~n892 ;
  assign y438 = ~n893 ;
  assign y439 = ~n894 ;
  assign y440 = ~1'b0 ;
  assign y441 = ~n896 ;
  assign y442 = n558 ;
  assign y443 = ~1'b0 ;
  assign y444 = ~n897 ;
  assign y445 = n806 ;
  assign y446 = ~1'b0 ;
  assign y447 = ~n259 ;
  assign y448 = ~1'b0 ;
  assign y449 = ~1'b0 ;
  assign y450 = ~n902 ;
  assign y451 = ~1'b0 ;
  assign y452 = ~1'b0 ;
  assign y453 = n165 ;
  assign y454 = ~1'b0 ;
  assign y455 = ~1'b0 ;
  assign y456 = n905 ;
  assign y457 = n908 ;
  assign y458 = ~n911 ;
  assign y459 = n912 ;
  assign y460 = ~n921 ;
  assign y461 = ~n924 ;
  assign y462 = n936 ;
  assign y463 = ~1'b0 ;
  assign y464 = n938 ;
  assign y465 = n939 ;
  assign y466 = ~1'b0 ;
  assign y467 = ~1'b0 ;
  assign y468 = ~n733 ;
  assign y469 = ~n945 ;
  assign y470 = ~n946 ;
  assign y471 = ~1'b0 ;
  assign y472 = n613 ;
  assign y473 = n949 ;
  assign y474 = ~1'b0 ;
  assign y475 = ~n950 ;
  assign y476 = ~1'b0 ;
  assign y477 = ~1'b0 ;
  assign y478 = n952 ;
  assign y479 = ~n956 ;
  assign y480 = ~n958 ;
  assign y481 = ~1'b0 ;
  assign y482 = ~1'b0 ;
  assign y483 = ~1'b0 ;
  assign y484 = ~n960 ;
  assign y485 = ~1'b0 ;
  assign y486 = ~n961 ;
  assign y487 = ~n969 ;
  assign y488 = n974 ;
  assign y489 = ~n975 ;
  assign y490 = ~n978 ;
  assign y491 = n981 ;
  assign y492 = n482 ;
  assign y493 = ~n983 ;
  assign y494 = n984 ;
  assign y495 = n985 ;
  assign y496 = ~1'b0 ;
  assign y497 = n307 ;
  assign y498 = ~1'b0 ;
  assign y499 = ~1'b0 ;
  assign y500 = ~n986 ;
  assign y501 = ~n988 ;
  assign y502 = ~1'b0 ;
  assign y503 = ~1'b0 ;
  assign y504 = ~1'b0 ;
  assign y505 = x77 ;
  assign y506 = ~1'b0 ;
  assign y507 = ~n989 ;
  assign y508 = ~1'b0 ;
  assign y509 = ~1'b0 ;
  assign y510 = n991 ;
  assign y511 = ~1'b0 ;
  assign y512 = ~n995 ;
  assign y513 = ~n307 ;
  assign y514 = ~1'b0 ;
  assign y515 = ~1'b0 ;
  assign y516 = ~1'b0 ;
  assign y517 = ~1'b0 ;
  assign y518 = ~1'b0 ;
  assign y519 = 1'b0 ;
  assign y520 = ~1'b0 ;
  assign y521 = ~n983 ;
  assign y522 = ~1'b0 ;
  assign y523 = n998 ;
  assign y524 = ~n1004 ;
  assign y525 = n1008 ;
  assign y526 = n926 ;
  assign y527 = n1012 ;
  assign y528 = ~x12 ;
  assign y529 = ~n1013 ;
  assign y530 = ~n1018 ;
  assign y531 = ~1'b0 ;
  assign y532 = ~x82 ;
  assign y533 = ~n1025 ;
  assign y534 = n1026 ;
  assign y535 = ~n1031 ;
  assign y536 = ~n1033 ;
  assign y537 = ~n1041 ;
  assign y538 = ~n1052 ;
  assign y539 = ~n1056 ;
  assign y540 = ~n1063 ;
  assign y541 = ~x75 ;
  assign y542 = ~n1067 ;
  assign y543 = ~n1072 ;
  assign y544 = n1077 ;
  assign y545 = n1079 ;
  assign y546 = n1082 ;
  assign y547 = ~n1084 ;
  assign y548 = 1'b0 ;
  assign y549 = n1087 ;
  assign y550 = ~1'b0 ;
  assign y551 = ~n1092 ;
  assign y552 = n1093 ;
  assign y553 = ~n1101 ;
  assign y554 = ~n1102 ;
  assign y555 = ~1'b0 ;
  assign y556 = n1103 ;
  assign y557 = ~1'b0 ;
  assign y558 = ~n1051 ;
  assign y559 = ~1'b0 ;
  assign y560 = ~n1105 ;
  assign y561 = ~n1106 ;
  assign y562 = ~n1107 ;
  assign y563 = ~n1116 ;
  assign y564 = ~n1118 ;
  assign y565 = n1122 ;
  assign y566 = n1124 ;
  assign y567 = ~n1126 ;
  assign y568 = ~1'b0 ;
  assign y569 = ~1'b0 ;
  assign y570 = ~1'b0 ;
  assign y571 = ~1'b0 ;
  assign y572 = ~n1129 ;
  assign y573 = ~1'b0 ;
  assign y574 = ~1'b0 ;
  assign y575 = ~1'b0 ;
  assign y576 = ~n1133 ;
  assign y577 = n1137 ;
  assign y578 = ~1'b0 ;
  assign y579 = n1139 ;
  assign y580 = ~1'b0 ;
  assign y581 = ~1'b0 ;
  assign y582 = ~n1141 ;
  assign y583 = ~n1144 ;
  assign y584 = ~1'b0 ;
  assign y585 = n1156 ;
  assign y586 = ~1'b0 ;
  assign y587 = ~n1158 ;
  assign y588 = n1160 ;
  assign y589 = ~x40 ;
  assign y590 = n1162 ;
  assign y591 = ~n1163 ;
  assign y592 = n1165 ;
  assign y593 = n1169 ;
  assign y594 = ~1'b0 ;
  assign y595 = ~n1172 ;
  assign y596 = ~1'b0 ;
  assign y597 = n1173 ;
  assign y598 = n1178 ;
  assign y599 = ~n1183 ;
  assign y600 = ~n1185 ;
  assign y601 = ~1'b0 ;
  assign y602 = n1188 ;
  assign y603 = ~1'b0 ;
  assign y604 = n1189 ;
  assign y605 = ~n1192 ;
  assign y606 = ~n1194 ;
  assign y607 = ~n1195 ;
  assign y608 = ~n1197 ;
  assign y609 = n1199 ;
  assign y610 = ~n1201 ;
  assign y611 = ~1'b0 ;
  assign y612 = n1202 ;
  assign y613 = n1203 ;
  assign y614 = ~1'b0 ;
  assign y615 = n1205 ;
  assign y616 = ~1'b0 ;
  assign y617 = ~1'b0 ;
  assign y618 = ~1'b0 ;
  assign y619 = ~n1207 ;
  assign y620 = ~n1208 ;
  assign y621 = n1211 ;
  assign y622 = ~n1219 ;
  assign y623 = ~1'b0 ;
  assign y624 = ~n1221 ;
  assign y625 = ~n1226 ;
  assign y626 = ~n1229 ;
  assign y627 = ~n1234 ;
  assign y628 = ~1'b0 ;
  assign y629 = ~n1235 ;
  assign y630 = n1236 ;
  assign y631 = ~n806 ;
  assign y632 = n1241 ;
  assign y633 = ~n1243 ;
  assign y634 = ~n1249 ;
  assign y635 = ~n1253 ;
  assign y636 = 1'b0 ;
  assign y637 = n1254 ;
  assign y638 = ~n1258 ;
  assign y639 = ~n427 ;
  assign y640 = 1'b0 ;
  assign y641 = ~n1265 ;
  assign y642 = ~1'b0 ;
  assign y643 = ~n1270 ;
  assign y644 = ~1'b0 ;
  assign y645 = n1273 ;
  assign y646 = ~n1274 ;
  assign y647 = ~n1277 ;
  assign y648 = n512 ;
  assign y649 = ~n1279 ;
  assign y650 = n1280 ;
  assign y651 = n1281 ;
  assign y652 = ~n1287 ;
  assign y653 = ~n1290 ;
  assign y654 = ~n1292 ;
  assign y655 = ~n1295 ;
  assign y656 = ~1'b0 ;
  assign y657 = ~n1298 ;
  assign y658 = ~1'b0 ;
  assign y659 = ~1'b0 ;
  assign y660 = n1299 ;
  assign y661 = ~n1301 ;
  assign y662 = n1302 ;
  assign y663 = n1303 ;
  assign y664 = n1308 ;
  assign y665 = ~1'b0 ;
  assign y666 = 1'b0 ;
  assign y667 = ~n1314 ;
  assign y668 = ~n1315 ;
  assign y669 = ~n1319 ;
  assign y670 = n1323 ;
  assign y671 = ~n1137 ;
  assign y672 = n1270 ;
  assign y673 = ~1'b0 ;
  assign y674 = ~1'b0 ;
  assign y675 = ~1'b0 ;
  assign y676 = ~1'b0 ;
  assign y677 = ~1'b0 ;
  assign y678 = ~1'b0 ;
  assign y679 = n1324 ;
  assign y680 = n323 ;
  assign y681 = n1325 ;
  assign y682 = n1334 ;
  assign y683 = n1221 ;
  assign y684 = ~n1340 ;
  assign y685 = ~n830 ;
  assign y686 = ~1'b0 ;
  assign y687 = ~n1348 ;
  assign y688 = ~1'b0 ;
  assign y689 = ~n1349 ;
  assign y690 = n1351 ;
  assign y691 = ~1'b0 ;
  assign y692 = n1352 ;
  assign y693 = n1355 ;
  assign y694 = ~1'b0 ;
  assign y695 = n1356 ;
  assign y696 = ~n1360 ;
  assign y697 = ~n1363 ;
  assign y698 = ~n544 ;
  assign y699 = ~1'b0 ;
  assign y700 = ~1'b0 ;
  assign y701 = ~n747 ;
  assign y702 = n1364 ;
  assign y703 = ~n1368 ;
  assign y704 = ~n1369 ;
  assign y705 = ~n1374 ;
  assign y706 = ~1'b0 ;
  assign y707 = n262 ;
  assign y708 = ~n1376 ;
  assign y709 = n1380 ;
  assign y710 = ~1'b0 ;
  assign y711 = n1381 ;
  assign y712 = ~1'b0 ;
  assign y713 = ~n1387 ;
  assign y714 = n1394 ;
  assign y715 = ~n1395 ;
  assign y716 = ~n1398 ;
  assign y717 = ~1'b0 ;
  assign y718 = ~1'b0 ;
  assign y719 = ~n1402 ;
  assign y720 = ~n1410 ;
  assign y721 = n1414 ;
  assign y722 = ~n1415 ;
  assign y723 = ~1'b0 ;
  assign y724 = ~n1416 ;
  assign y725 = ~n1419 ;
  assign y726 = n1420 ;
  assign y727 = ~n391 ;
  assign y728 = n978 ;
  assign y729 = n1425 ;
  assign y730 = ~1'b0 ;
  assign y731 = n1428 ;
  assign y732 = n1434 ;
  assign y733 = ~n1436 ;
  assign y734 = ~1'b0 ;
  assign y735 = ~n1437 ;
  assign y736 = ~1'b0 ;
  assign y737 = n1446 ;
  assign y738 = ~n1451 ;
  assign y739 = ~n1455 ;
  assign y740 = n1456 ;
  assign y741 = n1020 ;
  assign y742 = ~n1457 ;
  assign y743 = ~1'b0 ;
  assign y744 = ~n1461 ;
  assign y745 = ~1'b0 ;
  assign y746 = ~1'b0 ;
  assign y747 = ~n1463 ;
  assign y748 = ~1'b0 ;
  assign y749 = n1469 ;
  assign y750 = n1470 ;
  assign y751 = ~n1472 ;
  assign y752 = ~1'b0 ;
  assign y753 = ~n1474 ;
  assign y754 = n1475 ;
  assign y755 = n1477 ;
  assign y756 = n1478 ;
  assign y757 = n1480 ;
  assign y758 = ~n1482 ;
  assign y759 = n1484 ;
  assign y760 = ~1'b0 ;
  assign y761 = ~1'b0 ;
  assign y762 = ~n1485 ;
  assign y763 = ~n1487 ;
  assign y764 = ~1'b0 ;
  assign y765 = ~1'b0 ;
  assign y766 = ~n1493 ;
  assign y767 = n1495 ;
  assign y768 = ~n1496 ;
  assign y769 = n1497 ;
  assign y770 = ~n1498 ;
  assign y771 = ~1'b0 ;
  assign y772 = ~1'b0 ;
  assign y773 = n1499 ;
  assign y774 = n1502 ;
  assign y775 = ~n1513 ;
  assign y776 = ~1'b0 ;
  assign y777 = ~n1525 ;
  assign y778 = n1329 ;
  assign y779 = ~1'b0 ;
  assign y780 = ~n1532 ;
  assign y781 = ~n1534 ;
  assign y782 = ~n1536 ;
  assign y783 = n446 ;
  assign y784 = n1245 ;
  assign y785 = ~n1537 ;
  assign y786 = n1539 ;
  assign y787 = 1'b0 ;
  assign y788 = n1103 ;
  assign y789 = n1540 ;
  assign y790 = ~1'b0 ;
  assign y791 = 1'b0 ;
  assign y792 = n1542 ;
  assign y793 = ~n1543 ;
  assign y794 = ~n1545 ;
  assign y795 = n1547 ;
  assign y796 = ~1'b0 ;
  assign y797 = ~1'b0 ;
  assign y798 = ~n1554 ;
  assign y799 = ~n1561 ;
  assign y800 = n1564 ;
  assign y801 = n1566 ;
  assign y802 = ~1'b0 ;
  assign y803 = ~1'b0 ;
  assign y804 = ~n1569 ;
  assign y805 = ~n1572 ;
  assign y806 = ~1'b0 ;
  assign y807 = ~n1578 ;
  assign y808 = n1580 ;
  assign y809 = n1581 ;
  assign y810 = n1583 ;
  assign y811 = n1587 ;
  assign y812 = n1590 ;
  assign y813 = ~1'b0 ;
  assign y814 = ~n1592 ;
  assign y815 = n1534 ;
  assign y816 = n1595 ;
  assign y817 = n1602 ;
  assign y818 = ~n1608 ;
  assign y819 = ~1'b0 ;
  assign y820 = 1'b0 ;
  assign y821 = n1610 ;
  assign y822 = ~n1612 ;
  assign y823 = ~1'b0 ;
  assign y824 = ~n1613 ;
  assign y825 = ~1'b0 ;
  assign y826 = ~1'b0 ;
  assign y827 = ~n1616 ;
  assign y828 = ~n1622 ;
  assign y829 = n1624 ;
  assign y830 = ~1'b0 ;
  assign y831 = 1'b0 ;
  assign y832 = ~1'b0 ;
  assign y833 = ~1'b0 ;
  assign y834 = n1626 ;
  assign y835 = n1627 ;
  assign y836 = n1632 ;
  assign y837 = ~1'b0 ;
  assign y838 = ~n1636 ;
  assign y839 = n1639 ;
  assign y840 = ~1'b0 ;
  assign y841 = n1644 ;
  assign y842 = ~n1645 ;
  assign y843 = ~1'b0 ;
  assign y844 = ~n1648 ;
  assign y845 = ~1'b0 ;
  assign y846 = n1650 ;
  assign y847 = ~1'b0 ;
  assign y848 = ~n1651 ;
  assign y849 = n1652 ;
  assign y850 = ~1'b0 ;
  assign y851 = 1'b0 ;
  assign y852 = ~1'b0 ;
  assign y853 = n1662 ;
  assign y854 = ~n1664 ;
  assign y855 = ~1'b0 ;
  assign y856 = ~n1667 ;
  assign y857 = ~n1668 ;
  assign y858 = n1669 ;
  assign y859 = ~1'b0 ;
  assign y860 = n1673 ;
  assign y861 = n1674 ;
  assign y862 = ~n1675 ;
  assign y863 = ~1'b0 ;
  assign y864 = ~1'b0 ;
  assign y865 = ~1'b0 ;
  assign y866 = ~1'b0 ;
  assign y867 = ~1'b0 ;
  assign y868 = ~n636 ;
  assign y869 = 1'b0 ;
  assign y870 = ~n1677 ;
  assign y871 = ~n1680 ;
  assign y872 = n1681 ;
  assign y873 = n1685 ;
  assign y874 = ~n1688 ;
  assign y875 = n1692 ;
  assign y876 = n1693 ;
  assign y877 = ~n1703 ;
  assign y878 = n1704 ;
  assign y879 = ~n1707 ;
  assign y880 = ~1'b0 ;
  assign y881 = 1'b0 ;
  assign y882 = ~1'b0 ;
  assign y883 = n1710 ;
  assign y884 = n1713 ;
  assign y885 = n1716 ;
  assign y886 = ~n1720 ;
  assign y887 = ~1'b0 ;
  assign y888 = ~1'b0 ;
  assign y889 = ~n1722 ;
  assign y890 = ~n1724 ;
  assign y891 = ~1'b0 ;
  assign y892 = ~n1728 ;
  assign y893 = ~n1731 ;
  assign y894 = n1736 ;
  assign y895 = ~1'b0 ;
  assign y896 = ~n1738 ;
  assign y897 = ~1'b0 ;
  assign y898 = ~1'b0 ;
  assign y899 = ~1'b0 ;
  assign y900 = n1747 ;
  assign y901 = ~n1753 ;
  assign y902 = ~n1755 ;
  assign y903 = 1'b0 ;
  assign y904 = ~1'b0 ;
  assign y905 = ~n163 ;
  assign y906 = ~1'b0 ;
  assign y907 = ~1'b0 ;
  assign y908 = n1756 ;
  assign y909 = n1761 ;
  assign y910 = ~n1764 ;
  assign y911 = ~1'b0 ;
  assign y912 = ~1'b0 ;
  assign y913 = ~n1766 ;
  assign y914 = ~n1770 ;
  assign y915 = ~1'b0 ;
  assign y916 = n1534 ;
  assign y917 = ~1'b0 ;
  assign y918 = n1773 ;
  assign y919 = n1774 ;
  assign y920 = n1777 ;
  assign y921 = ~1'b0 ;
  assign y922 = n562 ;
  assign y923 = ~n1779 ;
  assign y924 = n1781 ;
  assign y925 = ~1'b0 ;
  assign y926 = ~n1782 ;
  assign y927 = ~n1498 ;
  assign y928 = n1784 ;
  assign y929 = ~n1789 ;
  assign y930 = n1790 ;
  assign y931 = ~n1805 ;
  assign y932 = ~n1807 ;
  assign y933 = ~n1808 ;
  assign y934 = ~n1030 ;
  assign y935 = ~n1811 ;
  assign y936 = ~n1814 ;
  assign y937 = n1816 ;
  assign y938 = n1817 ;
  assign y939 = ~1'b0 ;
  assign y940 = n1819 ;
  assign y941 = ~1'b0 ;
  assign y942 = ~1'b0 ;
  assign y943 = ~1'b0 ;
  assign y944 = n1823 ;
  assign y945 = ~1'b0 ;
  assign y946 = ~n1829 ;
  assign y947 = ~n1830 ;
  assign y948 = ~n1831 ;
  assign y949 = ~1'b0 ;
  assign y950 = ~n1833 ;
  assign y951 = ~1'b0 ;
  assign y952 = ~1'b0 ;
  assign y953 = ~n1835 ;
  assign y954 = n1839 ;
  assign y955 = ~1'b0 ;
  assign y956 = n1846 ;
  assign y957 = ~n1849 ;
  assign y958 = ~n1850 ;
  assign y959 = n1851 ;
  assign y960 = n1856 ;
  assign y961 = ~n1860 ;
  assign y962 = n1861 ;
  assign y963 = 1'b0 ;
  assign y964 = n1865 ;
  assign y965 = ~1'b0 ;
  assign y966 = n1866 ;
  assign y967 = ~n1868 ;
  assign y968 = ~n1664 ;
  assign y969 = ~n1537 ;
  assign y970 = ~1'b0 ;
  assign y971 = ~1'b0 ;
  assign y972 = ~1'b0 ;
  assign y973 = n1870 ;
  assign y974 = ~n1871 ;
  assign y975 = n1874 ;
  assign y976 = ~1'b0 ;
  assign y977 = n1877 ;
  assign y978 = n1878 ;
  assign y979 = ~1'b0 ;
  assign y980 = ~1'b0 ;
  assign y981 = n1883 ;
  assign y982 = ~n1891 ;
  assign y983 = ~n1892 ;
  assign y984 = n1894 ;
  assign y985 = ~n1897 ;
  assign y986 = ~n1898 ;
  assign y987 = n1899 ;
  assign y988 = ~n1904 ;
  assign y989 = ~1'b0 ;
  assign y990 = n1907 ;
  assign y991 = ~1'b0 ;
  assign y992 = ~1'b0 ;
  assign y993 = ~n1908 ;
  assign y994 = n1913 ;
  assign y995 = ~n1915 ;
  assign y996 = n1916 ;
  assign y997 = n1917 ;
  assign y998 = ~x62 ;
  assign y999 = ~1'b0 ;
  assign y1000 = ~1'b0 ;
  assign y1001 = n1918 ;
  assign y1002 = ~1'b0 ;
  assign y1003 = ~1'b0 ;
  assign y1004 = ~1'b0 ;
  assign y1005 = ~n1925 ;
  assign y1006 = ~n1930 ;
  assign y1007 = ~n1934 ;
  assign y1008 = n1935 ;
  assign y1009 = ~n1937 ;
  assign y1010 = ~n1945 ;
  assign y1011 = ~n1946 ;
  assign y1012 = ~1'b0 ;
  assign y1013 = n1947 ;
  assign y1014 = n1948 ;
  assign y1015 = n1951 ;
  assign y1016 = ~1'b0 ;
  assign y1017 = n1952 ;
  assign y1018 = ~n1954 ;
  assign y1019 = ~n1361 ;
  assign y1020 = ~1'b0 ;
  assign y1021 = ~n1808 ;
  assign y1022 = n1955 ;
  assign y1023 = ~1'b0 ;
  assign y1024 = ~n1957 ;
  assign y1025 = ~1'b0 ;
  assign y1026 = ~n1958 ;
  assign y1027 = ~n1961 ;
  assign y1028 = n1972 ;
  assign y1029 = ~n1975 ;
  assign y1030 = ~1'b0 ;
  assign y1031 = n1976 ;
  assign y1032 = ~n1126 ;
  assign y1033 = ~n1977 ;
  assign y1034 = ~n1979 ;
  assign y1035 = n1980 ;
  assign y1036 = ~n1981 ;
  assign y1037 = ~n1982 ;
  assign y1038 = ~1'b0 ;
  assign y1039 = ~1'b0 ;
  assign y1040 = ~n1985 ;
  assign y1041 = ~1'b0 ;
  assign y1042 = ~n1986 ;
  assign y1043 = ~n1987 ;
  assign y1044 = n1992 ;
  assign y1045 = ~1'b0 ;
  assign y1046 = ~n1993 ;
  assign y1047 = 1'b0 ;
  assign y1048 = ~1'b0 ;
  assign y1049 = ~n1996 ;
  assign y1050 = ~n1998 ;
  assign y1051 = n1999 ;
  assign y1052 = ~n315 ;
  assign y1053 = ~n2002 ;
  assign y1054 = ~n2003 ;
  assign y1055 = ~n983 ;
  assign y1056 = ~n2005 ;
  assign y1057 = n2006 ;
  assign y1058 = n2010 ;
  assign y1059 = ~1'b0 ;
  assign y1060 = n2012 ;
  assign y1061 = ~n2014 ;
  assign y1062 = ~n922 ;
  assign y1063 = 1'b0 ;
  assign y1064 = ~n2021 ;
  assign y1065 = n1651 ;
  assign y1066 = n2023 ;
  assign y1067 = ~1'b0 ;
  assign y1068 = ~n2034 ;
  assign y1069 = x60 ;
  assign y1070 = ~n2037 ;
  assign y1071 = ~n2038 ;
  assign y1072 = n2041 ;
  assign y1073 = ~n2044 ;
  assign y1074 = n2054 ;
  assign y1075 = ~n1875 ;
  assign y1076 = n1351 ;
  assign y1077 = n2055 ;
  assign y1078 = n2062 ;
  assign y1079 = ~1'b0 ;
  assign y1080 = n2070 ;
  assign y1081 = n2074 ;
  assign y1082 = ~1'b0 ;
  assign y1083 = 1'b0 ;
  assign y1084 = ~1'b0 ;
  assign y1085 = ~1'b0 ;
  assign y1086 = ~n2076 ;
  assign y1087 = n790 ;
  assign y1088 = ~n2086 ;
  assign y1089 = ~1'b0 ;
  assign y1090 = n2090 ;
  assign y1091 = n2094 ;
  assign y1092 = n2096 ;
  assign y1093 = ~1'b0 ;
  assign y1094 = n2099 ;
  assign y1095 = n2105 ;
  assign y1096 = n2109 ;
  assign y1097 = ~n2117 ;
  assign y1098 = ~n292 ;
  assign y1099 = ~1'b0 ;
  assign y1100 = ~1'b0 ;
  assign y1101 = n2122 ;
  assign y1102 = ~1'b0 ;
  assign y1103 = ~n2123 ;
  assign y1104 = ~1'b0 ;
  assign y1105 = n1548 ;
  assign y1106 = n2129 ;
  assign y1107 = n2137 ;
  assign y1108 = ~1'b0 ;
  assign y1109 = ~1'b0 ;
  assign y1110 = n2139 ;
  assign y1111 = ~n909 ;
  assign y1112 = ~n2142 ;
  assign y1113 = n2143 ;
  assign y1114 = ~1'b0 ;
  assign y1115 = 1'b0 ;
  assign y1116 = ~n2145 ;
  assign y1117 = ~1'b0 ;
  assign y1118 = ~n2146 ;
  assign y1119 = n2148 ;
  assign y1120 = n1724 ;
  assign y1121 = n825 ;
  assign y1122 = n2149 ;
  assign y1123 = ~n2153 ;
  assign y1124 = n2155 ;
  assign y1125 = n2163 ;
  assign y1126 = 1'b0 ;
  assign y1127 = ~1'b0 ;
  assign y1128 = ~1'b0 ;
  assign y1129 = ~1'b0 ;
  assign y1130 = ~n2165 ;
  assign y1131 = n2166 ;
  assign y1132 = ~n2168 ;
  assign y1133 = ~1'b0 ;
  assign y1134 = n2179 ;
  assign y1135 = ~n2181 ;
  assign y1136 = ~n811 ;
  assign y1137 = ~n2182 ;
  assign y1138 = ~n2183 ;
  assign y1139 = ~n2186 ;
  assign y1140 = ~n2190 ;
  assign y1141 = ~n2191 ;
  assign y1142 = n2193 ;
  assign y1143 = n430 ;
  assign y1144 = ~n2196 ;
  assign y1145 = n425 ;
  assign y1146 = ~1'b0 ;
  assign y1147 = ~n2200 ;
  assign y1148 = ~1'b0 ;
  assign y1149 = ~1'b0 ;
  assign y1150 = n2201 ;
  assign y1151 = ~n2206 ;
  assign y1152 = n2212 ;
  assign y1153 = ~1'b0 ;
  assign y1154 = n2213 ;
  assign y1155 = ~1'b0 ;
  assign y1156 = n2215 ;
  assign y1157 = ~1'b0 ;
  assign y1158 = n2218 ;
  assign y1159 = ~1'b0 ;
  assign y1160 = ~n2221 ;
  assign y1161 = n2222 ;
  assign y1162 = n2226 ;
  assign y1163 = ~1'b0 ;
  assign y1164 = ~n2229 ;
  assign y1165 = n2230 ;
  assign y1166 = ~1'b0 ;
  assign y1167 = ~n2233 ;
  assign y1168 = n2236 ;
  assign y1169 = ~1'b0 ;
  assign y1170 = ~n2240 ;
  assign y1171 = ~n2241 ;
  assign y1172 = ~n2242 ;
  assign y1173 = 1'b0 ;
  assign y1174 = ~n2245 ;
  assign y1175 = ~n2246 ;
  assign y1176 = n2250 ;
  assign y1177 = ~n2251 ;
  assign y1178 = n2256 ;
  assign y1179 = n2266 ;
  assign y1180 = n2268 ;
  assign y1181 = ~n2269 ;
  assign y1182 = ~n2271 ;
  assign y1183 = n2275 ;
  assign y1184 = n2276 ;
  assign y1185 = ~1'b0 ;
  assign y1186 = ~1'b0 ;
  assign y1187 = ~n2278 ;
  assign y1188 = n2279 ;
  assign y1189 = ~1'b0 ;
  assign y1190 = n2283 ;
  assign y1191 = n2285 ;
  assign y1192 = ~n2291 ;
  assign y1193 = 1'b0 ;
  assign y1194 = n2292 ;
  assign y1195 = ~n2295 ;
  assign y1196 = ~n2297 ;
  assign y1197 = n2303 ;
  assign y1198 = n2305 ;
  assign y1199 = n2308 ;
  assign y1200 = ~1'b0 ;
  assign y1201 = ~1'b0 ;
  assign y1202 = ~1'b0 ;
  assign y1203 = ~n2309 ;
  assign y1204 = ~1'b0 ;
  assign y1205 = n2312 ;
  assign y1206 = 1'b0 ;
  assign y1207 = n2313 ;
  assign y1208 = ~n2314 ;
  assign y1209 = ~n2318 ;
  assign y1210 = 1'b0 ;
  assign y1211 = n2319 ;
  assign y1212 = n2321 ;
  assign y1213 = ~n2322 ;
  assign y1214 = n2323 ;
  assign y1215 = ~1'b0 ;
  assign y1216 = n2324 ;
  assign y1217 = 1'b0 ;
  assign y1218 = ~n2329 ;
  assign y1219 = ~1'b0 ;
  assign y1220 = n2333 ;
  assign y1221 = n2337 ;
  assign y1222 = n1534 ;
  assign y1223 = ~1'b0 ;
  assign y1224 = ~n2340 ;
  assign y1225 = ~n2342 ;
  assign y1226 = n185 ;
  assign y1227 = ~n2343 ;
  assign y1228 = ~1'b0 ;
  assign y1229 = ~1'b0 ;
  assign y1230 = n2345 ;
  assign y1231 = ~1'b0 ;
  assign y1232 = n2347 ;
  assign y1233 = ~1'b0 ;
  assign y1234 = ~n2349 ;
  assign y1235 = ~1'b0 ;
  assign y1236 = ~n2351 ;
  assign y1237 = ~1'b0 ;
  assign y1238 = ~n2352 ;
  assign y1239 = ~1'b0 ;
  assign y1240 = n2358 ;
  assign y1241 = 1'b0 ;
  assign y1242 = n2364 ;
  assign y1243 = n2366 ;
  assign y1244 = ~n2367 ;
  assign y1245 = ~n2369 ;
  assign y1246 = ~n2371 ;
  assign y1247 = n2378 ;
  assign y1248 = ~n2384 ;
  assign y1249 = ~1'b0 ;
  assign y1250 = ~n2386 ;
  assign y1251 = n2395 ;
  assign y1252 = n2396 ;
  assign y1253 = ~1'b0 ;
  assign y1254 = ~1'b0 ;
  assign y1255 = n2398 ;
  assign y1256 = ~1'b0 ;
  assign y1257 = n2399 ;
  assign y1258 = ~1'b0 ;
  assign y1259 = ~1'b0 ;
  assign y1260 = ~1'b0 ;
  assign y1261 = ~1'b0 ;
  assign y1262 = ~1'b0 ;
  assign y1263 = ~1'b0 ;
  assign y1264 = n2400 ;
  assign y1265 = n2405 ;
  assign y1266 = ~1'b0 ;
  assign y1267 = ~1'b0 ;
  assign y1268 = ~1'b0 ;
  assign y1269 = ~1'b0 ;
  assign y1270 = n2408 ;
  assign y1271 = ~n485 ;
  assign y1272 = ~n2413 ;
  assign y1273 = ~n2415 ;
  assign y1274 = ~1'b0 ;
  assign y1275 = ~n2418 ;
  assign y1276 = n2422 ;
  assign y1277 = ~1'b0 ;
  assign y1278 = n1880 ;
  assign y1279 = n2426 ;
  assign y1280 = ~n2428 ;
  assign y1281 = n2433 ;
  assign y1282 = n2434 ;
  assign y1283 = ~1'b0 ;
  assign y1284 = ~n2438 ;
  assign y1285 = ~n2440 ;
  assign y1286 = ~1'b0 ;
  assign y1287 = ~1'b0 ;
  assign y1288 = n2441 ;
  assign y1289 = n2442 ;
  assign y1290 = n2443 ;
  assign y1291 = ~1'b0 ;
  assign y1292 = n1046 ;
  assign y1293 = n2445 ;
  assign y1294 = n2446 ;
  assign y1295 = n2450 ;
  assign y1296 = ~1'b0 ;
  assign y1297 = ~n2451 ;
  assign y1298 = n2452 ;
  assign y1299 = ~n2454 ;
  assign y1300 = ~n2458 ;
  assign y1301 = ~1'b0 ;
  assign y1302 = ~1'b0 ;
  assign y1303 = n2467 ;
  assign y1304 = ~1'b0 ;
  assign y1305 = n2468 ;
  assign y1306 = ~1'b0 ;
  assign y1307 = ~n2469 ;
  assign y1308 = ~n2470 ;
  assign y1309 = ~1'b0 ;
  assign y1310 = ~n2476 ;
  assign y1311 = n1443 ;
  assign y1312 = ~n2480 ;
  assign y1313 = n2482 ;
  assign y1314 = ~n2486 ;
  assign y1315 = ~n2490 ;
  assign y1316 = ~1'b0 ;
  assign y1317 = ~1'b0 ;
  assign y1318 = ~n2493 ;
  assign y1319 = n2496 ;
  assign y1320 = ~1'b0 ;
  assign y1321 = ~n2497 ;
  assign y1322 = ~1'b0 ;
  assign y1323 = ~n2499 ;
  assign y1324 = n2505 ;
  assign y1325 = n2506 ;
  assign y1326 = ~n2511 ;
  assign y1327 = ~n2516 ;
  assign y1328 = n2518 ;
  assign y1329 = n2521 ;
  assign y1330 = n2523 ;
  assign y1331 = ~n2525 ;
  assign y1332 = ~x87 ;
  assign y1333 = ~n2532 ;
  assign y1334 = n2541 ;
  assign y1335 = ~n2545 ;
  assign y1336 = ~1'b0 ;
  assign y1337 = ~n2546 ;
  assign y1338 = ~n2551 ;
  assign y1339 = n2552 ;
  assign y1340 = n2554 ;
  assign y1341 = ~1'b0 ;
  assign y1342 = ~n2555 ;
  assign y1343 = ~1'b0 ;
  assign y1344 = ~n2561 ;
  assign y1345 = ~1'b0 ;
  assign y1346 = ~n2565 ;
  assign y1347 = ~n2568 ;
  assign y1348 = ~n2569 ;
  assign y1349 = ~1'b0 ;
  assign y1350 = ~n2571 ;
  assign y1351 = n2575 ;
  assign y1352 = n2576 ;
  assign y1353 = n2579 ;
  assign y1354 = ~n2581 ;
  assign y1355 = ~n2592 ;
  assign y1356 = ~n2598 ;
  assign y1357 = n2600 ;
  assign y1358 = ~n2602 ;
  assign y1359 = n2603 ;
  assign y1360 = ~n2608 ;
  assign y1361 = x120 ;
  assign y1362 = n2610 ;
  assign y1363 = ~1'b0 ;
  assign y1364 = ~n2612 ;
  assign y1365 = n2614 ;
  assign y1366 = ~1'b0 ;
  assign y1367 = n2615 ;
  assign y1368 = n2620 ;
  assign y1369 = n2621 ;
  assign y1370 = ~1'b0 ;
  assign y1371 = ~n2624 ;
  assign y1372 = n1691 ;
  assign y1373 = ~n2626 ;
  assign y1374 = ~n2632 ;
  assign y1375 = ~n1784 ;
  assign y1376 = ~1'b0 ;
  assign y1377 = ~1'b0 ;
  assign y1378 = ~n2634 ;
  assign y1379 = ~n2637 ;
  assign y1380 = ~n2639 ;
  assign y1381 = ~1'b0 ;
  assign y1382 = n2641 ;
  assign y1383 = ~n2642 ;
  assign y1384 = ~n2643 ;
  assign y1385 = ~n2644 ;
  assign y1386 = n2647 ;
  assign y1387 = ~1'b0 ;
  assign y1388 = ~n2658 ;
  assign y1389 = n2659 ;
  assign y1390 = ~n2661 ;
  assign y1391 = ~n2666 ;
  assign y1392 = ~1'b0 ;
  assign y1393 = ~1'b0 ;
  assign y1394 = ~1'b0 ;
  assign y1395 = n2681 ;
  assign y1396 = n496 ;
  assign y1397 = ~1'b0 ;
  assign y1398 = n2689 ;
  assign y1399 = ~1'b0 ;
  assign y1400 = n2690 ;
  assign y1401 = n2691 ;
  assign y1402 = ~1'b0 ;
  assign y1403 = n2692 ;
  assign y1404 = ~n2693 ;
  assign y1405 = n2699 ;
  assign y1406 = n2702 ;
  assign y1407 = ~n2705 ;
  assign y1408 = ~1'b0 ;
  assign y1409 = ~n2716 ;
  assign y1410 = ~n2721 ;
  assign y1411 = ~1'b0 ;
  assign y1412 = ~n2733 ;
  assign y1413 = ~n2735 ;
  assign y1414 = n2738 ;
  assign y1415 = n2739 ;
  assign y1416 = ~1'b0 ;
  assign y1417 = ~1'b0 ;
  assign y1418 = ~1'b0 ;
  assign y1419 = x29 ;
  assign y1420 = ~n2745 ;
  assign y1421 = n2749 ;
  assign y1422 = ~1'b0 ;
  assign y1423 = 1'b0 ;
  assign y1424 = ~n2750 ;
  assign y1425 = n2756 ;
  assign y1426 = ~1'b0 ;
  assign y1427 = ~n2757 ;
  assign y1428 = ~n2759 ;
  assign y1429 = ~1'b0 ;
  assign y1430 = ~n2761 ;
  assign y1431 = ~1'b0 ;
  assign y1432 = ~1'b0 ;
  assign y1433 = ~1'b0 ;
  assign y1434 = ~1'b0 ;
  assign y1435 = ~1'b0 ;
  assign y1436 = n2770 ;
  assign y1437 = ~n2774 ;
  assign y1438 = ~n2775 ;
  assign y1439 = ~1'b0 ;
  assign y1440 = ~1'b0 ;
  assign y1441 = ~n2776 ;
  assign y1442 = n2777 ;
  assign y1443 = n2780 ;
  assign y1444 = n1315 ;
  assign y1445 = ~n1580 ;
  assign y1446 = x37 ;
  assign y1447 = ~n1329 ;
  assign y1448 = n2783 ;
  assign y1449 = ~1'b0 ;
  assign y1450 = n2786 ;
  assign y1451 = ~n2789 ;
  assign y1452 = n2792 ;
  assign y1453 = n2694 ;
  assign y1454 = ~1'b0 ;
  assign y1455 = n1782 ;
  assign y1456 = n2803 ;
  assign y1457 = n2804 ;
  assign y1458 = ~1'b0 ;
  assign y1459 = ~1'b0 ;
  assign y1460 = ~n2818 ;
  assign y1461 = ~n2819 ;
  assign y1462 = ~1'b0 ;
  assign y1463 = ~n2822 ;
  assign y1464 = ~1'b0 ;
  assign y1465 = n2824 ;
  assign y1466 = ~n2826 ;
  assign y1467 = ~1'b0 ;
  assign y1468 = ~n2827 ;
  assign y1469 = ~1'b0 ;
  assign y1470 = ~n2831 ;
  assign y1471 = ~n970 ;
  assign y1472 = ~n2833 ;
  assign y1473 = n2835 ;
  assign y1474 = ~n2838 ;
  assign y1475 = ~n2839 ;
  assign y1476 = ~n2842 ;
  assign y1477 = ~1'b0 ;
  assign y1478 = n2843 ;
  assign y1479 = n2849 ;
  assign y1480 = n2850 ;
  assign y1481 = ~n2855 ;
  assign y1482 = ~n2857 ;
  assign y1483 = n2858 ;
  assign y1484 = n2859 ;
  assign y1485 = n2866 ;
  assign y1486 = ~1'b0 ;
  assign y1487 = n704 ;
  assign y1488 = ~1'b0 ;
  assign y1489 = ~1'b0 ;
  assign y1490 = ~1'b0 ;
  assign y1491 = ~n2867 ;
  assign y1492 = ~n2872 ;
  assign y1493 = n2875 ;
  assign y1494 = ~1'b0 ;
  assign y1495 = n2815 ;
  assign y1496 = ~1'b0 ;
  assign y1497 = ~n2876 ;
  assign y1498 = n2879 ;
  assign y1499 = n2880 ;
  assign y1500 = n2881 ;
  assign y1501 = n2882 ;
  assign y1502 = n2884 ;
  assign y1503 = ~1'b0 ;
  assign y1504 = n2895 ;
  assign y1505 = ~n2896 ;
  assign y1506 = ~1'b0 ;
  assign y1507 = ~1'b0 ;
  assign y1508 = ~1'b0 ;
  assign y1509 = ~n2898 ;
  assign y1510 = ~n2899 ;
  assign y1511 = n2900 ;
  assign y1512 = ~1'b0 ;
  assign y1513 = ~n2903 ;
  assign y1514 = ~1'b0 ;
  assign y1515 = ~1'b0 ;
  assign y1516 = ~1'b0 ;
  assign y1517 = ~1'b0 ;
  assign y1518 = n2906 ;
  assign y1519 = n2907 ;
  assign y1520 = n2908 ;
  assign y1521 = n828 ;
  assign y1522 = ~n2913 ;
  assign y1523 = ~1'b0 ;
  assign y1524 = ~1'b0 ;
  assign y1525 = ~n2587 ;
  assign y1526 = n595 ;
  assign y1527 = n2915 ;
  assign y1528 = ~n2917 ;
  assign y1529 = ~1'b0 ;
  assign y1530 = n2919 ;
  assign y1531 = n2921 ;
  assign y1532 = n2924 ;
  assign y1533 = ~n2928 ;
  assign y1534 = ~1'b0 ;
  assign y1535 = n2931 ;
  assign y1536 = ~n2933 ;
  assign y1537 = ~n2936 ;
  assign y1538 = ~n2937 ;
  assign y1539 = ~1'b0 ;
  assign y1540 = n2938 ;
  assign y1541 = ~n2940 ;
  assign y1542 = ~1'b0 ;
  assign y1543 = ~n2941 ;
  assign y1544 = n2942 ;
  assign y1545 = ~n2943 ;
  assign y1546 = n2945 ;
  assign y1547 = ~n1487 ;
  assign y1548 = ~n2948 ;
  assign y1549 = n2949 ;
  assign y1550 = ~1'b0 ;
  assign y1551 = n2954 ;
  assign y1552 = ~n2955 ;
  assign y1553 = ~1'b0 ;
  assign y1554 = n2958 ;
  assign y1555 = n2959 ;
  assign y1556 = n2960 ;
  assign y1557 = n2966 ;
  assign y1558 = ~n2969 ;
  assign y1559 = n2971 ;
  assign y1560 = n2977 ;
  assign y1561 = n624 ;
  assign y1562 = ~n2983 ;
  assign y1563 = ~1'b0 ;
  assign y1564 = ~n2985 ;
  assign y1565 = ~1'b0 ;
  assign y1566 = ~1'b0 ;
  assign y1567 = ~n1037 ;
  assign y1568 = ~n2988 ;
  assign y1569 = ~n2989 ;
  assign y1570 = ~1'b0 ;
  assign y1571 = ~1'b0 ;
  assign y1572 = n2993 ;
  assign y1573 = n2995 ;
  assign y1574 = x85 ;
  assign y1575 = ~n2997 ;
  assign y1576 = n2998 ;
  assign y1577 = ~n3007 ;
  assign y1578 = n3015 ;
  assign y1579 = n3025 ;
  assign y1580 = ~1'b0 ;
  assign y1581 = ~n3027 ;
  assign y1582 = ~n3028 ;
  assign y1583 = ~1'b0 ;
  assign y1584 = ~n3031 ;
  assign y1585 = ~1'b0 ;
  assign y1586 = n373 ;
  assign y1587 = ~n3035 ;
  assign y1588 = ~n3037 ;
  assign y1589 = n3038 ;
  assign y1590 = ~1'b0 ;
  assign y1591 = n1419 ;
  assign y1592 = n3043 ;
  assign y1593 = ~1'b0 ;
  assign y1594 = ~1'b0 ;
  assign y1595 = n3046 ;
  assign y1596 = ~1'b0 ;
  assign y1597 = n3050 ;
  assign y1598 = ~n3053 ;
  assign y1599 = ~n3057 ;
  assign y1600 = n3060 ;
  assign y1601 = ~1'b0 ;
  assign y1602 = ~n3063 ;
  assign y1603 = n3066 ;
  assign y1604 = ~n3067 ;
  assign y1605 = ~1'b0 ;
  assign y1606 = ~n3068 ;
  assign y1607 = n3069 ;
  assign y1608 = ~n3071 ;
  assign y1609 = n3072 ;
  assign y1610 = ~1'b0 ;
  assign y1611 = ~n3075 ;
  assign y1612 = n3076 ;
  assign y1613 = ~1'b0 ;
  assign y1614 = ~1'b0 ;
  assign y1615 = ~1'b0 ;
  assign y1616 = n3077 ;
  assign y1617 = ~n3078 ;
  assign y1618 = n266 ;
  assign y1619 = n3079 ;
  assign y1620 = ~1'b0 ;
  assign y1621 = ~1'b0 ;
  assign y1622 = ~1'b0 ;
  assign y1623 = ~n3083 ;
  assign y1624 = n3087 ;
  assign y1625 = ~1'b0 ;
  assign y1626 = ~n3089 ;
  assign y1627 = n3094 ;
  assign y1628 = ~1'b0 ;
  assign y1629 = n3096 ;
  assign y1630 = ~1'b0 ;
  assign y1631 = ~n3097 ;
  assign y1632 = 1'b0 ;
  assign y1633 = n3098 ;
  assign y1634 = n3103 ;
  assign y1635 = ~n3104 ;
  assign y1636 = ~1'b0 ;
  assign y1637 = ~1'b0 ;
  assign y1638 = n3106 ;
  assign y1639 = ~1'b0 ;
  assign y1640 = n3108 ;
  assign y1641 = n3110 ;
  assign y1642 = ~1'b0 ;
  assign y1643 = ~1'b0 ;
  assign y1644 = ~1'b0 ;
  assign y1645 = n3112 ;
  assign y1646 = ~1'b0 ;
  assign y1647 = ~n3116 ;
  assign y1648 = ~n3118 ;
  assign y1649 = n237 ;
  assign y1650 = ~1'b0 ;
  assign y1651 = ~1'b0 ;
  assign y1652 = ~1'b0 ;
  assign y1653 = ~n3120 ;
  assign y1654 = ~1'b0 ;
  assign y1655 = ~1'b0 ;
  assign y1656 = ~n3121 ;
  assign y1657 = n3123 ;
  assign y1658 = n1251 ;
  assign y1659 = ~n3124 ;
  assign y1660 = ~n3126 ;
  assign y1661 = ~n3128 ;
  assign y1662 = ~n3135 ;
  assign y1663 = 1'b0 ;
  assign y1664 = ~1'b0 ;
  assign y1665 = n3136 ;
  assign y1666 = n3145 ;
  assign y1667 = ~1'b0 ;
  assign y1668 = n3147 ;
  assign y1669 = n3150 ;
  assign y1670 = ~1'b0 ;
  assign y1671 = 1'b0 ;
  assign y1672 = ~n3153 ;
  assign y1673 = n3156 ;
  assign y1674 = ~n3158 ;
  assign y1675 = ~1'b0 ;
  assign y1676 = ~n3163 ;
  assign y1677 = ~n3167 ;
  assign y1678 = ~n3170 ;
  assign y1679 = ~n3174 ;
  assign y1680 = ~n3176 ;
  assign y1681 = n3180 ;
  assign y1682 = ~n1630 ;
  assign y1683 = ~n3188 ;
  assign y1684 = n851 ;
  assign y1685 = ~n3191 ;
  assign y1686 = n3192 ;
  assign y1687 = ~n3194 ;
  assign y1688 = ~n3196 ;
  assign y1689 = ~1'b0 ;
  assign y1690 = ~1'b0 ;
  assign y1691 = n3198 ;
  assign y1692 = n3201 ;
  assign y1693 = ~n3203 ;
  assign y1694 = n3210 ;
  assign y1695 = ~n3213 ;
  assign y1696 = ~1'b0 ;
  assign y1697 = n3221 ;
  assign y1698 = ~1'b0 ;
  assign y1699 = ~n3223 ;
  assign y1700 = ~1'b0 ;
  assign y1701 = ~n3226 ;
  assign y1702 = ~1'b0 ;
  assign y1703 = ~n3228 ;
  assign y1704 = ~1'b0 ;
  assign y1705 = 1'b0 ;
  assign y1706 = ~n3229 ;
  assign y1707 = n3230 ;
  assign y1708 = ~n1758 ;
  assign y1709 = ~n221 ;
  assign y1710 = ~1'b0 ;
  assign y1711 = 1'b0 ;
  assign y1712 = ~n3231 ;
  assign y1713 = n3232 ;
  assign y1714 = ~1'b0 ;
  assign y1715 = n3236 ;
  assign y1716 = n1786 ;
  assign y1717 = n3237 ;
  assign y1718 = ~1'b0 ;
  assign y1719 = n932 ;
  assign y1720 = 1'b0 ;
  assign y1721 = n3149 ;
  assign y1722 = n189 ;
  assign y1723 = n3242 ;
  assign y1724 = n3244 ;
  assign y1725 = n2942 ;
  assign y1726 = ~n3247 ;
  assign y1727 = n3255 ;
  assign y1728 = ~1'b0 ;
  assign y1729 = ~1'b0 ;
  assign y1730 = n3264 ;
  assign y1731 = n3269 ;
  assign y1732 = ~n3270 ;
  assign y1733 = ~1'b0 ;
  assign y1734 = ~1'b0 ;
  assign y1735 = n753 ;
  assign y1736 = ~1'b0 ;
  assign y1737 = ~1'b0 ;
  assign y1738 = ~n3276 ;
  assign y1739 = n3278 ;
  assign y1740 = ~1'b0 ;
  assign y1741 = n3279 ;
  assign y1742 = ~n3281 ;
  assign y1743 = ~n3285 ;
  assign y1744 = ~1'b0 ;
  assign y1745 = ~1'b0 ;
  assign y1746 = ~1'b0 ;
  assign y1747 = ~n3290 ;
  assign y1748 = ~n3292 ;
  assign y1749 = ~n3293 ;
  assign y1750 = ~1'b0 ;
  assign y1751 = ~1'b0 ;
  assign y1752 = ~n3295 ;
  assign y1753 = ~1'b0 ;
  assign y1754 = ~n3298 ;
  assign y1755 = ~n3300 ;
  assign y1756 = ~n3302 ;
  assign y1757 = ~n3304 ;
  assign y1758 = n3307 ;
  assign y1759 = n3312 ;
  assign y1760 = ~n3318 ;
  assign y1761 = ~1'b0 ;
  assign y1762 = n3327 ;
  assign y1763 = n3328 ;
  assign y1764 = ~n3330 ;
  assign y1765 = ~1'b0 ;
  assign y1766 = ~1'b0 ;
  assign y1767 = ~n3338 ;
  assign y1768 = ~n2602 ;
  assign y1769 = ~1'b0 ;
  assign y1770 = n3340 ;
  assign y1771 = ~1'b0 ;
  assign y1772 = ~n2107 ;
  assign y1773 = ~1'b0 ;
  assign y1774 = n3344 ;
  assign y1775 = ~n3348 ;
  assign y1776 = ~n3356 ;
  assign y1777 = n3359 ;
  assign y1778 = ~n3363 ;
  assign y1779 = ~1'b0 ;
  assign y1780 = ~1'b0 ;
  assign y1781 = ~n3364 ;
  assign y1782 = ~1'b0 ;
  assign y1783 = ~1'b0 ;
  assign y1784 = ~1'b0 ;
  assign y1785 = ~n3373 ;
  assign y1786 = n3376 ;
  assign y1787 = n645 ;
  assign y1788 = n3377 ;
  assign y1789 = n3378 ;
  assign y1790 = n3379 ;
  assign y1791 = n3381 ;
  assign y1792 = ~n3382 ;
  assign y1793 = ~n1983 ;
  assign y1794 = n3388 ;
  assign y1795 = n3392 ;
  assign y1796 = ~1'b0 ;
  assign y1797 = ~1'b0 ;
  assign y1798 = ~1'b0 ;
  assign y1799 = ~1'b0 ;
  assign y1800 = n570 ;
  assign y1801 = ~1'b0 ;
  assign y1802 = ~n3396 ;
  assign y1803 = ~n3397 ;
  assign y1804 = n3400 ;
  assign y1805 = n3406 ;
  assign y1806 = ~n3407 ;
  assign y1807 = ~1'b0 ;
  assign y1808 = ~1'b0 ;
  assign y1809 = n3415 ;
  assign y1810 = n3428 ;
  assign y1811 = ~1'b0 ;
  assign y1812 = n3429 ;
  assign y1813 = ~n3430 ;
  assign y1814 = ~1'b0 ;
  assign y1815 = n3431 ;
  assign y1816 = ~n3432 ;
  assign y1817 = n3434 ;
  assign y1818 = n3436 ;
  assign y1819 = ~n3441 ;
  assign y1820 = ~n3443 ;
  assign y1821 = n3447 ;
  assign y1822 = ~1'b0 ;
  assign y1823 = n2923 ;
  assign y1824 = n3450 ;
  assign y1825 = ~1'b0 ;
  assign y1826 = ~1'b0 ;
  assign y1827 = n3452 ;
  assign y1828 = n3456 ;
  assign y1829 = n3461 ;
  assign y1830 = n3462 ;
  assign y1831 = ~n3468 ;
  assign y1832 = 1'b0 ;
  assign y1833 = n3473 ;
  assign y1834 = ~1'b0 ;
  assign y1835 = ~1'b0 ;
  assign y1836 = 1'b0 ;
  assign y1837 = ~1'b0 ;
  assign y1838 = ~n3475 ;
  assign y1839 = ~n3477 ;
  assign y1840 = ~n3479 ;
  assign y1841 = ~n3487 ;
  assign y1842 = n3488 ;
  assign y1843 = ~1'b0 ;
  assign y1844 = ~1'b0 ;
  assign y1845 = ~n1623 ;
  assign y1846 = ~1'b0 ;
  assign y1847 = n3489 ;
  assign y1848 = ~n3491 ;
  assign y1849 = n3494 ;
  assign y1850 = n3499 ;
  assign y1851 = ~n3502 ;
  assign y1852 = ~n3504 ;
  assign y1853 = ~1'b0 ;
  assign y1854 = n3505 ;
  assign y1855 = ~n3510 ;
  assign y1856 = n3518 ;
  assign y1857 = ~n3519 ;
  assign y1858 = n3523 ;
  assign y1859 = ~n3525 ;
  assign y1860 = ~n3526 ;
  assign y1861 = n3527 ;
  assign y1862 = ~x55 ;
  assign y1863 = n3532 ;
  assign y1864 = n1875 ;
  assign y1865 = ~1'b0 ;
  assign y1866 = ~1'b0 ;
  assign y1867 = n3534 ;
  assign y1868 = ~n3541 ;
  assign y1869 = ~1'b0 ;
  assign y1870 = n3547 ;
  assign y1871 = ~n3548 ;
  assign y1872 = ~n3552 ;
  assign y1873 = n3553 ;
  assign y1874 = ~n3557 ;
  assign y1875 = ~1'b0 ;
  assign y1876 = ~1'b0 ;
  assign y1877 = n3558 ;
  assign y1878 = ~n2602 ;
  assign y1879 = ~n3561 ;
  assign y1880 = ~n3507 ;
  assign y1881 = n3565 ;
  assign y1882 = ~n3569 ;
  assign y1883 = n3575 ;
  assign y1884 = n3577 ;
  assign y1885 = ~n3579 ;
  assign y1886 = ~1'b0 ;
  assign y1887 = n3580 ;
  assign y1888 = ~n3584 ;
  assign y1889 = ~n3585 ;
  assign y1890 = ~1'b0 ;
  assign y1891 = ~n3589 ;
  assign y1892 = ~1'b0 ;
  assign y1893 = ~x57 ;
  assign y1894 = ~1'b0 ;
  assign y1895 = ~1'b0 ;
  assign y1896 = ~n3595 ;
  assign y1897 = ~1'b0 ;
  assign y1898 = ~1'b0 ;
  assign y1899 = ~1'b0 ;
  assign y1900 = ~n3597 ;
  assign y1901 = ~1'b0 ;
  assign y1902 = n3599 ;
  assign y1903 = 1'b0 ;
  assign y1904 = ~n3602 ;
  assign y1905 = ~n3604 ;
  assign y1906 = n3605 ;
  assign y1907 = ~1'b0 ;
  assign y1908 = n3608 ;
  assign y1909 = ~1'b0 ;
  assign y1910 = n3610 ;
  assign y1911 = n3615 ;
  assign y1912 = ~1'b0 ;
  assign y1913 = n3619 ;
  assign y1914 = ~n3628 ;
  assign y1915 = ~n3262 ;
  assign y1916 = ~1'b0 ;
  assign y1917 = n3629 ;
  assign y1918 = ~n3630 ;
  assign y1919 = ~n3633 ;
  assign y1920 = n3634 ;
  assign y1921 = ~1'b0 ;
  assign y1922 = ~n3637 ;
  assign y1923 = ~n3650 ;
  assign y1924 = ~1'b0 ;
  assign y1925 = ~1'b0 ;
  assign y1926 = ~1'b0 ;
  assign y1927 = n296 ;
  assign y1928 = ~1'b0 ;
  assign y1929 = n3651 ;
  assign y1930 = ~1'b0 ;
  assign y1931 = ~1'b0 ;
  assign y1932 = ~1'b0 ;
  assign y1933 = ~n3655 ;
  assign y1934 = ~1'b0 ;
  assign y1935 = ~1'b0 ;
  assign y1936 = ~1'b0 ;
  assign y1937 = n3658 ;
  assign y1938 = ~1'b0 ;
  assign y1939 = ~1'b0 ;
  assign y1940 = ~n3661 ;
  assign y1941 = n3665 ;
  assign y1942 = ~n3669 ;
  assign y1943 = ~1'b0 ;
  assign y1944 = ~1'b0 ;
  assign y1945 = ~1'b0 ;
  assign y1946 = ~1'b0 ;
  assign y1947 = ~n3671 ;
  assign y1948 = ~n3672 ;
  assign y1949 = ~1'b0 ;
  assign y1950 = n3673 ;
  assign y1951 = ~n3674 ;
  assign y1952 = ~n3675 ;
  assign y1953 = ~n3677 ;
  assign y1954 = ~1'b0 ;
  assign y1955 = n183 ;
  assign y1956 = ~n3678 ;
  assign y1957 = ~1'b0 ;
  assign y1958 = ~1'b0 ;
  assign y1959 = ~1'b0 ;
  assign y1960 = ~n3680 ;
  assign y1961 = ~1'b0 ;
  assign y1962 = ~1'b0 ;
  assign y1963 = n707 ;
  assign y1964 = n3695 ;
  assign y1965 = n3696 ;
  assign y1966 = ~n3699 ;
  assign y1967 = n3700 ;
  assign y1968 = n3704 ;
  assign y1969 = ~1'b0 ;
  assign y1970 = ~1'b0 ;
  assign y1971 = ~n3707 ;
  assign y1972 = ~n3711 ;
  assign y1973 = ~1'b0 ;
  assign y1974 = ~1'b0 ;
  assign y1975 = ~1'b0 ;
  assign y1976 = n3712 ;
  assign y1977 = ~n3715 ;
  assign y1978 = ~1'b0 ;
  assign y1979 = 1'b0 ;
  assign y1980 = ~1'b0 ;
  assign y1981 = n3718 ;
  assign y1982 = n3721 ;
  assign y1983 = n3723 ;
  assign y1984 = ~n3725 ;
  assign y1985 = n3726 ;
  assign y1986 = n277 ;
  assign y1987 = ~1'b0 ;
  assign y1988 = ~1'b0 ;
  assign y1989 = ~1'b0 ;
  assign y1990 = ~1'b0 ;
  assign y1991 = n3728 ;
  assign y1992 = ~1'b0 ;
  assign y1993 = ~1'b0 ;
  assign y1994 = ~n3729 ;
  assign y1995 = n3730 ;
  assign y1996 = ~1'b0 ;
  assign y1997 = n3732 ;
  assign y1998 = n3734 ;
  assign y1999 = ~n3739 ;
  assign y2000 = ~n978 ;
  assign y2001 = n3740 ;
  assign y2002 = ~1'b0 ;
  assign y2003 = 1'b0 ;
  assign y2004 = ~n3744 ;
  assign y2005 = n3748 ;
  assign y2006 = ~n3749 ;
  assign y2007 = ~n3750 ;
  assign y2008 = n3753 ;
  assign y2009 = ~1'b0 ;
  assign y2010 = ~1'b0 ;
  assign y2011 = ~n3755 ;
  assign y2012 = n3758 ;
  assign y2013 = ~n305 ;
  assign y2014 = n3759 ;
  assign y2015 = ~n3762 ;
  assign y2016 = ~1'b0 ;
  assign y2017 = ~1'b0 ;
  assign y2018 = n3763 ;
  assign y2019 = ~n3769 ;
  assign y2020 = ~n3772 ;
  assign y2021 = ~n3773 ;
  assign y2022 = ~n3774 ;
  assign y2023 = n3776 ;
  assign y2024 = ~1'b0 ;
  assign y2025 = n3778 ;
  assign y2026 = ~n985 ;
  assign y2027 = ~n3780 ;
  assign y2028 = ~1'b0 ;
  assign y2029 = n3788 ;
  assign y2030 = 1'b0 ;
  assign y2031 = ~1'b0 ;
  assign y2032 = n3792 ;
  assign y2033 = ~1'b0 ;
  assign y2034 = ~1'b0 ;
  assign y2035 = n3793 ;
  assign y2036 = n3794 ;
  assign y2037 = n3795 ;
  assign y2038 = n3797 ;
  assign y2039 = ~1'b0 ;
  assign y2040 = n3800 ;
  assign y2041 = n3802 ;
  assign y2042 = ~1'b0 ;
  assign y2043 = n171 ;
  assign y2044 = n3803 ;
  assign y2045 = ~n806 ;
  assign y2046 = ~n2566 ;
  assign y2047 = ~n3770 ;
  assign y2048 = ~1'b0 ;
  assign y2049 = ~1'b0 ;
  assign y2050 = n3804 ;
  assign y2051 = n3813 ;
  assign y2052 = n3818 ;
  assign y2053 = n3821 ;
  assign y2054 = n3823 ;
  assign y2055 = ~1'b0 ;
  assign y2056 = n3828 ;
  assign y2057 = n3829 ;
  assign y2058 = ~1'b0 ;
  assign y2059 = ~n3831 ;
  assign y2060 = ~1'b0 ;
  assign y2061 = ~1'b0 ;
  assign y2062 = ~n3834 ;
  assign y2063 = n3836 ;
  assign y2064 = ~n3840 ;
  assign y2065 = ~n3844 ;
  assign y2066 = n3847 ;
  assign y2067 = ~1'b0 ;
  assign y2068 = n3853 ;
  assign y2069 = ~1'b0 ;
  assign y2070 = n3860 ;
  assign y2071 = ~1'b0 ;
  assign y2072 = ~n3861 ;
  assign y2073 = n3866 ;
  assign y2074 = n3868 ;
  assign y2075 = ~1'b0 ;
  assign y2076 = n3873 ;
  assign y2077 = ~n3875 ;
  assign y2078 = n1035 ;
  assign y2079 = ~1'b0 ;
  assign y2080 = n3877 ;
  assign y2081 = ~1'b0 ;
  assign y2082 = ~1'b0 ;
  assign y2083 = n3878 ;
  assign y2084 = ~n3882 ;
  assign y2085 = n3888 ;
  assign y2086 = ~n3891 ;
  assign y2087 = ~1'b0 ;
  assign y2088 = n3893 ;
  assign y2089 = ~1'b0 ;
  assign y2090 = ~1'b0 ;
  assign y2091 = ~1'b0 ;
  assign y2092 = n3897 ;
  assign y2093 = ~1'b0 ;
  assign y2094 = ~1'b0 ;
  assign y2095 = ~n3900 ;
  assign y2096 = n3902 ;
  assign y2097 = ~1'b0 ;
  assign y2098 = ~n3905 ;
  assign y2099 = ~1'b0 ;
  assign y2100 = ~n2427 ;
  assign y2101 = ~n1807 ;
  assign y2102 = ~n3906 ;
  assign y2103 = ~n3907 ;
  assign y2104 = ~n3908 ;
  assign y2105 = ~n3909 ;
  assign y2106 = n2313 ;
  assign y2107 = ~n3910 ;
  assign y2108 = ~1'b0 ;
  assign y2109 = ~1'b0 ;
  assign y2110 = ~n3915 ;
  assign y2111 = ~n3916 ;
  assign y2112 = ~n3917 ;
  assign y2113 = ~1'b0 ;
  assign y2114 = ~x2 ;
  assign y2115 = n3921 ;
  assign y2116 = n3922 ;
  assign y2117 = 1'b0 ;
  assign y2118 = 1'b0 ;
  assign y2119 = n3925 ;
  assign y2120 = ~n3927 ;
  assign y2121 = ~1'b0 ;
  assign y2122 = n3931 ;
  assign y2123 = n3934 ;
  assign y2124 = ~1'b0 ;
  assign y2125 = ~1'b0 ;
  assign y2126 = n3937 ;
  assign y2127 = ~1'b0 ;
  assign y2128 = ~n3944 ;
  assign y2129 = ~1'b0 ;
  assign y2130 = ~n3946 ;
  assign y2131 = ~1'b0 ;
  assign y2132 = n152 ;
  assign y2133 = n3948 ;
  assign y2134 = ~n3949 ;
  assign y2135 = ~1'b0 ;
  assign y2136 = ~1'b0 ;
  assign y2137 = ~n3953 ;
  assign y2138 = ~1'b0 ;
  assign y2139 = ~1'b0 ;
  assign y2140 = n3962 ;
  assign y2141 = n3966 ;
  assign y2142 = n3970 ;
  assign y2143 = n3973 ;
  assign y2144 = n3974 ;
  assign y2145 = n3975 ;
  assign y2146 = ~n3976 ;
  assign y2147 = ~n2087 ;
  assign y2148 = 1'b0 ;
  assign y2149 = ~n3977 ;
  assign y2150 = ~n3422 ;
  assign y2151 = ~n3978 ;
  assign y2152 = ~1'b0 ;
  assign y2153 = ~1'b0 ;
  assign y2154 = ~1'b0 ;
  assign y2155 = ~1'b0 ;
  assign y2156 = ~1'b0 ;
  assign y2157 = ~n806 ;
  assign y2158 = n3985 ;
  assign y2159 = ~1'b0 ;
  assign y2160 = ~1'b0 ;
  assign y2161 = ~1'b0 ;
  assign y2162 = ~1'b0 ;
  assign y2163 = ~n3987 ;
  assign y2164 = ~n3994 ;
  assign y2165 = ~1'b0 ;
  assign y2166 = n4001 ;
  assign y2167 = n4005 ;
  assign y2168 = ~n4011 ;
  assign y2169 = n4016 ;
  assign y2170 = n4027 ;
  assign y2171 = n4028 ;
  assign y2172 = ~1'b0 ;
  assign y2173 = ~1'b0 ;
  assign y2174 = ~n4029 ;
  assign y2175 = n4032 ;
  assign y2176 = n4034 ;
  assign y2177 = ~1'b0 ;
  assign y2178 = ~n4035 ;
  assign y2179 = ~n4038 ;
  assign y2180 = n4040 ;
  assign y2181 = ~n4042 ;
  assign y2182 = n4043 ;
  assign y2183 = ~1'b0 ;
  assign y2184 = ~n4047 ;
  assign y2185 = ~1'b0 ;
  assign y2186 = 1'b0 ;
  assign y2187 = ~n4048 ;
  assign y2188 = ~n4050 ;
  assign y2189 = n4054 ;
  assign y2190 = ~n4061 ;
  assign y2191 = n4064 ;
  assign y2192 = ~1'b0 ;
  assign y2193 = ~1'b0 ;
  assign y2194 = ~1'b0 ;
  assign y2195 = 1'b0 ;
  assign y2196 = ~n4069 ;
  assign y2197 = ~1'b0 ;
  assign y2198 = ~n4070 ;
  assign y2199 = ~1'b0 ;
  assign y2200 = ~1'b0 ;
  assign y2201 = ~1'b0 ;
  assign y2202 = ~n4071 ;
  assign y2203 = ~1'b0 ;
  assign y2204 = 1'b0 ;
  assign y2205 = n4072 ;
  assign y2206 = ~1'b0 ;
  assign y2207 = ~n4074 ;
  assign y2208 = ~n4078 ;
  assign y2209 = ~n4079 ;
  assign y2210 = ~n4081 ;
  assign y2211 = n4083 ;
  assign y2212 = n3878 ;
  assign y2213 = ~n4084 ;
  assign y2214 = n4087 ;
  assign y2215 = ~1'b0 ;
  assign y2216 = n4100 ;
  assign y2217 = ~1'b0 ;
  assign y2218 = ~n4107 ;
  assign y2219 = n4109 ;
  assign y2220 = n4112 ;
  assign y2221 = ~n4114 ;
  assign y2222 = 1'b0 ;
  assign y2223 = ~1'b0 ;
  assign y2224 = ~n4115 ;
  assign y2225 = n4118 ;
  assign y2226 = ~1'b0 ;
  assign y2227 = ~1'b0 ;
  assign y2228 = ~1'b0 ;
  assign y2229 = ~n4120 ;
  assign y2230 = ~1'b0 ;
  assign y2231 = ~1'b0 ;
  assign y2232 = ~n4122 ;
  assign y2233 = n4129 ;
  assign y2234 = n4133 ;
  assign y2235 = n4135 ;
  assign y2236 = ~x71 ;
  assign y2237 = n4139 ;
  assign y2238 = ~1'b0 ;
  assign y2239 = ~n4141 ;
  assign y2240 = ~n4144 ;
  assign y2241 = ~1'b0 ;
  assign y2242 = ~1'b0 ;
  assign y2243 = n4148 ;
  assign y2244 = ~n4150 ;
  assign y2245 = ~n4151 ;
  assign y2246 = ~n4155 ;
  assign y2247 = ~n4158 ;
  assign y2248 = ~1'b0 ;
  assign y2249 = ~n4167 ;
  assign y2250 = n4170 ;
  assign y2251 = ~1'b0 ;
  assign y2252 = ~1'b0 ;
  assign y2253 = ~1'b0 ;
  assign y2254 = n4173 ;
  assign y2255 = n1632 ;
  assign y2256 = ~1'b0 ;
  assign y2257 = ~1'b0 ;
  assign y2258 = ~n4181 ;
  assign y2259 = ~n4183 ;
  assign y2260 = n4186 ;
  assign y2261 = ~1'b0 ;
  assign y2262 = ~1'b0 ;
  assign y2263 = ~1'b0 ;
  assign y2264 = n4188 ;
  assign y2265 = ~n4189 ;
  assign y2266 = n4191 ;
  assign y2267 = ~n3074 ;
  assign y2268 = n4193 ;
  assign y2269 = ~1'b0 ;
  assign y2270 = ~1'b0 ;
  assign y2271 = ~1'b0 ;
  assign y2272 = ~n4200 ;
  assign y2273 = ~n432 ;
  assign y2274 = ~n4202 ;
  assign y2275 = ~n4210 ;
  assign y2276 = ~n4212 ;
  assign y2277 = ~n4213 ;
  assign y2278 = ~1'b0 ;
  assign y2279 = ~1'b0 ;
  assign y2280 = n4214 ;
  assign y2281 = n4215 ;
  assign y2282 = n4216 ;
  assign y2283 = 1'b0 ;
  assign y2284 = 1'b0 ;
  assign y2285 = ~n4217 ;
  assign y2286 = ~n4218 ;
  assign y2287 = n4219 ;
  assign y2288 = ~n4222 ;
  assign y2289 = n4227 ;
  assign y2290 = ~n895 ;
  assign y2291 = ~n4242 ;
  assign y2292 = n4244 ;
  assign y2293 = n4245 ;
  assign y2294 = ~n4247 ;
  assign y2295 = ~n4248 ;
  assign y2296 = ~1'b0 ;
  assign y2297 = ~n4249 ;
  assign y2298 = n4251 ;
  assign y2299 = ~1'b0 ;
  assign y2300 = ~n4252 ;
  assign y2301 = n4253 ;
  assign y2302 = ~1'b0 ;
  assign y2303 = ~1'b0 ;
  assign y2304 = n1491 ;
  assign y2305 = n4256 ;
  assign y2306 = ~n4259 ;
  assign y2307 = ~n4261 ;
  assign y2308 = n4265 ;
  assign y2309 = ~1'b0 ;
  assign y2310 = n4268 ;
  assign y2311 = ~n335 ;
  assign y2312 = ~1'b0 ;
  assign y2313 = n4269 ;
  assign y2314 = n2854 ;
  assign y2315 = n3870 ;
  assign y2316 = ~1'b0 ;
  assign y2317 = n4272 ;
  assign y2318 = 1'b0 ;
  assign y2319 = ~n4279 ;
  assign y2320 = ~1'b0 ;
  assign y2321 = ~1'b0 ;
  assign y2322 = ~n4282 ;
  assign y2323 = n4284 ;
  assign y2324 = ~n4288 ;
  assign y2325 = ~n4293 ;
  assign y2326 = ~1'b0 ;
  assign y2327 = 1'b0 ;
  assign y2328 = ~n4294 ;
  assign y2329 = ~n4300 ;
  assign y2330 = ~n4301 ;
  assign y2331 = ~1'b0 ;
  assign y2332 = n4304 ;
  assign y2333 = ~n3890 ;
  assign y2334 = ~n4306 ;
  assign y2335 = ~1'b0 ;
  assign y2336 = ~n4310 ;
  assign y2337 = n4312 ;
  assign y2338 = ~1'b0 ;
  assign y2339 = ~n4313 ;
  assign y2340 = 1'b0 ;
  assign y2341 = ~x11 ;
  assign y2342 = n4315 ;
  assign y2343 = ~n4318 ;
  assign y2344 = ~n4321 ;
  assign y2345 = ~1'b0 ;
  assign y2346 = ~1'b0 ;
  assign y2347 = n535 ;
  assign y2348 = n4322 ;
  assign y2349 = ~n4323 ;
  assign y2350 = n4328 ;
  assign y2351 = 1'b0 ;
  assign y2352 = n963 ;
  assign y2353 = n2383 ;
  assign y2354 = ~1'b0 ;
  assign y2355 = n4330 ;
  assign y2356 = n4334 ;
  assign y2357 = ~n3158 ;
  assign y2358 = n4336 ;
  assign y2359 = ~n4337 ;
  assign y2360 = ~1'b0 ;
  assign y2361 = n4338 ;
  assign y2362 = ~1'b0 ;
  assign y2363 = n4339 ;
  assign y2364 = n4340 ;
  assign y2365 = n4344 ;
  assign y2366 = n4345 ;
  assign y2367 = n4349 ;
  assign y2368 = ~1'b0 ;
  assign y2369 = ~1'b0 ;
  assign y2370 = n307 ;
  assign y2371 = ~n4350 ;
  assign y2372 = n4353 ;
  assign y2373 = ~1'b0 ;
  assign y2374 = n4354 ;
  assign y2375 = ~n339 ;
  assign y2376 = n4355 ;
  assign y2377 = ~n3339 ;
  assign y2378 = n4356 ;
  assign y2379 = ~n4361 ;
  assign y2380 = ~1'b0 ;
  assign y2381 = ~n4364 ;
  assign y2382 = ~n4366 ;
  assign y2383 = ~n4368 ;
  assign y2384 = n4372 ;
  assign y2385 = ~n667 ;
  assign y2386 = ~1'b0 ;
  assign y2387 = n4373 ;
  assign y2388 = n4375 ;
  assign y2389 = ~1'b0 ;
  assign y2390 = ~n4376 ;
  assign y2391 = ~n4377 ;
  assign y2392 = ~1'b0 ;
  assign y2393 = n4384 ;
  assign y2394 = n4388 ;
  assign y2395 = ~n4334 ;
  assign y2396 = ~1'b0 ;
  assign y2397 = n4390 ;
  assign y2398 = ~n2948 ;
  assign y2399 = n4391 ;
  assign y2400 = ~1'b0 ;
  assign y2401 = ~n2579 ;
  assign y2402 = ~1'b0 ;
  assign y2403 = ~n4397 ;
  assign y2404 = ~n4398 ;
  assign y2405 = n4410 ;
  assign y2406 = ~1'b0 ;
  assign y2407 = ~1'b0 ;
  assign y2408 = ~n4413 ;
  assign y2409 = ~n4415 ;
  assign y2410 = ~1'b0 ;
  assign y2411 = n4416 ;
  assign y2412 = n4419 ;
  assign y2413 = ~n4425 ;
  assign y2414 = n4429 ;
  assign y2415 = ~n4433 ;
  assign y2416 = n4434 ;
  assign y2417 = n4436 ;
  assign y2418 = n4438 ;
  assign y2419 = n4444 ;
  assign y2420 = ~1'b0 ;
  assign y2421 = n4445 ;
  assign y2422 = ~1'b0 ;
  assign y2423 = n4448 ;
  assign y2424 = ~1'b0 ;
  assign y2425 = n4462 ;
  assign y2426 = ~1'b0 ;
  assign y2427 = ~1'b0 ;
  assign y2428 = ~n4464 ;
  assign y2429 = ~n4465 ;
  assign y2430 = ~n4081 ;
  assign y2431 = ~n4471 ;
  assign y2432 = ~n4480 ;
  assign y2433 = ~n4482 ;
  assign y2434 = ~n4485 ;
  assign y2435 = 1'b0 ;
  assign y2436 = n4486 ;
  assign y2437 = ~n4493 ;
  assign y2438 = ~1'b0 ;
  assign y2439 = ~1'b0 ;
  assign y2440 = ~1'b0 ;
  assign y2441 = ~1'b0 ;
  assign y2442 = n4499 ;
  assign y2443 = ~n4501 ;
  assign y2444 = ~1'b0 ;
  assign y2445 = ~1'b0 ;
  assign y2446 = n4503 ;
  assign y2447 = ~n1491 ;
  assign y2448 = ~n4506 ;
  assign y2449 = ~1'b0 ;
  assign y2450 = ~1'b0 ;
  assign y2451 = n4507 ;
  assign y2452 = n4517 ;
  assign y2453 = n4520 ;
  assign y2454 = ~1'b0 ;
  assign y2455 = n4523 ;
  assign y2456 = ~1'b0 ;
  assign y2457 = ~n4527 ;
  assign y2458 = n4532 ;
  assign y2459 = n4549 ;
  assign y2460 = ~n4550 ;
  assign y2461 = ~n4553 ;
  assign y2462 = n4558 ;
  assign y2463 = n4560 ;
  assign y2464 = n4561 ;
  assign y2465 = n4564 ;
  assign y2466 = n4566 ;
  assign y2467 = n4567 ;
  assign y2468 = n1436 ;
  assign y2469 = ~n4568 ;
  assign y2470 = n4569 ;
  assign y2471 = n2019 ;
  assign y2472 = n4570 ;
  assign y2473 = ~1'b0 ;
  assign y2474 = ~n4572 ;
  assign y2475 = ~1'b0 ;
  assign y2476 = n4574 ;
  assign y2477 = ~n4579 ;
  assign y2478 = ~1'b0 ;
  assign y2479 = ~1'b0 ;
  assign y2480 = n4580 ;
  assign y2481 = ~n4585 ;
  assign y2482 = ~n4586 ;
  assign y2483 = ~1'b0 ;
  assign y2484 = n4589 ;
  assign y2485 = ~x46 ;
  assign y2486 = ~n4592 ;
  assign y2487 = ~1'b0 ;
  assign y2488 = n4598 ;
  assign y2489 = n4602 ;
  assign y2490 = ~n656 ;
  assign y2491 = n4603 ;
  assign y2492 = n4605 ;
  assign y2493 = ~n4610 ;
  assign y2494 = n4611 ;
  assign y2495 = n4612 ;
  assign y2496 = ~1'b0 ;
  assign y2497 = n4613 ;
  assign y2498 = ~1'b0 ;
  assign y2499 = ~n4615 ;
  assign y2500 = ~1'b0 ;
  assign y2501 = ~1'b0 ;
  assign y2502 = ~n4616 ;
  assign y2503 = n4618 ;
  assign y2504 = ~1'b0 ;
  assign y2505 = n4619 ;
  assign y2506 = n3482 ;
  assign y2507 = ~1'b0 ;
  assign y2508 = ~n4628 ;
  assign y2509 = n2808 ;
  assign y2510 = ~n4631 ;
  assign y2511 = n4632 ;
  assign y2512 = ~1'b0 ;
  assign y2513 = ~n4636 ;
  assign y2514 = ~n4639 ;
  assign y2515 = ~1'b0 ;
  assign y2516 = n4647 ;
  assign y2517 = n4648 ;
  assign y2518 = n4654 ;
  assign y2519 = ~n4656 ;
  assign y2520 = n4657 ;
  assign y2521 = ~n4660 ;
  assign y2522 = ~n4661 ;
  assign y2523 = ~1'b0 ;
  assign y2524 = ~1'b0 ;
  assign y2525 = n4662 ;
  assign y2526 = ~n4668 ;
  assign y2527 = ~1'b0 ;
  assign y2528 = n4669 ;
  assign y2529 = 1'b0 ;
  assign y2530 = ~1'b0 ;
  assign y2531 = ~1'b0 ;
  assign y2532 = n4673 ;
  assign y2533 = ~n4677 ;
  assign y2534 = ~n4683 ;
  assign y2535 = ~1'b0 ;
  assign y2536 = ~n3911 ;
  assign y2537 = n4685 ;
  assign y2538 = n4687 ;
  assign y2539 = ~1'b0 ;
  assign y2540 = ~n4689 ;
  assign y2541 = n4690 ;
  assign y2542 = ~1'b0 ;
  assign y2543 = n4691 ;
  assign y2544 = 1'b0 ;
  assign y2545 = ~n4692 ;
  assign y2546 = n4693 ;
  assign y2547 = n4699 ;
  assign y2548 = n4703 ;
  assign y2549 = ~n4705 ;
  assign y2550 = ~n4706 ;
  assign y2551 = n4707 ;
  assign y2552 = n4708 ;
  assign y2553 = n4711 ;
  assign y2554 = ~n4718 ;
  assign y2555 = ~1'b0 ;
  assign y2556 = ~1'b0 ;
  assign y2557 = n4720 ;
  assign y2558 = n4726 ;
  assign y2559 = 1'b0 ;
  assign y2560 = ~n4728 ;
  assign y2561 = ~1'b0 ;
  assign y2562 = ~1'b0 ;
  assign y2563 = ~1'b0 ;
  assign y2564 = ~n4730 ;
  assign y2565 = ~n4734 ;
  assign y2566 = n4735 ;
  assign y2567 = n4736 ;
  assign y2568 = ~1'b0 ;
  assign y2569 = n4742 ;
  assign y2570 = ~n4743 ;
  assign y2571 = ~n4745 ;
  assign y2572 = n4747 ;
  assign y2573 = n4752 ;
  assign y2574 = ~n1616 ;
  assign y2575 = n4755 ;
  assign y2576 = ~1'b0 ;
  assign y2577 = n4758 ;
  assign y2578 = n4759 ;
  assign y2579 = n4761 ;
  assign y2580 = 1'b0 ;
  assign y2581 = ~n4765 ;
  assign y2582 = ~n4768 ;
  assign y2583 = ~n4773 ;
  assign y2584 = ~1'b0 ;
  assign y2585 = ~n707 ;
  assign y2586 = ~1'b0 ;
  assign y2587 = ~n4775 ;
  assign y2588 = n4777 ;
  assign y2589 = ~1'b0 ;
  assign y2590 = ~1'b0 ;
  assign y2591 = ~1'b0 ;
  assign y2592 = ~1'b0 ;
  assign y2593 = ~1'b0 ;
  assign y2594 = n3717 ;
  assign y2595 = ~n4781 ;
  assign y2596 = ~1'b0 ;
  assign y2597 = n4784 ;
  assign y2598 = n4790 ;
  assign y2599 = ~1'b0 ;
  assign y2600 = ~n4791 ;
  assign y2601 = ~n4793 ;
  assign y2602 = n4797 ;
  assign y2603 = n4798 ;
  assign y2604 = ~1'b0 ;
  assign y2605 = n4802 ;
  assign y2606 = ~n4804 ;
  assign y2607 = ~1'b0 ;
  assign y2608 = ~n4806 ;
  assign y2609 = ~1'b0 ;
  assign y2610 = n4809 ;
  assign y2611 = ~n4811 ;
  assign y2612 = ~n2456 ;
  assign y2613 = n4296 ;
  assign y2614 = ~n4814 ;
  assign y2615 = n4817 ;
  assign y2616 = 1'b0 ;
  assign y2617 = ~1'b0 ;
  assign y2618 = n4819 ;
  assign y2619 = ~1'b0 ;
  assign y2620 = n4820 ;
  assign y2621 = ~1'b0 ;
  assign y2622 = n4823 ;
  assign y2623 = ~1'b0 ;
  assign y2624 = n4824 ;
  assign y2625 = ~n4825 ;
  assign y2626 = ~n4828 ;
  assign y2627 = ~n4830 ;
  assign y2628 = n4835 ;
  assign y2629 = n4838 ;
  assign y2630 = ~n4842 ;
  assign y2631 = ~n4843 ;
  assign y2632 = n4845 ;
  assign y2633 = n4850 ;
  assign y2634 = ~n4081 ;
  assign y2635 = ~n4851 ;
  assign y2636 = n4854 ;
  assign y2637 = n4856 ;
  assign y2638 = ~n1042 ;
  assign y2639 = ~1'b0 ;
  assign y2640 = n4857 ;
  assign y2641 = n4859 ;
  assign y2642 = n4860 ;
  assign y2643 = ~n4861 ;
  assign y2644 = ~1'b0 ;
  assign y2645 = ~1'b0 ;
  assign y2646 = ~1'b0 ;
  assign y2647 = ~n4865 ;
  assign y2648 = n4873 ;
  assign y2649 = n4877 ;
  assign y2650 = ~1'b0 ;
  assign y2651 = n4878 ;
  assign y2652 = ~1'b0 ;
  assign y2653 = n4882 ;
  assign y2654 = ~n4892 ;
  assign y2655 = ~1'b0 ;
  assign y2656 = ~n4893 ;
  assign y2657 = n4895 ;
  assign y2658 = n4898 ;
  assign y2659 = n4899 ;
  assign y2660 = ~n4906 ;
  assign y2661 = ~1'b0 ;
  assign y2662 = ~1'b0 ;
  assign y2663 = ~1'b0 ;
  assign y2664 = ~n4907 ;
  assign y2665 = ~n4910 ;
  assign y2666 = ~1'b0 ;
  assign y2667 = ~n4914 ;
  assign y2668 = n4915 ;
  assign y2669 = ~n4916 ;
  assign y2670 = ~n4920 ;
  assign y2671 = ~1'b0 ;
  assign y2672 = ~1'b0 ;
  assign y2673 = ~n4926 ;
  assign y2674 = ~n831 ;
  assign y2675 = ~1'b0 ;
  assign y2676 = n4928 ;
  assign y2677 = n4929 ;
  assign y2678 = ~n4933 ;
  assign y2679 = ~n4941 ;
  assign y2680 = n544 ;
  assign y2681 = n4942 ;
  assign y2682 = ~n4947 ;
  assign y2683 = n4948 ;
  assign y2684 = n529 ;
  assign y2685 = ~1'b0 ;
  assign y2686 = n4954 ;
  assign y2687 = ~1'b0 ;
  assign y2688 = n4346 ;
  assign y2689 = 1'b0 ;
  assign y2690 = ~n4956 ;
  assign y2691 = n4961 ;
  assign y2692 = ~n4964 ;
  assign y2693 = ~1'b0 ;
  assign y2694 = ~n4965 ;
  assign y2695 = n4966 ;
  assign y2696 = ~n4967 ;
  assign y2697 = ~n4968 ;
  assign y2698 = ~1'b0 ;
  assign y2699 = n4970 ;
  assign y2700 = n4974 ;
  assign y2701 = 1'b0 ;
  assign y2702 = ~n4978 ;
  assign y2703 = ~n4981 ;
  assign y2704 = n4990 ;
  assign y2705 = ~n4992 ;
  assign y2706 = ~n830 ;
  assign y2707 = ~1'b0 ;
  assign y2708 = ~n4995 ;
  assign y2709 = ~1'b0 ;
  assign y2710 = ~1'b0 ;
  assign y2711 = n2830 ;
  assign y2712 = ~n4996 ;
  assign y2713 = ~n2091 ;
  assign y2714 = ~1'b0 ;
  assign y2715 = n4998 ;
  assign y2716 = ~n5002 ;
  assign y2717 = ~n5003 ;
  assign y2718 = n5004 ;
  assign y2719 = ~1'b0 ;
  assign y2720 = ~n5007 ;
  assign y2721 = ~n5010 ;
  assign y2722 = ~n5011 ;
  assign y2723 = ~1'b0 ;
  assign y2724 = n5016 ;
  assign y2725 = ~1'b0 ;
  assign y2726 = n5018 ;
  assign y2727 = ~1'b0 ;
  assign y2728 = ~1'b0 ;
  assign y2729 = ~1'b0 ;
  assign y2730 = n5031 ;
  assign y2731 = ~n5036 ;
  assign y2732 = ~n5037 ;
  assign y2733 = 1'b0 ;
  assign y2734 = ~1'b0 ;
  assign y2735 = n5039 ;
  assign y2736 = ~1'b0 ;
  assign y2737 = n5040 ;
  assign y2738 = ~n5042 ;
  assign y2739 = ~n5048 ;
  assign y2740 = ~1'b0 ;
  assign y2741 = n5054 ;
  assign y2742 = n5057 ;
  assign y2743 = ~n5060 ;
  assign y2744 = n5065 ;
  assign y2745 = ~n5067 ;
  assign y2746 = ~n3852 ;
  assign y2747 = ~n5072 ;
  assign y2748 = ~n5074 ;
  assign y2749 = ~1'b0 ;
  assign y2750 = ~1'b0 ;
  assign y2751 = n5076 ;
  assign y2752 = ~1'b0 ;
  assign y2753 = ~n5085 ;
  assign y2754 = ~n5086 ;
  assign y2755 = 1'b0 ;
  assign y2756 = n5087 ;
  assign y2757 = n325 ;
  assign y2758 = x16 ;
  assign y2759 = ~n5090 ;
  assign y2760 = ~1'b0 ;
  assign y2761 = n5091 ;
  assign y2762 = n5093 ;
  assign y2763 = ~n5097 ;
  assign y2764 = ~n5098 ;
  assign y2765 = ~1'b0 ;
  assign y2766 = ~1'b0 ;
  assign y2767 = ~n5099 ;
  assign y2768 = ~1'b0 ;
  assign y2769 = ~1'b0 ;
  assign y2770 = ~n5101 ;
  assign y2771 = ~1'b0 ;
  assign y2772 = n3064 ;
  assign y2773 = ~1'b0 ;
  assign y2774 = ~n390 ;
  assign y2775 = ~1'b0 ;
  assign y2776 = ~1'b0 ;
  assign y2777 = n5102 ;
  assign y2778 = ~1'b0 ;
  assign y2779 = ~1'b0 ;
  assign y2780 = ~n5103 ;
  assign y2781 = ~1'b0 ;
  assign y2782 = ~n5105 ;
  assign y2783 = n5106 ;
  assign y2784 = n5110 ;
  assign y2785 = ~1'b0 ;
  assign y2786 = ~n5115 ;
  assign y2787 = 1'b0 ;
  assign y2788 = ~n5120 ;
  assign y2789 = ~n5121 ;
  assign y2790 = n5122 ;
  assign y2791 = n5123 ;
  assign y2792 = ~n3764 ;
  assign y2793 = ~1'b0 ;
  assign y2794 = n5127 ;
  assign y2795 = ~n5128 ;
  assign y2796 = ~1'b0 ;
  assign y2797 = ~1'b0 ;
  assign y2798 = ~1'b0 ;
  assign y2799 = n5130 ;
  assign y2800 = n5132 ;
  assign y2801 = ~1'b0 ;
  assign y2802 = ~1'b0 ;
  assign y2803 = ~1'b0 ;
  assign y2804 = ~1'b0 ;
  assign y2805 = ~1'b0 ;
  assign y2806 = ~1'b0 ;
  assign y2807 = n361 ;
  assign y2808 = ~n4958 ;
  assign y2809 = n5140 ;
  assign y2810 = n5143 ;
  assign y2811 = ~n4966 ;
  assign y2812 = n5152 ;
  assign y2813 = n5156 ;
  assign y2814 = ~n5158 ;
  assign y2815 = n5159 ;
  assign y2816 = ~1'b0 ;
  assign y2817 = ~1'b0 ;
  assign y2818 = ~n5059 ;
  assign y2819 = n5161 ;
  assign y2820 = n5168 ;
  assign y2821 = ~1'b0 ;
  assign y2822 = ~n5172 ;
  assign y2823 = n5176 ;
  assign y2824 = n5178 ;
  assign y2825 = ~1'b0 ;
  assign y2826 = ~n514 ;
  assign y2827 = 1'b0 ;
  assign y2828 = ~1'b0 ;
  assign y2829 = ~1'b0 ;
  assign y2830 = ~n5019 ;
  assign y2831 = ~1'b0 ;
  assign y2832 = n5179 ;
  assign y2833 = ~1'b0 ;
  assign y2834 = n5182 ;
  assign y2835 = n5184 ;
  assign y2836 = ~n3764 ;
  assign y2837 = n5193 ;
  assign y2838 = n5195 ;
  assign y2839 = ~n5196 ;
  assign y2840 = ~1'b0 ;
  assign y2841 = n5197 ;
  assign y2842 = ~n5198 ;
  assign y2843 = ~1'b0 ;
  assign y2844 = ~n3193 ;
  assign y2845 = ~1'b0 ;
  assign y2846 = ~1'b0 ;
  assign y2847 = n5200 ;
  assign y2848 = ~1'b0 ;
  assign y2849 = n5205 ;
  assign y2850 = n5211 ;
  assign y2851 = n5215 ;
  assign y2852 = n5217 ;
  assign y2853 = 1'b0 ;
  assign y2854 = ~1'b0 ;
  assign y2855 = ~1'b0 ;
  assign y2856 = ~n5219 ;
  assign y2857 = ~n5220 ;
  assign y2858 = ~n5226 ;
  assign y2859 = n5230 ;
  assign y2860 = ~1'b0 ;
  assign y2861 = ~n5231 ;
  assign y2862 = n5232 ;
  assign y2863 = ~n5233 ;
  assign y2864 = n5234 ;
  assign y2865 = 1'b0 ;
  assign y2866 = n5237 ;
  assign y2867 = ~1'b0 ;
  assign y2868 = ~n5240 ;
  assign y2869 = ~n5241 ;
  assign y2870 = ~1'b0 ;
  assign y2871 = n5242 ;
  assign y2872 = n5243 ;
  assign y2873 = ~1'b0 ;
  assign y2874 = ~1'b0 ;
  assign y2875 = n5245 ;
  assign y2876 = ~n5246 ;
  assign y2877 = ~n5247 ;
  assign y2878 = ~1'b0 ;
  assign y2879 = n5248 ;
  assign y2880 = ~n5249 ;
  assign y2881 = ~1'b0 ;
  assign y2882 = n5251 ;
  assign y2883 = ~1'b0 ;
  assign y2884 = n5252 ;
  assign y2885 = ~n5253 ;
  assign y2886 = n5254 ;
  assign y2887 = ~1'b0 ;
  assign y2888 = ~n5257 ;
  assign y2889 = n5258 ;
  assign y2890 = ~n5259 ;
  assign y2891 = ~1'b0 ;
  assign y2892 = n5263 ;
  assign y2893 = n5268 ;
  assign y2894 = ~n5271 ;
  assign y2895 = n5273 ;
  assign y2896 = ~1'b0 ;
  assign y2897 = n5278 ;
  assign y2898 = ~1'b0 ;
  assign y2899 = ~1'b0 ;
  assign y2900 = 1'b0 ;
  assign y2901 = ~n5280 ;
  assign y2902 = ~n5282 ;
  assign y2903 = ~n1423 ;
  assign y2904 = ~1'b0 ;
  assign y2905 = 1'b0 ;
  assign y2906 = n5283 ;
  assign y2907 = ~1'b0 ;
  assign y2908 = ~n5290 ;
  assign y2909 = ~1'b0 ;
  assign y2910 = ~n5292 ;
  assign y2911 = ~1'b0 ;
  assign y2912 = ~n5297 ;
  assign y2913 = ~n5300 ;
  assign y2914 = ~n5302 ;
  assign y2915 = ~1'b0 ;
  assign y2916 = n5308 ;
  assign y2917 = ~n3272 ;
  assign y2918 = n5309 ;
  assign y2919 = n5310 ;
  assign y2920 = n5313 ;
  assign y2921 = ~1'b0 ;
  assign y2922 = ~1'b0 ;
  assign y2923 = ~1'b0 ;
  assign y2924 = ~n5315 ;
  assign y2925 = ~n5318 ;
  assign y2926 = n5320 ;
  assign y2927 = ~n5321 ;
  assign y2928 = ~1'b0 ;
  assign y2929 = ~n5324 ;
  assign y2930 = n5328 ;
  assign y2931 = ~n2585 ;
  assign y2932 = n5329 ;
  assign y2933 = n5332 ;
  assign y2934 = ~1'b0 ;
  assign y2935 = n5333 ;
  assign y2936 = ~1'b0 ;
  assign y2937 = ~1'b0 ;
  assign y2938 = ~n5337 ;
  assign y2939 = ~1'b0 ;
  assign y2940 = n5341 ;
  assign y2941 = n724 ;
  assign y2942 = ~1'b0 ;
  assign y2943 = ~n5346 ;
  assign y2944 = n5347 ;
  assign y2945 = ~1'b0 ;
  assign y2946 = n5349 ;
  assign y2947 = ~n5356 ;
  assign y2948 = n5358 ;
  assign y2949 = n5360 ;
  assign y2950 = ~1'b0 ;
  assign y2951 = ~n5361 ;
  assign y2952 = n5363 ;
  assign y2953 = ~n5372 ;
  assign y2954 = ~n5373 ;
  assign y2955 = ~n5377 ;
  assign y2956 = ~1'b0 ;
  assign y2957 = n5378 ;
  assign y2958 = n5387 ;
  assign y2959 = ~n5388 ;
  assign y2960 = ~n5390 ;
  assign y2961 = ~n5392 ;
  assign y2962 = n5397 ;
  assign y2963 = ~n5399 ;
  assign y2964 = ~n5400 ;
  assign y2965 = ~1'b0 ;
  assign y2966 = ~1'b0 ;
  assign y2967 = n5404 ;
  assign y2968 = n5410 ;
  assign y2969 = n5369 ;
  assign y2970 = n5411 ;
  assign y2971 = ~n5414 ;
  assign y2972 = x124 ;
  assign y2973 = ~1'b0 ;
  assign y2974 = n5415 ;
  assign y2975 = ~n5417 ;
  assign y2976 = ~1'b0 ;
  assign y2977 = ~n5420 ;
  assign y2978 = ~1'b0 ;
  assign y2979 = ~1'b0 ;
  assign y2980 = ~1'b0 ;
  assign y2981 = n5424 ;
  assign y2982 = n5429 ;
  assign y2983 = ~1'b0 ;
  assign y2984 = ~n5430 ;
  assign y2985 = n5432 ;
  assign y2986 = ~1'b0 ;
  assign y2987 = ~n1487 ;
  assign y2988 = ~n5436 ;
  assign y2989 = ~1'b0 ;
  assign y2990 = n5437 ;
  assign y2991 = n5438 ;
  assign y2992 = n5439 ;
  assign y2993 = n5440 ;
  assign y2994 = ~n5445 ;
  assign y2995 = ~n5450 ;
  assign y2996 = ~1'b0 ;
  assign y2997 = n5451 ;
  assign y2998 = ~n5460 ;
  assign y2999 = ~1'b0 ;
  assign y3000 = ~1'b0 ;
  assign y3001 = ~1'b0 ;
  assign y3002 = ~n5463 ;
  assign y3003 = ~1'b0 ;
  assign y3004 = ~n5464 ;
  assign y3005 = n5466 ;
  assign y3006 = 1'b0 ;
  assign y3007 = ~1'b0 ;
  assign y3008 = n5467 ;
  assign y3009 = ~n1133 ;
  assign y3010 = ~n5470 ;
  assign y3011 = n5475 ;
  assign y3012 = ~1'b0 ;
  assign y3013 = n5476 ;
  assign y3014 = n5479 ;
  assign y3015 = ~n5482 ;
  assign y3016 = n5483 ;
  assign y3017 = n3906 ;
  assign y3018 = ~1'b0 ;
  assign y3019 = n5486 ;
  assign y3020 = ~n1179 ;
  assign y3021 = ~1'b0 ;
  assign y3022 = n5491 ;
  assign y3023 = n5492 ;
  assign y3024 = ~n5510 ;
  assign y3025 = ~n5516 ;
  assign y3026 = ~1'b0 ;
  assign y3027 = n5517 ;
  assign y3028 = ~1'b0 ;
  assign y3029 = ~1'b0 ;
  assign y3030 = ~n5524 ;
  assign y3031 = n5526 ;
  assign y3032 = n1891 ;
  assign y3033 = ~1'b0 ;
  assign y3034 = n5528 ;
  assign y3035 = ~1'b0 ;
  assign y3036 = ~n5534 ;
  assign y3037 = ~1'b0 ;
  assign y3038 = ~1'b0 ;
  assign y3039 = ~n5536 ;
  assign y3040 = ~1'b0 ;
  assign y3041 = ~n5537 ;
  assign y3042 = ~n5540 ;
  assign y3043 = n211 ;
  assign y3044 = 1'b0 ;
  assign y3045 = n5541 ;
  assign y3046 = ~1'b0 ;
  assign y3047 = 1'b0 ;
  assign y3048 = n5549 ;
  assign y3049 = ~n5550 ;
  assign y3050 = ~n3934 ;
  assign y3051 = n358 ;
  assign y3052 = n2878 ;
  assign y3053 = n5552 ;
  assign y3054 = n5555 ;
  assign y3055 = n5556 ;
  assign y3056 = n5558 ;
  assign y3057 = ~1'b0 ;
  assign y3058 = n5559 ;
  assign y3059 = ~1'b0 ;
  assign y3060 = ~n5560 ;
  assign y3061 = 1'b0 ;
  assign y3062 = ~1'b0 ;
  assign y3063 = n5562 ;
  assign y3064 = ~1'b0 ;
  assign y3065 = ~1'b0 ;
  assign y3066 = ~n5566 ;
  assign y3067 = ~1'b0 ;
  assign y3068 = ~1'b0 ;
  assign y3069 = ~n5572 ;
  assign y3070 = ~1'b0 ;
  assign y3071 = ~n5573 ;
  assign y3072 = ~n5574 ;
  assign y3073 = n5575 ;
  assign y3074 = n1685 ;
  assign y3075 = ~n5579 ;
  assign y3076 = ~n5580 ;
  assign y3077 = n5583 ;
  assign y3078 = ~1'b0 ;
  assign y3079 = ~n5584 ;
  assign y3080 = ~n5588 ;
  assign y3081 = ~1'b0 ;
  assign y3082 = n5589 ;
  assign y3083 = ~n5590 ;
  assign y3084 = ~1'b0 ;
  assign y3085 = ~n5593 ;
  assign y3086 = n5594 ;
  assign y3087 = ~n5600 ;
  assign y3088 = ~n5605 ;
  assign y3089 = n5606 ;
  assign y3090 = n5608 ;
  assign y3091 = n5613 ;
  assign y3092 = ~n5615 ;
  assign y3093 = ~1'b0 ;
  assign y3094 = ~1'b0 ;
  assign y3095 = ~1'b0 ;
  assign y3096 = ~n5622 ;
  assign y3097 = n5623 ;
  assign y3098 = 1'b0 ;
  assign y3099 = ~n5629 ;
  assign y3100 = n5634 ;
  assign y3101 = ~n5638 ;
  assign y3102 = n5642 ;
  assign y3103 = ~1'b0 ;
  assign y3104 = ~1'b0 ;
  assign y3105 = 1'b0 ;
  assign y3106 = n5643 ;
  assign y3107 = ~n5648 ;
  assign y3108 = n5649 ;
  assign y3109 = n5651 ;
  assign y3110 = ~1'b0 ;
  assign y3111 = ~1'b0 ;
  assign y3112 = ~1'b0 ;
  assign y3113 = ~1'b0 ;
  assign y3114 = ~1'b0 ;
  assign y3115 = n5653 ;
  assign y3116 = n5654 ;
  assign y3117 = n5658 ;
  assign y3118 = ~1'b0 ;
  assign y3119 = ~1'b0 ;
  assign y3120 = n5532 ;
  assign y3121 = ~1'b0 ;
  assign y3122 = n5659 ;
  assign y3123 = n5661 ;
  assign y3124 = n5258 ;
  assign y3125 = ~n5663 ;
  assign y3126 = n5667 ;
  assign y3127 = ~n5672 ;
  assign y3128 = ~n5676 ;
  assign y3129 = ~1'b0 ;
  assign y3130 = ~n5683 ;
  assign y3131 = ~n5685 ;
  assign y3132 = ~n5687 ;
  assign y3133 = ~1'b0 ;
  assign y3134 = n5691 ;
  assign y3135 = ~1'b0 ;
  assign y3136 = ~1'b0 ;
  assign y3137 = ~n4350 ;
  assign y3138 = ~n3415 ;
  assign y3139 = n5692 ;
  assign y3140 = ~n5693 ;
  assign y3141 = ~n5698 ;
  assign y3142 = n5700 ;
  assign y3143 = n5705 ;
  assign y3144 = ~n5709 ;
  assign y3145 = ~1'b0 ;
  assign y3146 = n5713 ;
  assign y3147 = n5716 ;
  assign y3148 = ~n5718 ;
  assign y3149 = ~n5720 ;
  assign y3150 = ~n5722 ;
  assign y3151 = n5726 ;
  assign y3152 = ~n3780 ;
  assign y3153 = n5727 ;
  assign y3154 = ~n5729 ;
  assign y3155 = ~n5732 ;
  assign y3156 = n5733 ;
  assign y3157 = n5745 ;
  assign y3158 = ~n5746 ;
  assign y3159 = n5753 ;
  assign y3160 = ~1'b0 ;
  assign y3161 = ~1'b0 ;
  assign y3162 = ~n5755 ;
  assign y3163 = ~n5757 ;
  assign y3164 = n5758 ;
  assign y3165 = ~n5760 ;
  assign y3166 = n5761 ;
  assign y3167 = ~1'b0 ;
  assign y3168 = ~n4589 ;
  assign y3169 = ~n5763 ;
  assign y3170 = n5764 ;
  assign y3171 = ~n2978 ;
  assign y3172 = ~n5768 ;
  assign y3173 = n5771 ;
  assign y3174 = 1'b0 ;
  assign y3175 = ~1'b0 ;
  assign y3176 = n5778 ;
  assign y3177 = ~n5779 ;
  assign y3178 = ~n5782 ;
  assign y3179 = ~1'b0 ;
  assign y3180 = ~1'b0 ;
  assign y3181 = ~n5787 ;
  assign y3182 = n5791 ;
  assign y3183 = ~1'b0 ;
  assign y3184 = ~1'b0 ;
  assign y3185 = n5794 ;
  assign y3186 = n5796 ;
  assign y3187 = n5801 ;
  assign y3188 = ~n5804 ;
  assign y3189 = ~1'b0 ;
  assign y3190 = ~n5807 ;
  assign y3191 = ~1'b0 ;
  assign y3192 = ~n5809 ;
  assign y3193 = ~1'b0 ;
  assign y3194 = ~n5814 ;
  assign y3195 = n5817 ;
  assign y3196 = ~1'b0 ;
  assign y3197 = n5821 ;
  assign y3198 = n5822 ;
  assign y3199 = ~1'b0 ;
  assign y3200 = ~n5826 ;
  assign y3201 = ~n5834 ;
  assign y3202 = ~n5836 ;
  assign y3203 = n5837 ;
  assign y3204 = ~1'b0 ;
  assign y3205 = ~1'b0 ;
  assign y3206 = n5838 ;
  assign y3207 = ~1'b0 ;
  assign y3208 = ~1'b0 ;
  assign y3209 = n5840 ;
  assign y3210 = ~1'b0 ;
  assign y3211 = ~1'b0 ;
  assign y3212 = n5842 ;
  assign y3213 = n5854 ;
  assign y3214 = ~n5855 ;
  assign y3215 = n5857 ;
  assign y3216 = n5862 ;
  assign y3217 = ~n5865 ;
  assign y3218 = ~1'b0 ;
  assign y3219 = ~1'b0 ;
  assign y3220 = ~1'b0 ;
  assign y3221 = n3426 ;
  assign y3222 = n5866 ;
  assign y3223 = ~n728 ;
  assign y3224 = n5867 ;
  assign y3225 = ~n5871 ;
  assign y3226 = ~n5874 ;
  assign y3227 = ~n5875 ;
  assign y3228 = ~n5876 ;
  assign y3229 = n5878 ;
  assign y3230 = ~1'b0 ;
  assign y3231 = ~1'b0 ;
  assign y3232 = ~n5880 ;
  assign y3233 = ~1'b0 ;
  assign y3234 = ~n5882 ;
  assign y3235 = ~1'b0 ;
  assign y3236 = ~1'b0 ;
  assign y3237 = n5887 ;
  assign y3238 = n5889 ;
  assign y3239 = n5890 ;
  assign y3240 = ~1'b0 ;
  assign y3241 = ~n5891 ;
  assign y3242 = n5894 ;
  assign y3243 = ~n5897 ;
  assign y3244 = ~1'b0 ;
  assign y3245 = ~n5900 ;
  assign y3246 = ~n5903 ;
  assign y3247 = ~1'b0 ;
  assign y3248 = ~1'b0 ;
  assign y3249 = n5904 ;
  assign y3250 = n5909 ;
  assign y3251 = n356 ;
  assign y3252 = n5912 ;
  assign y3253 = ~n5918 ;
  assign y3254 = ~n5920 ;
  assign y3255 = n5923 ;
  assign y3256 = n5924 ;
  assign y3257 = ~1'b0 ;
  assign y3258 = ~1'b0 ;
  assign y3259 = n5926 ;
  assign y3260 = ~n5931 ;
  assign y3261 = ~n2570 ;
  assign y3262 = n5933 ;
  assign y3263 = ~1'b0 ;
  assign y3264 = n5935 ;
  assign y3265 = ~n221 ;
  assign y3266 = n5938 ;
  assign y3267 = ~1'b0 ;
  assign y3268 = ~n5943 ;
  assign y3269 = ~1'b0 ;
  assign y3270 = ~1'b0 ;
  assign y3271 = n5944 ;
  assign y3272 = ~n5946 ;
  assign y3273 = n5947 ;
  assign y3274 = ~1'b0 ;
  assign y3275 = ~1'b0 ;
  assign y3276 = ~n5950 ;
  assign y3277 = ~1'b0 ;
  assign y3278 = 1'b0 ;
  assign y3279 = ~1'b0 ;
  assign y3280 = ~1'b0 ;
  assign y3281 = ~n5951 ;
  assign y3282 = ~1'b0 ;
  assign y3283 = ~1'b0 ;
  assign y3284 = n5956 ;
  assign y3285 = ~n5958 ;
  assign y3286 = ~n5965 ;
  assign y3287 = ~n5966 ;
  assign y3288 = ~n5973 ;
  assign y3289 = n5974 ;
  assign y3290 = ~1'b0 ;
  assign y3291 = ~1'b0 ;
  assign y3292 = ~1'b0 ;
  assign y3293 = n5975 ;
  assign y3294 = ~n5977 ;
  assign y3295 = ~1'b0 ;
  assign y3296 = n5979 ;
  assign y3297 = ~1'b0 ;
  assign y3298 = ~n5980 ;
  assign y3299 = ~n5981 ;
  assign y3300 = ~1'b0 ;
  assign y3301 = ~1'b0 ;
  assign y3302 = n5984 ;
  assign y3303 = n5986 ;
  assign y3304 = ~1'b0 ;
  assign y3305 = ~1'b0 ;
  assign y3306 = ~n5996 ;
  assign y3307 = ~n6001 ;
  assign y3308 = ~1'b0 ;
  assign y3309 = ~n6004 ;
  assign y3310 = n6012 ;
  assign y3311 = ~n6016 ;
  assign y3312 = 1'b0 ;
  assign y3313 = ~n6017 ;
  assign y3314 = ~n6018 ;
  assign y3315 = ~n6019 ;
  assign y3316 = ~n6020 ;
  assign y3317 = ~1'b0 ;
  assign y3318 = n6023 ;
  assign y3319 = n6027 ;
  assign y3320 = n6030 ;
  assign y3321 = 1'b0 ;
  assign y3322 = 1'b0 ;
  assign y3323 = ~1'b0 ;
  assign y3324 = n6036 ;
  assign y3325 = ~1'b0 ;
  assign y3326 = n6041 ;
  assign y3327 = n3407 ;
  assign y3328 = ~1'b0 ;
  assign y3329 = n6045 ;
  assign y3330 = n6046 ;
  assign y3331 = ~1'b0 ;
  assign y3332 = 1'b0 ;
  assign y3333 = x77 ;
  assign y3334 = n6047 ;
  assign y3335 = ~1'b0 ;
  assign y3336 = ~n4190 ;
  assign y3337 = ~1'b0 ;
  assign y3338 = n6050 ;
  assign y3339 = n6054 ;
  assign y3340 = n2073 ;
  assign y3341 = n6057 ;
  assign y3342 = ~n3979 ;
  assign y3343 = ~n6062 ;
  assign y3344 = ~n6064 ;
  assign y3345 = ~x37 ;
  assign y3346 = n6067 ;
  assign y3347 = ~1'b0 ;
  assign y3348 = ~1'b0 ;
  assign y3349 = ~1'b0 ;
  assign y3350 = ~1'b0 ;
  assign y3351 = ~n6069 ;
  assign y3352 = n6070 ;
  assign y3353 = ~n6071 ;
  assign y3354 = n6075 ;
  assign y3355 = ~n6080 ;
  assign y3356 = ~n6083 ;
  assign y3357 = ~1'b0 ;
  assign y3358 = ~n6084 ;
  assign y3359 = ~1'b0 ;
  assign y3360 = ~n6086 ;
  assign y3361 = ~1'b0 ;
  assign y3362 = ~1'b0 ;
  assign y3363 = n6089 ;
  assign y3364 = ~1'b0 ;
  assign y3365 = ~1'b0 ;
  assign y3366 = n6091 ;
  assign y3367 = ~1'b0 ;
  assign y3368 = ~1'b0 ;
  assign y3369 = ~n4304 ;
  assign y3370 = n6092 ;
  assign y3371 = n6094 ;
  assign y3372 = n6096 ;
  assign y3373 = ~n6101 ;
  assign y3374 = ~1'b0 ;
  assign y3375 = ~1'b0 ;
  assign y3376 = ~n6102 ;
  assign y3377 = ~1'b0 ;
  assign y3378 = ~1'b0 ;
  assign y3379 = x84 ;
  assign y3380 = n6106 ;
  assign y3381 = ~n1162 ;
  assign y3382 = n6108 ;
  assign y3383 = ~1'b0 ;
  assign y3384 = n6112 ;
  assign y3385 = ~1'b0 ;
  assign y3386 = n2291 ;
  assign y3387 = ~1'b0 ;
  assign y3388 = ~n6114 ;
  assign y3389 = ~n6116 ;
  assign y3390 = ~1'b0 ;
  assign y3391 = ~1'b0 ;
  assign y3392 = ~1'b0 ;
  assign y3393 = ~1'b0 ;
  assign y3394 = ~n6117 ;
  assign y3395 = ~1'b0 ;
  assign y3396 = ~n6121 ;
  assign y3397 = ~n6129 ;
  assign y3398 = n4005 ;
  assign y3399 = ~n3172 ;
  assign y3400 = 1'b0 ;
  assign y3401 = ~n6057 ;
  assign y3402 = n6131 ;
  assign y3403 = ~n6132 ;
  assign y3404 = ~1'b0 ;
  assign y3405 = ~n6142 ;
  assign y3406 = ~n6144 ;
  assign y3407 = ~1'b0 ;
  assign y3408 = n6147 ;
  assign y3409 = ~n5704 ;
  assign y3410 = n6149 ;
  assign y3411 = n6153 ;
  assign y3412 = ~n6155 ;
  assign y3413 = ~1'b0 ;
  assign y3414 = ~1'b0 ;
  assign y3415 = 1'b0 ;
  assign y3416 = n6159 ;
  assign y3417 = n6162 ;
  assign y3418 = n4366 ;
  assign y3419 = ~1'b0 ;
  assign y3420 = n6164 ;
  assign y3421 = ~1'b0 ;
  assign y3422 = ~n6166 ;
  assign y3423 = ~n6171 ;
  assign y3424 = ~n6175 ;
  assign y3425 = ~n6178 ;
  assign y3426 = ~n6186 ;
  assign y3427 = ~1'b0 ;
  assign y3428 = n5280 ;
  assign y3429 = ~1'b0 ;
  assign y3430 = 1'b0 ;
  assign y3431 = ~n6188 ;
  assign y3432 = ~n6192 ;
  assign y3433 = n6114 ;
  assign y3434 = ~1'b0 ;
  assign y3435 = ~1'b0 ;
  assign y3436 = ~1'b0 ;
  assign y3437 = n6193 ;
  assign y3438 = n6197 ;
  assign y3439 = ~1'b0 ;
  assign y3440 = ~n6206 ;
  assign y3441 = ~n6207 ;
  assign y3442 = n6208 ;
  assign y3443 = n6211 ;
  assign y3444 = n6212 ;
  assign y3445 = n6217 ;
  assign y3446 = 1'b0 ;
  assign y3447 = n6220 ;
  assign y3448 = ~1'b0 ;
  assign y3449 = 1'b0 ;
  assign y3450 = ~1'b0 ;
  assign y3451 = ~1'b0 ;
  assign y3452 = ~n6222 ;
  assign y3453 = ~1'b0 ;
  assign y3454 = ~n5442 ;
  assign y3455 = n6223 ;
  assign y3456 = ~1'b0 ;
  assign y3457 = n6224 ;
  assign y3458 = n6226 ;
  assign y3459 = n6227 ;
  assign y3460 = ~1'b0 ;
  assign y3461 = n6233 ;
  assign y3462 = n6236 ;
  assign y3463 = n6237 ;
  assign y3464 = ~n5347 ;
  assign y3465 = n6239 ;
  assign y3466 = n6240 ;
  assign y3467 = ~1'b0 ;
  assign y3468 = 1'b0 ;
  assign y3469 = n6241 ;
  assign y3470 = 1'b0 ;
  assign y3471 = ~1'b0 ;
  assign y3472 = ~n6242 ;
  assign y3473 = ~1'b0 ;
  assign y3474 = n6247 ;
  assign y3475 = ~1'b0 ;
  assign y3476 = ~n6251 ;
  assign y3477 = ~1'b0 ;
  assign y3478 = ~1'b0 ;
  assign y3479 = ~1'b0 ;
  assign y3480 = ~1'b0 ;
  assign y3481 = ~1'b0 ;
  assign y3482 = ~n6256 ;
  assign y3483 = n3286 ;
  assign y3484 = n6259 ;
  assign y3485 = ~n6260 ;
  assign y3486 = n6261 ;
  assign y3487 = n6263 ;
  assign y3488 = n6268 ;
  assign y3489 = n6270 ;
  assign y3490 = ~1'b0 ;
  assign y3491 = ~n6272 ;
  assign y3492 = n6278 ;
  assign y3493 = ~1'b0 ;
  assign y3494 = ~1'b0 ;
  assign y3495 = ~n6281 ;
  assign y3496 = ~1'b0 ;
  assign y3497 = n272 ;
  assign y3498 = n6283 ;
  assign y3499 = ~n6286 ;
  assign y3500 = ~n6288 ;
  assign y3501 = ~1'b0 ;
  assign y3502 = n6294 ;
  assign y3503 = n6299 ;
  assign y3504 = ~1'b0 ;
  assign y3505 = ~1'b0 ;
  assign y3506 = ~1'b0 ;
  assign y3507 = n6306 ;
  assign y3508 = n6307 ;
  assign y3509 = n6309 ;
  assign y3510 = n6313 ;
  assign y3511 = ~1'b0 ;
  assign y3512 = ~n6317 ;
  assign y3513 = n6318 ;
  assign y3514 = n6319 ;
  assign y3515 = ~1'b0 ;
  assign y3516 = n1281 ;
  assign y3517 = ~1'b0 ;
  assign y3518 = ~n6320 ;
  assign y3519 = ~n6321 ;
  assign y3520 = ~1'b0 ;
  assign y3521 = ~n6322 ;
  assign y3522 = ~n6324 ;
  assign y3523 = ~n6328 ;
  assign y3524 = ~1'b0 ;
  assign y3525 = ~1'b0 ;
  assign y3526 = ~1'b0 ;
  assign y3527 = n5801 ;
  assign y3528 = ~1'b0 ;
  assign y3529 = ~1'b0 ;
  assign y3530 = ~n6330 ;
  assign y3531 = ~n6335 ;
  assign y3532 = n6336 ;
  assign y3533 = n4081 ;
  assign y3534 = n6340 ;
  assign y3535 = ~1'b0 ;
  assign y3536 = ~1'b0 ;
  assign y3537 = n6341 ;
  assign y3538 = n6350 ;
  assign y3539 = ~n6357 ;
  assign y3540 = ~n6358 ;
  assign y3541 = n6360 ;
  assign y3542 = n6361 ;
  assign y3543 = ~1'b0 ;
  assign y3544 = ~n6362 ;
  assign y3545 = n6366 ;
  assign y3546 = ~n2775 ;
  assign y3547 = 1'b0 ;
  assign y3548 = ~n6370 ;
  assign y3549 = ~1'b0 ;
  assign y3550 = ~n1335 ;
  assign y3551 = ~n6373 ;
  assign y3552 = n6377 ;
  assign y3553 = n6385 ;
  assign y3554 = n4804 ;
  assign y3555 = ~n6388 ;
  assign y3556 = ~1'b0 ;
  assign y3557 = ~n6389 ;
  assign y3558 = 1'b0 ;
  assign y3559 = ~n6391 ;
  assign y3560 = ~n6393 ;
  assign y3561 = n6394 ;
  assign y3562 = ~1'b0 ;
  assign y3563 = n6401 ;
  assign y3564 = ~n6402 ;
  assign y3565 = ~n6404 ;
  assign y3566 = ~1'b0 ;
  assign y3567 = ~n6406 ;
  assign y3568 = n6408 ;
  assign y3569 = ~n6414 ;
  assign y3570 = ~n6418 ;
  assign y3571 = ~n6419 ;
  assign y3572 = ~1'b0 ;
  assign y3573 = n6422 ;
  assign y3574 = ~n6425 ;
  assign y3575 = ~1'b0 ;
  assign y3576 = n6427 ;
  assign y3577 = ~x12 ;
  assign y3578 = ~1'b0 ;
  assign y3579 = ~n6428 ;
  assign y3580 = ~1'b0 ;
  assign y3581 = ~n6429 ;
  assign y3582 = ~1'b0 ;
  assign y3583 = ~1'b0 ;
  assign y3584 = ~1'b0 ;
  assign y3585 = ~n6432 ;
  assign y3586 = ~n6433 ;
  assign y3587 = ~n6436 ;
  assign y3588 = ~n6441 ;
  assign y3589 = ~1'b0 ;
  assign y3590 = n3494 ;
  assign y3591 = ~n6442 ;
  assign y3592 = n6444 ;
  assign y3593 = n6445 ;
  assign y3594 = n6448 ;
  assign y3595 = n6449 ;
  assign y3596 = ~1'b0 ;
  assign y3597 = 1'b0 ;
  assign y3598 = ~n6455 ;
  assign y3599 = n6457 ;
  assign y3600 = ~1'b0 ;
  assign y3601 = ~n6467 ;
  assign y3602 = ~n6469 ;
  assign y3603 = ~1'b0 ;
  assign y3604 = ~1'b0 ;
  assign y3605 = ~1'b0 ;
  assign y3606 = n6470 ;
  assign y3607 = ~1'b0 ;
  assign y3608 = ~n6471 ;
  assign y3609 = n568 ;
  assign y3610 = ~n5367 ;
  assign y3611 = ~1'b0 ;
  assign y3612 = ~n4900 ;
  assign y3613 = n4833 ;
  assign y3614 = ~1'b0 ;
  assign y3615 = ~n6482 ;
  assign y3616 = n6485 ;
  assign y3617 = n6486 ;
  assign y3618 = n6492 ;
  assign y3619 = ~1'b0 ;
  assign y3620 = ~n6493 ;
  assign y3621 = n6494 ;
  assign y3622 = ~n6495 ;
  assign y3623 = n6496 ;
  assign y3624 = ~1'b0 ;
  assign y3625 = ~1'b0 ;
  assign y3626 = n6497 ;
  assign y3627 = n2819 ;
  assign y3628 = ~1'b0 ;
  assign y3629 = n6505 ;
  assign y3630 = ~n6507 ;
  assign y3631 = n6508 ;
  assign y3632 = ~n6509 ;
  assign y3633 = n6512 ;
  assign y3634 = n6517 ;
  assign y3635 = ~1'b0 ;
  assign y3636 = ~n6520 ;
  assign y3637 = n6525 ;
  assign y3638 = ~1'b0 ;
  assign y3639 = ~n6527 ;
  assign y3640 = n6530 ;
  assign y3641 = ~n1116 ;
  assign y3642 = n6533 ;
  assign y3643 = ~1'b0 ;
  assign y3644 = n6539 ;
  assign y3645 = ~1'b0 ;
  assign y3646 = ~1'b0 ;
  assign y3647 = ~n4318 ;
  assign y3648 = ~n6542 ;
  assign y3649 = ~1'b0 ;
  assign y3650 = n6549 ;
  assign y3651 = ~n6554 ;
  assign y3652 = ~n6555 ;
  assign y3653 = ~1'b0 ;
  assign y3654 = ~n6557 ;
  assign y3655 = n6559 ;
  assign y3656 = n6562 ;
  assign y3657 = ~1'b0 ;
  assign y3658 = n6563 ;
  assign y3659 = n6159 ;
  assign y3660 = n4117 ;
  assign y3661 = n6564 ;
  assign y3662 = n6566 ;
  assign y3663 = ~n4648 ;
  assign y3664 = 1'b0 ;
  assign y3665 = ~1'b0 ;
  assign y3666 = ~1'b0 ;
  assign y3667 = ~n6569 ;
  assign y3668 = n6575 ;
  assign y3669 = n3295 ;
  assign y3670 = ~n6578 ;
  assign y3671 = n6581 ;
  assign y3672 = 1'b0 ;
  assign y3673 = ~n6582 ;
  assign y3674 = ~1'b0 ;
  assign y3675 = ~1'b0 ;
  assign y3676 = n5324 ;
  assign y3677 = 1'b0 ;
  assign y3678 = 1'b0 ;
  assign y3679 = n6583 ;
  assign y3680 = ~1'b0 ;
  assign y3681 = ~n6587 ;
  assign y3682 = ~1'b0 ;
  assign y3683 = ~1'b0 ;
  assign y3684 = ~n6589 ;
  assign y3685 = ~n4760 ;
  assign y3686 = ~1'b0 ;
  assign y3687 = ~n1669 ;
  assign y3688 = ~n6590 ;
  assign y3689 = n6596 ;
  assign y3690 = n6598 ;
  assign y3691 = n6601 ;
  assign y3692 = n6605 ;
  assign y3693 = ~n6608 ;
  assign y3694 = n6612 ;
  assign y3695 = ~1'b0 ;
  assign y3696 = ~1'b0 ;
  assign y3697 = ~1'b0 ;
  assign y3698 = ~1'b0 ;
  assign y3699 = ~n6614 ;
  assign y3700 = ~1'b0 ;
  assign y3701 = ~1'b0 ;
  assign y3702 = ~n6618 ;
  assign y3703 = ~1'b0 ;
  assign y3704 = ~n6621 ;
  assign y3705 = n6623 ;
  assign y3706 = ~n6626 ;
  assign y3707 = n6629 ;
  assign y3708 = ~n6632 ;
  assign y3709 = ~1'b0 ;
  assign y3710 = ~n6636 ;
  assign y3711 = ~n6643 ;
  assign y3712 = ~1'b0 ;
  assign y3713 = n503 ;
  assign y3714 = n6644 ;
  assign y3715 = ~n6646 ;
  assign y3716 = ~n6649 ;
  assign y3717 = n6652 ;
  assign y3718 = ~n6654 ;
  assign y3719 = n6664 ;
  assign y3720 = ~1'b0 ;
  assign y3721 = ~1'b0 ;
  assign y3722 = ~n4600 ;
  assign y3723 = n6667 ;
  assign y3724 = n6670 ;
  assign y3725 = n6673 ;
  assign y3726 = ~n6675 ;
  assign y3727 = ~1'b0 ;
  assign y3728 = ~n6679 ;
  assign y3729 = ~n6685 ;
  assign y3730 = n1880 ;
  assign y3731 = n6687 ;
  assign y3732 = n6690 ;
  assign y3733 = n6692 ;
  assign y3734 = n6242 ;
  assign y3735 = ~n1181 ;
  assign y3736 = 1'b0 ;
  assign y3737 = ~1'b0 ;
  assign y3738 = ~n6698 ;
  assign y3739 = ~1'b0 ;
  assign y3740 = ~n6703 ;
  assign y3741 = ~n1637 ;
  assign y3742 = ~n6708 ;
  assign y3743 = ~n6710 ;
  assign y3744 = ~1'b0 ;
  assign y3745 = ~n6711 ;
  assign y3746 = ~n6719 ;
  assign y3747 = ~n6721 ;
  assign y3748 = ~n4578 ;
  assign y3749 = ~n2310 ;
  assign y3750 = ~n5885 ;
  assign y3751 = n6725 ;
  assign y3752 = ~1'b0 ;
  assign y3753 = ~1'b0 ;
  assign y3754 = n6726 ;
  assign y3755 = n6728 ;
  assign y3756 = ~1'b0 ;
  assign y3757 = ~n6730 ;
  assign y3758 = ~1'b0 ;
  assign y3759 = ~1'b0 ;
  assign y3760 = n6731 ;
  assign y3761 = n6732 ;
  assign y3762 = n6734 ;
  assign y3763 = ~1'b0 ;
  assign y3764 = ~n3667 ;
  assign y3765 = ~n6735 ;
  assign y3766 = ~1'b0 ;
  assign y3767 = ~n6736 ;
  assign y3768 = 1'b0 ;
  assign y3769 = n6738 ;
  assign y3770 = n6744 ;
  assign y3771 = n6746 ;
  assign y3772 = ~1'b0 ;
  assign y3773 = ~n6747 ;
  assign y3774 = ~n6753 ;
  assign y3775 = n6757 ;
  assign y3776 = ~1'b0 ;
  assign y3777 = ~1'b0 ;
  assign y3778 = ~n6764 ;
  assign y3779 = ~1'b0 ;
  assign y3780 = n6769 ;
  assign y3781 = n6773 ;
  assign y3782 = ~n6776 ;
  assign y3783 = ~n6780 ;
  assign y3784 = 1'b0 ;
  assign y3785 = ~n6782 ;
  assign y3786 = n6783 ;
  assign y3787 = n6786 ;
  assign y3788 = ~1'b0 ;
  assign y3789 = ~1'b0 ;
  assign y3790 = ~n6787 ;
  assign y3791 = ~1'b0 ;
  assign y3792 = ~n6788 ;
  assign y3793 = ~n6790 ;
  assign y3794 = n6792 ;
  assign y3795 = n6793 ;
  assign y3796 = ~n6794 ;
  assign y3797 = ~1'b0 ;
  assign y3798 = n6796 ;
  assign y3799 = ~1'b0 ;
  assign y3800 = ~n6799 ;
  assign y3801 = n6803 ;
  assign y3802 = ~1'b0 ;
  assign y3803 = ~n6811 ;
  assign y3804 = ~1'b0 ;
  assign y3805 = ~n1764 ;
  assign y3806 = n6813 ;
  assign y3807 = n6816 ;
  assign y3808 = ~1'b0 ;
  assign y3809 = ~1'b0 ;
  assign y3810 = ~1'b0 ;
  assign y3811 = ~1'b0 ;
  assign y3812 = ~1'b0 ;
  assign y3813 = ~1'b0 ;
  assign y3814 = n6531 ;
  assign y3815 = ~n6817 ;
  assign y3816 = ~1'b0 ;
  assign y3817 = ~1'b0 ;
  assign y3818 = n6822 ;
  assign y3819 = n1786 ;
  assign y3820 = ~1'b0 ;
  assign y3821 = n6825 ;
  assign y3822 = ~n6827 ;
  assign y3823 = ~n3824 ;
  assign y3824 = ~n6831 ;
  assign y3825 = ~n307 ;
  assign y3826 = ~n6832 ;
  assign y3827 = n6833 ;
  assign y3828 = ~1'b0 ;
  assign y3829 = ~n6835 ;
  assign y3830 = 1'b0 ;
  assign y3831 = n6451 ;
  assign y3832 = ~1'b0 ;
  assign y3833 = ~1'b0 ;
  assign y3834 = ~1'b0 ;
  assign y3835 = n6837 ;
  assign y3836 = ~1'b0 ;
  assign y3837 = n6840 ;
  assign y3838 = ~1'b0 ;
  assign y3839 = ~n6842 ;
  assign y3840 = ~1'b0 ;
  assign y3841 = ~n6846 ;
  assign y3842 = ~1'b0 ;
  assign y3843 = ~n6856 ;
  assign y3844 = ~1'b0 ;
  assign y3845 = ~n6859 ;
  assign y3846 = n2792 ;
  assign y3847 = n6860 ;
  assign y3848 = n6866 ;
  assign y3849 = 1'b0 ;
  assign y3850 = n6873 ;
  assign y3851 = ~1'b0 ;
  assign y3852 = ~n6874 ;
  assign y3853 = ~n6876 ;
  assign y3854 = ~1'b0 ;
  assign y3855 = ~n6877 ;
  assign y3856 = ~n6878 ;
  assign y3857 = n6881 ;
  assign y3858 = n6883 ;
  assign y3859 = ~n6891 ;
  assign y3860 = n6897 ;
  assign y3861 = n6901 ;
  assign y3862 = ~n6902 ;
  assign y3863 = n6904 ;
  assign y3864 = n6905 ;
  assign y3865 = ~n6908 ;
  assign y3866 = ~n6912 ;
  assign y3867 = ~1'b0 ;
  assign y3868 = ~n6917 ;
  assign y3869 = n6919 ;
  assign y3870 = n6922 ;
  assign y3871 = ~1'b0 ;
  assign y3872 = ~1'b0 ;
  assign y3873 = ~1'b0 ;
  assign y3874 = n6926 ;
  assign y3875 = ~1'b0 ;
  assign y3876 = ~1'b0 ;
  assign y3877 = ~1'b0 ;
  assign y3878 = ~1'b0 ;
  assign y3879 = n6928 ;
  assign y3880 = ~n6930 ;
  assign y3881 = ~1'b0 ;
  assign y3882 = ~1'b0 ;
  assign y3883 = n6933 ;
  assign y3884 = ~n6937 ;
  assign y3885 = ~1'b0 ;
  assign y3886 = ~1'b0 ;
  assign y3887 = ~n877 ;
  assign y3888 = ~1'b0 ;
  assign y3889 = 1'b0 ;
  assign y3890 = ~1'b0 ;
  assign y3891 = ~n6939 ;
  assign y3892 = ~1'b0 ;
  assign y3893 = ~n6940 ;
  assign y3894 = ~1'b0 ;
  assign y3895 = n6942 ;
  assign y3896 = ~1'b0 ;
  assign y3897 = ~1'b0 ;
  assign y3898 = n3369 ;
  assign y3899 = ~1'b0 ;
  assign y3900 = n6943 ;
  assign y3901 = ~1'b0 ;
  assign y3902 = n3763 ;
  assign y3903 = ~1'b0 ;
  assign y3904 = ~n6948 ;
  assign y3905 = n6954 ;
  assign y3906 = ~n4564 ;
  assign y3907 = ~n6957 ;
  assign y3908 = n6961 ;
  assign y3909 = n6962 ;
  assign y3910 = ~n6964 ;
  assign y3911 = ~n6969 ;
  assign y3912 = n6971 ;
  assign y3913 = ~n6972 ;
  assign y3914 = ~1'b0 ;
  assign y3915 = ~n6975 ;
  assign y3916 = ~1'b0 ;
  assign y3917 = n6980 ;
  assign y3918 = ~n6983 ;
  assign y3919 = n6984 ;
  assign y3920 = n6985 ;
  assign y3921 = ~1'b0 ;
  assign y3922 = n6987 ;
  assign y3923 = ~1'b0 ;
  assign y3924 = ~n5103 ;
  assign y3925 = ~1'b0 ;
  assign y3926 = ~n6988 ;
  assign y3927 = ~n6990 ;
  assign y3928 = ~1'b0 ;
  assign y3929 = ~n6994 ;
  assign y3930 = n6995 ;
  assign y3931 = ~n6998 ;
  assign y3932 = ~n7000 ;
  assign y3933 = n7001 ;
  assign y3934 = ~1'b0 ;
  assign y3935 = ~1'b0 ;
  assign y3936 = ~n7002 ;
  assign y3937 = ~1'b0 ;
  assign y3938 = ~n7006 ;
  assign y3939 = ~n7011 ;
  assign y3940 = ~1'b0 ;
  assign y3941 = n7015 ;
  assign y3942 = ~n7020 ;
  assign y3943 = n7031 ;
  assign y3944 = n7040 ;
  assign y3945 = ~1'b0 ;
  assign y3946 = ~1'b0 ;
  assign y3947 = n7044 ;
  assign y3948 = ~n7046 ;
  assign y3949 = ~n7047 ;
  assign y3950 = ~n7050 ;
  assign y3951 = n7054 ;
  assign y3952 = ~1'b0 ;
  assign y3953 = n7057 ;
  assign y3954 = n7060 ;
  assign y3955 = ~n7062 ;
  assign y3956 = n7069 ;
  assign y3957 = n7073 ;
  assign y3958 = ~1'b0 ;
  assign y3959 = ~n7078 ;
  assign y3960 = n7079 ;
  assign y3961 = ~n7082 ;
  assign y3962 = n7089 ;
  assign y3963 = n6760 ;
  assign y3964 = ~n7090 ;
  assign y3965 = ~1'b0 ;
  assign y3966 = ~n7094 ;
  assign y3967 = n7095 ;
  assign y3968 = ~n894 ;
  assign y3969 = ~1'b0 ;
  assign y3970 = n6915 ;
  assign y3971 = n7096 ;
  assign y3972 = ~n7100 ;
  assign y3973 = ~n7102 ;
  assign y3974 = n7104 ;
  assign y3975 = n7105 ;
  assign y3976 = ~n6578 ;
  assign y3977 = n7107 ;
  assign y3978 = n7109 ;
  assign y3979 = ~n7110 ;
  assign y3980 = ~1'b0 ;
  assign y3981 = n7111 ;
  assign y3982 = ~n7124 ;
  assign y3983 = ~n7125 ;
  assign y3984 = ~n2198 ;
  assign y3985 = ~1'b0 ;
  assign y3986 = n934 ;
  assign y3987 = ~n6321 ;
  assign y3988 = n7128 ;
  assign y3989 = ~n7129 ;
  assign y3990 = n7138 ;
  assign y3991 = ~n7139 ;
  assign y3992 = ~n7141 ;
  assign y3993 = ~1'b0 ;
  assign y3994 = ~1'b0 ;
  assign y3995 = ~n7142 ;
  assign y3996 = n7143 ;
  assign y3997 = ~n7155 ;
  assign y3998 = ~n7156 ;
  assign y3999 = ~1'b0 ;
  assign y4000 = ~n7157 ;
  assign y4001 = ~1'b0 ;
  assign y4002 = ~1'b0 ;
  assign y4003 = ~n7163 ;
  assign y4004 = n7166 ;
  assign y4005 = ~1'b0 ;
  assign y4006 = ~1'b0 ;
  assign y4007 = ~n7167 ;
  assign y4008 = ~n7168 ;
  assign y4009 = n7170 ;
  assign y4010 = ~n7172 ;
  assign y4011 = 1'b0 ;
  assign y4012 = n7176 ;
  assign y4013 = ~1'b0 ;
  assign y4014 = ~1'b0 ;
  assign y4015 = ~1'b0 ;
  assign y4016 = ~1'b0 ;
  assign y4017 = n7179 ;
  assign y4018 = ~n7180 ;
  assign y4019 = ~1'b0 ;
  assign y4020 = ~1'b0 ;
  assign y4021 = ~1'b0 ;
  assign y4022 = ~n7184 ;
  assign y4023 = 1'b0 ;
  assign y4024 = n7185 ;
  assign y4025 = ~n7186 ;
  assign y4026 = n7188 ;
  assign y4027 = n7190 ;
  assign y4028 = ~1'b0 ;
  assign y4029 = ~1'b0 ;
  assign y4030 = n7193 ;
  assign y4031 = ~n7194 ;
  assign y4032 = ~n7196 ;
  assign y4033 = ~n3615 ;
  assign y4034 = n7199 ;
  assign y4035 = ~n7202 ;
  assign y4036 = ~1'b0 ;
  assign y4037 = n7204 ;
  assign y4038 = 1'b0 ;
  assign y4039 = ~n7208 ;
  assign y4040 = ~1'b0 ;
  assign y4041 = ~1'b0 ;
  assign y4042 = ~1'b0 ;
  assign y4043 = ~n7211 ;
  assign y4044 = n7212 ;
  assign y4045 = x54 ;
  assign y4046 = ~n7213 ;
  assign y4047 = n7215 ;
  assign y4048 = n7216 ;
  assign y4049 = ~1'b0 ;
  assign y4050 = n7217 ;
  assign y4051 = ~1'b0 ;
  assign y4052 = 1'b0 ;
  assign y4053 = n7219 ;
  assign y4054 = ~n7221 ;
  assign y4055 = ~n7222 ;
  assign y4056 = ~n7226 ;
  assign y4057 = ~1'b0 ;
  assign y4058 = ~1'b0 ;
  assign y4059 = ~1'b0 ;
  assign y4060 = ~1'b0 ;
  assign y4061 = ~1'b0 ;
  assign y4062 = n7227 ;
  assign y4063 = ~n7229 ;
  assign y4064 = x107 ;
  assign y4065 = ~1'b0 ;
  assign y4066 = ~1'b0 ;
  assign y4067 = n7230 ;
  assign y4068 = ~1'b0 ;
  assign y4069 = ~n7233 ;
  assign y4070 = ~n7236 ;
  assign y4071 = n7239 ;
  assign y4072 = n7244 ;
  assign y4073 = ~1'b0 ;
  assign y4074 = ~n7245 ;
  assign y4075 = n7246 ;
  assign y4076 = ~n7249 ;
  assign y4077 = ~n7250 ;
  assign y4078 = ~n7253 ;
  assign y4079 = ~n7257 ;
  assign y4080 = n7262 ;
  assign y4081 = ~n5552 ;
  assign y4082 = n7263 ;
  assign y4083 = ~1'b0 ;
  assign y4084 = ~1'b0 ;
  assign y4085 = ~n7265 ;
  assign y4086 = ~1'b0 ;
  assign y4087 = n7266 ;
  assign y4088 = n7269 ;
  assign y4089 = ~1'b0 ;
  assign y4090 = ~n7271 ;
  assign y4091 = ~n7273 ;
  assign y4092 = n7275 ;
  assign y4093 = ~1'b0 ;
  assign y4094 = ~n7276 ;
  assign y4095 = n7277 ;
  assign y4096 = ~n7278 ;
  assign y4097 = n7280 ;
  assign y4098 = ~1'b0 ;
  assign y4099 = ~n7283 ;
  assign y4100 = n7284 ;
  assign y4101 = ~1'b0 ;
  assign y4102 = 1'b0 ;
  assign y4103 = 1'b0 ;
  assign y4104 = ~n7285 ;
  assign y4105 = n7287 ;
  assign y4106 = 1'b0 ;
  assign y4107 = ~1'b0 ;
  assign y4108 = ~n7293 ;
  assign y4109 = ~1'b0 ;
  assign y4110 = n7296 ;
  assign y4111 = n7299 ;
  assign y4112 = ~1'b0 ;
  assign y4113 = ~n7300 ;
  assign y4114 = ~n7302 ;
  assign y4115 = ~n7303 ;
  assign y4116 = n7305 ;
  assign y4117 = ~1'b0 ;
  assign y4118 = ~1'b0 ;
  assign y4119 = n7306 ;
  assign y4120 = ~n1762 ;
  assign y4121 = ~1'b0 ;
  assign y4122 = ~n7307 ;
  assign y4123 = ~1'b0 ;
  assign y4124 = ~1'b0 ;
  assign y4125 = ~1'b0 ;
  assign y4126 = n7308 ;
  assign y4127 = ~1'b0 ;
  assign y4128 = ~n2885 ;
  assign y4129 = ~1'b0 ;
  assign y4130 = ~1'b0 ;
  assign y4131 = ~n7310 ;
  assign y4132 = ~1'b0 ;
  assign y4133 = ~n7334 ;
  assign y4134 = ~1'b0 ;
  assign y4135 = ~1'b0 ;
  assign y4136 = n7337 ;
  assign y4137 = ~n7339 ;
  assign y4138 = ~n7343 ;
  assign y4139 = ~1'b0 ;
  assign y4140 = ~1'b0 ;
  assign y4141 = ~n7345 ;
  assign y4142 = ~n7348 ;
  assign y4143 = ~1'b0 ;
  assign y4144 = ~1'b0 ;
  assign y4145 = n7350 ;
  assign y4146 = n7358 ;
  assign y4147 = 1'b0 ;
  assign y4148 = ~1'b0 ;
  assign y4149 = n7360 ;
  assign y4150 = n7361 ;
  assign y4151 = ~n7362 ;
  assign y4152 = n7367 ;
  assign y4153 = ~1'b0 ;
  assign y4154 = ~1'b0 ;
  assign y4155 = ~n7368 ;
  assign y4156 = n7369 ;
  assign y4157 = n7370 ;
  assign y4158 = ~n7371 ;
  assign y4159 = ~1'b0 ;
  assign y4160 = ~1'b0 ;
  assign y4161 = ~1'b0 ;
  assign y4162 = ~n7372 ;
  assign y4163 = ~n2944 ;
  assign y4164 = ~n7375 ;
  assign y4165 = 1'b0 ;
  assign y4166 = ~n7376 ;
  assign y4167 = ~1'b0 ;
  assign y4168 = ~1'b0 ;
  assign y4169 = ~1'b0 ;
  assign y4170 = ~1'b0 ;
  assign y4171 = ~1'b0 ;
  assign y4172 = ~1'b0 ;
  assign y4173 = ~1'b0 ;
  assign y4174 = n6371 ;
  assign y4175 = ~1'b0 ;
  assign y4176 = ~1'b0 ;
  assign y4177 = ~1'b0 ;
  assign y4178 = ~n5748 ;
  assign y4179 = ~1'b0 ;
  assign y4180 = n7378 ;
  assign y4181 = n7381 ;
  assign y4182 = ~n7383 ;
  assign y4183 = n7389 ;
  assign y4184 = ~1'b0 ;
  assign y4185 = ~n7397 ;
  assign y4186 = n7404 ;
  assign y4187 = n7408 ;
  assign y4188 = ~1'b0 ;
  assign y4189 = ~1'b0 ;
  assign y4190 = ~1'b0 ;
  assign y4191 = ~n7416 ;
  assign y4192 = ~1'b0 ;
  assign y4193 = n5501 ;
  assign y4194 = ~n7418 ;
  assign y4195 = ~n7421 ;
  assign y4196 = ~n7423 ;
  assign y4197 = ~1'b0 ;
  assign y4198 = ~n5720 ;
  assign y4199 = ~1'b0 ;
  assign y4200 = ~n7424 ;
  assign y4201 = ~n7432 ;
  assign y4202 = ~1'b0 ;
  assign y4203 = ~n3415 ;
  assign y4204 = ~n7436 ;
  assign y4205 = ~n7440 ;
  assign y4206 = ~1'b0 ;
  assign y4207 = n7441 ;
  assign y4208 = ~n7445 ;
  assign y4209 = ~1'b0 ;
  assign y4210 = ~1'b0 ;
  assign y4211 = n7446 ;
  assign y4212 = ~n7454 ;
  assign y4213 = n7456 ;
  assign y4214 = ~n7457 ;
  assign y4215 = n7459 ;
  assign y4216 = ~1'b0 ;
  assign y4217 = ~1'b0 ;
  assign y4218 = ~1'b0 ;
  assign y4219 = ~1'b0 ;
  assign y4220 = ~1'b0 ;
  assign y4221 = ~n7467 ;
  assign y4222 = n7468 ;
  assign y4223 = ~n7469 ;
  assign y4224 = ~1'b0 ;
  assign y4225 = ~1'b0 ;
  assign y4226 = ~n390 ;
  assign y4227 = ~1'b0 ;
  assign y4228 = n7474 ;
  assign y4229 = ~1'b0 ;
  assign y4230 = n4571 ;
  assign y4231 = ~1'b0 ;
  assign y4232 = n7475 ;
  assign y4233 = ~1'b0 ;
  assign y4234 = n3251 ;
  assign y4235 = ~n7476 ;
  assign y4236 = ~1'b0 ;
  assign y4237 = ~1'b0 ;
  assign y4238 = ~n7478 ;
  assign y4239 = n7479 ;
  assign y4240 = ~1'b0 ;
  assign y4241 = ~n7487 ;
  assign y4242 = ~1'b0 ;
  assign y4243 = ~n3454 ;
  assign y4244 = n7488 ;
  assign y4245 = ~n7490 ;
  assign y4246 = n7492 ;
  assign y4247 = ~1'b0 ;
  assign y4248 = n7495 ;
  assign y4249 = ~n7497 ;
  assign y4250 = ~n7505 ;
  assign y4251 = ~1'b0 ;
  assign y4252 = n7506 ;
  assign y4253 = n7512 ;
  assign y4254 = ~1'b0 ;
  assign y4255 = n7519 ;
  assign y4256 = 1'b0 ;
  assign y4257 = n7522 ;
  assign y4258 = ~n7523 ;
  assign y4259 = n985 ;
  assign y4260 = ~n7524 ;
  assign y4261 = n7525 ;
  assign y4262 = n7527 ;
  assign y4263 = ~n7529 ;
  assign y4264 = ~1'b0 ;
  assign y4265 = ~1'b0 ;
  assign y4266 = n7531 ;
  assign y4267 = ~n7535 ;
  assign y4268 = ~1'b0 ;
  assign y4269 = n7536 ;
  assign y4270 = ~n7543 ;
  assign y4271 = ~1'b0 ;
  assign y4272 = n7544 ;
  assign y4273 = n7545 ;
  assign y4274 = ~1'b0 ;
  assign y4275 = n7547 ;
  assign y4276 = n7549 ;
  assign y4277 = n7550 ;
  assign y4278 = n7556 ;
  assign y4279 = ~n7558 ;
  assign y4280 = n7567 ;
  assign y4281 = n7574 ;
  assign y4282 = ~1'b0 ;
  assign y4283 = ~n7576 ;
  assign y4284 = ~n7584 ;
  assign y4285 = n7592 ;
  assign y4286 = ~n6829 ;
  assign y4287 = ~1'b0 ;
  assign y4288 = n825 ;
  assign y4289 = n7593 ;
  assign y4290 = ~1'b0 ;
  assign y4291 = n7597 ;
  assign y4292 = ~1'b0 ;
  assign y4293 = n7598 ;
  assign y4294 = ~n7600 ;
  assign y4295 = ~n7601 ;
  assign y4296 = ~n6051 ;
  assign y4297 = ~1'b0 ;
  assign y4298 = ~1'b0 ;
  assign y4299 = ~n7602 ;
  assign y4300 = n7608 ;
  assign y4301 = n7612 ;
  assign y4302 = ~1'b0 ;
  assign y4303 = n1910 ;
  assign y4304 = n7613 ;
  assign y4305 = ~n7616 ;
  assign y4306 = ~n7622 ;
  assign y4307 = n7626 ;
  assign y4308 = n7629 ;
  assign y4309 = ~1'b0 ;
  assign y4310 = n7633 ;
  assign y4311 = ~1'b0 ;
  assign y4312 = ~n7637 ;
  assign y4313 = ~1'b0 ;
  assign y4314 = ~n4876 ;
  assign y4315 = ~n7639 ;
  assign y4316 = ~n7640 ;
  assign y4317 = 1'b0 ;
  assign y4318 = ~1'b0 ;
  assign y4319 = ~n7641 ;
  assign y4320 = 1'b0 ;
  assign y4321 = ~n6890 ;
  assign y4322 = ~1'b0 ;
  assign y4323 = n2315 ;
  assign y4324 = ~n7643 ;
  assign y4325 = ~n7644 ;
  assign y4326 = ~n7646 ;
  assign y4327 = ~1'b0 ;
  assign y4328 = n7648 ;
  assign y4329 = n5434 ;
  assign y4330 = 1'b0 ;
  assign y4331 = ~1'b0 ;
  assign y4332 = n7652 ;
  assign y4333 = ~n7653 ;
  assign y4334 = ~n7657 ;
  assign y4335 = n7658 ;
  assign y4336 = ~1'b0 ;
  assign y4337 = ~n7659 ;
  assign y4338 = ~n7660 ;
  assign y4339 = ~n7662 ;
  assign y4340 = n7666 ;
  assign y4341 = ~n7668 ;
  assign y4342 = ~1'b0 ;
  assign y4343 = ~n3066 ;
  assign y4344 = ~1'b0 ;
  assign y4345 = ~n7670 ;
  assign y4346 = n7675 ;
  assign y4347 = ~n7678 ;
  assign y4348 = ~1'b0 ;
  assign y4349 = n7679 ;
  assign y4350 = n7686 ;
  assign y4351 = ~1'b0 ;
  assign y4352 = ~n7692 ;
  assign y4353 = n7695 ;
  assign y4354 = ~1'b0 ;
  assign y4355 = ~n7697 ;
  assign y4356 = ~1'b0 ;
  assign y4357 = ~n7703 ;
  assign y4358 = n7704 ;
  assign y4359 = ~1'b0 ;
  assign y4360 = n7705 ;
  assign y4361 = ~1'b0 ;
  assign y4362 = ~1'b0 ;
  assign y4363 = 1'b0 ;
  assign y4364 = ~1'b0 ;
  assign y4365 = ~n7706 ;
  assign y4366 = ~1'b0 ;
  assign y4367 = n7707 ;
  assign y4368 = ~1'b0 ;
  assign y4369 = ~n7708 ;
  assign y4370 = n7709 ;
  assign y4371 = ~1'b0 ;
  assign y4372 = n1899 ;
  assign y4373 = ~1'b0 ;
  assign y4374 = n7712 ;
  assign y4375 = n7716 ;
  assign y4376 = n7719 ;
  assign y4377 = ~1'b0 ;
  assign y4378 = 1'b0 ;
  assign y4379 = n7721 ;
  assign y4380 = 1'b0 ;
  assign y4381 = n7723 ;
  assign y4382 = n5223 ;
  assign y4383 = ~1'b0 ;
  assign y4384 = ~n7724 ;
  assign y4385 = ~n5152 ;
  assign y4386 = n7725 ;
  assign y4387 = ~n7727 ;
  assign y4388 = n7729 ;
  assign y4389 = n7731 ;
  assign y4390 = ~n7732 ;
  assign y4391 = n7733 ;
  assign y4392 = ~n7740 ;
  assign y4393 = ~n3544 ;
  assign y4394 = 1'b0 ;
  assign y4395 = n7741 ;
  assign y4396 = ~n7744 ;
  assign y4397 = ~n7749 ;
  assign y4398 = n7750 ;
  assign y4399 = n7753 ;
  assign y4400 = n7755 ;
  assign y4401 = n7758 ;
  assign y4402 = n7762 ;
  assign y4403 = ~n7763 ;
  assign y4404 = ~n7764 ;
  assign y4405 = ~1'b0 ;
  assign y4406 = n7766 ;
  assign y4407 = n5120 ;
  assign y4408 = ~n7767 ;
  assign y4409 = n7769 ;
  assign y4410 = n7770 ;
  assign y4411 = ~n7773 ;
  assign y4412 = n7777 ;
  assign y4413 = ~1'b0 ;
  assign y4414 = ~1'b0 ;
  assign y4415 = ~1'b0 ;
  assign y4416 = n7780 ;
  assign y4417 = n7784 ;
  assign y4418 = n7788 ;
  assign y4419 = n7791 ;
  assign y4420 = ~n7792 ;
  assign y4421 = n7793 ;
  assign y4422 = n7794 ;
  assign y4423 = n1880 ;
  assign y4424 = ~n7795 ;
  assign y4425 = ~n7796 ;
  assign y4426 = n7801 ;
  assign y4427 = ~n5293 ;
  assign y4428 = n7803 ;
  assign y4429 = ~1'b0 ;
  assign y4430 = ~n7809 ;
  assign y4431 = ~n7810 ;
  assign y4432 = ~n7812 ;
  assign y4433 = n7815 ;
  assign y4434 = ~1'b0 ;
  assign y4435 = ~n7816 ;
  assign y4436 = ~n1548 ;
  assign y4437 = n7819 ;
  assign y4438 = ~n7834 ;
  assign y4439 = ~n2897 ;
  assign y4440 = ~n7835 ;
  assign y4441 = ~n7836 ;
  assign y4442 = n3445 ;
  assign y4443 = n6901 ;
  assign y4444 = ~1'b0 ;
  assign y4445 = ~1'b0 ;
  assign y4446 = n7845 ;
  assign y4447 = ~n7851 ;
  assign y4448 = n2043 ;
  assign y4449 = n7853 ;
  assign y4450 = ~1'b0 ;
  assign y4451 = n7855 ;
  assign y4452 = ~n7857 ;
  assign y4453 = n7864 ;
  assign y4454 = ~1'b0 ;
  assign y4455 = n7867 ;
  assign y4456 = ~1'b0 ;
  assign y4457 = n7868 ;
  assign y4458 = ~n7873 ;
  assign y4459 = ~n7874 ;
  assign y4460 = n7879 ;
  assign y4461 = ~n7886 ;
  assign y4462 = n7888 ;
  assign y4463 = ~1'b0 ;
  assign y4464 = ~1'b0 ;
  assign y4465 = ~n7889 ;
  assign y4466 = ~n7892 ;
  assign y4467 = ~n7896 ;
  assign y4468 = ~n7898 ;
  assign y4469 = ~1'b0 ;
  assign y4470 = n7900 ;
  assign y4471 = n7902 ;
  assign y4472 = n7904 ;
  assign y4473 = ~1'b0 ;
  assign y4474 = ~1'b0 ;
  assign y4475 = ~n7905 ;
  assign y4476 = ~n7913 ;
  assign y4477 = ~n5652 ;
  assign y4478 = ~n7915 ;
  assign y4479 = ~1'b0 ;
  assign y4480 = ~n7922 ;
  assign y4481 = ~n7924 ;
  assign y4482 = ~1'b0 ;
  assign y4483 = n2505 ;
  assign y4484 = ~1'b0 ;
  assign y4485 = n7925 ;
  assign y4486 = ~n7926 ;
  assign y4487 = ~n7927 ;
  assign y4488 = ~n7929 ;
  assign y4489 = n7930 ;
  assign y4490 = ~n7932 ;
  assign y4491 = ~n7933 ;
  assign y4492 = ~1'b0 ;
  assign y4493 = ~n7934 ;
  assign y4494 = ~n5239 ;
  assign y4495 = ~1'b0 ;
  assign y4496 = ~1'b0 ;
  assign y4497 = ~1'b0 ;
  assign y4498 = ~n7935 ;
  assign y4499 = n7936 ;
  assign y4500 = ~n6495 ;
  assign y4501 = ~n7938 ;
  assign y4502 = ~n7940 ;
  assign y4503 = n7941 ;
  assign y4504 = n7943 ;
  assign y4505 = ~n7944 ;
  assign y4506 = n7948 ;
  assign y4507 = n7951 ;
  assign y4508 = ~1'b0 ;
  assign y4509 = ~n7952 ;
  assign y4510 = n7956 ;
  assign y4511 = ~1'b0 ;
  assign y4512 = n7957 ;
  assign y4513 = n7961 ;
  assign y4514 = ~1'b0 ;
  assign y4515 = ~1'b0 ;
  assign y4516 = ~n7963 ;
  assign y4517 = ~1'b0 ;
  assign y4518 = ~1'b0 ;
  assign y4519 = ~n7965 ;
  assign y4520 = ~1'b0 ;
  assign y4521 = ~1'b0 ;
  assign y4522 = ~1'b0 ;
  assign y4523 = n7967 ;
  assign y4524 = n7968 ;
  assign y4525 = ~n7970 ;
  assign y4526 = ~n5222 ;
  assign y4527 = n7971 ;
  assign y4528 = n7974 ;
  assign y4529 = ~n7976 ;
  assign y4530 = ~1'b0 ;
  assign y4531 = ~n7978 ;
  assign y4532 = n7986 ;
  assign y4533 = ~1'b0 ;
  assign y4534 = ~1'b0 ;
  assign y4535 = n7987 ;
  assign y4536 = n5018 ;
  assign y4537 = n7991 ;
  assign y4538 = ~1'b0 ;
  assign y4539 = ~1'b0 ;
  assign y4540 = ~1'b0 ;
  assign y4541 = n7995 ;
  assign y4542 = ~n7996 ;
  assign y4543 = n7801 ;
  assign y4544 = ~n7999 ;
  assign y4545 = ~n8007 ;
  assign y4546 = ~1'b0 ;
  assign y4547 = ~1'b0 ;
  assign y4548 = 1'b0 ;
  assign y4549 = ~n8008 ;
  assign y4550 = ~1'b0 ;
  assign y4551 = ~n8011 ;
  assign y4552 = n8014 ;
  assign y4553 = n8019 ;
  assign y4554 = ~1'b0 ;
  assign y4555 = n8020 ;
  assign y4556 = n8024 ;
  assign y4557 = n8026 ;
  assign y4558 = ~1'b0 ;
  assign y4559 = ~1'b0 ;
  assign y4560 = ~n8029 ;
  assign y4561 = ~1'b0 ;
  assign y4562 = ~n8032 ;
  assign y4563 = ~n8033 ;
  assign y4564 = n8034 ;
  assign y4565 = ~n8037 ;
  assign y4566 = n8040 ;
  assign y4567 = n8043 ;
  assign y4568 = n6326 ;
  assign y4569 = n8046 ;
  assign y4570 = n8048 ;
  assign y4571 = ~1'b0 ;
  assign y4572 = ~1'b0 ;
  assign y4573 = n8050 ;
  assign y4574 = n3672 ;
  assign y4575 = n8054 ;
  assign y4576 = n8055 ;
  assign y4577 = ~1'b0 ;
  assign y4578 = ~n8056 ;
  assign y4579 = n8064 ;
  assign y4580 = n8065 ;
  assign y4581 = ~n8069 ;
  assign y4582 = n2818 ;
  assign y4583 = ~1'b0 ;
  assign y4584 = ~n8077 ;
  assign y4585 = ~n8078 ;
  assign y4586 = ~n8080 ;
  assign y4587 = n8084 ;
  assign y4588 = ~n8087 ;
  assign y4589 = 1'b0 ;
  assign y4590 = ~n8088 ;
  assign y4591 = ~1'b0 ;
  assign y4592 = ~1'b0 ;
  assign y4593 = ~1'b0 ;
  assign y4594 = n781 ;
  assign y4595 = n8090 ;
  assign y4596 = n8092 ;
  assign y4597 = n8096 ;
  assign y4598 = ~1'b0 ;
  assign y4599 = ~n8098 ;
  assign y4600 = ~1'b0 ;
  assign y4601 = ~n8102 ;
  assign y4602 = n4274 ;
  assign y4603 = ~1'b0 ;
  assign y4604 = ~1'b0 ;
  assign y4605 = ~1'b0 ;
  assign y4606 = ~1'b0 ;
  assign y4607 = ~1'b0 ;
  assign y4608 = ~n8107 ;
  assign y4609 = ~n8110 ;
  assign y4610 = n8112 ;
  assign y4611 = ~1'b0 ;
  assign y4612 = ~1'b0 ;
  assign y4613 = 1'b0 ;
  assign y4614 = ~n8115 ;
  assign y4615 = n8116 ;
  assign y4616 = ~n8117 ;
  assign y4617 = ~n8118 ;
  assign y4618 = ~n6992 ;
  assign y4619 = n8120 ;
  assign y4620 = ~n1601 ;
  assign y4621 = ~1'b0 ;
  assign y4622 = ~n8121 ;
  assign y4623 = 1'b0 ;
  assign y4624 = n8124 ;
  assign y4625 = ~n8125 ;
  assign y4626 = ~1'b0 ;
  assign y4627 = ~n2981 ;
  assign y4628 = n8126 ;
  assign y4629 = n8131 ;
  assign y4630 = n8133 ;
  assign y4631 = ~1'b0 ;
  assign y4632 = ~n8136 ;
  assign y4633 = ~1'b0 ;
  assign y4634 = n1772 ;
  assign y4635 = n8138 ;
  assign y4636 = n8144 ;
  assign y4637 = n8146 ;
  assign y4638 = ~1'b0 ;
  assign y4639 = n8154 ;
  assign y4640 = n1880 ;
  assign y4641 = ~n8155 ;
  assign y4642 = ~n8160 ;
  assign y4643 = ~n8163 ;
  assign y4644 = n8164 ;
  assign y4645 = ~1'b0 ;
  assign y4646 = n8169 ;
  assign y4647 = ~n8170 ;
  assign y4648 = n8173 ;
  assign y4649 = n8175 ;
  assign y4650 = n8176 ;
  assign y4651 = ~n8178 ;
  assign y4652 = ~n8182 ;
  assign y4653 = ~n8183 ;
  assign y4654 = ~n8185 ;
  assign y4655 = ~n8186 ;
  assign y4656 = ~1'b0 ;
  assign y4657 = n8190 ;
  assign y4658 = ~1'b0 ;
  assign y4659 = n6874 ;
  assign y4660 = 1'b0 ;
  assign y4661 = 1'b0 ;
  assign y4662 = ~n8192 ;
  assign y4663 = ~1'b0 ;
  assign y4664 = n8194 ;
  assign y4665 = ~n3829 ;
  assign y4666 = 1'b0 ;
  assign y4667 = ~1'b0 ;
  assign y4668 = ~1'b0 ;
  assign y4669 = n8198 ;
  assign y4670 = n8199 ;
  assign y4671 = ~1'b0 ;
  assign y4672 = n3120 ;
  assign y4673 = n8200 ;
  assign y4674 = ~1'b0 ;
  assign y4675 = ~1'b0 ;
  assign y4676 = ~n8203 ;
  assign y4677 = ~1'b0 ;
  assign y4678 = ~n8204 ;
  assign y4679 = x11 ;
  assign y4680 = ~1'b0 ;
  assign y4681 = n8209 ;
  assign y4682 = ~n8216 ;
  assign y4683 = ~1'b0 ;
  assign y4684 = ~1'b0 ;
  assign y4685 = n8218 ;
  assign y4686 = n1655 ;
  assign y4687 = ~x12 ;
  assign y4688 = n8219 ;
  assign y4689 = ~1'b0 ;
  assign y4690 = ~1'b0 ;
  assign y4691 = ~1'b0 ;
  assign y4692 = ~n2155 ;
  assign y4693 = n8224 ;
  assign y4694 = ~n8225 ;
  assign y4695 = 1'b0 ;
  assign y4696 = n8230 ;
  assign y4697 = ~1'b0 ;
  assign y4698 = ~1'b0 ;
  assign y4699 = ~1'b0 ;
  assign y4700 = n8232 ;
  assign y4701 = n4598 ;
  assign y4702 = ~n8237 ;
  assign y4703 = ~n8246 ;
  assign y4704 = n8247 ;
  assign y4705 = ~1'b0 ;
  assign y4706 = ~1'b0 ;
  assign y4707 = n8250 ;
  assign y4708 = ~1'b0 ;
  assign y4709 = ~1'b0 ;
  assign y4710 = ~1'b0 ;
  assign y4711 = ~n7364 ;
  assign y4712 = ~n8251 ;
  assign y4713 = ~n8253 ;
  assign y4714 = n8254 ;
  assign y4715 = ~n8259 ;
  assign y4716 = 1'b0 ;
  assign y4717 = ~n8261 ;
  assign y4718 = ~1'b0 ;
  assign y4719 = ~1'b0 ;
  assign y4720 = n8262 ;
  assign y4721 = n8265 ;
  assign y4722 = ~n7543 ;
  assign y4723 = ~1'b0 ;
  assign y4724 = ~n5089 ;
  assign y4725 = ~1'b0 ;
  assign y4726 = ~n8268 ;
  assign y4727 = n8270 ;
  assign y4728 = ~n8274 ;
  assign y4729 = ~n8280 ;
  assign y4730 = n8282 ;
  assign y4731 = ~n1932 ;
  assign y4732 = ~1'b0 ;
  assign y4733 = ~1'b0 ;
  assign y4734 = n8284 ;
  assign y4735 = ~n8285 ;
  assign y4736 = n3144 ;
  assign y4737 = n8288 ;
  assign y4738 = n8289 ;
  assign y4739 = ~1'b0 ;
  assign y4740 = ~1'b0 ;
  assign y4741 = n8292 ;
  assign y4742 = n8295 ;
  assign y4743 = ~n8300 ;
  assign y4744 = n8304 ;
  assign y4745 = ~n8306 ;
  assign y4746 = n8307 ;
  assign y4747 = ~n8309 ;
  assign y4748 = ~1'b0 ;
  assign y4749 = ~1'b0 ;
  assign y4750 = n8310 ;
  assign y4751 = n8314 ;
  assign y4752 = ~1'b0 ;
  assign y4753 = ~n8315 ;
  assign y4754 = 1'b0 ;
  assign y4755 = ~n8318 ;
  assign y4756 = ~1'b0 ;
  assign y4757 = n3947 ;
  assign y4758 = n1554 ;
  assign y4759 = n8320 ;
  assign y4760 = ~1'b0 ;
  assign y4761 = ~1'b0 ;
  assign y4762 = ~n8327 ;
  assign y4763 = ~1'b0 ;
  assign y4764 = n3195 ;
  assign y4765 = n8330 ;
  assign y4766 = ~1'b0 ;
  assign y4767 = ~n8332 ;
  assign y4768 = n8333 ;
  assign y4769 = ~n8338 ;
  assign y4770 = n8342 ;
  assign y4771 = ~n8343 ;
  assign y4772 = ~n8345 ;
  assign y4773 = n8347 ;
  assign y4774 = n8350 ;
  assign y4775 = ~n1256 ;
  assign y4776 = n8358 ;
  assign y4777 = ~n8360 ;
  assign y4778 = n8362 ;
  assign y4779 = n8363 ;
  assign y4780 = ~1'b0 ;
  assign y4781 = n8368 ;
  assign y4782 = n8369 ;
  assign y4783 = ~n8370 ;
  assign y4784 = ~1'b0 ;
  assign y4785 = ~1'b0 ;
  assign y4786 = ~1'b0 ;
  assign y4787 = ~1'b0 ;
  assign y4788 = ~n8371 ;
  assign y4789 = 1'b0 ;
  assign y4790 = ~1'b0 ;
  assign y4791 = ~x55 ;
  assign y4792 = n8374 ;
  assign y4793 = ~n8376 ;
  assign y4794 = ~1'b0 ;
  assign y4795 = n8377 ;
  assign y4796 = ~n8379 ;
  assign y4797 = 1'b0 ;
  assign y4798 = ~n8385 ;
  assign y4799 = n8387 ;
  assign y4800 = ~n7694 ;
  assign y4801 = ~1'b0 ;
  assign y4802 = ~1'b0 ;
  assign y4803 = ~1'b0 ;
  assign y4804 = ~n8389 ;
  assign y4805 = n7726 ;
  assign y4806 = n8390 ;
  assign y4807 = ~n8392 ;
  assign y4808 = ~n1356 ;
  assign y4809 = ~1'b0 ;
  assign y4810 = ~1'b0 ;
  assign y4811 = ~n8393 ;
  assign y4812 = ~n8395 ;
  assign y4813 = n8397 ;
  assign y4814 = n8398 ;
  assign y4815 = 1'b0 ;
  assign y4816 = ~1'b0 ;
  assign y4817 = ~n8404 ;
  assign y4818 = ~n8409 ;
  assign y4819 = ~n8411 ;
  assign y4820 = ~1'b0 ;
  assign y4821 = ~1'b0 ;
  assign y4822 = n8413 ;
  assign y4823 = ~n8414 ;
  assign y4824 = ~1'b0 ;
  assign y4825 = n8418 ;
  assign y4826 = n8419 ;
  assign y4827 = ~n8423 ;
  assign y4828 = n4895 ;
  assign y4829 = n8429 ;
  assign y4830 = ~n558 ;
  assign y4831 = n8430 ;
  assign y4832 = n8431 ;
  assign y4833 = ~1'b0 ;
  assign y4834 = ~n8433 ;
  assign y4835 = ~1'b0 ;
  assign y4836 = ~1'b0 ;
  assign y4837 = n8436 ;
  assign y4838 = ~1'b0 ;
  assign y4839 = ~n8437 ;
  assign y4840 = ~n8439 ;
  assign y4841 = ~1'b0 ;
  assign y4842 = x62 ;
  assign y4843 = ~n8440 ;
  assign y4844 = n8441 ;
  assign y4845 = n8445 ;
  assign y4846 = ~n8446 ;
  assign y4847 = n8447 ;
  assign y4848 = ~1'b0 ;
  assign y4849 = ~n8452 ;
  assign y4850 = n8454 ;
  assign y4851 = ~n8456 ;
  assign y4852 = ~1'b0 ;
  assign y4853 = ~1'b0 ;
  assign y4854 = x85 ;
  assign y4855 = n8458 ;
  assign y4856 = ~n8461 ;
  assign y4857 = ~n8462 ;
  assign y4858 = ~n1480 ;
  assign y4859 = ~n8463 ;
  assign y4860 = n8464 ;
  assign y4861 = ~n8472 ;
  assign y4862 = ~n544 ;
  assign y4863 = ~n8474 ;
  assign y4864 = 1'b0 ;
  assign y4865 = n8476 ;
  assign y4866 = ~n8486 ;
  assign y4867 = ~n8490 ;
  assign y4868 = n8491 ;
  assign y4869 = ~1'b0 ;
  assign y4870 = ~1'b0 ;
  assign y4871 = ~n8492 ;
  assign y4872 = ~n3900 ;
  assign y4873 = ~1'b0 ;
  assign y4874 = ~1'b0 ;
  assign y4875 = ~n2056 ;
  assign y4876 = ~1'b0 ;
  assign y4877 = ~n8494 ;
  assign y4878 = n8504 ;
  assign y4879 = n8506 ;
  assign y4880 = ~n8510 ;
  assign y4881 = ~n8511 ;
  assign y4882 = ~1'b0 ;
  assign y4883 = ~n8513 ;
  assign y4884 = ~n868 ;
  assign y4885 = ~1'b0 ;
  assign y4886 = ~1'b0 ;
  assign y4887 = n8517 ;
  assign y4888 = ~1'b0 ;
  assign y4889 = n8518 ;
  assign y4890 = ~1'b0 ;
  assign y4891 = ~n8519 ;
  assign y4892 = ~n8520 ;
  assign y4893 = ~1'b0 ;
  assign y4894 = ~n8522 ;
  assign y4895 = ~n983 ;
  assign y4896 = ~1'b0 ;
  assign y4897 = ~1'b0 ;
  assign y4898 = n3019 ;
  assign y4899 = n8524 ;
  assign y4900 = n8526 ;
  assign y4901 = ~1'b0 ;
  assign y4902 = n8530 ;
  assign y4903 = n8533 ;
  assign y4904 = ~n8535 ;
  assign y4905 = n8536 ;
  assign y4906 = n8564 ;
  assign y4907 = ~n8567 ;
  assign y4908 = n8570 ;
  assign y4909 = ~1'b0 ;
  assign y4910 = n8577 ;
  assign y4911 = ~1'b0 ;
  assign y4912 = n4224 ;
  assign y4913 = n8578 ;
  assign y4914 = ~n2811 ;
  assign y4915 = ~1'b0 ;
  assign y4916 = ~n8580 ;
  assign y4917 = n8581 ;
  assign y4918 = n8582 ;
  assign y4919 = n8584 ;
  assign y4920 = n8585 ;
  assign y4921 = ~1'b0 ;
  assign y4922 = n8587 ;
  assign y4923 = ~n8592 ;
  assign y4924 = ~n8594 ;
  assign y4925 = n891 ;
  assign y4926 = n2436 ;
  assign y4927 = 1'b0 ;
  assign y4928 = ~1'b0 ;
  assign y4929 = ~n8595 ;
  assign y4930 = ~n8596 ;
  assign y4931 = ~1'b0 ;
  assign y4932 = n8597 ;
  assign y4933 = n8599 ;
  assign y4934 = ~1'b0 ;
  assign y4935 = ~1'b0 ;
  assign y4936 = n8604 ;
  assign y4937 = ~n8605 ;
  assign y4938 = ~1'b0 ;
  assign y4939 = ~n8610 ;
  assign y4940 = ~n8613 ;
  assign y4941 = n8623 ;
  assign y4942 = n8624 ;
  assign y4943 = 1'b0 ;
  assign y4944 = n8628 ;
  assign y4945 = ~1'b0 ;
  assign y4946 = n8633 ;
  assign y4947 = 1'b0 ;
  assign y4948 = ~1'b0 ;
  assign y4949 = ~1'b0 ;
  assign y4950 = ~1'b0 ;
  assign y4951 = ~n8635 ;
  assign y4952 = n8638 ;
  assign y4953 = ~n8642 ;
  assign y4954 = ~1'b0 ;
  assign y4955 = n8643 ;
  assign y4956 = ~1'b0 ;
  assign y4957 = ~1'b0 ;
  assign y4958 = n7841 ;
  assign y4959 = ~1'b0 ;
  assign y4960 = ~n8644 ;
  assign y4961 = ~1'b0 ;
  assign y4962 = ~n8646 ;
  assign y4963 = n8649 ;
  assign y4964 = n8653 ;
  assign y4965 = n8657 ;
  assign y4966 = 1'b0 ;
  assign y4967 = n8664 ;
  assign y4968 = ~n8665 ;
  assign y4969 = ~n8666 ;
  assign y4970 = ~1'b0 ;
  assign y4971 = ~1'b0 ;
  assign y4972 = ~n8667 ;
  assign y4973 = ~1'b0 ;
  assign y4974 = ~1'b0 ;
  assign y4975 = ~n8671 ;
  assign y4976 = ~n8675 ;
  assign y4977 = ~1'b0 ;
  assign y4978 = ~1'b0 ;
  assign y4979 = n8681 ;
  assign y4980 = n8683 ;
  assign y4981 = ~n8684 ;
  assign y4982 = n4819 ;
  assign y4983 = ~n8687 ;
  assign y4984 = n8694 ;
  assign y4985 = n8698 ;
  assign y4986 = n8701 ;
  assign y4987 = n8708 ;
  assign y4988 = ~n8710 ;
  assign y4989 = ~n8711 ;
  assign y4990 = n8713 ;
  assign y4991 = ~n8716 ;
  assign y4992 = n8721 ;
  assign y4993 = ~1'b0 ;
  assign y4994 = ~n8723 ;
  assign y4995 = n8724 ;
  assign y4996 = ~n8725 ;
  assign y4997 = ~1'b0 ;
  assign y4998 = n181 ;
  assign y4999 = ~n8726 ;
  assign y5000 = n8728 ;
  assign y5001 = ~n8737 ;
  assign y5002 = ~1'b0 ;
  assign y5003 = ~n8740 ;
  assign y5004 = ~n8743 ;
  assign y5005 = ~n8744 ;
  assign y5006 = n8746 ;
  assign y5007 = n8751 ;
  assign y5008 = n8754 ;
  assign y5009 = n8759 ;
  assign y5010 = ~n8770 ;
  assign y5011 = ~n8772 ;
  assign y5012 = ~1'b0 ;
  assign y5013 = ~n8776 ;
  assign y5014 = ~1'b0 ;
  assign y5015 = ~n2745 ;
  assign y5016 = ~n8777 ;
  assign y5017 = 1'b0 ;
  assign y5018 = ~1'b0 ;
  assign y5019 = ~n8781 ;
  assign y5020 = n6523 ;
  assign y5021 = ~1'b0 ;
  assign y5022 = n8793 ;
  assign y5023 = n8794 ;
  assign y5024 = ~n8795 ;
  assign y5025 = ~n8796 ;
  assign y5026 = n8803 ;
  assign y5027 = ~n1815 ;
  assign y5028 = n8804 ;
  assign y5029 = ~n8807 ;
  assign y5030 = ~1'b0 ;
  assign y5031 = ~1'b0 ;
  assign y5032 = ~1'b0 ;
  assign y5033 = ~n5977 ;
  assign y5034 = n8811 ;
  assign y5035 = ~1'b0 ;
  assign y5036 = n8814 ;
  assign y5037 = n8816 ;
  assign y5038 = ~1'b0 ;
  assign y5039 = ~n8818 ;
  assign y5040 = ~n8820 ;
  assign y5041 = ~1'b0 ;
  assign y5042 = ~1'b0 ;
  assign y5043 = ~n8829 ;
  assign y5044 = ~1'b0 ;
  assign y5045 = ~1'b0 ;
  assign y5046 = ~1'b0 ;
  assign y5047 = ~1'b0 ;
  assign y5048 = n4253 ;
  assign y5049 = ~1'b0 ;
  assign y5050 = 1'b0 ;
  assign y5051 = n8832 ;
  assign y5052 = 1'b0 ;
  assign y5053 = ~n8833 ;
  assign y5054 = n8837 ;
  assign y5055 = ~n8840 ;
  assign y5056 = ~n8843 ;
  assign y5057 = n8365 ;
  assign y5058 = ~1'b0 ;
  assign y5059 = ~n8846 ;
  assign y5060 = n8849 ;
  assign y5061 = ~n8851 ;
  assign y5062 = ~1'b0 ;
  assign y5063 = n8852 ;
  assign y5064 = ~n8854 ;
  assign y5065 = ~1'b0 ;
  assign y5066 = n8857 ;
  assign y5067 = ~1'b0 ;
  assign y5068 = n8862 ;
  assign y5069 = ~n8863 ;
  assign y5070 = ~1'b0 ;
  assign y5071 = n8867 ;
  assign y5072 = ~1'b0 ;
  assign y5073 = n8869 ;
  assign y5074 = ~1'b0 ;
  assign y5075 = ~n8871 ;
  assign y5076 = ~n8873 ;
  assign y5077 = n8875 ;
  assign y5078 = ~1'b0 ;
  assign y5079 = n8879 ;
  assign y5080 = n8880 ;
  assign y5081 = n3320 ;
  assign y5082 = ~1'b0 ;
  assign y5083 = n8883 ;
  assign y5084 = ~1'b0 ;
  assign y5085 = ~n8887 ;
  assign y5086 = ~1'b0 ;
  assign y5087 = n8889 ;
  assign y5088 = ~n8891 ;
  assign y5089 = ~n8894 ;
  assign y5090 = ~1'b0 ;
  assign y5091 = ~1'b0 ;
  assign y5092 = ~n8900 ;
  assign y5093 = n8902 ;
  assign y5094 = n8903 ;
  assign y5095 = ~1'b0 ;
  assign y5096 = n8905 ;
  assign y5097 = ~1'b0 ;
  assign y5098 = ~1'b0 ;
  assign y5099 = ~n8907 ;
  assign y5100 = n8910 ;
  assign y5101 = ~n8914 ;
  assign y5102 = n1281 ;
  assign y5103 = ~n8916 ;
  assign y5104 = ~1'b0 ;
  assign y5105 = n8918 ;
  assign y5106 = ~1'b0 ;
  assign y5107 = n8922 ;
  assign y5108 = n8930 ;
  assign y5109 = ~1'b0 ;
  assign y5110 = ~1'b0 ;
  assign y5111 = ~n8931 ;
  assign y5112 = ~1'b0 ;
  assign y5113 = ~1'b0 ;
  assign y5114 = n8936 ;
  assign y5115 = ~1'b0 ;
  assign y5116 = ~n8938 ;
  assign y5117 = n8941 ;
  assign y5118 = n8942 ;
  assign y5119 = ~n8951 ;
  assign y5120 = ~n512 ;
  assign y5121 = ~n8952 ;
  assign y5122 = ~1'b0 ;
  assign y5123 = ~1'b0 ;
  assign y5124 = n8956 ;
  assign y5125 = n8958 ;
  assign y5126 = ~n8959 ;
  assign y5127 = ~1'b0 ;
  assign y5128 = n8963 ;
  assign y5129 = ~1'b0 ;
  assign y5130 = ~n2182 ;
  assign y5131 = ~n8968 ;
  assign y5132 = ~n8970 ;
  assign y5133 = ~n8972 ;
  assign y5134 = n8973 ;
  assign y5135 = ~1'b0 ;
  assign y5136 = n8975 ;
  assign y5137 = n8978 ;
  assign y5138 = ~n8983 ;
  assign y5139 = ~1'b0 ;
  assign y5140 = n8984 ;
  assign y5141 = n8985 ;
  assign y5142 = ~n8986 ;
  assign y5143 = n8987 ;
  assign y5144 = ~n8989 ;
  assign y5145 = 1'b0 ;
  assign y5146 = n8992 ;
  assign y5147 = ~1'b0 ;
  assign y5148 = ~n8993 ;
  assign y5149 = ~n8997 ;
  assign y5150 = ~n8999 ;
  assign y5151 = ~1'b0 ;
  assign y5152 = n9001 ;
  assign y5153 = ~1'b0 ;
  assign y5154 = ~n9011 ;
  assign y5155 = ~n9013 ;
  assign y5156 = 1'b0 ;
  assign y5157 = ~1'b0 ;
  assign y5158 = ~1'b0 ;
  assign y5159 = ~1'b0 ;
  assign y5160 = ~1'b0 ;
  assign y5161 = ~1'b0 ;
  assign y5162 = ~1'b0 ;
  assign y5163 = ~n9014 ;
  assign y5164 = ~x123 ;
  assign y5165 = n9015 ;
  assign y5166 = ~1'b0 ;
  assign y5167 = n9016 ;
  assign y5168 = n6401 ;
  assign y5169 = ~n9021 ;
  assign y5170 = 1'b0 ;
  assign y5171 = ~n9022 ;
  assign y5172 = ~1'b0 ;
  assign y5173 = ~1'b0 ;
  assign y5174 = ~1'b0 ;
  assign y5175 = n1441 ;
  assign y5176 = ~n9024 ;
  assign y5177 = ~1'b0 ;
  assign y5178 = n9028 ;
  assign y5179 = ~n4497 ;
  assign y5180 = ~1'b0 ;
  assign y5181 = n9030 ;
  assign y5182 = ~n9034 ;
  assign y5183 = n9035 ;
  assign y5184 = n6064 ;
  assign y5185 = ~n9036 ;
  assign y5186 = ~1'b0 ;
  assign y5187 = ~n9038 ;
  assign y5188 = ~n9040 ;
  assign y5189 = n9050 ;
  assign y5190 = ~1'b0 ;
  assign y5191 = ~n9051 ;
  assign y5192 = n9053 ;
  assign y5193 = ~1'b0 ;
  assign y5194 = ~1'b0 ;
  assign y5195 = n9056 ;
  assign y5196 = ~1'b0 ;
  assign y5197 = n9058 ;
  assign y5198 = ~n5584 ;
  assign y5199 = ~1'b0 ;
  assign y5200 = n9059 ;
  assign y5201 = ~1'b0 ;
  assign y5202 = ~n9060 ;
  assign y5203 = ~n9064 ;
  assign y5204 = ~n9066 ;
  assign y5205 = n9068 ;
  assign y5206 = n9070 ;
  assign y5207 = ~n9071 ;
  assign y5208 = ~1'b0 ;
  assign y5209 = ~1'b0 ;
  assign y5210 = n835 ;
  assign y5211 = n9076 ;
  assign y5212 = ~1'b0 ;
  assign y5213 = n9079 ;
  assign y5214 = ~n9083 ;
  assign y5215 = ~1'b0 ;
  assign y5216 = n9087 ;
  assign y5217 = n9088 ;
  assign y5218 = n9089 ;
  assign y5219 = ~1'b0 ;
  assign y5220 = n9093 ;
  assign y5221 = n9098 ;
  assign y5222 = ~n9108 ;
  assign y5223 = ~n889 ;
  assign y5224 = ~n8972 ;
  assign y5225 = ~1'b0 ;
  assign y5226 = ~1'b0 ;
  assign y5227 = ~n9109 ;
  assign y5228 = ~1'b0 ;
  assign y5229 = ~1'b0 ;
  assign y5230 = n3137 ;
  assign y5231 = ~n9111 ;
  assign y5232 = n9116 ;
  assign y5233 = n9118 ;
  assign y5234 = 1'b0 ;
  assign y5235 = ~n9119 ;
  assign y5236 = ~n9122 ;
  assign y5237 = ~1'b0 ;
  assign y5238 = ~n9126 ;
  assign y5239 = n1317 ;
  assign y5240 = ~n9128 ;
  assign y5241 = ~n9129 ;
  assign y5242 = ~1'b0 ;
  assign y5243 = ~1'b0 ;
  assign y5244 = n9135 ;
  assign y5245 = n9136 ;
  assign y5246 = ~1'b0 ;
  assign y5247 = n9139 ;
  assign y5248 = n9142 ;
  assign y5249 = n288 ;
  assign y5250 = n9145 ;
  assign y5251 = n9146 ;
  assign y5252 = ~1'b0 ;
  assign y5253 = ~n9149 ;
  assign y5254 = n9150 ;
  assign y5255 = ~1'b0 ;
  assign y5256 = ~1'b0 ;
  assign y5257 = ~1'b0 ;
  assign y5258 = n9152 ;
  assign y5259 = 1'b0 ;
  assign y5260 = ~1'b0 ;
  assign y5261 = ~n9156 ;
  assign y5262 = n528 ;
  assign y5263 = ~1'b0 ;
  assign y5264 = ~1'b0 ;
  assign y5265 = n9158 ;
  assign y5266 = ~x54 ;
  assign y5267 = ~1'b0 ;
  assign y5268 = n9161 ;
  assign y5269 = ~n9165 ;
  assign y5270 = ~1'b0 ;
  assign y5271 = n9166 ;
  assign y5272 = ~1'b0 ;
  assign y5273 = ~n9168 ;
  assign y5274 = n9169 ;
  assign y5275 = ~1'b0 ;
  assign y5276 = ~1'b0 ;
  assign y5277 = ~1'b0 ;
  assign y5278 = n9172 ;
  assign y5279 = ~n9178 ;
  assign y5280 = n9179 ;
  assign y5281 = n9183 ;
  assign y5282 = ~n9185 ;
  assign y5283 = ~1'b0 ;
  assign y5284 = ~1'b0 ;
  assign y5285 = n8737 ;
  assign y5286 = ~n2896 ;
  assign y5287 = n2715 ;
  assign y5288 = ~n9186 ;
  assign y5289 = ~n9187 ;
  assign y5290 = n9190 ;
  assign y5291 = ~n9197 ;
  assign y5292 = ~n9198 ;
  assign y5293 = n9205 ;
  assign y5294 = n9207 ;
  assign y5295 = ~1'b0 ;
  assign y5296 = ~1'b0 ;
  assign y5297 = ~1'b0 ;
  assign y5298 = n9208 ;
  assign y5299 = ~n9213 ;
  assign y5300 = n9214 ;
  assign y5301 = n9215 ;
  assign y5302 = ~n9220 ;
  assign y5303 = n9224 ;
  assign y5304 = ~1'b0 ;
  assign y5305 = n9047 ;
  assign y5306 = n9226 ;
  assign y5307 = ~n9227 ;
  assign y5308 = ~n9237 ;
  assign y5309 = n5159 ;
  assign y5310 = ~n9239 ;
  assign y5311 = n9245 ;
  assign y5312 = n9247 ;
  assign y5313 = ~1'b0 ;
  assign y5314 = ~1'b0 ;
  assign y5315 = ~n9250 ;
  assign y5316 = n9251 ;
  assign y5317 = ~n9254 ;
  assign y5318 = n1180 ;
  assign y5319 = ~n9256 ;
  assign y5320 = ~1'b0 ;
  assign y5321 = ~n9257 ;
  assign y5322 = n9258 ;
  assign y5323 = n9259 ;
  assign y5324 = ~1'b0 ;
  assign y5325 = n9262 ;
  assign y5326 = n9265 ;
  assign y5327 = ~n9266 ;
  assign y5328 = ~1'b0 ;
  assign y5329 = n9267 ;
  assign y5330 = ~1'b0 ;
  assign y5331 = ~1'b0 ;
  assign y5332 = ~n9268 ;
  assign y5333 = n9270 ;
  assign y5334 = ~n9273 ;
  assign y5335 = n9275 ;
  assign y5336 = ~n9277 ;
  assign y5337 = ~n9279 ;
  assign y5338 = n9280 ;
  assign y5339 = n9281 ;
  assign y5340 = ~1'b0 ;
  assign y5341 = ~n9286 ;
  assign y5342 = ~1'b0 ;
  assign y5343 = n9288 ;
  assign y5344 = n6607 ;
  assign y5345 = n9292 ;
  assign y5346 = ~1'b0 ;
  assign y5347 = ~1'b0 ;
  assign y5348 = 1'b0 ;
  assign y5349 = n9294 ;
  assign y5350 = ~1'b0 ;
  assign y5351 = ~1'b0 ;
  assign y5352 = ~n9299 ;
  assign y5353 = ~n9300 ;
  assign y5354 = ~n9302 ;
  assign y5355 = ~1'b0 ;
  assign y5356 = ~n9305 ;
  assign y5357 = n9310 ;
  assign y5358 = ~1'b0 ;
  assign y5359 = ~n9311 ;
  assign y5360 = ~n2906 ;
  assign y5361 = ~n9312 ;
  assign y5362 = n9313 ;
  assign y5363 = n9321 ;
  assign y5364 = n9322 ;
  assign y5365 = ~1'b0 ;
  assign y5366 = ~1'b0 ;
  assign y5367 = ~1'b0 ;
  assign y5368 = ~1'b0 ;
  assign y5369 = ~n9324 ;
  assign y5370 = ~n9326 ;
  assign y5371 = ~n9332 ;
  assign y5372 = ~1'b0 ;
  assign y5373 = ~1'b0 ;
  assign y5374 = n9338 ;
  assign y5375 = n8220 ;
  assign y5376 = ~1'b0 ;
  assign y5377 = n9341 ;
  assign y5378 = ~1'b0 ;
  assign y5379 = ~n9343 ;
  assign y5380 = ~1'b0 ;
  assign y5381 = ~n7256 ;
  assign y5382 = ~n9344 ;
  assign y5383 = n9347 ;
  assign y5384 = ~1'b0 ;
  assign y5385 = ~n9349 ;
  assign y5386 = 1'b0 ;
  assign y5387 = ~n9353 ;
  assign y5388 = ~1'b0 ;
  assign y5389 = ~1'b0 ;
  assign y5390 = ~1'b0 ;
  assign y5391 = ~1'b0 ;
  assign y5392 = ~n9354 ;
  assign y5393 = ~n9355 ;
  assign y5394 = n9356 ;
  assign y5395 = ~1'b0 ;
  assign y5396 = n9364 ;
  assign y5397 = n9365 ;
  assign y5398 = ~n9374 ;
  assign y5399 = ~1'b0 ;
  assign y5400 = ~n3363 ;
  assign y5401 = ~n9376 ;
  assign y5402 = n9378 ;
  assign y5403 = ~1'b0 ;
  assign y5404 = n9335 ;
  assign y5405 = ~n6994 ;
  assign y5406 = ~1'b0 ;
  assign y5407 = n9380 ;
  assign y5408 = ~n9386 ;
  assign y5409 = n9387 ;
  assign y5410 = ~n9393 ;
  assign y5411 = ~1'b0 ;
  assign y5412 = ~1'b0 ;
  assign y5413 = ~1'b0 ;
  assign y5414 = n9397 ;
  assign y5415 = ~n9399 ;
  assign y5416 = ~1'b0 ;
  assign y5417 = ~1'b0 ;
  assign y5418 = ~1'b0 ;
  assign y5419 = ~1'b0 ;
  assign y5420 = ~1'b0 ;
  assign y5421 = ~1'b0 ;
  assign y5422 = 1'b0 ;
  assign y5423 = n9411 ;
  assign y5424 = n9412 ;
  assign y5425 = ~1'b0 ;
  assign y5426 = ~n9413 ;
  assign y5427 = ~1'b0 ;
  assign y5428 = ~1'b0 ;
  assign y5429 = ~1'b0 ;
  assign y5430 = 1'b0 ;
  assign y5431 = n9414 ;
  assign y5432 = n9415 ;
  assign y5433 = ~n562 ;
  assign y5434 = n9418 ;
  assign y5435 = n9419 ;
  assign y5436 = n9422 ;
  assign y5437 = ~n9423 ;
  assign y5438 = n5363 ;
  assign y5439 = ~n9424 ;
  assign y5440 = ~1'b0 ;
  assign y5441 = n8936 ;
  assign y5442 = ~n9429 ;
  assign y5443 = n9437 ;
  assign y5444 = ~1'b0 ;
  assign y5445 = ~n9439 ;
  assign y5446 = n9442 ;
  assign y5447 = ~n9444 ;
  assign y5448 = n9446 ;
  assign y5449 = ~1'b0 ;
  assign y5450 = 1'b0 ;
  assign y5451 = ~1'b0 ;
  assign y5452 = ~n9447 ;
  assign y5453 = ~1'b0 ;
  assign y5454 = n2203 ;
  assign y5455 = 1'b0 ;
  assign y5456 = ~1'b0 ;
  assign y5457 = n9448 ;
  assign y5458 = ~1'b0 ;
  assign y5459 = ~1'b0 ;
  assign y5460 = ~n9449 ;
  assign y5461 = n9450 ;
  assign y5462 = ~1'b0 ;
  assign y5463 = ~n9452 ;
  assign y5464 = ~1'b0 ;
  assign y5465 = ~n2542 ;
  assign y5466 = ~n9455 ;
  assign y5467 = ~1'b0 ;
  assign y5468 = ~n9461 ;
  assign y5469 = ~n2792 ;
  assign y5470 = n9462 ;
  assign y5471 = ~n9470 ;
  assign y5472 = n9473 ;
  assign y5473 = ~1'b0 ;
  assign y5474 = ~n9474 ;
  assign y5475 = 1'b0 ;
  assign y5476 = ~n9475 ;
  assign y5477 = n9479 ;
  assign y5478 = 1'b0 ;
  assign y5479 = n9481 ;
  assign y5480 = ~1'b0 ;
  assign y5481 = ~1'b0 ;
  assign y5482 = n9482 ;
  assign y5483 = n9487 ;
  assign y5484 = n9494 ;
  assign y5485 = n4157 ;
  assign y5486 = ~1'b0 ;
  assign y5487 = n9495 ;
  assign y5488 = ~n9501 ;
  assign y5489 = ~1'b0 ;
  assign y5490 = n9502 ;
  assign y5491 = n9503 ;
  assign y5492 = ~1'b0 ;
  assign y5493 = n9506 ;
  assign y5494 = ~1'b0 ;
  assign y5495 = n9508 ;
  assign y5496 = ~1'b0 ;
  assign y5497 = n9511 ;
  assign y5498 = ~1'b0 ;
  assign y5499 = n9512 ;
  assign y5500 = n9514 ;
  assign y5501 = ~n9517 ;
  assign y5502 = ~n9519 ;
  assign y5503 = ~1'b0 ;
  assign y5504 = 1'b0 ;
  assign y5505 = ~n6268 ;
  assign y5506 = n9520 ;
  assign y5507 = n9523 ;
  assign y5508 = ~n9526 ;
  assign y5509 = ~1'b0 ;
  assign y5510 = ~1'b0 ;
  assign y5511 = ~1'b0 ;
  assign y5512 = ~1'b0 ;
  assign y5513 = n9530 ;
  assign y5514 = ~n1329 ;
  assign y5515 = n9531 ;
  assign y5516 = n9533 ;
  assign y5517 = ~n9534 ;
  assign y5518 = ~1'b0 ;
  assign y5519 = n9536 ;
  assign y5520 = ~1'b0 ;
  assign y5521 = ~n9542 ;
  assign y5522 = n9544 ;
  assign y5523 = n9547 ;
  assign y5524 = ~1'b0 ;
  assign y5525 = n4364 ;
  assign y5526 = n9548 ;
  assign y5527 = ~n3521 ;
  assign y5528 = ~n9549 ;
  assign y5529 = ~1'b0 ;
  assign y5530 = n9553 ;
  assign y5531 = ~1'b0 ;
  assign y5532 = n9554 ;
  assign y5533 = ~1'b0 ;
  assign y5534 = ~1'b0 ;
  assign y5535 = n9556 ;
  assign y5536 = ~n9559 ;
  assign y5537 = 1'b0 ;
  assign y5538 = n9560 ;
  assign y5539 = ~n9569 ;
  assign y5540 = ~n9571 ;
  assign y5541 = ~n9572 ;
  assign y5542 = n9574 ;
  assign y5543 = n9575 ;
  assign y5544 = ~n9576 ;
  assign y5545 = ~1'b0 ;
  assign y5546 = ~n8185 ;
  assign y5547 = n9585 ;
  assign y5548 = ~1'b0 ;
  assign y5549 = ~n9586 ;
  assign y5550 = ~1'b0 ;
  assign y5551 = ~n9590 ;
  assign y5552 = ~n9592 ;
  assign y5553 = n9594 ;
  assign y5554 = ~1'b0 ;
  assign y5555 = ~1'b0 ;
  assign y5556 = ~n9596 ;
  assign y5557 = ~1'b0 ;
  assign y5558 = 1'b0 ;
  assign y5559 = ~n9604 ;
  assign y5560 = n9606 ;
  assign y5561 = ~1'b0 ;
  assign y5562 = ~1'b0 ;
  assign y5563 = ~n9608 ;
  assign y5564 = ~1'b0 ;
  assign y5565 = ~1'b0 ;
  assign y5566 = ~1'b0 ;
  assign y5567 = n9609 ;
  assign y5568 = ~1'b0 ;
  assign y5569 = n9612 ;
  assign y5570 = n9614 ;
  assign y5571 = ~n9615 ;
  assign y5572 = ~n9617 ;
  assign y5573 = n9618 ;
  assign y5574 = ~n9620 ;
  assign y5575 = n9623 ;
  assign y5576 = ~n9624 ;
  assign y5577 = n9626 ;
  assign y5578 = n9628 ;
  assign y5579 = n9629 ;
  assign y5580 = ~n9630 ;
  assign y5581 = ~n9641 ;
  assign y5582 = ~1'b0 ;
  assign y5583 = n9648 ;
  assign y5584 = n9653 ;
  assign y5585 = ~n9657 ;
  assign y5586 = ~1'b0 ;
  assign y5587 = n9658 ;
  assign y5588 = ~1'b0 ;
  assign y5589 = ~1'b0 ;
  assign y5590 = n9660 ;
  assign y5591 = ~1'b0 ;
  assign y5592 = n7563 ;
  assign y5593 = n9668 ;
  assign y5594 = n9670 ;
  assign y5595 = ~1'b0 ;
  assign y5596 = n9671 ;
  assign y5597 = ~n8224 ;
  assign y5598 = ~1'b0 ;
  assign y5599 = n9672 ;
  assign y5600 = ~1'b0 ;
  assign y5601 = n8496 ;
  assign y5602 = n9675 ;
  assign y5603 = n729 ;
  assign y5604 = n9676 ;
  assign y5605 = n9677 ;
  assign y5606 = ~n9680 ;
  assign y5607 = n9681 ;
  assign y5608 = n9299 ;
  assign y5609 = n9683 ;
  assign y5610 = n9684 ;
  assign y5611 = n9690 ;
  assign y5612 = n9695 ;
  assign y5613 = ~n9697 ;
  assign y5614 = ~1'b0 ;
  assign y5615 = ~n9704 ;
  assign y5616 = ~n3947 ;
  assign y5617 = ~1'b0 ;
  assign y5618 = ~n9706 ;
  assign y5619 = n9708 ;
  assign y5620 = ~1'b0 ;
  assign y5621 = ~n9709 ;
  assign y5622 = n9710 ;
  assign y5623 = ~n9711 ;
  assign y5624 = ~1'b0 ;
  assign y5625 = ~n9716 ;
  assign y5626 = ~1'b0 ;
  assign y5627 = ~n6959 ;
  assign y5628 = n504 ;
  assign y5629 = n9717 ;
  assign y5630 = ~n9718 ;
  assign y5631 = ~1'b0 ;
  assign y5632 = ~n9719 ;
  assign y5633 = ~1'b0 ;
  assign y5634 = ~1'b0 ;
  assign y5635 = n9725 ;
  assign y5636 = ~n9732 ;
  assign y5637 = ~n9736 ;
  assign y5638 = ~1'b0 ;
  assign y5639 = ~n9737 ;
  assign y5640 = ~n9745 ;
  assign y5641 = 1'b0 ;
  assign y5642 = ~1'b0 ;
  assign y5643 = ~1'b0 ;
  assign y5644 = ~1'b0 ;
  assign y5645 = ~n9746 ;
  assign y5646 = n9749 ;
  assign y5647 = 1'b0 ;
  assign y5648 = n9751 ;
  assign y5649 = n9753 ;
  assign y5650 = ~n9761 ;
  assign y5651 = ~1'b0 ;
  assign y5652 = ~n9766 ;
  assign y5653 = ~n9775 ;
  assign y5654 = n9777 ;
  assign y5655 = n9779 ;
  assign y5656 = ~n9782 ;
  assign y5657 = n9785 ;
  assign y5658 = n9789 ;
  assign y5659 = n9795 ;
  assign y5660 = ~n9798 ;
  assign y5661 = n9799 ;
  assign y5662 = ~n2340 ;
  assign y5663 = n3226 ;
  assign y5664 = n9800 ;
  assign y5665 = ~n9805 ;
  assign y5666 = ~1'b0 ;
  assign y5667 = ~n9806 ;
  assign y5668 = ~n9808 ;
  assign y5669 = ~n9811 ;
  assign y5670 = ~1'b0 ;
  assign y5671 = ~1'b0 ;
  assign y5672 = ~1'b0 ;
  assign y5673 = ~n5910 ;
  assign y5674 = ~n9816 ;
  assign y5675 = ~n4265 ;
  assign y5676 = n9822 ;
  assign y5677 = ~n9823 ;
  assign y5678 = n9826 ;
  assign y5679 = n9827 ;
  assign y5680 = ~n9828 ;
  assign y5681 = n9831 ;
  assign y5682 = ~n9833 ;
  assign y5683 = ~1'b0 ;
  assign y5684 = n9836 ;
  assign y5685 = n9838 ;
  assign y5686 = ~1'b0 ;
  assign y5687 = n550 ;
  assign y5688 = ~n1001 ;
  assign y5689 = n9839 ;
  assign y5690 = ~n9840 ;
  assign y5691 = n9845 ;
  assign y5692 = ~1'b0 ;
  assign y5693 = n9846 ;
  assign y5694 = n9848 ;
  assign y5695 = n9850 ;
  assign y5696 = ~n9851 ;
  assign y5697 = n9852 ;
  assign y5698 = ~n9853 ;
  assign y5699 = ~1'b0 ;
  assign y5700 = n9854 ;
  assign y5701 = ~1'b0 ;
  assign y5702 = ~1'b0 ;
  assign y5703 = ~1'b0 ;
  assign y5704 = ~1'b0 ;
  assign y5705 = n9856 ;
  assign y5706 = ~n9859 ;
  assign y5707 = ~n9863 ;
  assign y5708 = n9865 ;
  assign y5709 = n9866 ;
  assign y5710 = n9867 ;
  assign y5711 = ~n9869 ;
  assign y5712 = ~1'b0 ;
  assign y5713 = ~1'b0 ;
  assign y5714 = n9870 ;
  assign y5715 = ~n9874 ;
  assign y5716 = ~n9877 ;
  assign y5717 = ~1'b0 ;
  assign y5718 = ~n9887 ;
  assign y5719 = ~n9891 ;
  assign y5720 = ~n1862 ;
  assign y5721 = n9892 ;
  assign y5722 = ~1'b0 ;
  assign y5723 = n9894 ;
  assign y5724 = ~n9895 ;
  assign y5725 = n9896 ;
  assign y5726 = n579 ;
  assign y5727 = ~n9897 ;
  assign y5728 = ~n6575 ;
  assign y5729 = n3166 ;
  assign y5730 = 1'b0 ;
  assign y5731 = ~n9901 ;
  assign y5732 = ~1'b0 ;
  assign y5733 = ~1'b0 ;
  assign y5734 = ~1'b0 ;
  assign y5735 = ~1'b0 ;
  assign y5736 = ~1'b0 ;
  assign y5737 = ~x36 ;
  assign y5738 = ~1'b0 ;
  assign y5739 = ~n9903 ;
  assign y5740 = ~n9906 ;
  assign y5741 = ~1'b0 ;
  assign y5742 = ~n9911 ;
  assign y5743 = ~1'b0 ;
  assign y5744 = n8762 ;
  assign y5745 = ~1'b0 ;
  assign y5746 = n9914 ;
  assign y5747 = ~1'b0 ;
  assign y5748 = ~n9915 ;
  assign y5749 = ~n9916 ;
  assign y5750 = ~1'b0 ;
  assign y5751 = n9919 ;
  assign y5752 = ~n9924 ;
  assign y5753 = ~n9928 ;
  assign y5754 = ~n9938 ;
  assign y5755 = ~n8824 ;
  assign y5756 = ~1'b0 ;
  assign y5757 = n9940 ;
  assign y5758 = n9946 ;
  assign y5759 = ~1'b0 ;
  assign y5760 = ~n9947 ;
  assign y5761 = ~n9952 ;
  assign y5762 = ~1'b0 ;
  assign y5763 = ~1'b0 ;
  assign y5764 = ~n9954 ;
  assign y5765 = n9959 ;
  assign y5766 = 1'b0 ;
  assign y5767 = ~n9961 ;
  assign y5768 = ~n9962 ;
  assign y5769 = n9979 ;
  assign y5770 = ~n9981 ;
  assign y5771 = ~1'b0 ;
  assign y5772 = ~1'b0 ;
  assign y5773 = n6393 ;
  assign y5774 = ~1'b0 ;
  assign y5775 = ~1'b0 ;
  assign y5776 = n9988 ;
  assign y5777 = n9990 ;
  assign y5778 = ~1'b0 ;
  assign y5779 = n6313 ;
  assign y5780 = ~1'b0 ;
  assign y5781 = ~n2459 ;
  assign y5782 = n9992 ;
  assign y5783 = n9997 ;
  assign y5784 = ~1'b0 ;
  assign y5785 = ~n10006 ;
  assign y5786 = ~1'b0 ;
  assign y5787 = n10011 ;
  assign y5788 = 1'b0 ;
  assign y5789 = ~n10015 ;
  assign y5790 = ~1'b0 ;
  assign y5791 = ~1'b0 ;
  assign y5792 = ~n10016 ;
  assign y5793 = ~n10020 ;
  assign y5794 = n10021 ;
  assign y5795 = ~n10022 ;
  assign y5796 = n10024 ;
  assign y5797 = ~n10026 ;
  assign y5798 = ~n10027 ;
  assign y5799 = n5223 ;
  assign y5800 = ~n10029 ;
  assign y5801 = ~n10031 ;
  assign y5802 = n4648 ;
  assign y5803 = ~n8872 ;
  assign y5804 = n10042 ;
  assign y5805 = ~1'b0 ;
  assign y5806 = ~1'b0 ;
  assign y5807 = ~1'b0 ;
  assign y5808 = ~1'b0 ;
  assign y5809 = ~n5688 ;
  assign y5810 = 1'b0 ;
  assign y5811 = ~1'b0 ;
  assign y5812 = n6727 ;
  assign y5813 = ~1'b0 ;
  assign y5814 = ~n10045 ;
  assign y5815 = ~1'b0 ;
  assign y5816 = ~n10046 ;
  assign y5817 = ~n10047 ;
  assign y5818 = n10048 ;
  assign y5819 = n629 ;
  assign y5820 = n183 ;
  assign y5821 = ~n10049 ;
  assign y5822 = n10051 ;
  assign y5823 = ~n10054 ;
  assign y5824 = ~n10055 ;
  assign y5825 = n4028 ;
  assign y5826 = ~n10058 ;
  assign y5827 = n9381 ;
  assign y5828 = n10063 ;
  assign y5829 = ~n10065 ;
  assign y5830 = ~n10068 ;
  assign y5831 = ~n10069 ;
  assign y5832 = ~1'b0 ;
  assign y5833 = 1'b0 ;
  assign y5834 = ~1'b0 ;
  assign y5835 = n1645 ;
  assign y5836 = n10072 ;
  assign y5837 = ~n10074 ;
  assign y5838 = ~1'b0 ;
  assign y5839 = ~n9572 ;
  assign y5840 = ~n10076 ;
  assign y5841 = ~n10077 ;
  assign y5842 = n10078 ;
  assign y5843 = ~n10079 ;
  assign y5844 = ~n10080 ;
  assign y5845 = ~n10081 ;
  assign y5846 = ~1'b0 ;
  assign y5847 = n10083 ;
  assign y5848 = ~1'b0 ;
  assign y5849 = n10086 ;
  assign y5850 = ~n10089 ;
  assign y5851 = ~1'b0 ;
  assign y5852 = n10091 ;
  assign y5853 = ~1'b0 ;
  assign y5854 = ~1'b0 ;
  assign y5855 = 1'b0 ;
  assign y5856 = ~n10095 ;
  assign y5857 = ~1'b0 ;
  assign y5858 = ~1'b0 ;
  assign y5859 = ~n10096 ;
  assign y5860 = ~1'b0 ;
  assign y5861 = n10098 ;
  assign y5862 = ~n10099 ;
  assign y5863 = ~n10118 ;
  assign y5864 = ~n7242 ;
  assign y5865 = ~1'b0 ;
  assign y5866 = ~n10120 ;
  assign y5867 = n10121 ;
  assign y5868 = ~1'b0 ;
  assign y5869 = ~n10125 ;
  assign y5870 = ~n10126 ;
  assign y5871 = ~n10128 ;
  assign y5872 = ~n10132 ;
  assign y5873 = 1'b0 ;
  assign y5874 = ~1'b0 ;
  assign y5875 = ~n10134 ;
  assign y5876 = 1'b0 ;
  assign y5877 = ~1'b0 ;
  assign y5878 = ~1'b0 ;
  assign y5879 = ~n10136 ;
  assign y5880 = 1'b0 ;
  assign y5881 = ~1'b0 ;
  assign y5882 = ~n10139 ;
  assign y5883 = ~n10141 ;
  assign y5884 = n10142 ;
  assign y5885 = n10144 ;
  assign y5886 = ~1'b0 ;
  assign y5887 = n10149 ;
  assign y5888 = ~1'b0 ;
  assign y5889 = n2420 ;
  assign y5890 = ~1'b0 ;
  assign y5891 = n10151 ;
  assign y5892 = ~1'b0 ;
  assign y5893 = ~n10153 ;
  assign y5894 = ~1'b0 ;
  assign y5895 = ~n10156 ;
  assign y5896 = ~n10157 ;
  assign y5897 = ~1'b0 ;
  assign y5898 = ~n10158 ;
  assign y5899 = ~n10160 ;
  assign y5900 = ~n10165 ;
  assign y5901 = ~n4376 ;
  assign y5902 = ~n10166 ;
  assign y5903 = ~1'b0 ;
  assign y5904 = ~1'b0 ;
  assign y5905 = ~n10170 ;
  assign y5906 = n10172 ;
  assign y5907 = n10177 ;
  assign y5908 = ~n704 ;
  assign y5909 = ~n10178 ;
  assign y5910 = ~1'b0 ;
  assign y5911 = n10179 ;
  assign y5912 = ~1'b0 ;
  assign y5913 = ~n2322 ;
  assign y5914 = n10183 ;
  assign y5915 = n10184 ;
  assign y5916 = ~n10187 ;
  assign y5917 = ~1'b0 ;
  assign y5918 = n6563 ;
  assign y5919 = ~1'b0 ;
  assign y5920 = n10189 ;
  assign y5921 = ~n10190 ;
  assign y5922 = ~1'b0 ;
  assign y5923 = ~n10191 ;
  assign y5924 = n10192 ;
  assign y5925 = ~n10195 ;
  assign y5926 = ~n10197 ;
  assign y5927 = n10199 ;
  assign y5928 = ~n10203 ;
  assign y5929 = ~n10212 ;
  assign y5930 = ~1'b0 ;
  assign y5931 = n10213 ;
  assign y5932 = 1'b0 ;
  assign y5933 = ~n10216 ;
  assign y5934 = x125 ;
  assign y5935 = ~1'b0 ;
  assign y5936 = ~1'b0 ;
  assign y5937 = n10217 ;
  assign y5938 = ~1'b0 ;
  assign y5939 = ~n10225 ;
  assign y5940 = ~1'b0 ;
  assign y5941 = ~1'b0 ;
  assign y5942 = ~n2932 ;
  assign y5943 = ~1'b0 ;
  assign y5944 = ~n10227 ;
  assign y5945 = ~1'b0 ;
  assign y5946 = 1'b0 ;
  assign y5947 = n10230 ;
  assign y5948 = n10231 ;
  assign y5949 = 1'b0 ;
  assign y5950 = n10237 ;
  assign y5951 = ~n10241 ;
  assign y5952 = n10242 ;
  assign y5953 = ~1'b0 ;
  assign y5954 = ~1'b0 ;
  assign y5955 = ~n10243 ;
  assign y5956 = ~n10245 ;
  assign y5957 = ~n10247 ;
  assign y5958 = 1'b0 ;
  assign y5959 = n10250 ;
  assign y5960 = ~n10255 ;
  assign y5961 = n10257 ;
  assign y5962 = n10261 ;
  assign y5963 = ~n10262 ;
  assign y5964 = ~n10265 ;
  assign y5965 = n10266 ;
  assign y5966 = ~n10268 ;
  assign y5967 = ~n10277 ;
  assign y5968 = x18 ;
  assign y5969 = n10278 ;
  assign y5970 = n10281 ;
  assign y5971 = ~1'b0 ;
  assign y5972 = ~1'b0 ;
  assign y5973 = n10282 ;
  assign y5974 = ~n10283 ;
  assign y5975 = ~n10284 ;
  assign y5976 = ~n10285 ;
  assign y5977 = ~1'b0 ;
  assign y5978 = n1116 ;
  assign y5979 = ~n10287 ;
  assign y5980 = ~1'b0 ;
  assign y5981 = n10292 ;
  assign y5982 = ~n10293 ;
  assign y5983 = ~1'b0 ;
  assign y5984 = ~1'b0 ;
  assign y5985 = ~1'b0 ;
  assign y5986 = ~1'b0 ;
  assign y5987 = ~n10295 ;
  assign y5988 = ~1'b0 ;
  assign y5989 = ~n10296 ;
  assign y5990 = ~1'b0 ;
  assign y5991 = ~n10297 ;
  assign y5992 = ~1'b0 ;
  assign y5993 = ~n10301 ;
  assign y5994 = ~1'b0 ;
  assign y5995 = n10302 ;
  assign y5996 = ~1'b0 ;
  assign y5997 = ~n10303 ;
  assign y5998 = n10304 ;
  assign y5999 = ~1'b0 ;
  assign y6000 = ~n6718 ;
  assign y6001 = ~1'b0 ;
  assign y6002 = ~1'b0 ;
  assign y6003 = n10305 ;
  assign y6004 = n10308 ;
  assign y6005 = n10311 ;
  assign y6006 = ~1'b0 ;
  assign y6007 = ~1'b0 ;
  assign y6008 = n10315 ;
  assign y6009 = n2093 ;
  assign y6010 = ~n10318 ;
  assign y6011 = n10319 ;
  assign y6012 = ~1'b0 ;
  assign y6013 = ~1'b0 ;
  assign y6014 = n10323 ;
  assign y6015 = ~1'b0 ;
  assign y6016 = n10324 ;
  assign y6017 = n10328 ;
  assign y6018 = ~n10331 ;
  assign y6019 = ~1'b0 ;
  assign y6020 = n10336 ;
  assign y6021 = n10343 ;
  assign y6022 = n10350 ;
  assign y6023 = ~1'b0 ;
  assign y6024 = ~1'b0 ;
  assign y6025 = ~1'b0 ;
  assign y6026 = ~1'b0 ;
  assign y6027 = n10354 ;
  assign y6028 = n5023 ;
  assign y6029 = ~1'b0 ;
  assign y6030 = ~n10356 ;
  assign y6031 = x84 ;
  assign y6032 = n10357 ;
  assign y6033 = ~1'b0 ;
  assign y6034 = ~1'b0 ;
  assign y6035 = ~n10359 ;
  assign y6036 = n10361 ;
  assign y6037 = n10367 ;
  assign y6038 = ~1'b0 ;
  assign y6039 = ~n10375 ;
  assign y6040 = ~1'b0 ;
  assign y6041 = ~1'b0 ;
  assign y6042 = ~n2785 ;
  assign y6043 = n10377 ;
  assign y6044 = ~n10378 ;
  assign y6045 = n10381 ;
  assign y6046 = ~1'b0 ;
  assign y6047 = ~1'b0 ;
  assign y6048 = ~n10382 ;
  assign y6049 = n10387 ;
  assign y6050 = n10392 ;
  assign y6051 = ~1'b0 ;
  assign y6052 = ~1'b0 ;
  assign y6053 = ~n10398 ;
  assign y6054 = ~1'b0 ;
  assign y6055 = ~n10400 ;
  assign y6056 = n10405 ;
  assign y6057 = n10408 ;
  assign y6058 = n10411 ;
  assign y6059 = n10412 ;
  assign y6060 = 1'b0 ;
  assign y6061 = ~n409 ;
  assign y6062 = ~n10414 ;
  assign y6063 = n10417 ;
  assign y6064 = ~1'b0 ;
  assign y6065 = ~1'b0 ;
  assign y6066 = ~1'b0 ;
  assign y6067 = ~n10419 ;
  assign y6068 = ~n10420 ;
  assign y6069 = ~1'b0 ;
  assign y6070 = ~n10422 ;
  assign y6071 = n10423 ;
  assign y6072 = 1'b0 ;
  assign y6073 = n10424 ;
  assign y6074 = ~n10429 ;
  assign y6075 = ~1'b0 ;
  assign y6076 = n10431 ;
  assign y6077 = ~n10432 ;
  assign y6078 = ~1'b0 ;
  assign y6079 = n10435 ;
  assign y6080 = ~n10436 ;
  assign y6081 = ~n10438 ;
  assign y6082 = ~n10441 ;
  assign y6083 = ~1'b0 ;
  assign y6084 = ~1'b0 ;
  assign y6085 = ~n10442 ;
  assign y6086 = ~n10446 ;
  assign y6087 = n10448 ;
  assign y6088 = ~n10453 ;
  assign y6089 = ~n10456 ;
  assign y6090 = ~1'b0 ;
  assign y6091 = ~n10461 ;
  assign y6092 = ~n10462 ;
  assign y6093 = ~1'b0 ;
  assign y6094 = n10463 ;
  assign y6095 = n10466 ;
  assign y6096 = n10468 ;
  assign y6097 = ~1'b0 ;
  assign y6098 = ~n10470 ;
  assign y6099 = n10471 ;
  assign y6100 = ~1'b0 ;
  assign y6101 = ~n10474 ;
  assign y6102 = n3050 ;
  assign y6103 = ~1'b0 ;
  assign y6104 = n10478 ;
  assign y6105 = n9719 ;
  assign y6106 = ~n1329 ;
  assign y6107 = ~1'b0 ;
  assign y6108 = ~1'b0 ;
  assign y6109 = n10479 ;
  assign y6110 = ~1'b0 ;
  assign y6111 = ~n10482 ;
  assign y6112 = ~1'b0 ;
  assign y6113 = ~n10483 ;
  assign y6114 = n10486 ;
  assign y6115 = ~n10489 ;
  assign y6116 = ~1'b0 ;
  assign y6117 = ~1'b0 ;
  assign y6118 = ~n10492 ;
  assign y6119 = n10493 ;
  assign y6120 = ~n877 ;
  assign y6121 = ~n520 ;
  assign y6122 = ~n10496 ;
  assign y6123 = ~1'b0 ;
  assign y6124 = ~1'b0 ;
  assign y6125 = ~1'b0 ;
  assign y6126 = 1'b0 ;
  assign y6127 = n10497 ;
  assign y6128 = n1905 ;
  assign y6129 = n10498 ;
  assign y6130 = ~n10499 ;
  assign y6131 = ~n10500 ;
  assign y6132 = n3868 ;
  assign y6133 = ~n10507 ;
  assign y6134 = ~1'b0 ;
  assign y6135 = ~n10513 ;
  assign y6136 = 1'b0 ;
  assign y6137 = ~n10514 ;
  assign y6138 = n10518 ;
  assign y6139 = ~n10519 ;
  assign y6140 = ~n10521 ;
  assign y6141 = ~1'b0 ;
  assign y6142 = n10523 ;
  assign y6143 = n10524 ;
  assign y6144 = 1'b0 ;
  assign y6145 = n10527 ;
  assign y6146 = ~1'b0 ;
  assign y6147 = ~1'b0 ;
  assign y6148 = n10529 ;
  assign y6149 = ~n10534 ;
  assign y6150 = ~n10537 ;
  assign y6151 = ~n10543 ;
  assign y6152 = ~n10551 ;
  assign y6153 = ~n10552 ;
  assign y6154 = ~1'b0 ;
  assign y6155 = 1'b0 ;
  assign y6156 = ~n10553 ;
  assign y6157 = n10554 ;
  assign y6158 = ~1'b0 ;
  assign y6159 = 1'b0 ;
  assign y6160 = 1'b0 ;
  assign y6161 = 1'b0 ;
  assign y6162 = ~1'b0 ;
  assign y6163 = ~n10555 ;
  assign y6164 = ~n10556 ;
  assign y6165 = ~1'b0 ;
  assign y6166 = ~1'b0 ;
  assign y6167 = ~n10558 ;
  assign y6168 = ~n10559 ;
  assign y6169 = ~n10560 ;
  assign y6170 = ~n10565 ;
  assign y6171 = n10566 ;
  assign y6172 = n10568 ;
  assign y6173 = ~1'b0 ;
  assign y6174 = n10571 ;
  assign y6175 = ~1'b0 ;
  assign y6176 = ~1'b0 ;
  assign y6177 = ~1'b0 ;
  assign y6178 = ~1'b0 ;
  assign y6179 = ~n3587 ;
  assign y6180 = n10572 ;
  assign y6181 = ~1'b0 ;
  assign y6182 = ~n10147 ;
  assign y6183 = ~n10576 ;
  assign y6184 = ~1'b0 ;
  assign y6185 = ~n10589 ;
  assign y6186 = ~1'b0 ;
  assign y6187 = n10595 ;
  assign y6188 = n10597 ;
  assign y6189 = n10598 ;
  assign y6190 = ~1'b0 ;
  assign y6191 = ~1'b0 ;
  assign y6192 = ~1'b0 ;
  assign y6193 = n9315 ;
  assign y6194 = n10599 ;
  assign y6195 = n10600 ;
  assign y6196 = n10604 ;
  assign y6197 = ~n10605 ;
  assign y6198 = ~1'b0 ;
  assign y6199 = ~n10616 ;
  assign y6200 = n10617 ;
  assign y6201 = ~1'b0 ;
  assign y6202 = ~1'b0 ;
  assign y6203 = ~1'b0 ;
  assign y6204 = ~1'b0 ;
  assign y6205 = ~n5028 ;
  assign y6206 = ~1'b0 ;
  assign y6207 = n10618 ;
  assign y6208 = n10619 ;
  assign y6209 = n10621 ;
  assign y6210 = n10624 ;
  assign y6211 = ~1'b0 ;
  assign y6212 = ~n10628 ;
  assign y6213 = n10630 ;
  assign y6214 = ~n10635 ;
  assign y6215 = ~1'b0 ;
  assign y6216 = ~n10636 ;
  assign y6217 = ~n10641 ;
  assign y6218 = ~n10642 ;
  assign y6219 = ~1'b0 ;
  assign y6220 = ~n10644 ;
  assign y6221 = ~1'b0 ;
  assign y6222 = ~n10659 ;
  assign y6223 = ~1'b0 ;
  assign y6224 = ~n10660 ;
  assign y6225 = ~1'b0 ;
  assign y6226 = n10662 ;
  assign y6227 = ~1'b0 ;
  assign y6228 = n10663 ;
  assign y6229 = ~1'b0 ;
  assign y6230 = ~1'b0 ;
  assign y6231 = ~1'b0 ;
  assign y6232 = ~n10665 ;
  assign y6233 = ~n8861 ;
  assign y6234 = ~n10666 ;
  assign y6235 = n10669 ;
  assign y6236 = n10671 ;
  assign y6237 = n10679 ;
  assign y6238 = ~1'b0 ;
  assign y6239 = n10681 ;
  assign y6240 = ~n10682 ;
  assign y6241 = ~1'b0 ;
  assign y6242 = n6667 ;
  assign y6243 = ~1'b0 ;
  assign y6244 = ~n10684 ;
  assign y6245 = ~n10686 ;
  assign y6246 = ~1'b0 ;
  assign y6247 = 1'b0 ;
  assign y6248 = n10690 ;
  assign y6249 = ~1'b0 ;
  assign y6250 = ~1'b0 ;
  assign y6251 = ~1'b0 ;
  assign y6252 = ~n10696 ;
  assign y6253 = n10698 ;
  assign y6254 = n7695 ;
  assign y6255 = n10699 ;
  assign y6256 = n10703 ;
  assign y6257 = ~n10704 ;
  assign y6258 = ~n7509 ;
  assign y6259 = n10707 ;
  assign y6260 = ~n10708 ;
  assign y6261 = ~n10709 ;
  assign y6262 = ~1'b0 ;
  assign y6263 = ~n4087 ;
  assign y6264 = ~n1932 ;
  assign y6265 = ~1'b0 ;
  assign y6266 = ~1'b0 ;
  assign y6267 = ~1'b0 ;
  assign y6268 = ~1'b0 ;
  assign y6269 = ~n10710 ;
  assign y6270 = ~1'b0 ;
  assign y6271 = ~n10712 ;
  assign y6272 = ~1'b0 ;
  assign y6273 = ~1'b0 ;
  assign y6274 = ~1'b0 ;
  assign y6275 = n10715 ;
  assign y6276 = n10716 ;
  assign y6277 = ~n4252 ;
  assign y6278 = n10718 ;
  assign y6279 = 1'b0 ;
  assign y6280 = ~n10721 ;
  assign y6281 = n10725 ;
  assign y6282 = ~1'b0 ;
  assign y6283 = ~n10728 ;
  assign y6284 = n10747 ;
  assign y6285 = n10748 ;
  assign y6286 = ~1'b0 ;
  assign y6287 = ~1'b0 ;
  assign y6288 = ~n10750 ;
  assign y6289 = ~n10499 ;
  assign y6290 = n10754 ;
  assign y6291 = ~1'b0 ;
  assign y6292 = ~n10758 ;
  assign y6293 = 1'b0 ;
  assign y6294 = ~1'b0 ;
  assign y6295 = n10759 ;
  assign y6296 = ~n10760 ;
  assign y6297 = n10761 ;
  assign y6298 = n10765 ;
  assign y6299 = ~n10769 ;
  assign y6300 = n10771 ;
  assign y6301 = n4682 ;
  assign y6302 = ~n10774 ;
  assign y6303 = ~n10776 ;
  assign y6304 = ~n10788 ;
  assign y6305 = 1'b0 ;
  assign y6306 = ~1'b0 ;
  assign y6307 = ~1'b0 ;
  assign y6308 = ~n3436 ;
  assign y6309 = ~n10789 ;
  assign y6310 = n10790 ;
  assign y6311 = n10795 ;
  assign y6312 = n10797 ;
  assign y6313 = ~n10799 ;
  assign y6314 = ~n10800 ;
  assign y6315 = n10802 ;
  assign y6316 = ~1'b0 ;
  assign y6317 = ~1'b0 ;
  assign y6318 = n10803 ;
  assign y6319 = n10805 ;
  assign y6320 = n10806 ;
  assign y6321 = ~n3428 ;
  assign y6322 = ~1'b0 ;
  assign y6323 = ~n10810 ;
  assign y6324 = n5418 ;
  assign y6325 = 1'b0 ;
  assign y6326 = ~1'b0 ;
  assign y6327 = ~1'b0 ;
  assign y6328 = n10813 ;
  assign y6329 = ~n10815 ;
  assign y6330 = ~n10820 ;
  assign y6331 = ~1'b0 ;
  assign y6332 = ~1'b0 ;
  assign y6333 = n10825 ;
  assign y6334 = 1'b0 ;
  assign y6335 = n10827 ;
  assign y6336 = n10832 ;
  assign y6337 = ~n10835 ;
  assign y6338 = ~1'b0 ;
  assign y6339 = ~1'b0 ;
  assign y6340 = n10836 ;
  assign y6341 = n10841 ;
  assign y6342 = ~1'b0 ;
  assign y6343 = ~1'b0 ;
  assign y6344 = n10843 ;
  assign y6345 = n10847 ;
  assign y6346 = n10848 ;
  assign y6347 = ~1'b0 ;
  assign y6348 = n10849 ;
  assign y6349 = 1'b0 ;
  assign y6350 = ~n10853 ;
  assign y6351 = ~n10856 ;
  assign y6352 = n10857 ;
  assign y6353 = ~n10858 ;
  assign y6354 = n10859 ;
  assign y6355 = n10860 ;
  assign y6356 = ~1'b0 ;
  assign y6357 = ~n10861 ;
  assign y6358 = ~n10863 ;
  assign y6359 = x102 ;
  assign y6360 = ~1'b0 ;
  assign y6361 = ~1'b0 ;
  assign y6362 = ~1'b0 ;
  assign y6363 = n10866 ;
  assign y6364 = ~n10867 ;
  assign y6365 = n10868 ;
  assign y6366 = ~n10869 ;
  assign y6367 = ~1'b0 ;
  assign y6368 = n10874 ;
  assign y6369 = ~n10876 ;
  assign y6370 = ~1'b0 ;
  assign y6371 = n10881 ;
  assign y6372 = n10886 ;
  assign y6373 = ~n10889 ;
  assign y6374 = n10890 ;
  assign y6375 = ~n5526 ;
  assign y6376 = n6102 ;
  assign y6377 = ~1'b0 ;
  assign y6378 = ~1'b0 ;
  assign y6379 = n10891 ;
  assign y6380 = ~1'b0 ;
  assign y6381 = ~1'b0 ;
  assign y6382 = ~1'b0 ;
  assign y6383 = ~n10895 ;
  assign y6384 = ~n10896 ;
  assign y6385 = ~n10899 ;
  assign y6386 = ~n10901 ;
  assign y6387 = ~1'b0 ;
  assign y6388 = n10903 ;
  assign y6389 = n10905 ;
  assign y6390 = n134 ;
  assign y6391 = ~n10909 ;
  assign y6392 = n1784 ;
  assign y6393 = n10912 ;
  assign y6394 = ~1'b0 ;
  assign y6395 = n10913 ;
  assign y6396 = ~1'b0 ;
  assign y6397 = ~n10914 ;
  assign y6398 = ~n10916 ;
  assign y6399 = ~n10922 ;
  assign y6400 = n10925 ;
  assign y6401 = ~1'b0 ;
  assign y6402 = n10927 ;
  assign y6403 = ~n10929 ;
  assign y6404 = ~1'b0 ;
  assign y6405 = ~1'b0 ;
  assign y6406 = ~n10934 ;
  assign y6407 = n10935 ;
  assign y6408 = ~1'b0 ;
  assign y6409 = ~n10936 ;
  assign y6410 = ~n9254 ;
  assign y6411 = ~1'b0 ;
  assign y6412 = ~1'b0 ;
  assign y6413 = n10943 ;
  assign y6414 = n10944 ;
  assign y6415 = ~1'b0 ;
  assign y6416 = ~1'b0 ;
  assign y6417 = ~n10947 ;
  assign y6418 = ~n10948 ;
  assign y6419 = ~1'b0 ;
  assign y6420 = ~n10949 ;
  assign y6421 = n10951 ;
  assign y6422 = n10952 ;
  assign y6423 = ~n963 ;
  assign y6424 = ~1'b0 ;
  assign y6425 = n10954 ;
  assign y6426 = n10955 ;
  assign y6427 = n10956 ;
  assign y6428 = ~n10957 ;
  assign y6429 = ~1'b0 ;
  assign y6430 = ~1'b0 ;
  assign y6431 = ~1'b0 ;
  assign y6432 = ~1'b0 ;
  assign y6433 = n10961 ;
  assign y6434 = ~1'b0 ;
  assign y6435 = n5395 ;
  assign y6436 = ~n10967 ;
  assign y6437 = ~n10968 ;
  assign y6438 = ~n10970 ;
  assign y6439 = ~n10971 ;
  assign y6440 = ~1'b0 ;
  assign y6441 = n10972 ;
  assign y6442 = ~n10978 ;
  assign y6443 = 1'b0 ;
  assign y6444 = ~n10980 ;
  assign y6445 = n10985 ;
  assign y6446 = n10986 ;
  assign y6447 = ~n10995 ;
  assign y6448 = ~1'b0 ;
  assign y6449 = n10997 ;
  assign y6450 = n10998 ;
  assign y6451 = n10999 ;
  assign y6452 = n11001 ;
  assign y6453 = ~n11008 ;
  assign y6454 = ~n11009 ;
  assign y6455 = ~n11010 ;
  assign y6456 = ~n11012 ;
  assign y6457 = ~n11016 ;
  assign y6458 = n11017 ;
  assign y6459 = ~n11019 ;
  assign y6460 = 1'b0 ;
  assign y6461 = ~1'b0 ;
  assign y6462 = ~1'b0 ;
  assign y6463 = ~n11021 ;
  assign y6464 = ~n11023 ;
  assign y6465 = ~x15 ;
  assign y6466 = n11025 ;
  assign y6467 = ~1'b0 ;
  assign y6468 = ~1'b0 ;
  assign y6469 = ~n11030 ;
  assign y6470 = ~1'b0 ;
  assign y6471 = ~1'b0 ;
  assign y6472 = 1'b0 ;
  assign y6473 = ~1'b0 ;
  assign y6474 = n11031 ;
  assign y6475 = ~n11034 ;
  assign y6476 = ~n11037 ;
  assign y6477 = ~n11038 ;
  assign y6478 = ~1'b0 ;
  assign y6479 = ~n11040 ;
  assign y6480 = ~n11041 ;
  assign y6481 = ~n806 ;
  assign y6482 = ~n11043 ;
  assign y6483 = n11044 ;
  assign y6484 = ~1'b0 ;
  assign y6485 = 1'b0 ;
  assign y6486 = ~1'b0 ;
  assign y6487 = ~1'b0 ;
  assign y6488 = n11051 ;
  assign y6489 = n7185 ;
  assign y6490 = n11052 ;
  assign y6491 = n11053 ;
  assign y6492 = ~1'b0 ;
  assign y6493 = ~n11054 ;
  assign y6494 = ~n11066 ;
  assign y6495 = ~1'b0 ;
  assign y6496 = n11067 ;
  assign y6497 = ~1'b0 ;
  assign y6498 = ~1'b0 ;
  assign y6499 = ~1'b0 ;
  assign y6500 = 1'b0 ;
  assign y6501 = n5783 ;
  assign y6502 = n11068 ;
  assign y6503 = ~1'b0 ;
  assign y6504 = ~n11069 ;
  assign y6505 = ~n11070 ;
  assign y6506 = n11071 ;
  assign y6507 = ~n11073 ;
  assign y6508 = ~1'b0 ;
  assign y6509 = ~1'b0 ;
  assign y6510 = n11077 ;
  assign y6511 = n11084 ;
  assign y6512 = n11085 ;
  assign y6513 = ~1'b0 ;
  assign y6514 = ~n11088 ;
  assign y6515 = ~1'b0 ;
  assign y6516 = ~1'b0 ;
  assign y6517 = n3278 ;
  assign y6518 = n11091 ;
  assign y6519 = ~1'b0 ;
  assign y6520 = ~1'b0 ;
  assign y6521 = ~1'b0 ;
  assign y6522 = n11096 ;
  assign y6523 = ~1'b0 ;
  assign y6524 = ~1'b0 ;
  assign y6525 = ~1'b0 ;
  assign y6526 = n11099 ;
  assign y6527 = ~n11100 ;
  assign y6528 = n1916 ;
  assign y6529 = ~n11102 ;
  assign y6530 = ~1'b0 ;
  assign y6531 = n11106 ;
  assign y6532 = n11107 ;
  assign y6533 = ~1'b0 ;
  assign y6534 = ~n1169 ;
  assign y6535 = ~n11108 ;
  assign y6536 = n11110 ;
  assign y6537 = ~1'b0 ;
  assign y6538 = ~1'b0 ;
  assign y6539 = ~n11114 ;
  assign y6540 = n11115 ;
  assign y6541 = ~n11118 ;
  assign y6542 = ~1'b0 ;
  assign y6543 = ~n11119 ;
  assign y6544 = ~n11121 ;
  assign y6545 = ~n11122 ;
  assign y6546 = n11123 ;
  assign y6547 = ~n11127 ;
  assign y6548 = ~1'b0 ;
  assign y6549 = n11128 ;
  assign y6550 = ~n11131 ;
  assign y6551 = ~n11134 ;
  assign y6552 = ~n11139 ;
  assign y6553 = ~1'b0 ;
  assign y6554 = ~n11141 ;
  assign y6555 = n11142 ;
  assign y6556 = ~n11146 ;
  assign y6557 = ~1'b0 ;
  assign y6558 = n11149 ;
  assign y6559 = ~1'b0 ;
  assign y6560 = ~n11150 ;
  assign y6561 = ~n11153 ;
  assign y6562 = n11156 ;
  assign y6563 = ~1'b0 ;
  assign y6564 = n11157 ;
  assign y6565 = ~1'b0 ;
  assign y6566 = ~1'b0 ;
  assign y6567 = ~1'b0 ;
  assign y6568 = n11158 ;
  assign y6569 = ~1'b0 ;
  assign y6570 = n11161 ;
  assign y6571 = 1'b0 ;
  assign y6572 = ~1'b0 ;
  assign y6573 = ~n11165 ;
  assign y6574 = ~1'b0 ;
  assign y6575 = n11166 ;
  assign y6576 = n11168 ;
  assign y6577 = ~n11170 ;
  assign y6578 = n11173 ;
  assign y6579 = ~1'b0 ;
  assign y6580 = ~1'b0 ;
  assign y6581 = ~n11174 ;
  assign y6582 = n808 ;
  assign y6583 = n11175 ;
  assign y6584 = ~n11178 ;
  assign y6585 = ~n11181 ;
  assign y6586 = ~1'b0 ;
  assign y6587 = n11183 ;
  assign y6588 = n11185 ;
  assign y6589 = ~1'b0 ;
  assign y6590 = n11190 ;
  assign y6591 = ~1'b0 ;
  assign y6592 = x0 ;
  assign y6593 = ~1'b0 ;
  assign y6594 = ~n11193 ;
  assign y6595 = ~n11197 ;
  assign y6596 = ~1'b0 ;
  assign y6597 = n11198 ;
  assign y6598 = ~n11202 ;
  assign y6599 = n2602 ;
  assign y6600 = ~n11205 ;
  assign y6601 = ~1'b0 ;
  assign y6602 = n11207 ;
  assign y6603 = ~n11208 ;
  assign y6604 = ~n5855 ;
  assign y6605 = n3667 ;
  assign y6606 = ~n11209 ;
  assign y6607 = ~n11210 ;
  assign y6608 = n10675 ;
  assign y6609 = ~n11212 ;
  assign y6610 = n11222 ;
  assign y6611 = ~n11223 ;
  assign y6612 = ~1'b0 ;
  assign y6613 = ~1'b0 ;
  assign y6614 = ~1'b0 ;
  assign y6615 = n11226 ;
  assign y6616 = ~1'b0 ;
  assign y6617 = ~n11233 ;
  assign y6618 = n4731 ;
  assign y6619 = ~1'b0 ;
  assign y6620 = ~n1812 ;
  assign y6621 = n11236 ;
  assign y6622 = ~n11237 ;
  assign y6623 = ~n2602 ;
  assign y6624 = ~1'b0 ;
  assign y6625 = ~n11241 ;
  assign y6626 = ~1'b0 ;
  assign y6627 = n11243 ;
  assign y6628 = n11244 ;
  assign y6629 = ~n11247 ;
  assign y6630 = n11248 ;
  assign y6631 = 1'b0 ;
  assign y6632 = n7365 ;
  assign y6633 = ~1'b0 ;
  assign y6634 = 1'b0 ;
  assign y6635 = n11254 ;
  assign y6636 = n11259 ;
  assign y6637 = n11260 ;
  assign y6638 = ~1'b0 ;
  assign y6639 = ~1'b0 ;
  assign y6640 = n11266 ;
  assign y6641 = ~1'b0 ;
  assign y6642 = n11268 ;
  assign y6643 = ~n11271 ;
  assign y6644 = ~1'b0 ;
  assign y6645 = n11273 ;
  assign y6646 = n11275 ;
  assign y6647 = n879 ;
  assign y6648 = ~n11279 ;
  assign y6649 = ~1'b0 ;
  assign y6650 = ~n11280 ;
  assign y6651 = ~1'b0 ;
  assign y6652 = ~1'b0 ;
  assign y6653 = ~1'b0 ;
  assign y6654 = ~1'b0 ;
  assign y6655 = ~n11283 ;
  assign y6656 = ~n11284 ;
  assign y6657 = n11286 ;
  assign y6658 = n11290 ;
  assign y6659 = n11291 ;
  assign y6660 = ~1'b0 ;
  assign y6661 = n11296 ;
  assign y6662 = n11298 ;
  assign y6663 = ~n11300 ;
  assign y6664 = ~1'b0 ;
  assign y6665 = n11303 ;
  assign y6666 = n11305 ;
  assign y6667 = ~n11307 ;
  assign y6668 = n11312 ;
  assign y6669 = ~1'b0 ;
  assign y6670 = n11314 ;
  assign y6671 = 1'b0 ;
  assign y6672 = ~n11315 ;
  assign y6673 = ~n4911 ;
  assign y6674 = ~n11316 ;
  assign y6675 = n693 ;
  assign y6676 = ~n4326 ;
  assign y6677 = ~n11319 ;
  assign y6678 = n11324 ;
  assign y6679 = n11325 ;
  assign y6680 = n11327 ;
  assign y6681 = ~1'b0 ;
  assign y6682 = ~1'b0 ;
  assign y6683 = ~1'b0 ;
  assign y6684 = ~n11331 ;
  assign y6685 = ~n11332 ;
  assign y6686 = ~n2839 ;
  assign y6687 = ~n11339 ;
  assign y6688 = ~n11341 ;
  assign y6689 = ~n11342 ;
  assign y6690 = ~n11346 ;
  assign y6691 = ~n11347 ;
  assign y6692 = ~1'b0 ;
  assign y6693 = ~n408 ;
  assign y6694 = n8838 ;
  assign y6695 = n11349 ;
  assign y6696 = ~1'b0 ;
  assign y6697 = 1'b0 ;
  assign y6698 = ~n11351 ;
  assign y6699 = ~1'b0 ;
  assign y6700 = ~n11354 ;
  assign y6701 = ~n11355 ;
  assign y6702 = n11356 ;
  assign y6703 = ~1'b0 ;
  assign y6704 = n11357 ;
  assign y6705 = ~n11358 ;
  assign y6706 = n11360 ;
  assign y6707 = ~n11362 ;
  assign y6708 = ~1'b0 ;
  assign y6709 = ~1'b0 ;
  assign y6710 = ~1'b0 ;
  assign y6711 = ~n11363 ;
  assign y6712 = ~n5839 ;
  assign y6713 = n11367 ;
  assign y6714 = ~1'b0 ;
  assign y6715 = ~n5960 ;
  assign y6716 = 1'b0 ;
  assign y6717 = ~n11368 ;
  assign y6718 = ~1'b0 ;
  assign y6719 = n11369 ;
  assign y6720 = n11372 ;
  assign y6721 = ~n11373 ;
  assign y6722 = ~n11374 ;
  assign y6723 = ~n11375 ;
  assign y6724 = ~1'b0 ;
  assign y6725 = n11378 ;
  assign y6726 = x13 ;
  assign y6727 = ~n11384 ;
  assign y6728 = n5613 ;
  assign y6729 = ~n11385 ;
  assign y6730 = n7986 ;
  assign y6731 = n11389 ;
  assign y6732 = n3872 ;
  assign y6733 = ~1'b0 ;
  assign y6734 = ~n11391 ;
  assign y6735 = ~n11392 ;
  assign y6736 = n11393 ;
  assign y6737 = n11396 ;
  assign y6738 = n11400 ;
  assign y6739 = ~n11404 ;
  assign y6740 = n11406 ;
  assign y6741 = ~n11409 ;
  assign y6742 = ~n11412 ;
  assign y6743 = n11415 ;
  assign y6744 = ~n11418 ;
  assign y6745 = n11432 ;
  assign y6746 = ~1'b0 ;
  assign y6747 = ~n11435 ;
  assign y6748 = ~n11436 ;
  assign y6749 = ~1'b0 ;
  assign y6750 = ~1'b0 ;
  assign y6751 = n2592 ;
  assign y6752 = ~1'b0 ;
  assign y6753 = n11437 ;
  assign y6754 = n11438 ;
  assign y6755 = ~n11440 ;
  assign y6756 = n11444 ;
  assign y6757 = ~n11446 ;
  assign y6758 = ~n11458 ;
  assign y6759 = ~n11461 ;
  assign y6760 = ~n11466 ;
  assign y6761 = n11468 ;
  assign y6762 = ~1'b0 ;
  assign y6763 = ~n11469 ;
  assign y6764 = ~1'b0 ;
  assign y6765 = ~1'b0 ;
  assign y6766 = ~1'b0 ;
  assign y6767 = ~n11471 ;
  assign y6768 = n11472 ;
  assign y6769 = ~1'b0 ;
  assign y6770 = ~n5802 ;
  assign y6771 = n11482 ;
  assign y6772 = n11489 ;
  assign y6773 = ~n11491 ;
  assign y6774 = n11498 ;
  assign y6775 = ~1'b0 ;
  assign y6776 = ~n11501 ;
  assign y6777 = ~1'b0 ;
  assign y6778 = ~n11503 ;
  assign y6779 = n11507 ;
  assign y6780 = ~1'b0 ;
  assign y6781 = ~n11508 ;
  assign y6782 = x72 ;
  assign y6783 = ~n11511 ;
  assign y6784 = n11513 ;
  assign y6785 = ~1'b0 ;
  assign y6786 = ~n11517 ;
  assign y6787 = n11519 ;
  assign y6788 = n11520 ;
  assign y6789 = n11522 ;
  assign y6790 = ~n11523 ;
  assign y6791 = n11537 ;
  assign y6792 = 1'b0 ;
  assign y6793 = ~n11539 ;
  assign y6794 = ~n11541 ;
  assign y6795 = ~1'b0 ;
  assign y6796 = n11542 ;
  assign y6797 = ~n11543 ;
  assign y6798 = ~n11546 ;
  assign y6799 = ~n11547 ;
  assign y6800 = ~n11548 ;
  assign y6801 = n4098 ;
  assign y6802 = ~1'b0 ;
  assign y6803 = n11550 ;
  assign y6804 = ~1'b0 ;
  assign y6805 = n8005 ;
  assign y6806 = ~n11553 ;
  assign y6807 = ~n11556 ;
  assign y6808 = ~1'b0 ;
  assign y6809 = ~n11557 ;
  assign y6810 = ~n11559 ;
  assign y6811 = 1'b0 ;
  assign y6812 = n11560 ;
  assign y6813 = ~1'b0 ;
  assign y6814 = ~1'b0 ;
  assign y6815 = ~1'b0 ;
  assign y6816 = ~1'b0 ;
  assign y6817 = n11561 ;
  assign y6818 = ~n5014 ;
  assign y6819 = ~n11564 ;
  assign y6820 = n3078 ;
  assign y6821 = ~n3324 ;
  assign y6822 = ~n11566 ;
  assign y6823 = n2709 ;
  assign y6824 = n11570 ;
  assign y6825 = ~n11576 ;
  assign y6826 = 1'b0 ;
  assign y6827 = n11577 ;
  assign y6828 = n11580 ;
  assign y6829 = ~1'b0 ;
  assign y6830 = ~1'b0 ;
  assign y6831 = n11582 ;
  assign y6832 = ~n11584 ;
  assign y6833 = ~1'b0 ;
  assign y6834 = ~n11586 ;
  assign y6835 = n11587 ;
  assign y6836 = ~1'b0 ;
  assign y6837 = ~n11588 ;
  assign y6838 = ~n11589 ;
  assign y6839 = n11590 ;
  assign y6840 = ~n11598 ;
  assign y6841 = ~1'b0 ;
  assign y6842 = n11599 ;
  assign y6843 = n11603 ;
  assign y6844 = n11605 ;
  assign y6845 = n11608 ;
  assign y6846 = n11609 ;
  assign y6847 = ~n11614 ;
  assign y6848 = ~1'b0 ;
  assign y6849 = 1'b0 ;
  assign y6850 = ~1'b0 ;
  assign y6851 = ~n11615 ;
  assign y6852 = 1'b0 ;
  assign y6853 = ~n11616 ;
  assign y6854 = n11622 ;
  assign y6855 = n11626 ;
  assign y6856 = ~n11628 ;
  assign y6857 = ~n11630 ;
  assign y6858 = n11634 ;
  assign y6859 = n11635 ;
  assign y6860 = ~n11636 ;
  assign y6861 = n11637 ;
  assign y6862 = ~1'b0 ;
  assign y6863 = n11652 ;
  assign y6864 = ~1'b0 ;
  assign y6865 = ~n11653 ;
  assign y6866 = ~n11654 ;
  assign y6867 = ~n11661 ;
  assign y6868 = n11663 ;
  assign y6869 = ~1'b0 ;
  assign y6870 = ~1'b0 ;
  assign y6871 = ~1'b0 ;
  assign y6872 = n11668 ;
  assign y6873 = n11669 ;
  assign y6874 = n11673 ;
  assign y6875 = ~n11674 ;
  assign y6876 = ~1'b0 ;
  assign y6877 = n11678 ;
  assign y6878 = ~1'b0 ;
  assign y6879 = ~n11683 ;
  assign y6880 = ~1'b0 ;
  assign y6881 = n11684 ;
  assign y6882 = ~n11686 ;
  assign y6883 = 1'b0 ;
  assign y6884 = ~n11691 ;
  assign y6885 = n11696 ;
  assign y6886 = ~1'b0 ;
  assign y6887 = n134 ;
  assign y6888 = 1'b0 ;
  assign y6889 = ~1'b0 ;
  assign y6890 = n11698 ;
  assign y6891 = ~n11700 ;
  assign y6892 = n11701 ;
  assign y6893 = ~1'b0 ;
  assign y6894 = ~n11703 ;
  assign y6895 = ~n11704 ;
  assign y6896 = n11705 ;
  assign y6897 = ~n11707 ;
  assign y6898 = n11711 ;
  assign y6899 = ~n11712 ;
  assign y6900 = n11713 ;
  assign y6901 = n11715 ;
  assign y6902 = n11717 ;
  assign y6903 = ~1'b0 ;
  assign y6904 = ~n11720 ;
  assign y6905 = n11723 ;
  assign y6906 = ~n11726 ;
  assign y6907 = n3483 ;
  assign y6908 = n7476 ;
  assign y6909 = ~n11731 ;
  assign y6910 = ~n6644 ;
  assign y6911 = ~n11732 ;
  assign y6912 = n11733 ;
  assign y6913 = ~n11737 ;
  assign y6914 = ~1'b0 ;
  assign y6915 = ~1'b0 ;
  assign y6916 = ~1'b0 ;
  assign y6917 = ~1'b0 ;
  assign y6918 = ~n11739 ;
  assign y6919 = ~1'b0 ;
  assign y6920 = n11740 ;
  assign y6921 = ~1'b0 ;
  assign y6922 = ~n11741 ;
  assign y6923 = ~n11743 ;
  assign y6924 = 1'b0 ;
  assign y6925 = n11744 ;
  assign y6926 = ~1'b0 ;
  assign y6927 = ~n11746 ;
  assign y6928 = n11750 ;
  assign y6929 = ~n11756 ;
  assign y6930 = ~n11758 ;
  assign y6931 = ~n11759 ;
  assign y6932 = ~1'b0 ;
  assign y6933 = ~n11761 ;
  assign y6934 = ~1'b0 ;
  assign y6935 = ~n8441 ;
  assign y6936 = ~n11762 ;
  assign y6937 = n11763 ;
  assign y6938 = ~1'b0 ;
  assign y6939 = ~n11767 ;
  assign y6940 = ~n11770 ;
  assign y6941 = ~n11771 ;
  assign y6942 = n11774 ;
  assign y6943 = ~1'b0 ;
  assign y6944 = ~1'b0 ;
  assign y6945 = ~n11775 ;
  assign y6946 = n11777 ;
  assign y6947 = ~1'b0 ;
  assign y6948 = ~n11778 ;
  assign y6949 = n11779 ;
  assign y6950 = ~n11780 ;
  assign y6951 = ~n11782 ;
  assign y6952 = n8363 ;
  assign y6953 = n11784 ;
  assign y6954 = ~1'b0 ;
  assign y6955 = ~1'b0 ;
  assign y6956 = n11786 ;
  assign y6957 = n7804 ;
  assign y6958 = ~n11788 ;
  assign y6959 = ~n11790 ;
  assign y6960 = ~n11792 ;
  assign y6961 = ~n11794 ;
  assign y6962 = ~n11795 ;
  assign y6963 = n11797 ;
  assign y6964 = ~1'b0 ;
  assign y6965 = ~1'b0 ;
  assign y6966 = n11798 ;
  assign y6967 = ~n11799 ;
  assign y6968 = n11802 ;
  assign y6969 = n11804 ;
  assign y6970 = ~1'b0 ;
  assign y6971 = ~1'b0 ;
  assign y6972 = ~1'b0 ;
  assign y6973 = ~1'b0 ;
  assign y6974 = n11807 ;
  assign y6975 = ~1'b0 ;
  assign y6976 = n11809 ;
  assign y6977 = ~1'b0 ;
  assign y6978 = ~1'b0 ;
  assign y6979 = ~1'b0 ;
  assign y6980 = ~n11810 ;
  assign y6981 = ~n11811 ;
  assign y6982 = ~1'b0 ;
  assign y6983 = ~n11813 ;
  assign y6984 = ~1'b0 ;
  assign y6985 = ~n7435 ;
  assign y6986 = n1010 ;
  assign y6987 = ~n11814 ;
  assign y6988 = ~1'b0 ;
  assign y6989 = ~n11815 ;
  assign y6990 = ~1'b0 ;
  assign y6991 = n11816 ;
  assign y6992 = ~1'b0 ;
  assign y6993 = ~1'b0 ;
  assign y6994 = ~1'b0 ;
  assign y6995 = n11818 ;
  assign y6996 = ~n11819 ;
  assign y6997 = n11823 ;
  assign y6998 = ~1'b0 ;
  assign y6999 = ~1'b0 ;
  assign y7000 = ~n11824 ;
  assign y7001 = n11828 ;
  assign y7002 = ~1'b0 ;
  assign y7003 = ~1'b0 ;
  assign y7004 = 1'b0 ;
  assign y7005 = ~1'b0 ;
  assign y7006 = n11829 ;
  assign y7007 = n809 ;
  assign y7008 = ~1'b0 ;
  assign y7009 = ~n11831 ;
  assign y7010 = ~n1724 ;
  assign y7011 = ~1'b0 ;
  assign y7012 = ~1'b0 ;
  assign y7013 = n11833 ;
  assign y7014 = ~n11836 ;
  assign y7015 = n11124 ;
  assign y7016 = ~n11837 ;
  assign y7017 = ~1'b0 ;
  assign y7018 = ~1'b0 ;
  assign y7019 = n11840 ;
  assign y7020 = ~1'b0 ;
  assign y7021 = n11843 ;
  assign y7022 = n11844 ;
  assign y7023 = ~1'b0 ;
  assign y7024 = ~n882 ;
  assign y7025 = ~1'b0 ;
  assign y7026 = n11848 ;
  assign y7027 = n3064 ;
  assign y7028 = ~n11851 ;
  assign y7029 = ~1'b0 ;
  assign y7030 = ~n3426 ;
  assign y7031 = n11854 ;
  assign y7032 = ~n11857 ;
  assign y7033 = n11858 ;
  assign y7034 = ~n9285 ;
  assign y7035 = ~n11861 ;
  assign y7036 = ~1'b0 ;
  assign y7037 = n11862 ;
  assign y7038 = ~1'b0 ;
  assign y7039 = n11863 ;
  assign y7040 = n11864 ;
  assign y7041 = n11865 ;
  assign y7042 = ~1'b0 ;
  assign y7043 = n11866 ;
  assign y7044 = n11868 ;
  assign y7045 = ~1'b0 ;
  assign y7046 = n3795 ;
  assign y7047 = n11877 ;
  assign y7048 = ~1'b0 ;
  assign y7049 = ~1'b0 ;
  assign y7050 = ~n11880 ;
  assign y7051 = n11881 ;
  assign y7052 = n9490 ;
  assign y7053 = n8244 ;
  assign y7054 = n11882 ;
  assign y7055 = ~1'b0 ;
  assign y7056 = 1'b0 ;
  assign y7057 = n11885 ;
  assign y7058 = ~1'b0 ;
  assign y7059 = ~1'b0 ;
  assign y7060 = n7454 ;
  assign y7061 = n11887 ;
  assign y7062 = ~1'b0 ;
  assign y7063 = n11894 ;
  assign y7064 = n11896 ;
  assign y7065 = n11898 ;
  assign y7066 = ~n10453 ;
  assign y7067 = ~1'b0 ;
  assign y7068 = ~1'b0 ;
  assign y7069 = ~1'b0 ;
  assign y7070 = n11900 ;
  assign y7071 = ~1'b0 ;
  assign y7072 = n11902 ;
  assign y7073 = ~n11904 ;
  assign y7074 = ~1'b0 ;
  assign y7075 = ~1'b0 ;
  assign y7076 = n11906 ;
  assign y7077 = ~1'b0 ;
  assign y7078 = n11909 ;
  assign y7079 = ~n6144 ;
  assign y7080 = ~1'b0 ;
  assign y7081 = ~1'b0 ;
  assign y7082 = ~n7364 ;
  assign y7083 = n11913 ;
  assign y7084 = x73 ;
  assign y7085 = 1'b0 ;
  assign y7086 = n11914 ;
  assign y7087 = n11917 ;
  assign y7088 = n11918 ;
  assign y7089 = 1'b0 ;
  assign y7090 = ~1'b0 ;
  assign y7091 = n11920 ;
  assign y7092 = ~1'b0 ;
  assign y7093 = ~n11921 ;
  assign y7094 = ~1'b0 ;
  assign y7095 = ~n11922 ;
  assign y7096 = ~1'b0 ;
  assign y7097 = ~1'b0 ;
  assign y7098 = ~n11925 ;
  assign y7099 = ~1'b0 ;
  assign y7100 = 1'b0 ;
  assign y7101 = ~1'b0 ;
  assign y7102 = ~n11928 ;
  assign y7103 = n11931 ;
  assign y7104 = n11933 ;
  assign y7105 = ~n11936 ;
  assign y7106 = ~n11938 ;
  assign y7107 = ~n11941 ;
  assign y7108 = n11943 ;
  assign y7109 = n11947 ;
  assign y7110 = ~n11948 ;
  assign y7111 = ~n11952 ;
  assign y7112 = ~1'b0 ;
  assign y7113 = n11959 ;
  assign y7114 = ~1'b0 ;
  assign y7115 = ~1'b0 ;
  assign y7116 = n5448 ;
  assign y7117 = n11960 ;
  assign y7118 = ~1'b0 ;
  assign y7119 = ~1'b0 ;
  assign y7120 = ~1'b0 ;
  assign y7121 = ~1'b0 ;
  assign y7122 = ~1'b0 ;
  assign y7123 = n11961 ;
  assign y7124 = ~n11962 ;
  assign y7125 = ~1'b0 ;
  assign y7126 = ~n1402 ;
  assign y7127 = ~1'b0 ;
  assign y7128 = ~n11964 ;
  assign y7129 = ~n11965 ;
  assign y7130 = ~1'b0 ;
  assign y7131 = n11967 ;
  assign y7132 = ~1'b0 ;
  assign y7133 = ~n11968 ;
  assign y7134 = ~1'b0 ;
  assign y7135 = ~n11972 ;
  assign y7136 = n11974 ;
  assign y7137 = ~n11977 ;
  assign y7138 = n11978 ;
  assign y7139 = ~n11979 ;
  assign y7140 = ~n11984 ;
  assign y7141 = ~n4366 ;
  assign y7142 = 1'b0 ;
  assign y7143 = ~1'b0 ;
  assign y7144 = 1'b0 ;
  assign y7145 = ~1'b0 ;
  assign y7146 = ~1'b0 ;
  assign y7147 = ~1'b0 ;
  assign y7148 = ~1'b0 ;
  assign y7149 = n11987 ;
  assign y7150 = n4954 ;
  assign y7151 = ~1'b0 ;
  assign y7152 = ~n11988 ;
  assign y7153 = ~1'b0 ;
  assign y7154 = n11990 ;
  assign y7155 = ~n1212 ;
  assign y7156 = n11992 ;
  assign y7157 = ~1'b0 ;
  assign y7158 = n11996 ;
  assign y7159 = ~n11999 ;
  assign y7160 = ~n12001 ;
  assign y7161 = ~n12003 ;
  assign y7162 = n5685 ;
  assign y7163 = ~1'b0 ;
  assign y7164 = ~n12004 ;
  assign y7165 = ~n12006 ;
  assign y7166 = n12007 ;
  assign y7167 = ~1'b0 ;
  assign y7168 = n12010 ;
  assign y7169 = n12011 ;
  assign y7170 = n890 ;
  assign y7171 = ~1'b0 ;
  assign y7172 = ~n12013 ;
  assign y7173 = ~n2775 ;
  assign y7174 = ~n12014 ;
  assign y7175 = n12017 ;
  assign y7176 = ~1'b0 ;
  assign y7177 = ~n4697 ;
  assign y7178 = ~1'b0 ;
  assign y7179 = ~n12020 ;
  assign y7180 = n10548 ;
  assign y7181 = ~n12021 ;
  assign y7182 = ~n12023 ;
  assign y7183 = ~1'b0 ;
  assign y7184 = ~n12029 ;
  assign y7185 = ~1'b0 ;
  assign y7186 = 1'b0 ;
  assign y7187 = n12032 ;
  assign y7188 = ~n12033 ;
  assign y7189 = 1'b0 ;
  assign y7190 = ~n12040 ;
  assign y7191 = n12043 ;
  assign y7192 = ~1'b0 ;
  assign y7193 = n12044 ;
  assign y7194 = ~1'b0 ;
  assign y7195 = ~n12050 ;
  assign y7196 = ~1'b0 ;
  assign y7197 = n12057 ;
  assign y7198 = ~n12060 ;
  assign y7199 = ~n12063 ;
  assign y7200 = ~1'b0 ;
  assign y7201 = n12064 ;
  assign y7202 = n12066 ;
  assign y7203 = 1'b0 ;
  assign y7204 = n12071 ;
  assign y7205 = ~n12072 ;
  assign y7206 = ~n1867 ;
  assign y7207 = ~1'b0 ;
  assign y7208 = n12073 ;
  assign y7209 = n12076 ;
  assign y7210 = n12082 ;
  assign y7211 = ~1'b0 ;
  assign y7212 = ~1'b0 ;
  assign y7213 = ~n7799 ;
  assign y7214 = n8511 ;
  assign y7215 = ~1'b0 ;
  assign y7216 = n12084 ;
  assign y7217 = ~n12088 ;
  assign y7218 = ~1'b0 ;
  assign y7219 = 1'b0 ;
  assign y7220 = ~1'b0 ;
  assign y7221 = n12093 ;
  assign y7222 = n12095 ;
  assign y7223 = ~1'b0 ;
  assign y7224 = ~n12098 ;
  assign y7225 = ~n12100 ;
  assign y7226 = ~n12101 ;
  assign y7227 = ~1'b0 ;
  assign y7228 = ~n12104 ;
  assign y7229 = ~1'b0 ;
  assign y7230 = ~1'b0 ;
  assign y7231 = ~n272 ;
  assign y7232 = ~n12108 ;
  assign y7233 = ~1'b0 ;
  assign y7234 = ~n12115 ;
  assign y7235 = ~n12117 ;
  assign y7236 = ~1'b0 ;
  assign y7237 = 1'b0 ;
  assign y7238 = ~1'b0 ;
  assign y7239 = ~n12118 ;
  assign y7240 = ~n12122 ;
  assign y7241 = ~1'b0 ;
  assign y7242 = n12124 ;
  assign y7243 = ~1'b0 ;
  assign y7244 = n12125 ;
  assign y7245 = 1'b0 ;
  assign y7246 = ~n12128 ;
  assign y7247 = ~n12132 ;
  assign y7248 = ~1'b0 ;
  assign y7249 = n2040 ;
  assign y7250 = ~n3041 ;
  assign y7251 = ~n12134 ;
  assign y7252 = ~n12138 ;
  assign y7253 = ~1'b0 ;
  assign y7254 = ~1'b0 ;
  assign y7255 = ~n1579 ;
  assign y7256 = n12139 ;
  assign y7257 = ~n2936 ;
  assign y7258 = ~n12140 ;
  assign y7259 = n12142 ;
  assign y7260 = n6436 ;
  assign y7261 = ~n12145 ;
  assign y7262 = ~n12147 ;
  assign y7263 = n12148 ;
  assign y7264 = ~1'b0 ;
  assign y7265 = ~1'b0 ;
  assign y7266 = n12149 ;
  assign y7267 = ~n12151 ;
  assign y7268 = n11164 ;
  assign y7269 = ~1'b0 ;
  assign y7270 = ~n12156 ;
  assign y7271 = n11051 ;
  assign y7272 = ~1'b0 ;
  assign y7273 = ~n12157 ;
  assign y7274 = ~n12159 ;
  assign y7275 = ~1'b0 ;
  assign y7276 = ~1'b0 ;
  assign y7277 = ~n6735 ;
  assign y7278 = n10443 ;
  assign y7279 = ~n8322 ;
  assign y7280 = n12161 ;
  assign y7281 = ~n12164 ;
  assign y7282 = n12166 ;
  assign y7283 = n12171 ;
  assign y7284 = ~1'b0 ;
  assign y7285 = ~n12174 ;
  assign y7286 = ~n12179 ;
  assign y7287 = ~1'b0 ;
  assign y7288 = n12181 ;
  assign y7289 = 1'b0 ;
  assign y7290 = ~1'b0 ;
  assign y7291 = ~1'b0 ;
  assign y7292 = ~n12182 ;
  assign y7293 = ~n12183 ;
  assign y7294 = n6759 ;
  assign y7295 = ~1'b0 ;
  assign y7296 = ~1'b0 ;
  assign y7297 = n12184 ;
  assign y7298 = n12186 ;
  assign y7299 = n12187 ;
  assign y7300 = ~n10724 ;
  assign y7301 = ~n12189 ;
  assign y7302 = 1'b0 ;
  assign y7303 = ~1'b0 ;
  assign y7304 = 1'b0 ;
  assign y7305 = ~n12191 ;
  assign y7306 = ~n1238 ;
  assign y7307 = ~1'b0 ;
  assign y7308 = ~1'b0 ;
  assign y7309 = ~n5096 ;
  assign y7310 = n998 ;
  assign y7311 = ~1'b0 ;
  assign y7312 = ~n886 ;
  assign y7313 = ~1'b0 ;
  assign y7314 = 1'b0 ;
  assign y7315 = n12194 ;
  assign y7316 = ~1'b0 ;
  assign y7317 = n12195 ;
  assign y7318 = ~1'b0 ;
  assign y7319 = ~n12196 ;
  assign y7320 = ~n12197 ;
  assign y7321 = ~1'b0 ;
  assign y7322 = n12198 ;
  assign y7323 = n12202 ;
  assign y7324 = ~n12206 ;
  assign y7325 = ~1'b0 ;
  assign y7326 = n12209 ;
  assign y7327 = ~1'b0 ;
  assign y7328 = ~n12217 ;
  assign y7329 = n12218 ;
  assign y7330 = ~1'b0 ;
  assign y7331 = ~1'b0 ;
  assign y7332 = n12225 ;
  assign y7333 = ~1'b0 ;
  assign y7334 = n12228 ;
  assign y7335 = n12229 ;
  assign y7336 = ~1'b0 ;
  assign y7337 = n12232 ;
  assign y7338 = ~n12238 ;
  assign y7339 = ~n7169 ;
  assign y7340 = ~1'b0 ;
  assign y7341 = ~1'b0 ;
  assign y7342 = ~n12240 ;
  assign y7343 = ~n12241 ;
  assign y7344 = ~n12247 ;
  assign y7345 = ~n12248 ;
  assign y7346 = ~n12249 ;
  assign y7347 = ~1'b0 ;
  assign y7348 = ~1'b0 ;
  assign y7349 = n12250 ;
  assign y7350 = ~1'b0 ;
  assign y7351 = n12252 ;
  assign y7352 = ~n12257 ;
  assign y7353 = 1'b0 ;
  assign y7354 = ~n12258 ;
  assign y7355 = ~n10172 ;
  assign y7356 = ~n8596 ;
  assign y7357 = ~1'b0 ;
  assign y7358 = ~n12260 ;
  assign y7359 = ~n8535 ;
  assign y7360 = ~1'b0 ;
  assign y7361 = ~1'b0 ;
  assign y7362 = ~n12261 ;
  assign y7363 = ~n12262 ;
  assign y7364 = ~n5068 ;
  assign y7365 = ~n12264 ;
  assign y7366 = ~1'b0 ;
  assign y7367 = n12266 ;
  assign y7368 = n12268 ;
  assign y7369 = ~n12269 ;
  assign y7370 = ~n2271 ;
  assign y7371 = n12272 ;
  assign y7372 = ~n891 ;
  assign y7373 = ~1'b0 ;
  assign y7374 = ~1'b0 ;
  assign y7375 = ~1'b0 ;
  assign y7376 = ~n12277 ;
  assign y7377 = ~1'b0 ;
  assign y7378 = n12279 ;
  assign y7379 = ~n12281 ;
  assign y7380 = n12283 ;
  assign y7381 = n12287 ;
  assign y7382 = ~n12288 ;
  assign y7383 = n12298 ;
  assign y7384 = n12302 ;
  assign y7385 = ~1'b0 ;
  assign y7386 = n12304 ;
  assign y7387 = ~n12306 ;
  assign y7388 = n7944 ;
  assign y7389 = n12309 ;
  assign y7390 = ~1'b0 ;
  assign y7391 = n12312 ;
  assign y7392 = ~1'b0 ;
  assign y7393 = ~n12317 ;
  assign y7394 = ~n12319 ;
  assign y7395 = 1'b0 ;
  assign y7396 = ~n12321 ;
  assign y7397 = n12323 ;
  assign y7398 = ~1'b0 ;
  assign y7399 = ~1'b0 ;
  assign y7400 = ~n12326 ;
  assign y7401 = ~n12327 ;
  assign y7402 = ~1'b0 ;
  assign y7403 = ~1'b0 ;
  assign y7404 = n12336 ;
  assign y7405 = n12337 ;
  assign y7406 = ~n2636 ;
  assign y7407 = n12338 ;
  assign y7408 = ~1'b0 ;
  assign y7409 = ~1'b0 ;
  assign y7410 = ~1'b0 ;
  assign y7411 = n12340 ;
  assign y7412 = n10847 ;
  assign y7413 = 1'b0 ;
  assign y7414 = ~n12342 ;
  assign y7415 = ~1'b0 ;
  assign y7416 = 1'b0 ;
  assign y7417 = n3491 ;
  assign y7418 = ~n12344 ;
  assign y7419 = n12345 ;
  assign y7420 = ~1'b0 ;
  assign y7421 = ~1'b0 ;
  assign y7422 = ~n12346 ;
  assign y7423 = ~1'b0 ;
  assign y7424 = n12347 ;
  assign y7425 = ~n12349 ;
  assign y7426 = ~n12353 ;
  assign y7427 = n12354 ;
  assign y7428 = ~n4259 ;
  assign y7429 = n12355 ;
  assign y7430 = ~1'b0 ;
  assign y7431 = n8725 ;
  assign y7432 = ~1'b0 ;
  assign y7433 = n12357 ;
  assign y7434 = ~n12360 ;
  assign y7435 = ~n12361 ;
  assign y7436 = ~n12363 ;
  assign y7437 = ~n12368 ;
  assign y7438 = ~1'b0 ;
  assign y7439 = ~n12370 ;
  assign y7440 = ~1'b0 ;
  assign y7441 = ~1'b0 ;
  assign y7442 = n12371 ;
  assign y7443 = ~n12372 ;
  assign y7444 = ~1'b0 ;
  assign y7445 = n12375 ;
  assign y7446 = ~1'b0 ;
  assign y7447 = ~1'b0 ;
  assign y7448 = x111 ;
  assign y7449 = ~1'b0 ;
  assign y7450 = ~n12377 ;
  assign y7451 = ~n12380 ;
  assign y7452 = n868 ;
  assign y7453 = n12381 ;
  assign y7454 = ~1'b0 ;
  assign y7455 = ~n4630 ;
  assign y7456 = ~n12387 ;
  assign y7457 = ~n12388 ;
  assign y7458 = ~n12391 ;
  assign y7459 = ~n4560 ;
  assign y7460 = 1'b0 ;
  assign y7461 = n12393 ;
  assign y7462 = ~1'b0 ;
  assign y7463 = ~1'b0 ;
  assign y7464 = ~n6757 ;
  assign y7465 = ~1'b0 ;
  assign y7466 = ~1'b0 ;
  assign y7467 = ~1'b0 ;
  assign y7468 = ~1'b0 ;
  assign y7469 = n12394 ;
  assign y7470 = n12396 ;
  assign y7471 = 1'b0 ;
  assign y7472 = ~n12397 ;
  assign y7473 = ~1'b0 ;
  assign y7474 = ~1'b0 ;
  assign y7475 = n3697 ;
  assign y7476 = ~n12399 ;
  assign y7477 = ~n12400 ;
  assign y7478 = ~1'b0 ;
  assign y7479 = ~n12404 ;
  assign y7480 = ~n9797 ;
  assign y7481 = ~n12405 ;
  assign y7482 = ~1'b0 ;
  assign y7483 = n12406 ;
  assign y7484 = n12407 ;
  assign y7485 = n12411 ;
  assign y7486 = 1'b0 ;
  assign y7487 = ~n12412 ;
  assign y7488 = n12414 ;
  assign y7489 = n12347 ;
  assign y7490 = ~n12416 ;
  assign y7491 = n12417 ;
  assign y7492 = 1'b0 ;
  assign y7493 = ~1'b0 ;
  assign y7494 = ~1'b0 ;
  assign y7495 = ~1'b0 ;
  assign y7496 = n2094 ;
  assign y7497 = ~1'b0 ;
  assign y7498 = n12418 ;
  assign y7499 = ~n12428 ;
  assign y7500 = ~1'b0 ;
  assign y7501 = ~1'b0 ;
  assign y7502 = ~1'b0 ;
  assign y7503 = n424 ;
  assign y7504 = ~n12430 ;
  assign y7505 = 1'b0 ;
  assign y7506 = ~n12433 ;
  assign y7507 = n12434 ;
  assign y7508 = n12436 ;
  assign y7509 = n12439 ;
  assign y7510 = ~1'b0 ;
  assign y7511 = n10840 ;
  assign y7512 = ~n12440 ;
  assign y7513 = n640 ;
  assign y7514 = ~n12442 ;
  assign y7515 = ~1'b0 ;
  assign y7516 = ~1'b0 ;
  assign y7517 = ~1'b0 ;
  assign y7518 = n12443 ;
  assign y7519 = ~n12444 ;
  assign y7520 = n12446 ;
  assign y7521 = ~1'b0 ;
  assign y7522 = ~n12447 ;
  assign y7523 = n8737 ;
  assign y7524 = n12452 ;
  assign y7525 = n12455 ;
  assign y7526 = n12456 ;
  assign y7527 = ~1'b0 ;
  assign y7528 = ~n12457 ;
  assign y7529 = ~n12458 ;
  assign y7530 = n12462 ;
  assign y7531 = ~1'b0 ;
  assign y7532 = n12464 ;
  assign y7533 = n12467 ;
  assign y7534 = n12474 ;
  assign y7535 = ~1'b0 ;
  assign y7536 = ~n12476 ;
  assign y7537 = ~n12477 ;
  assign y7538 = n12482 ;
  assign y7539 = n12484 ;
  assign y7540 = ~1'b0 ;
  assign y7541 = ~1'b0 ;
  assign y7542 = ~1'b0 ;
  assign y7543 = ~1'b0 ;
  assign y7544 = ~1'b0 ;
  assign y7545 = ~n12486 ;
  assign y7546 = n12488 ;
  assign y7547 = ~1'b0 ;
  assign y7548 = ~1'b0 ;
  assign y7549 = ~n12497 ;
  assign y7550 = ~n12499 ;
  assign y7551 = ~n12502 ;
  assign y7552 = ~1'b0 ;
  assign y7553 = ~n12503 ;
  assign y7554 = n12504 ;
  assign y7555 = ~1'b0 ;
  assign y7556 = ~n12512 ;
  assign y7557 = ~1'b0 ;
  assign y7558 = n12513 ;
  assign y7559 = 1'b0 ;
  assign y7560 = n12515 ;
  assign y7561 = n1724 ;
  assign y7562 = ~1'b0 ;
  assign y7563 = ~n12517 ;
  assign y7564 = ~1'b0 ;
  assign y7565 = 1'b0 ;
  assign y7566 = 1'b0 ;
  assign y7567 = n11423 ;
  assign y7568 = n12519 ;
  assign y7569 = ~n12525 ;
  assign y7570 = ~n12527 ;
  assign y7571 = n12529 ;
  assign y7572 = ~n12532 ;
  assign y7573 = n12535 ;
  assign y7574 = 1'b0 ;
  assign y7575 = n12537 ;
  assign y7576 = n616 ;
  assign y7577 = ~1'b0 ;
  assign y7578 = 1'b0 ;
  assign y7579 = ~1'b0 ;
  assign y7580 = n12539 ;
  assign y7581 = ~1'b0 ;
  assign y7582 = n12543 ;
  assign y7583 = n12548 ;
  assign y7584 = ~1'b0 ;
  assign y7585 = 1'b0 ;
  assign y7586 = n12549 ;
  assign y7587 = n12551 ;
  assign y7588 = ~1'b0 ;
  assign y7589 = ~n12553 ;
  assign y7590 = n12556 ;
  assign y7591 = n12564 ;
  assign y7592 = ~1'b0 ;
  assign y7593 = n12566 ;
  assign y7594 = 1'b0 ;
  assign y7595 = ~n12571 ;
  assign y7596 = ~n12572 ;
  assign y7597 = n12573 ;
  assign y7598 = ~n12574 ;
  assign y7599 = ~n12579 ;
  assign y7600 = ~1'b0 ;
  assign y7601 = n12580 ;
  assign y7602 = ~1'b0 ;
  assign y7603 = n12581 ;
  assign y7604 = 1'b0 ;
  assign y7605 = ~n12587 ;
  assign y7606 = ~n12589 ;
  assign y7607 = ~n12590 ;
  assign y7608 = n12597 ;
  assign y7609 = n12599 ;
  assign y7610 = 1'b0 ;
  assign y7611 = 1'b0 ;
  assign y7612 = ~1'b0 ;
  assign y7613 = ~1'b0 ;
  assign y7614 = ~1'b0 ;
  assign y7615 = ~1'b0 ;
  assign y7616 = n12600 ;
  assign y7617 = n12603 ;
  assign y7618 = n12605 ;
  assign y7619 = ~1'b0 ;
  assign y7620 = ~1'b0 ;
  assign y7621 = 1'b0 ;
  assign y7622 = n12611 ;
  assign y7623 = n12614 ;
  assign y7624 = n12617 ;
  assign y7625 = ~1'b0 ;
  assign y7626 = ~1'b0 ;
  assign y7627 = n12619 ;
  assign y7628 = ~1'b0 ;
  assign y7629 = n12621 ;
  assign y7630 = n12622 ;
  assign y7631 = ~1'b0 ;
  assign y7632 = n12624 ;
  assign y7633 = n12633 ;
  assign y7634 = n12634 ;
  assign y7635 = n12635 ;
  assign y7636 = n12637 ;
  assign y7637 = n12639 ;
  assign y7638 = n12643 ;
  assign y7639 = n12644 ;
  assign y7640 = ~n12648 ;
  assign y7641 = n12651 ;
  assign y7642 = ~1'b0 ;
  assign y7643 = n12652 ;
  assign y7644 = ~1'b0 ;
  assign y7645 = ~1'b0 ;
  assign y7646 = ~n9285 ;
  assign y7647 = ~1'b0 ;
  assign y7648 = ~n12654 ;
  assign y7649 = ~1'b0 ;
  assign y7650 = ~1'b0 ;
  assign y7651 = ~1'b0 ;
  assign y7652 = ~n12656 ;
  assign y7653 = n12658 ;
  assign y7654 = n12662 ;
  assign y7655 = n12665 ;
  assign y7656 = ~1'b0 ;
  assign y7657 = n12667 ;
  assign y7658 = ~1'b0 ;
  assign y7659 = ~1'b0 ;
  assign y7660 = ~1'b0 ;
  assign y7661 = ~n12670 ;
  assign y7662 = n12671 ;
  assign y7663 = ~n5455 ;
  assign y7664 = ~1'b0 ;
  assign y7665 = n11203 ;
  assign y7666 = ~1'b0 ;
  assign y7667 = ~1'b0 ;
  assign y7668 = ~n12672 ;
  assign y7669 = n1166 ;
  assign y7670 = n12676 ;
  assign y7671 = ~1'b0 ;
  assign y7672 = n12677 ;
  assign y7673 = n12678 ;
  assign y7674 = n12686 ;
  assign y7675 = n12687 ;
  assign y7676 = ~1'b0 ;
  assign y7677 = ~1'b0 ;
  assign y7678 = n12689 ;
  assign y7679 = ~n12692 ;
  assign y7680 = n12694 ;
  assign y7681 = ~n12699 ;
  assign y7682 = ~1'b0 ;
  assign y7683 = ~1'b0 ;
  assign y7684 = ~n12705 ;
  assign y7685 = ~n12707 ;
  assign y7686 = ~1'b0 ;
  assign y7687 = n12708 ;
  assign y7688 = ~n12710 ;
  assign y7689 = n12712 ;
  assign y7690 = ~1'b0 ;
  assign y7691 = ~n12713 ;
  assign y7692 = n12714 ;
  assign y7693 = ~1'b0 ;
  assign y7694 = ~n1704 ;
  assign y7695 = ~n12716 ;
  assign y7696 = ~n12718 ;
  assign y7697 = n12723 ;
  assign y7698 = n9609 ;
  assign y7699 = n12063 ;
  assign y7700 = ~1'b0 ;
  assign y7701 = n12725 ;
  assign y7702 = n12728 ;
  assign y7703 = ~1'b0 ;
  assign y7704 = ~1'b0 ;
  assign y7705 = ~1'b0 ;
  assign y7706 = ~1'b0 ;
  assign y7707 = n12730 ;
  assign y7708 = ~n12731 ;
  assign y7709 = ~n12733 ;
  assign y7710 = n12738 ;
  assign y7711 = ~1'b0 ;
  assign y7712 = n12740 ;
  assign y7713 = ~n12744 ;
  assign y7714 = ~1'b0 ;
  assign y7715 = n12746 ;
  assign y7716 = ~1'b0 ;
  assign y7717 = ~n12750 ;
  assign y7718 = ~1'b0 ;
  assign y7719 = ~1'b0 ;
  assign y7720 = ~n12753 ;
  assign y7721 = ~1'b0 ;
  assign y7722 = n12756 ;
  assign y7723 = n12759 ;
  assign y7724 = ~1'b0 ;
  assign y7725 = ~n12767 ;
  assign y7726 = n12769 ;
  assign y7727 = ~n12770 ;
  assign y7728 = n12771 ;
  assign y7729 = ~1'b0 ;
  assign y7730 = n12774 ;
  assign y7731 = n12782 ;
  assign y7732 = n12783 ;
  assign y7733 = ~n12784 ;
  assign y7734 = ~n12785 ;
  assign y7735 = ~1'b0 ;
  assign y7736 = n12787 ;
  assign y7737 = ~1'b0 ;
  assign y7738 = ~1'b0 ;
  assign y7739 = ~1'b0 ;
  assign y7740 = ~1'b0 ;
  assign y7741 = ~1'b0 ;
  assign y7742 = ~1'b0 ;
  assign y7743 = ~1'b0 ;
  assign y7744 = ~1'b0 ;
  assign y7745 = ~1'b0 ;
  assign y7746 = ~n12795 ;
  assign y7747 = ~1'b0 ;
  assign y7748 = ~n436 ;
  assign y7749 = ~n518 ;
  assign y7750 = 1'b0 ;
  assign y7751 = n12796 ;
  assign y7752 = 1'b0 ;
  assign y7753 = ~n12797 ;
  assign y7754 = ~n12801 ;
  assign y7755 = ~n12802 ;
  assign y7756 = n12807 ;
  assign y7757 = ~1'b0 ;
  assign y7758 = ~n12809 ;
  assign y7759 = ~n8590 ;
  assign y7760 = ~n3651 ;
  assign y7761 = ~n12810 ;
  assign y7762 = ~1'b0 ;
  assign y7763 = n12812 ;
  assign y7764 = ~n12813 ;
  assign y7765 = n12816 ;
  assign y7766 = n12819 ;
  assign y7767 = ~n12822 ;
  assign y7768 = ~1'b0 ;
  assign y7769 = ~n12823 ;
  assign y7770 = ~n12827 ;
  assign y7771 = ~n1203 ;
  assign y7772 = ~n12832 ;
  assign y7773 = 1'b0 ;
  assign y7774 = ~n12838 ;
  assign y7775 = ~1'b0 ;
  assign y7776 = n12839 ;
  assign y7777 = ~n10067 ;
  assign y7778 = ~1'b0 ;
  assign y7779 = n12843 ;
  assign y7780 = ~1'b0 ;
  assign y7781 = n12846 ;
  assign y7782 = n12850 ;
  assign y7783 = ~n12851 ;
  assign y7784 = ~1'b0 ;
  assign y7785 = ~n12852 ;
  assign y7786 = n12853 ;
  assign y7787 = ~1'b0 ;
  assign y7788 = ~1'b0 ;
  assign y7789 = ~1'b0 ;
  assign y7790 = ~n12857 ;
  assign y7791 = ~n12863 ;
  assign y7792 = n12864 ;
  assign y7793 = n12865 ;
  assign y7794 = n12869 ;
  assign y7795 = ~1'b0 ;
  assign y7796 = ~1'b0 ;
  assign y7797 = ~n12870 ;
  assign y7798 = n1629 ;
  assign y7799 = n12871 ;
  assign y7800 = ~n12873 ;
  assign y7801 = n12874 ;
  assign y7802 = ~n12877 ;
  assign y7803 = n12880 ;
  assign y7804 = n12884 ;
  assign y7805 = n3064 ;
  assign y7806 = n12743 ;
  assign y7807 = ~1'b0 ;
  assign y7808 = n12886 ;
  assign y7809 = n12889 ;
  assign y7810 = 1'b0 ;
  assign y7811 = ~1'b0 ;
  assign y7812 = ~n12890 ;
  assign y7813 = ~n12891 ;
  assign y7814 = ~1'b0 ;
  assign y7815 = ~n12895 ;
  assign y7816 = ~n12897 ;
  assign y7817 = 1'b0 ;
  assign y7818 = ~n2981 ;
  assign y7819 = n12900 ;
  assign y7820 = ~n12901 ;
  assign y7821 = n12903 ;
  assign y7822 = ~n12904 ;
  assign y7823 = ~n12907 ;
  assign y7824 = ~n12910 ;
  assign y7825 = ~1'b0 ;
  assign y7826 = ~1'b0 ;
  assign y7827 = n12911 ;
  assign y7828 = n12915 ;
  assign y7829 = ~1'b0 ;
  assign y7830 = ~1'b0 ;
  assign y7831 = ~n12918 ;
  assign y7832 = ~n12927 ;
  assign y7833 = n2325 ;
  assign y7834 = ~1'b0 ;
  assign y7835 = ~1'b0 ;
  assign y7836 = ~1'b0 ;
  assign y7837 = ~1'b0 ;
  assign y7838 = n12928 ;
  assign y7839 = ~1'b0 ;
  assign y7840 = ~1'b0 ;
  assign y7841 = ~1'b0 ;
  assign y7842 = n12929 ;
  assign y7843 = n10866 ;
  assign y7844 = ~1'b0 ;
  assign y7845 = ~n12930 ;
  assign y7846 = n12932 ;
  assign y7847 = n12935 ;
  assign y7848 = n12936 ;
  assign y7849 = ~n12940 ;
  assign y7850 = 1'b0 ;
  assign y7851 = ~n12942 ;
  assign y7852 = ~n1432 ;
  assign y7853 = n12944 ;
  assign y7854 = n10317 ;
  assign y7855 = n12951 ;
  assign y7856 = ~1'b0 ;
  assign y7857 = ~1'b0 ;
  assign y7858 = ~1'b0 ;
  assign y7859 = ~n12952 ;
  assign y7860 = ~1'b0 ;
  assign y7861 = n12956 ;
  assign y7862 = n12958 ;
  assign y7863 = ~n12962 ;
  assign y7864 = ~1'b0 ;
  assign y7865 = ~n12966 ;
  assign y7866 = ~n12968 ;
  assign y7867 = n12974 ;
  assign y7868 = n12975 ;
  assign y7869 = n12976 ;
  assign y7870 = ~1'b0 ;
  assign y7871 = n12978 ;
  assign y7872 = ~1'b0 ;
  assign y7873 = n12980 ;
  assign y7874 = ~n12982 ;
  assign y7875 = n12983 ;
  assign y7876 = ~1'b0 ;
  assign y7877 = ~n12987 ;
  assign y7878 = n12989 ;
  assign y7879 = ~n12990 ;
  assign y7880 = ~n12992 ;
  assign y7881 = ~1'b0 ;
  assign y7882 = ~1'b0 ;
  assign y7883 = n12993 ;
  assign y7884 = n12994 ;
  assign y7885 = ~1'b0 ;
  assign y7886 = ~n12996 ;
  assign y7887 = n12997 ;
  assign y7888 = n12999 ;
  assign y7889 = ~1'b0 ;
  assign y7890 = n13001 ;
  assign y7891 = ~n13005 ;
  assign y7892 = ~1'b0 ;
  assign y7893 = ~n13009 ;
  assign y7894 = n13012 ;
  assign y7895 = ~n13017 ;
  assign y7896 = n13020 ;
  assign y7897 = n13021 ;
  assign y7898 = ~n10518 ;
  assign y7899 = ~1'b0 ;
  assign y7900 = ~n13024 ;
  assign y7901 = ~n6371 ;
  assign y7902 = ~1'b0 ;
  assign y7903 = ~n13027 ;
  assign y7904 = ~n10482 ;
  assign y7905 = ~1'b0 ;
  assign y7906 = ~n13029 ;
  assign y7907 = ~n13037 ;
  assign y7908 = ~n872 ;
  assign y7909 = ~1'b0 ;
  assign y7910 = n13038 ;
  assign y7911 = n13040 ;
  assign y7912 = n13041 ;
  assign y7913 = n13043 ;
  assign y7914 = ~n13045 ;
  assign y7915 = ~n13048 ;
  assign y7916 = ~n13051 ;
  assign y7917 = n13057 ;
  assign y7918 = ~n13060 ;
  assign y7919 = n13063 ;
  assign y7920 = n13065 ;
  assign y7921 = n13067 ;
  assign y7922 = ~1'b0 ;
  assign y7923 = ~1'b0 ;
  assign y7924 = ~n7223 ;
  assign y7925 = ~n13070 ;
  assign y7926 = ~1'b0 ;
  assign y7927 = ~n13074 ;
  assign y7928 = ~n6369 ;
  assign y7929 = ~1'b0 ;
  assign y7930 = ~n13076 ;
  assign y7931 = ~n13078 ;
  assign y7932 = n13079 ;
  assign y7933 = ~n13082 ;
  assign y7934 = n13084 ;
  assign y7935 = n6357 ;
  assign y7936 = n13086 ;
  assign y7937 = ~1'b0 ;
  assign y7938 = n13088 ;
  assign y7939 = n13090 ;
  assign y7940 = n13091 ;
  assign y7941 = n13093 ;
  assign y7942 = 1'b0 ;
  assign y7943 = n13094 ;
  assign y7944 = ~1'b0 ;
  assign y7945 = ~n13096 ;
  assign y7946 = ~1'b0 ;
  assign y7947 = ~n9483 ;
  assign y7948 = ~n13097 ;
  assign y7949 = n13102 ;
  assign y7950 = ~n13105 ;
  assign y7951 = 1'b0 ;
  assign y7952 = ~1'b0 ;
  assign y7953 = ~n13107 ;
  assign y7954 = ~n13108 ;
  assign y7955 = n13110 ;
  assign y7956 = ~n13113 ;
  assign y7957 = ~1'b0 ;
  assign y7958 = ~n13115 ;
  assign y7959 = n5564 ;
  assign y7960 = ~1'b0 ;
  assign y7961 = n13116 ;
  assign y7962 = 1'b0 ;
  assign y7963 = n428 ;
  assign y7964 = n13117 ;
  assign y7965 = ~1'b0 ;
  assign y7966 = n13118 ;
  assign y7967 = ~n13119 ;
  assign y7968 = ~1'b0 ;
  assign y7969 = n13120 ;
  assign y7970 = ~n13121 ;
  assign y7971 = n13126 ;
  assign y7972 = n13128 ;
  assign y7973 = ~1'b0 ;
  assign y7974 = ~1'b0 ;
  assign y7975 = ~1'b0 ;
  assign y7976 = n6022 ;
  assign y7977 = ~n13135 ;
  assign y7978 = n10785 ;
  assign y7979 = ~n13139 ;
  assign y7980 = n13141 ;
  assign y7981 = ~n13145 ;
  assign y7982 = n13146 ;
  assign y7983 = ~n13147 ;
  assign y7984 = ~1'b0 ;
  assign y7985 = ~1'b0 ;
  assign y7986 = n13148 ;
  assign y7987 = ~n13149 ;
  assign y7988 = ~1'b0 ;
  assign y7989 = n13152 ;
  assign y7990 = n13153 ;
  assign y7991 = ~n13157 ;
  assign y7992 = ~n13161 ;
  assign y7993 = n13162 ;
  assign y7994 = ~n13163 ;
  assign y7995 = ~n13166 ;
  assign y7996 = ~n13167 ;
  assign y7997 = ~n13168 ;
  assign y7998 = ~n13174 ;
  assign y7999 = ~1'b0 ;
  assign y8000 = ~n13176 ;
  assign y8001 = n13181 ;
  assign y8002 = ~1'b0 ;
  assign y8003 = ~1'b0 ;
  assign y8004 = ~1'b0 ;
  assign y8005 = ~n13185 ;
  assign y8006 = ~1'b0 ;
  assign y8007 = n1624 ;
  assign y8008 = n13187 ;
  assign y8009 = ~1'b0 ;
  assign y8010 = ~1'b0 ;
  assign y8011 = ~n11411 ;
  assign y8012 = ~n13192 ;
  assign y8013 = n13193 ;
  assign y8014 = ~1'b0 ;
  assign y8015 = n13197 ;
  assign y8016 = ~1'b0 ;
  assign y8017 = ~1'b0 ;
  assign y8018 = ~1'b0 ;
  assign y8019 = ~n13198 ;
  assign y8020 = n13200 ;
  assign y8021 = n13201 ;
  assign y8022 = ~n10573 ;
  assign y8023 = ~1'b0 ;
  assign y8024 = ~1'b0 ;
  assign y8025 = n13202 ;
  assign y8026 = n13203 ;
  assign y8027 = ~1'b0 ;
  assign y8028 = ~n13209 ;
  assign y8029 = n13211 ;
  assign y8030 = ~1'b0 ;
  assign y8031 = ~n13213 ;
  assign y8032 = ~n13216 ;
  assign y8033 = ~1'b0 ;
  assign y8034 = ~1'b0 ;
  assign y8035 = ~1'b0 ;
  assign y8036 = ~n13220 ;
  assign y8037 = n4980 ;
  assign y8038 = n13222 ;
  assign y8039 = n12083 ;
  assign y8040 = n13229 ;
  assign y8041 = ~n13231 ;
  assign y8042 = n7127 ;
  assign y8043 = ~1'b0 ;
  assign y8044 = ~n13233 ;
  assign y8045 = ~1'b0 ;
  assign y8046 = ~n13234 ;
  assign y8047 = n13239 ;
  assign y8048 = n2257 ;
  assign y8049 = ~1'b0 ;
  assign y8050 = ~n13240 ;
  assign y8051 = ~1'b0 ;
  assign y8052 = ~1'b0 ;
  assign y8053 = ~n13241 ;
  assign y8054 = ~1'b0 ;
  assign y8055 = ~n13242 ;
  assign y8056 = n13243 ;
  assign y8057 = n13244 ;
  assign y8058 = ~1'b0 ;
  assign y8059 = n7926 ;
  assign y8060 = n13247 ;
  assign y8061 = n13248 ;
  assign y8062 = 1'b0 ;
  assign y8063 = n13250 ;
  assign y8064 = ~n13251 ;
  assign y8065 = ~1'b0 ;
  assign y8066 = ~n13254 ;
  assign y8067 = ~n2400 ;
  assign y8068 = ~1'b0 ;
  assign y8069 = ~n13255 ;
  assign y8070 = ~1'b0 ;
  assign y8071 = ~1'b0 ;
  assign y8072 = ~n6932 ;
  assign y8073 = ~1'b0 ;
  assign y8074 = ~1'b0 ;
  assign y8075 = ~1'b0 ;
  assign y8076 = n13257 ;
  assign y8077 = ~1'b0 ;
  assign y8078 = ~n294 ;
  assign y8079 = ~1'b0 ;
  assign y8080 = ~1'b0 ;
  assign y8081 = ~n13260 ;
  assign y8082 = ~n13261 ;
  assign y8083 = ~1'b0 ;
  assign y8084 = n13262 ;
  assign y8085 = ~n13265 ;
  assign y8086 = 1'b0 ;
  assign y8087 = ~1'b0 ;
  assign y8088 = ~1'b0 ;
  assign y8089 = ~x108 ;
  assign y8090 = ~1'b0 ;
  assign y8091 = n4582 ;
  assign y8092 = ~n11185 ;
  assign y8093 = ~n13266 ;
  assign y8094 = 1'b0 ;
  assign y8095 = ~n13271 ;
  assign y8096 = ~n13274 ;
  assign y8097 = ~1'b0 ;
  assign y8098 = ~1'b0 ;
  assign y8099 = n13275 ;
  assign y8100 = n13277 ;
  assign y8101 = ~n13279 ;
  assign y8102 = ~1'b0 ;
  assign y8103 = ~n4252 ;
  assign y8104 = ~1'b0 ;
  assign y8105 = n13280 ;
  assign y8106 = ~1'b0 ;
  assign y8107 = n13282 ;
  assign y8108 = ~n7607 ;
  assign y8109 = ~1'b0 ;
  assign y8110 = ~1'b0 ;
  assign y8111 = ~n13286 ;
  assign y8112 = ~1'b0 ;
  assign y8113 = 1'b0 ;
  assign y8114 = ~n13289 ;
  assign y8115 = ~n13291 ;
  assign y8116 = ~1'b0 ;
  assign y8117 = ~n1329 ;
  assign y8118 = ~1'b0 ;
  assign y8119 = n13292 ;
  assign y8120 = n13295 ;
  assign y8121 = ~1'b0 ;
  assign y8122 = ~n13298 ;
  assign y8123 = n10911 ;
  assign y8124 = ~1'b0 ;
  assign y8125 = ~1'b0 ;
  assign y8126 = ~n13299 ;
  assign y8127 = ~1'b0 ;
  assign y8128 = n13300 ;
  assign y8129 = ~n13301 ;
  assign y8130 = n13302 ;
  assign y8131 = ~1'b0 ;
  assign y8132 = ~n13303 ;
  assign y8133 = ~1'b0 ;
  assign y8134 = 1'b0 ;
  assign y8135 = ~n13304 ;
  assign y8136 = n13305 ;
  assign y8137 = n13307 ;
  assign y8138 = ~1'b0 ;
  assign y8139 = n7997 ;
  assign y8140 = ~1'b0 ;
  assign y8141 = ~n13310 ;
  assign y8142 = ~1'b0 ;
  assign y8143 = ~n13313 ;
  assign y8144 = ~n13316 ;
  assign y8145 = n4748 ;
  assign y8146 = n13319 ;
  assign y8147 = n13320 ;
  assign y8148 = ~1'b0 ;
  assign y8149 = ~1'b0 ;
  assign y8150 = ~1'b0 ;
  assign y8151 = n13321 ;
  assign y8152 = ~1'b0 ;
  assign y8153 = n13323 ;
  assign y8154 = ~1'b0 ;
  assign y8155 = n3904 ;
  assign y8156 = n13326 ;
  assign y8157 = n13328 ;
  assign y8158 = ~n10006 ;
  assign y8159 = ~n13331 ;
  assign y8160 = ~n13332 ;
  assign y8161 = n13352 ;
  assign y8162 = n13358 ;
  assign y8163 = n13360 ;
  assign y8164 = ~n13361 ;
  assign y8165 = ~n13362 ;
  assign y8166 = ~1'b0 ;
  assign y8167 = ~n13365 ;
  assign y8168 = ~1'b0 ;
  assign y8169 = 1'b0 ;
  assign y8170 = ~n13367 ;
  assign y8171 = n13370 ;
  assign y8172 = ~n13371 ;
  assign y8173 = ~1'b0 ;
  assign y8174 = n13372 ;
  assign y8175 = ~1'b0 ;
  assign y8176 = n13374 ;
  assign y8177 = n13385 ;
  assign y8178 = ~n13390 ;
  assign y8179 = n13392 ;
  assign y8180 = ~n13394 ;
  assign y8181 = n11785 ;
  assign y8182 = ~1'b0 ;
  assign y8183 = ~n13397 ;
  assign y8184 = ~1'b0 ;
  assign y8185 = ~n3454 ;
  assign y8186 = ~1'b0 ;
  assign y8187 = ~1'b0 ;
  assign y8188 = n13399 ;
  assign y8189 = ~n361 ;
  assign y8190 = n13402 ;
  assign y8191 = ~1'b0 ;
  assign y8192 = ~n13415 ;
  assign y8193 = ~1'b0 ;
  assign y8194 = ~1'b0 ;
  assign y8195 = ~1'b0 ;
  assign y8196 = ~n13416 ;
  assign y8197 = ~1'b0 ;
  assign y8198 = n13422 ;
  assign y8199 = n13423 ;
  assign y8200 = n13425 ;
  assign y8201 = ~n13428 ;
  assign y8202 = ~1'b0 ;
  assign y8203 = ~1'b0 ;
  assign y8204 = ~n13433 ;
  assign y8205 = ~1'b0 ;
  assign y8206 = n11175 ;
  assign y8207 = ~n13434 ;
  assign y8208 = ~1'b0 ;
  assign y8209 = ~1'b0 ;
  assign y8210 = ~n13436 ;
  assign y8211 = ~1'b0 ;
  assign y8212 = ~1'b0 ;
  assign y8213 = ~n13438 ;
  assign y8214 = ~n802 ;
  assign y8215 = ~n13440 ;
  assign y8216 = ~n567 ;
  assign y8217 = ~1'b0 ;
  assign y8218 = ~1'b0 ;
  assign y8219 = ~n13442 ;
  assign y8220 = ~n13444 ;
  assign y8221 = ~n5282 ;
  assign y8222 = ~n8909 ;
  assign y8223 = n13446 ;
  assign y8224 = n6180 ;
  assign y8225 = n13448 ;
  assign y8226 = n13449 ;
  assign y8227 = n13451 ;
  assign y8228 = ~1'b0 ;
  assign y8229 = n13452 ;
  assign y8230 = n13453 ;
  assign y8231 = n10292 ;
  assign y8232 = ~n1031 ;
  assign y8233 = ~n13454 ;
  assign y8234 = ~n13463 ;
  assign y8235 = ~n13467 ;
  assign y8236 = ~n13469 ;
  assign y8237 = n13470 ;
  assign y8238 = n10312 ;
  assign y8239 = ~n5054 ;
  assign y8240 = n13471 ;
  assign y8241 = ~n13473 ;
  assign y8242 = ~1'b0 ;
  assign y8243 = ~n13477 ;
  assign y8244 = ~n13479 ;
  assign y8245 = ~1'b0 ;
  assign y8246 = ~1'b0 ;
  assign y8247 = ~n13480 ;
  assign y8248 = ~1'b0 ;
  assign y8249 = ~1'b0 ;
  assign y8250 = n13483 ;
  assign y8251 = n13484 ;
  assign y8252 = ~n13486 ;
  assign y8253 = ~1'b0 ;
  assign y8254 = ~1'b0 ;
  assign y8255 = ~n13487 ;
  assign y8256 = ~n13492 ;
  assign y8257 = ~n13493 ;
  assign y8258 = ~1'b0 ;
  assign y8259 = ~1'b0 ;
  assign y8260 = 1'b0 ;
  assign y8261 = n13495 ;
  assign y8262 = n13488 ;
  assign y8263 = n13496 ;
  assign y8264 = ~1'b0 ;
  assign y8265 = ~1'b0 ;
  assign y8266 = ~1'b0 ;
  assign y8267 = ~n13498 ;
  assign y8268 = ~n13502 ;
  assign y8269 = ~n424 ;
  assign y8270 = n13504 ;
  assign y8271 = n8629 ;
  assign y8272 = n13505 ;
  assign y8273 = ~1'b0 ;
  assign y8274 = n13507 ;
  assign y8275 = ~n13508 ;
  assign y8276 = ~n13510 ;
  assign y8277 = ~1'b0 ;
  assign y8278 = n13512 ;
  assign y8279 = ~n13514 ;
  assign y8280 = ~n13516 ;
  assign y8281 = n13518 ;
  assign y8282 = ~1'b0 ;
  assign y8283 = ~1'b0 ;
  assign y8284 = ~n13519 ;
  assign y8285 = n13520 ;
  assign y8286 = ~1'b0 ;
  assign y8287 = ~n13521 ;
  assign y8288 = ~1'b0 ;
  assign y8289 = ~1'b0 ;
  assign y8290 = ~1'b0 ;
  assign y8291 = ~1'b0 ;
  assign y8292 = n13522 ;
  assign y8293 = ~1'b0 ;
  assign y8294 = n13525 ;
  assign y8295 = 1'b0 ;
  assign y8296 = ~n13527 ;
  assign y8297 = 1'b0 ;
  assign y8298 = ~1'b0 ;
  assign y8299 = ~n290 ;
  assign y8300 = n13533 ;
  assign y8301 = n13542 ;
  assign y8302 = n13546 ;
  assign y8303 = ~1'b0 ;
  assign y8304 = ~n9176 ;
  assign y8305 = n13549 ;
  assign y8306 = ~1'b0 ;
  assign y8307 = ~n13550 ;
  assign y8308 = n2999 ;
  assign y8309 = ~1'b0 ;
  assign y8310 = n13554 ;
  assign y8311 = ~n13557 ;
  assign y8312 = ~1'b0 ;
  assign y8313 = ~n13558 ;
  assign y8314 = ~n13562 ;
  assign y8315 = 1'b0 ;
  assign y8316 = ~n13564 ;
  assign y8317 = ~n13567 ;
  assign y8318 = ~1'b0 ;
  assign y8319 = ~1'b0 ;
  assign y8320 = ~1'b0 ;
  assign y8321 = ~1'b0 ;
  assign y8322 = ~n13568 ;
  assign y8323 = ~1'b0 ;
  assign y8324 = ~n13569 ;
  assign y8325 = ~n13579 ;
  assign y8326 = ~1'b0 ;
  assign y8327 = ~1'b0 ;
  assign y8328 = ~n13583 ;
  assign y8329 = n13585 ;
  assign y8330 = n5708 ;
  assign y8331 = n13589 ;
  assign y8332 = ~1'b0 ;
  assign y8333 = ~1'b0 ;
  assign y8334 = ~1'b0 ;
  assign y8335 = ~1'b0 ;
  assign y8336 = ~n13590 ;
  assign y8337 = ~1'b0 ;
  assign y8338 = ~n13592 ;
  assign y8339 = ~1'b0 ;
  assign y8340 = n7361 ;
  assign y8341 = ~n5327 ;
  assign y8342 = ~n13595 ;
  assign y8343 = ~1'b0 ;
  assign y8344 = n11710 ;
  assign y8345 = ~n13596 ;
  assign y8346 = ~n13598 ;
  assign y8347 = x97 ;
  assign y8348 = n13600 ;
  assign y8349 = ~n13601 ;
  assign y8350 = n13603 ;
  assign y8351 = ~n2718 ;
  assign y8352 = n13614 ;
  assign y8353 = n13621 ;
  assign y8354 = ~1'b0 ;
  assign y8355 = ~n13624 ;
  assign y8356 = ~1'b0 ;
  assign y8357 = ~1'b0 ;
  assign y8358 = ~n13625 ;
  assign y8359 = ~1'b0 ;
  assign y8360 = ~n13627 ;
  assign y8361 = ~n13628 ;
  assign y8362 = ~1'b0 ;
  assign y8363 = ~1'b0 ;
  assign y8364 = n13630 ;
  assign y8365 = n13631 ;
  assign y8366 = n13636 ;
  assign y8367 = n11782 ;
  assign y8368 = ~1'b0 ;
  assign y8369 = ~1'b0 ;
  assign y8370 = n13637 ;
  assign y8371 = ~n13641 ;
  assign y8372 = n13643 ;
  assign y8373 = ~n13645 ;
  assign y8374 = ~1'b0 ;
  assign y8375 = ~1'b0 ;
  assign y8376 = n3708 ;
  assign y8377 = n13648 ;
  assign y8378 = ~1'b0 ;
  assign y8379 = n8046 ;
  assign y8380 = ~1'b0 ;
  assign y8381 = 1'b0 ;
  assign y8382 = x49 ;
  assign y8383 = 1'b0 ;
  assign y8384 = n13651 ;
  assign y8385 = ~1'b0 ;
  assign y8386 = n13653 ;
  assign y8387 = n13656 ;
  assign y8388 = n13657 ;
  assign y8389 = ~n13658 ;
  assign y8390 = n6642 ;
  assign y8391 = ~n13659 ;
  assign y8392 = n13660 ;
  assign y8393 = ~n13661 ;
  assign y8394 = ~n13663 ;
  assign y8395 = ~1'b0 ;
  assign y8396 = ~n13664 ;
  assign y8397 = ~1'b0 ;
  assign y8398 = n13667 ;
  assign y8399 = n13668 ;
  assign y8400 = ~1'b0 ;
  assign y8401 = ~n13671 ;
  assign y8402 = ~1'b0 ;
  assign y8403 = n13673 ;
  assign y8404 = ~n13675 ;
  assign y8405 = ~n13678 ;
  assign y8406 = n13680 ;
  assign y8407 = ~n13681 ;
  assign y8408 = n13683 ;
  assign y8409 = ~1'b0 ;
  assign y8410 = ~1'b0 ;
  assign y8411 = n13034 ;
  assign y8412 = ~n13688 ;
  assign y8413 = ~1'b0 ;
  assign y8414 = ~1'b0 ;
  assign y8415 = n13690 ;
  assign y8416 = n13691 ;
  assign y8417 = ~n13693 ;
  assign y8418 = ~n13696 ;
  assign y8419 = n13698 ;
  assign y8420 = ~n5663 ;
  assign y8421 = ~n13704 ;
  assign y8422 = 1'b0 ;
  assign y8423 = x115 ;
  assign y8424 = ~n13706 ;
  assign y8425 = ~1'b0 ;
  assign y8426 = ~n13709 ;
  assign y8427 = ~n13714 ;
  assign y8428 = n13719 ;
  assign y8429 = ~n13723 ;
  assign y8430 = ~n4298 ;
  assign y8431 = n13724 ;
  assign y8432 = ~n13730 ;
  assign y8433 = n13731 ;
  assign y8434 = ~n13733 ;
  assign y8435 = ~1'b0 ;
  assign y8436 = ~n13734 ;
  assign y8437 = ~1'b0 ;
  assign y8438 = n13738 ;
  assign y8439 = n13739 ;
  assign y8440 = n2091 ;
  assign y8441 = 1'b0 ;
  assign y8442 = ~1'b0 ;
  assign y8443 = ~n13741 ;
  assign y8444 = ~n2213 ;
  assign y8445 = ~n13742 ;
  assign y8446 = n13744 ;
  assign y8447 = ~n13747 ;
  assign y8448 = n13752 ;
  assign y8449 = ~n13759 ;
  assign y8450 = ~n13763 ;
  assign y8451 = ~1'b0 ;
  assign y8452 = ~1'b0 ;
  assign y8453 = n13769 ;
  assign y8454 = n457 ;
  assign y8455 = ~1'b0 ;
  assign y8456 = n13774 ;
  assign y8457 = n13777 ;
  assign y8458 = n5120 ;
  assign y8459 = ~n13780 ;
  assign y8460 = 1'b0 ;
  assign y8461 = n13781 ;
  assign y8462 = n13783 ;
  assign y8463 = ~1'b0 ;
  assign y8464 = ~n13785 ;
  assign y8465 = ~1'b0 ;
  assign y8466 = n13787 ;
  assign y8467 = ~n13794 ;
  assign y8468 = 1'b0 ;
  assign y8469 = 1'b0 ;
  assign y8470 = 1'b0 ;
  assign y8471 = n13798 ;
  assign y8472 = ~n13800 ;
  assign y8473 = n5352 ;
  assign y8474 = n8706 ;
  assign y8475 = ~1'b0 ;
  assign y8476 = ~1'b0 ;
  assign y8477 = ~n13805 ;
  assign y8478 = n6780 ;
  assign y8479 = n13809 ;
  assign y8480 = ~1'b0 ;
  assign y8481 = 1'b0 ;
  assign y8482 = ~n2503 ;
  assign y8483 = ~n13813 ;
  assign y8484 = ~1'b0 ;
  assign y8485 = n13815 ;
  assign y8486 = ~n13816 ;
  assign y8487 = ~1'b0 ;
  assign y8488 = ~1'b0 ;
  assign y8489 = ~1'b0 ;
  assign y8490 = ~n2831 ;
  assign y8491 = ~1'b0 ;
  assign y8492 = ~1'b0 ;
  assign y8493 = ~n13821 ;
  assign y8494 = ~1'b0 ;
  assign y8495 = n13822 ;
  assign y8496 = n7785 ;
  assign y8497 = n1037 ;
  assign y8498 = ~n13823 ;
  assign y8499 = n13824 ;
  assign y8500 = n8807 ;
  assign y8501 = ~1'b0 ;
  assign y8502 = ~1'b0 ;
  assign y8503 = ~n13826 ;
  assign y8504 = ~1'b0 ;
  assign y8505 = ~1'b0 ;
  assign y8506 = ~n13829 ;
  assign y8507 = n13831 ;
  assign y8508 = n13832 ;
  assign y8509 = ~1'b0 ;
  assign y8510 = ~1'b0 ;
  assign y8511 = n13833 ;
  assign y8512 = n13837 ;
  assign y8513 = ~n13839 ;
  assign y8514 = n13840 ;
  assign y8515 = ~n13844 ;
  assign y8516 = n13846 ;
  assign y8517 = ~n13849 ;
  assign y8518 = ~n13853 ;
  assign y8519 = ~1'b0 ;
  assign y8520 = n13854 ;
  assign y8521 = ~n3189 ;
  assign y8522 = n13856 ;
  assign y8523 = ~1'b0 ;
  assign y8524 = ~1'b0 ;
  assign y8525 = ~1'b0 ;
  assign y8526 = ~1'b0 ;
  assign y8527 = ~n13859 ;
  assign y8528 = ~1'b0 ;
  assign y8529 = ~1'b0 ;
  assign y8530 = n13861 ;
  assign y8531 = ~n13871 ;
  assign y8532 = ~1'b0 ;
  assign y8533 = ~n13872 ;
  assign y8534 = ~1'b0 ;
  assign y8535 = n13873 ;
  assign y8536 = ~1'b0 ;
  assign y8537 = ~n13876 ;
  assign y8538 = ~1'b0 ;
  assign y8539 = 1'b0 ;
  assign y8540 = ~n13878 ;
  assign y8541 = ~n13880 ;
  assign y8542 = ~1'b0 ;
  assign y8543 = 1'b0 ;
  assign y8544 = ~1'b0 ;
  assign y8545 = ~1'b0 ;
  assign y8546 = ~1'b0 ;
  assign y8547 = ~n13888 ;
  assign y8548 = ~1'b0 ;
  assign y8549 = ~1'b0 ;
  assign y8550 = ~n13893 ;
  assign y8551 = ~n13896 ;
  assign y8552 = ~n8496 ;
  assign y8553 = ~n13897 ;
  assign y8554 = ~1'b0 ;
  assign y8555 = ~1'b0 ;
  assign y8556 = n13900 ;
  assign y8557 = n13901 ;
  assign y8558 = n13903 ;
  assign y8559 = n13907 ;
  assign y8560 = n13908 ;
  assign y8561 = ~n13909 ;
  assign y8562 = ~n13910 ;
  assign y8563 = ~1'b0 ;
  assign y8564 = n13912 ;
  assign y8565 = ~1'b0 ;
  assign y8566 = n5417 ;
  assign y8567 = ~1'b0 ;
  assign y8568 = ~n13918 ;
  assign y8569 = ~n13919 ;
  assign y8570 = ~n13922 ;
  assign y8571 = n13925 ;
  assign y8572 = ~n13927 ;
  assign y8573 = n8235 ;
  assign y8574 = n13932 ;
  assign y8575 = ~n13935 ;
  assign y8576 = n13937 ;
  assign y8577 = n13938 ;
  assign y8578 = ~n4654 ;
  assign y8579 = ~n13939 ;
  assign y8580 = ~1'b0 ;
  assign y8581 = n13940 ;
  assign y8582 = ~1'b0 ;
  assign y8583 = ~n13942 ;
  assign y8584 = ~1'b0 ;
  assign y8585 = ~1'b0 ;
  assign y8586 = ~n13945 ;
  assign y8587 = ~n13947 ;
  assign y8588 = ~n13948 ;
  assign y8589 = n3196 ;
  assign y8590 = ~1'b0 ;
  assign y8591 = ~n13949 ;
  assign y8592 = ~n13950 ;
  assign y8593 = n13957 ;
  assign y8594 = ~1'b0 ;
  assign y8595 = ~n13959 ;
  assign y8596 = ~1'b0 ;
  assign y8597 = n5142 ;
  assign y8598 = n13961 ;
  assign y8599 = ~n13964 ;
  assign y8600 = ~n13968 ;
  assign y8601 = ~1'b0 ;
  assign y8602 = ~n3477 ;
  assign y8603 = ~1'b0 ;
  assign y8604 = ~1'b0 ;
  assign y8605 = ~1'b0 ;
  assign y8606 = ~n13970 ;
  assign y8607 = ~n297 ;
  assign y8608 = n13973 ;
  assign y8609 = n13978 ;
  assign y8610 = ~n13980 ;
  assign y8611 = ~n13987 ;
  assign y8612 = n13988 ;
  assign y8613 = ~1'b0 ;
  assign y8614 = n13990 ;
  assign y8615 = n1188 ;
  assign y8616 = ~n13991 ;
  assign y8617 = ~1'b0 ;
  assign y8618 = ~1'b0 ;
  assign y8619 = ~n13995 ;
  assign y8620 = ~n13999 ;
  assign y8621 = 1'b0 ;
  assign y8622 = ~n14000 ;
  assign y8623 = ~n14001 ;
  assign y8624 = ~n14003 ;
  assign y8625 = ~1'b0 ;
  assign y8626 = n14010 ;
  assign y8627 = ~n14012 ;
  assign y8628 = n14013 ;
  assign y8629 = n14020 ;
  assign y8630 = ~n14021 ;
  assign y8631 = n14026 ;
  assign y8632 = ~n14027 ;
  assign y8633 = ~n14030 ;
  assign y8634 = n14033 ;
  assign y8635 = ~1'b0 ;
  assign y8636 = ~n14035 ;
  assign y8637 = ~1'b0 ;
  assign y8638 = ~n14036 ;
  assign y8639 = ~n14041 ;
  assign y8640 = ~1'b0 ;
  assign y8641 = ~1'b0 ;
  assign y8642 = ~1'b0 ;
  assign y8643 = 1'b0 ;
  assign y8644 = ~n14042 ;
  assign y8645 = ~n14049 ;
  assign y8646 = ~1'b0 ;
  assign y8647 = ~1'b0 ;
  assign y8648 = ~n14051 ;
  assign y8649 = ~n6370 ;
  assign y8650 = ~1'b0 ;
  assign y8651 = n14054 ;
  assign y8652 = ~1'b0 ;
  assign y8653 = n14060 ;
  assign y8654 = n8773 ;
  assign y8655 = ~n14064 ;
  assign y8656 = ~n14066 ;
  assign y8657 = ~n14067 ;
  assign y8658 = ~n14069 ;
  assign y8659 = n8958 ;
  assign y8660 = ~n5007 ;
  assign y8661 = ~n14070 ;
  assign y8662 = ~1'b0 ;
  assign y8663 = ~1'b0 ;
  assign y8664 = n14071 ;
  assign y8665 = ~n14072 ;
  assign y8666 = ~1'b0 ;
  assign y8667 = ~1'b0 ;
  assign y8668 = n14077 ;
  assign y8669 = ~1'b0 ;
  assign y8670 = ~1'b0 ;
  assign y8671 = ~n14078 ;
  assign y8672 = ~n12275 ;
  assign y8673 = ~1'b0 ;
  assign y8674 = ~1'b0 ;
  assign y8675 = ~1'b0 ;
  assign y8676 = ~n14081 ;
  assign y8677 = n3230 ;
  assign y8678 = n13096 ;
  assign y8679 = n12262 ;
  assign y8680 = n14082 ;
  assign y8681 = ~n14084 ;
  assign y8682 = 1'b0 ;
  assign y8683 = ~n14089 ;
  assign y8684 = ~n14091 ;
  assign y8685 = ~1'b0 ;
  assign y8686 = ~n14093 ;
  assign y8687 = ~n14094 ;
  assign y8688 = 1'b0 ;
  assign y8689 = ~n14097 ;
  assign y8690 = n14098 ;
  assign y8691 = ~n14107 ;
  assign y8692 = ~1'b0 ;
  assign y8693 = ~1'b0 ;
  assign y8694 = n14108 ;
  assign y8695 = ~n14111 ;
  assign y8696 = ~1'b0 ;
  assign y8697 = n13447 ;
  assign y8698 = ~n14114 ;
  assign y8699 = ~1'b0 ;
  assign y8700 = ~n14116 ;
  assign y8701 = ~n13376 ;
  assign y8702 = ~n14117 ;
  assign y8703 = n14120 ;
  assign y8704 = 1'b0 ;
  assign y8705 = ~n14121 ;
  assign y8706 = n14124 ;
  assign y8707 = ~1'b0 ;
  assign y8708 = ~n14125 ;
  assign y8709 = ~1'b0 ;
  assign y8710 = n14126 ;
  assign y8711 = ~1'b0 ;
  assign y8712 = n14130 ;
  assign y8713 = ~n14131 ;
  assign y8714 = ~n7726 ;
  assign y8715 = n11569 ;
  assign y8716 = ~1'b0 ;
  assign y8717 = ~n7994 ;
  assign y8718 = ~1'b0 ;
  assign y8719 = ~n14133 ;
  assign y8720 = 1'b0 ;
  assign y8721 = ~n14137 ;
  assign y8722 = ~1'b0 ;
  assign y8723 = ~n14139 ;
  assign y8724 = n14142 ;
  assign y8725 = ~n14144 ;
  assign y8726 = ~n14146 ;
  assign y8727 = n14151 ;
  assign y8728 = ~n14153 ;
  assign y8729 = ~1'b0 ;
  assign y8730 = n14154 ;
  assign y8731 = n14155 ;
  assign y8732 = n14158 ;
  assign y8733 = ~1'b0 ;
  assign y8734 = n14159 ;
  assign y8735 = n14160 ;
  assign y8736 = ~n14161 ;
  assign y8737 = n14162 ;
  assign y8738 = ~1'b0 ;
  assign y8739 = ~n14166 ;
  assign y8740 = ~1'b0 ;
  assign y8741 = ~n14168 ;
  assign y8742 = n14169 ;
  assign y8743 = n14170 ;
  assign y8744 = ~n14172 ;
  assign y8745 = n14174 ;
  assign y8746 = n14175 ;
  assign y8747 = ~n14177 ;
  assign y8748 = n14178 ;
  assign y8749 = ~1'b0 ;
  assign y8750 = n14180 ;
  assign y8751 = n820 ;
  assign y8752 = ~1'b0 ;
  assign y8753 = n14181 ;
  assign y8754 = n14185 ;
  assign y8755 = ~1'b0 ;
  assign y8756 = ~n2673 ;
  assign y8757 = ~1'b0 ;
  assign y8758 = n14186 ;
  assign y8759 = ~1'b0 ;
  assign y8760 = ~n14187 ;
  assign y8761 = ~1'b0 ;
  assign y8762 = n14190 ;
  assign y8763 = ~n14191 ;
  assign y8764 = n14193 ;
  assign y8765 = ~1'b0 ;
  assign y8766 = ~1'b0 ;
  assign y8767 = ~1'b0 ;
  assign y8768 = ~1'b0 ;
  assign y8769 = ~1'b0 ;
  assign y8770 = ~n14195 ;
  assign y8771 = ~n14198 ;
  assign y8772 = n14207 ;
  assign y8773 = ~n14209 ;
  assign y8774 = n14212 ;
  assign y8775 = ~1'b0 ;
  assign y8776 = n14214 ;
  assign y8777 = ~n14216 ;
  assign y8778 = ~n14218 ;
  assign y8779 = ~1'b0 ;
  assign y8780 = 1'b0 ;
  assign y8781 = ~n14220 ;
  assign y8782 = n9252 ;
  assign y8783 = ~n14223 ;
  assign y8784 = ~1'b0 ;
  assign y8785 = n14230 ;
  assign y8786 = n14231 ;
  assign y8787 = ~n14233 ;
  assign y8788 = ~1'b0 ;
  assign y8789 = n14235 ;
  assign y8790 = n14237 ;
  assign y8791 = ~n14244 ;
  assign y8792 = ~n1432 ;
  assign y8793 = ~1'b0 ;
  assign y8794 = ~1'b0 ;
  assign y8795 = n14245 ;
  assign y8796 = n14248 ;
  assign y8797 = ~1'b0 ;
  assign y8798 = n14253 ;
  assign y8799 = n14254 ;
  assign y8800 = n10922 ;
  assign y8801 = ~n14256 ;
  assign y8802 = ~1'b0 ;
  assign y8803 = n14257 ;
  assign y8804 = n14258 ;
  assign y8805 = n14262 ;
  assign y8806 = ~n14263 ;
  assign y8807 = 1'b0 ;
  assign y8808 = 1'b0 ;
  assign y8809 = ~1'b0 ;
  assign y8810 = ~1'b0 ;
  assign y8811 = ~1'b0 ;
  assign y8812 = n14265 ;
  assign y8813 = ~1'b0 ;
  assign y8814 = ~1'b0 ;
  assign y8815 = n14267 ;
  assign y8816 = ~1'b0 ;
  assign y8817 = ~n14268 ;
  assign y8818 = ~1'b0 ;
  assign y8819 = n14274 ;
  assign y8820 = n10556 ;
  assign y8821 = n14277 ;
  assign y8822 = ~1'b0 ;
  assign y8823 = ~n14280 ;
  assign y8824 = ~1'b0 ;
  assign y8825 = ~1'b0 ;
  assign y8826 = ~1'b0 ;
  assign y8827 = n14281 ;
  assign y8828 = n14282 ;
  assign y8829 = ~n14283 ;
  assign y8830 = ~n14284 ;
  assign y8831 = n4998 ;
  assign y8832 = n14286 ;
  assign y8833 = n14289 ;
  assign y8834 = ~1'b0 ;
  assign y8835 = ~1'b0 ;
  assign y8836 = ~n5417 ;
  assign y8837 = n14293 ;
  assign y8838 = n14297 ;
  assign y8839 = ~1'b0 ;
  assign y8840 = n14300 ;
  assign y8841 = ~1'b0 ;
  assign y8842 = ~1'b0 ;
  assign y8843 = ~n14303 ;
  assign y8844 = ~1'b0 ;
  assign y8845 = ~n9492 ;
  assign y8846 = n14307 ;
  assign y8847 = ~1'b0 ;
  assign y8848 = n14313 ;
  assign y8849 = ~1'b0 ;
  assign y8850 = ~n14315 ;
  assign y8851 = n5985 ;
  assign y8852 = n14316 ;
  assign y8853 = n14318 ;
  assign y8854 = ~n7244 ;
  assign y8855 = ~n2178 ;
  assign y8856 = 1'b0 ;
  assign y8857 = ~n14321 ;
  assign y8858 = ~1'b0 ;
  assign y8859 = ~1'b0 ;
  assign y8860 = n14323 ;
  assign y8861 = ~1'b0 ;
  assign y8862 = n14324 ;
  assign y8863 = ~n14330 ;
  assign y8864 = n14331 ;
  assign y8865 = n14333 ;
  assign y8866 = ~n14335 ;
  assign y8867 = n14337 ;
  assign y8868 = n14338 ;
  assign y8869 = n14340 ;
  assign y8870 = n14342 ;
  assign y8871 = ~n14343 ;
  assign y8872 = n9096 ;
  assign y8873 = n14344 ;
  assign y8874 = n14346 ;
  assign y8875 = n6626 ;
  assign y8876 = n14347 ;
  assign y8877 = 1'b0 ;
  assign y8878 = ~n4664 ;
  assign y8879 = 1'b0 ;
  assign y8880 = n9726 ;
  assign y8881 = n7529 ;
  assign y8882 = ~1'b0 ;
  assign y8883 = ~1'b0 ;
  assign y8884 = ~1'b0 ;
  assign y8885 = ~n14350 ;
  assign y8886 = ~n14353 ;
  assign y8887 = ~1'b0 ;
  assign y8888 = n14354 ;
  assign y8889 = ~1'b0 ;
  assign y8890 = ~n14356 ;
  assign y8891 = n14359 ;
  assign y8892 = 1'b0 ;
  assign y8893 = n14360 ;
  assign y8894 = n14361 ;
  assign y8895 = n13903 ;
  assign y8896 = ~n14362 ;
  assign y8897 = n6918 ;
  assign y8898 = ~n14365 ;
  assign y8899 = ~n14372 ;
  assign y8900 = n14376 ;
  assign y8901 = ~1'b0 ;
  assign y8902 = ~n14378 ;
  assign y8903 = 1'b0 ;
  assign y8904 = ~1'b0 ;
  assign y8905 = n14379 ;
  assign y8906 = ~n14381 ;
  assign y8907 = ~n3585 ;
  assign y8908 = ~1'b0 ;
  assign y8909 = ~n7959 ;
  assign y8910 = ~n14382 ;
  assign y8911 = ~n14385 ;
  assign y8912 = ~1'b0 ;
  assign y8913 = ~1'b0 ;
  assign y8914 = n14387 ;
  assign y8915 = n14390 ;
  assign y8916 = n10392 ;
  assign y8917 = ~1'b0 ;
  assign y8918 = ~1'b0 ;
  assign y8919 = n14392 ;
  assign y8920 = n14398 ;
  assign y8921 = 1'b0 ;
  assign y8922 = ~n14399 ;
  assign y8923 = n14408 ;
  assign y8924 = ~n14409 ;
  assign y8925 = 1'b0 ;
  assign y8926 = ~n14410 ;
  assign y8927 = ~n11889 ;
  assign y8928 = ~1'b0 ;
  assign y8929 = ~1'b0 ;
  assign y8930 = ~1'b0 ;
  assign y8931 = ~n14411 ;
  assign y8932 = ~n8737 ;
  assign y8933 = n14414 ;
  assign y8934 = ~1'b0 ;
  assign y8935 = n14415 ;
  assign y8936 = ~n14417 ;
  assign y8937 = n14418 ;
  assign y8938 = n14420 ;
  assign y8939 = ~1'b0 ;
  assign y8940 = ~n14425 ;
  assign y8941 = ~n12156 ;
  assign y8942 = ~n14426 ;
  assign y8943 = n14428 ;
  assign y8944 = n12408 ;
  assign y8945 = n14431 ;
  assign y8946 = ~1'b0 ;
  assign y8947 = ~1'b0 ;
  assign y8948 = ~1'b0 ;
  assign y8949 = 1'b0 ;
  assign y8950 = n10968 ;
  assign y8951 = ~n14432 ;
  assign y8952 = n14436 ;
  assign y8953 = n14438 ;
  assign y8954 = n13376 ;
  assign y8955 = ~n14439 ;
  assign y8956 = ~1'b0 ;
  assign y8957 = ~1'b0 ;
  assign y8958 = ~1'b0 ;
  assign y8959 = ~1'b0 ;
  assign y8960 = ~1'b0 ;
  assign y8961 = n10611 ;
  assign y8962 = ~1'b0 ;
  assign y8963 = n14442 ;
  assign y8964 = n14443 ;
  assign y8965 = n14446 ;
  assign y8966 = n14447 ;
  assign y8967 = ~1'b0 ;
  assign y8968 = ~1'b0 ;
  assign y8969 = n14463 ;
  assign y8970 = n14464 ;
  assign y8971 = ~n14466 ;
  assign y8972 = 1'b0 ;
  assign y8973 = ~1'b0 ;
  assign y8974 = n12234 ;
  assign y8975 = n14469 ;
  assign y8976 = n14473 ;
  assign y8977 = n14475 ;
  assign y8978 = ~1'b0 ;
  assign y8979 = ~n14477 ;
  assign y8980 = ~1'b0 ;
  assign y8981 = ~1'b0 ;
  assign y8982 = ~1'b0 ;
  assign y8983 = ~1'b0 ;
  assign y8984 = ~1'b0 ;
  assign y8985 = ~1'b0 ;
  assign y8986 = ~n14480 ;
  assign y8987 = ~n14489 ;
  assign y8988 = ~1'b0 ;
  assign y8989 = n14491 ;
  assign y8990 = ~n7718 ;
  assign y8991 = ~1'b0 ;
  assign y8992 = ~n10793 ;
  assign y8993 = ~n14120 ;
  assign y8994 = ~1'b0 ;
  assign y8995 = ~1'b0 ;
  assign y8996 = n6011 ;
  assign y8997 = n14496 ;
  assign y8998 = ~n14498 ;
  assign y8999 = ~n14499 ;
  assign y9000 = 1'b0 ;
  assign y9001 = ~n316 ;
  assign y9002 = ~n14500 ;
  assign y9003 = ~n14501 ;
  assign y9004 = ~1'b0 ;
  assign y9005 = ~n14502 ;
  assign y9006 = ~n14504 ;
  assign y9007 = n14510 ;
  assign y9008 = ~1'b0 ;
  assign y9009 = n6671 ;
  assign y9010 = ~n14511 ;
  assign y9011 = n14512 ;
  assign y9012 = ~1'b0 ;
  assign y9013 = ~1'b0 ;
  assign y9014 = ~n14514 ;
  assign y9015 = n14515 ;
  assign y9016 = ~1'b0 ;
  assign y9017 = n14532 ;
  assign y9018 = ~1'b0 ;
  assign y9019 = n14533 ;
  assign y9020 = ~n14534 ;
  assign y9021 = ~n14537 ;
  assign y9022 = ~n14538 ;
  assign y9023 = ~1'b0 ;
  assign y9024 = n14539 ;
  assign y9025 = n14540 ;
  assign y9026 = ~1'b0 ;
  assign y9027 = n14541 ;
  assign y9028 = n14547 ;
  assign y9029 = n14549 ;
  assign y9030 = ~n14554 ;
  assign y9031 = ~n14555 ;
  assign y9032 = n14556 ;
  assign y9033 = ~1'b0 ;
  assign y9034 = ~n14557 ;
  assign y9035 = n14558 ;
  assign y9036 = n14560 ;
  assign y9037 = n14562 ;
  assign y9038 = ~n14564 ;
  assign y9039 = ~n14569 ;
  assign y9040 = ~1'b0 ;
  assign y9041 = ~n2756 ;
  assign y9042 = ~n14575 ;
  assign y9043 = ~n4971 ;
  assign y9044 = ~n14580 ;
  assign y9045 = ~n14583 ;
  assign y9046 = ~n14585 ;
  assign y9047 = ~n14588 ;
  assign y9048 = ~n14591 ;
  assign y9049 = n14593 ;
  assign y9050 = ~1'b0 ;
  assign y9051 = ~n14598 ;
  assign y9052 = n14600 ;
  assign y9053 = ~1'b0 ;
  assign y9054 = ~n14603 ;
  assign y9055 = ~n14604 ;
  assign y9056 = ~1'b0 ;
  assign y9057 = n14606 ;
  assign y9058 = ~n14609 ;
  assign y9059 = ~n14611 ;
  assign y9060 = n14612 ;
  assign y9061 = n14613 ;
  assign y9062 = ~1'b0 ;
  assign y9063 = ~n14619 ;
  assign y9064 = ~1'b0 ;
  assign y9065 = n14621 ;
  assign y9066 = n14626 ;
  assign y9067 = ~n10485 ;
  assign y9068 = ~n14629 ;
  assign y9069 = ~n14632 ;
  assign y9070 = n14636 ;
  assign y9071 = ~1'b0 ;
  assign y9072 = ~1'b0 ;
  assign y9073 = ~1'b0 ;
  assign y9074 = ~n14637 ;
  assign y9075 = ~n14638 ;
  assign y9076 = n14639 ;
  assign y9077 = ~n2966 ;
  assign y9078 = ~1'b0 ;
  assign y9079 = n14642 ;
  assign y9080 = ~1'b0 ;
  assign y9081 = n14644 ;
  assign y9082 = n14646 ;
  assign y9083 = ~1'b0 ;
  assign y9084 = n14648 ;
  assign y9085 = 1'b0 ;
  assign y9086 = ~1'b0 ;
  assign y9087 = n11442 ;
  assign y9088 = n14650 ;
  assign y9089 = ~n9488 ;
  assign y9090 = ~n14652 ;
  assign y9091 = n14655 ;
  assign y9092 = n14657 ;
  assign y9093 = ~1'b0 ;
  assign y9094 = ~1'b0 ;
  assign y9095 = n14658 ;
  assign y9096 = ~1'b0 ;
  assign y9097 = ~1'b0 ;
  assign y9098 = ~1'b0 ;
  assign y9099 = ~n3494 ;
  assign y9100 = ~n14660 ;
  assign y9101 = n14662 ;
  assign y9102 = n14664 ;
  assign y9103 = ~n4505 ;
  assign y9104 = ~1'b0 ;
  assign y9105 = ~1'b0 ;
  assign y9106 = n14666 ;
  assign y9107 = ~n14673 ;
  assign y9108 = ~n14676 ;
  assign y9109 = ~1'b0 ;
  assign y9110 = ~n14677 ;
  assign y9111 = ~1'b0 ;
  assign y9112 = ~n14678 ;
  assign y9113 = ~1'b0 ;
  assign y9114 = ~n11051 ;
  assign y9115 = ~n14679 ;
  assign y9116 = ~1'b0 ;
  assign y9117 = n14686 ;
  assign y9118 = n14691 ;
  assign y9119 = ~1'b0 ;
  assign y9120 = ~n14696 ;
  assign y9121 = ~n14697 ;
  assign y9122 = ~n14704 ;
  assign y9123 = ~n14707 ;
  assign y9124 = n14711 ;
  assign y9125 = ~1'b0 ;
  assign y9126 = n14712 ;
  assign y9127 = ~1'b0 ;
  assign y9128 = 1'b0 ;
  assign y9129 = ~1'b0 ;
  assign y9130 = n14714 ;
  assign y9131 = n14716 ;
  assign y9132 = ~n14720 ;
  assign y9133 = ~1'b0 ;
  assign y9134 = ~n14722 ;
  assign y9135 = n14723 ;
  assign y9136 = ~1'b0 ;
  assign y9137 = ~1'b0 ;
  assign y9138 = ~1'b0 ;
  assign y9139 = ~n14726 ;
  assign y9140 = ~n14728 ;
  assign y9141 = ~1'b0 ;
  assign y9142 = n14729 ;
  assign y9143 = n14731 ;
  assign y9144 = ~1'b0 ;
  assign y9145 = n14736 ;
  assign y9146 = ~n14737 ;
  assign y9147 = ~n14742 ;
  assign y9148 = ~n14749 ;
  assign y9149 = ~n14751 ;
  assign y9150 = ~1'b0 ;
  assign y9151 = ~n14752 ;
  assign y9152 = n14753 ;
  assign y9153 = n14759 ;
  assign y9154 = ~n14760 ;
  assign y9155 = ~1'b0 ;
  assign y9156 = n14763 ;
  assign y9157 = ~n14764 ;
  assign y9158 = ~n14766 ;
  assign y9159 = ~n3398 ;
  assign y9160 = n14767 ;
  assign y9161 = 1'b0 ;
  assign y9162 = ~n14772 ;
  assign y9163 = ~1'b0 ;
  assign y9164 = ~1'b0 ;
  assign y9165 = n14774 ;
  assign y9166 = ~1'b0 ;
  assign y9167 = ~n14782 ;
  assign y9168 = n14785 ;
  assign y9169 = 1'b0 ;
  assign y9170 = n14786 ;
  assign y9171 = ~1'b0 ;
  assign y9172 = ~1'b0 ;
  assign y9173 = 1'b0 ;
  assign y9174 = ~n14787 ;
  assign y9175 = ~n4241 ;
  assign y9176 = ~n9412 ;
  assign y9177 = ~1'b0 ;
  assign y9178 = ~1'b0 ;
  assign y9179 = ~n14788 ;
  assign y9180 = n14791 ;
  assign y9181 = n14795 ;
  assign y9182 = ~1'b0 ;
  assign y9183 = ~n10386 ;
  assign y9184 = n173 ;
  assign y9185 = ~n14797 ;
  assign y9186 = ~n14798 ;
  assign y9187 = n14799 ;
  assign y9188 = ~1'b0 ;
  assign y9189 = ~n14800 ;
  assign y9190 = ~1'b0 ;
  assign y9191 = ~1'b0 ;
  assign y9192 = ~1'b0 ;
  assign y9193 = ~1'b0 ;
  assign y9194 = n14801 ;
  assign y9195 = ~1'b0 ;
  assign y9196 = ~1'b0 ;
  assign y9197 = ~1'b0 ;
  assign y9198 = ~1'b0 ;
  assign y9199 = n14809 ;
  assign y9200 = ~n14814 ;
  assign y9201 = ~1'b0 ;
  assign y9202 = ~n14816 ;
  assign y9203 = ~n13693 ;
  assign y9204 = n14818 ;
  assign y9205 = n14821 ;
  assign y9206 = ~1'b0 ;
  assign y9207 = ~n14822 ;
  assign y9208 = n14823 ;
  assign y9209 = ~1'b0 ;
  assign y9210 = ~n14824 ;
  assign y9211 = ~n14825 ;
  assign y9212 = ~1'b0 ;
  assign y9213 = ~n14826 ;
  assign y9214 = n14830 ;
  assign y9215 = n14834 ;
  assign y9216 = ~1'b0 ;
  assign y9217 = n14835 ;
  assign y9218 = ~1'b0 ;
  assign y9219 = ~1'b0 ;
  assign y9220 = ~1'b0 ;
  assign y9221 = n14841 ;
  assign y9222 = n14842 ;
  assign y9223 = n14843 ;
  assign y9224 = ~n2255 ;
  assign y9225 = ~n14844 ;
  assign y9226 = n14845 ;
  assign y9227 = ~1'b0 ;
  assign y9228 = n5819 ;
  assign y9229 = n14847 ;
  assign y9230 = ~1'b0 ;
  assign y9231 = n14848 ;
  assign y9232 = n14849 ;
  assign y9233 = 1'b0 ;
  assign y9234 = 1'b0 ;
  assign y9235 = ~n14851 ;
  assign y9236 = n14853 ;
  assign y9237 = ~n14854 ;
  assign y9238 = ~1'b0 ;
  assign y9239 = ~1'b0 ;
  assign y9240 = ~1'b0 ;
  assign y9241 = ~n14855 ;
  assign y9242 = ~1'b0 ;
  assign y9243 = ~n14856 ;
  assign y9244 = ~n14863 ;
  assign y9245 = n14866 ;
  assign y9246 = n14869 ;
  assign y9247 = ~n14873 ;
  assign y9248 = n14874 ;
  assign y9249 = n14876 ;
  assign y9250 = ~1'b0 ;
  assign y9251 = n14878 ;
  assign y9252 = n14880 ;
  assign y9253 = ~1'b0 ;
  assign y9254 = ~1'b0 ;
  assign y9255 = ~1'b0 ;
  assign y9256 = ~1'b0 ;
  assign y9257 = ~n14882 ;
  assign y9258 = ~1'b0 ;
  assign y9259 = ~n14884 ;
  assign y9260 = ~1'b0 ;
  assign y9261 = ~n14891 ;
  assign y9262 = ~1'b0 ;
  assign y9263 = ~n14895 ;
  assign y9264 = n7803 ;
  assign y9265 = n14896 ;
  assign y9266 = ~n14908 ;
  assign y9267 = ~1'b0 ;
  assign y9268 = ~n14909 ;
  assign y9269 = ~n14911 ;
  assign y9270 = ~1'b0 ;
  assign y9271 = n14916 ;
  assign y9272 = ~n14917 ;
  assign y9273 = ~1'b0 ;
  assign y9274 = ~n14919 ;
  assign y9275 = n14920 ;
  assign y9276 = ~n3210 ;
  assign y9277 = ~n14921 ;
  assign y9278 = 1'b0 ;
  assign y9279 = n211 ;
  assign y9280 = n14923 ;
  assign y9281 = ~n3256 ;
  assign y9282 = ~1'b0 ;
  assign y9283 = n14924 ;
  assign y9284 = ~1'b0 ;
  assign y9285 = ~n14927 ;
  assign y9286 = ~n14931 ;
  assign y9287 = ~n14935 ;
  assign y9288 = ~1'b0 ;
  assign y9289 = ~1'b0 ;
  assign y9290 = ~n3805 ;
  assign y9291 = n11116 ;
  assign y9292 = ~1'b0 ;
  assign y9293 = 1'b0 ;
  assign y9294 = ~1'b0 ;
  assign y9295 = n14937 ;
  assign y9296 = ~n14939 ;
  assign y9297 = n14946 ;
  assign y9298 = ~n14949 ;
  assign y9299 = ~n14953 ;
  assign y9300 = n14954 ;
  assign y9301 = n14955 ;
  assign y9302 = ~1'b0 ;
  assign y9303 = ~n14956 ;
  assign y9304 = ~n14962 ;
  assign y9305 = ~1'b0 ;
  assign y9306 = ~n14963 ;
  assign y9307 = ~n14964 ;
  assign y9308 = ~1'b0 ;
  assign y9309 = n14968 ;
  assign y9310 = ~n14971 ;
  assign y9311 = ~n14973 ;
  assign y9312 = ~n14976 ;
  assign y9313 = 1'b0 ;
  assign y9314 = ~1'b0 ;
  assign y9315 = ~1'b0 ;
  assign y9316 = n14977 ;
  assign y9317 = ~1'b0 ;
  assign y9318 = ~1'b0 ;
  assign y9319 = ~1'b0 ;
  assign y9320 = ~n14982 ;
  assign y9321 = n14985 ;
  assign y9322 = n14986 ;
  assign y9323 = ~1'b0 ;
  assign y9324 = ~1'b0 ;
  assign y9325 = ~1'b0 ;
  assign y9326 = ~n14989 ;
  assign y9327 = n14992 ;
  assign y9328 = ~1'b0 ;
  assign y9329 = ~n14997 ;
  assign y9330 = 1'b0 ;
  assign y9331 = ~n14999 ;
  assign y9332 = ~n15000 ;
  assign y9333 = ~n15007 ;
  assign y9334 = n15008 ;
  assign y9335 = ~1'b0 ;
  assign y9336 = ~1'b0 ;
  assign y9337 = ~n15009 ;
  assign y9338 = ~n15013 ;
  assign y9339 = n4929 ;
  assign y9340 = ~1'b0 ;
  assign y9341 = ~n15014 ;
  assign y9342 = ~n15016 ;
  assign y9343 = n15018 ;
  assign y9344 = ~1'b0 ;
  assign y9345 = ~n5913 ;
  assign y9346 = ~n15020 ;
  assign y9347 = n15022 ;
  assign y9348 = n15023 ;
  assign y9349 = 1'b0 ;
  assign y9350 = n15025 ;
  assign y9351 = ~n15033 ;
  assign y9352 = ~n15036 ;
  assign y9353 = n15038 ;
  assign y9354 = n14842 ;
  assign y9355 = ~n15043 ;
  assign y9356 = n15044 ;
  assign y9357 = n15046 ;
  assign y9358 = n15047 ;
  assign y9359 = n15049 ;
  assign y9360 = ~1'b0 ;
  assign y9361 = ~n1848 ;
  assign y9362 = n15050 ;
  assign y9363 = ~n15060 ;
  assign y9364 = ~1'b0 ;
  assign y9365 = n15063 ;
  assign y9366 = ~n15065 ;
  assign y9367 = ~1'b0 ;
  assign y9368 = n15067 ;
  assign y9369 = ~n15068 ;
  assign y9370 = ~1'b0 ;
  assign y9371 = ~n15077 ;
  assign y9372 = ~1'b0 ;
  assign y9373 = ~1'b0 ;
  assign y9374 = ~n15079 ;
  assign y9375 = n15082 ;
  assign y9376 = ~1'b0 ;
  assign y9377 = ~n15085 ;
  assign y9378 = ~1'b0 ;
  assign y9379 = ~1'b0 ;
  assign y9380 = ~1'b0 ;
  assign y9381 = ~1'b0 ;
  assign y9382 = ~1'b0 ;
  assign y9383 = n15089 ;
  assign y9384 = n15093 ;
  assign y9385 = ~n15094 ;
  assign y9386 = n15098 ;
  assign y9387 = n15099 ;
  assign y9388 = n15100 ;
  assign y9389 = ~1'b0 ;
  assign y9390 = 1'b0 ;
  assign y9391 = ~1'b0 ;
  assign y9392 = ~n15104 ;
  assign y9393 = ~n15105 ;
  assign y9394 = ~1'b0 ;
  assign y9395 = ~1'b0 ;
  assign y9396 = n444 ;
  assign y9397 = ~1'b0 ;
  assign y9398 = ~n15110 ;
  assign y9399 = ~n15111 ;
  assign y9400 = ~n15114 ;
  assign y9401 = ~n15115 ;
  assign y9402 = ~n15118 ;
  assign y9403 = n15121 ;
  assign y9404 = ~n15122 ;
  assign y9405 = ~1'b0 ;
  assign y9406 = ~n15123 ;
  assign y9407 = ~1'b0 ;
  assign y9408 = n15124 ;
  assign y9409 = ~1'b0 ;
  assign y9410 = ~1'b0 ;
  assign y9411 = n5214 ;
  assign y9412 = ~1'b0 ;
  assign y9413 = ~n11464 ;
  assign y9414 = n15125 ;
  assign y9415 = n571 ;
  assign y9416 = n11846 ;
  assign y9417 = n15127 ;
  assign y9418 = n15129 ;
  assign y9419 = ~1'b0 ;
  assign y9420 = ~n15130 ;
  assign y9421 = ~n15133 ;
  assign y9422 = ~1'b0 ;
  assign y9423 = ~n15139 ;
  assign y9424 = ~n15141 ;
  assign y9425 = ~n15142 ;
  assign y9426 = ~n15148 ;
  assign y9427 = n15151 ;
  assign y9428 = ~1'b0 ;
  assign y9429 = ~n15153 ;
  assign y9430 = ~n15155 ;
  assign y9431 = n15157 ;
  assign y9432 = ~n15160 ;
  assign y9433 = n15161 ;
  assign y9434 = ~n15162 ;
  assign y9435 = n15164 ;
  assign y9436 = ~n5367 ;
  assign y9437 = n15166 ;
  assign y9438 = n15168 ;
  assign y9439 = ~n15169 ;
  assign y9440 = ~n15171 ;
  assign y9441 = ~n15173 ;
  assign y9442 = ~n15175 ;
  assign y9443 = ~1'b0 ;
  assign y9444 = ~n15178 ;
  assign y9445 = ~n15180 ;
  assign y9446 = n15183 ;
  assign y9447 = ~1'b0 ;
  assign y9448 = n15185 ;
  assign y9449 = ~1'b0 ;
  assign y9450 = n15186 ;
  assign y9451 = ~1'b0 ;
  assign y9452 = n15190 ;
  assign y9453 = ~n15191 ;
  assign y9454 = n846 ;
  assign y9455 = n15194 ;
  assign y9456 = n15196 ;
  assign y9457 = ~n15203 ;
  assign y9458 = ~1'b0 ;
  assign y9459 = n15204 ;
  assign y9460 = ~1'b0 ;
  assign y9461 = ~n15209 ;
  assign y9462 = n15211 ;
  assign y9463 = 1'b0 ;
  assign y9464 = 1'b0 ;
  assign y9465 = ~n15213 ;
  assign y9466 = 1'b0 ;
  assign y9467 = ~n15214 ;
  assign y9468 = ~1'b0 ;
  assign y9469 = ~1'b0 ;
  assign y9470 = x63 ;
  assign y9471 = ~1'b0 ;
  assign y9472 = ~1'b0 ;
  assign y9473 = ~1'b0 ;
  assign y9474 = n2481 ;
  assign y9475 = n15215 ;
  assign y9476 = ~1'b0 ;
  assign y9477 = n15217 ;
  assign y9478 = ~1'b0 ;
  assign y9479 = ~1'b0 ;
  assign y9480 = n15227 ;
  assign y9481 = ~1'b0 ;
  assign y9482 = ~n15229 ;
  assign y9483 = n15234 ;
  assign y9484 = n15238 ;
  assign y9485 = n15242 ;
  assign y9486 = ~1'b0 ;
  assign y9487 = ~1'b0 ;
  assign y9488 = ~1'b0 ;
  assign y9489 = 1'b0 ;
  assign y9490 = n15245 ;
  assign y9491 = n15246 ;
  assign y9492 = ~1'b0 ;
  assign y9493 = n15248 ;
  assign y9494 = n15251 ;
  assign y9495 = n15256 ;
  assign y9496 = ~1'b0 ;
  assign y9497 = ~1'b0 ;
  assign y9498 = n15261 ;
  assign y9499 = n15264 ;
  assign y9500 = n15265 ;
  assign y9501 = n15266 ;
  assign y9502 = ~1'b0 ;
  assign y9503 = ~n15270 ;
  assign y9504 = ~1'b0 ;
  assign y9505 = ~1'b0 ;
  assign y9506 = n5687 ;
  assign y9507 = ~n15271 ;
  assign y9508 = n15274 ;
  assign y9509 = ~1'b0 ;
  assign y9510 = ~1'b0 ;
  assign y9511 = n15276 ;
  assign y9512 = ~1'b0 ;
  assign y9513 = n15278 ;
  assign y9514 = n15283 ;
  assign y9515 = ~n15284 ;
  assign y9516 = ~1'b0 ;
  assign y9517 = n15285 ;
  assign y9518 = ~n15286 ;
  assign y9519 = ~1'b0 ;
  assign y9520 = n15288 ;
  assign y9521 = n15291 ;
  assign y9522 = ~1'b0 ;
  assign y9523 = ~n15292 ;
  assign y9524 = ~1'b0 ;
  assign y9525 = ~1'b0 ;
  assign y9526 = n15294 ;
  assign y9527 = ~n15298 ;
  assign y9528 = ~n15299 ;
  assign y9529 = n10530 ;
  assign y9530 = ~n15300 ;
  assign y9531 = ~n13909 ;
  assign y9532 = ~n15303 ;
  assign y9533 = ~n15304 ;
  assign y9534 = ~1'b0 ;
  assign y9535 = ~n15305 ;
  assign y9536 = ~1'b0 ;
  assign y9537 = ~1'b0 ;
  assign y9538 = n1724 ;
  assign y9539 = ~1'b0 ;
  assign y9540 = n15307 ;
  assign y9541 = ~n15311 ;
  assign y9542 = n11856 ;
  assign y9543 = ~1'b0 ;
  assign y9544 = ~n15317 ;
  assign y9545 = n15318 ;
  assign y9546 = n9047 ;
  assign y9547 = n15320 ;
  assign y9548 = ~n15322 ;
  assign y9549 = n15324 ;
  assign y9550 = n15326 ;
  assign y9551 = ~1'b0 ;
  assign y9552 = ~1'b0 ;
  assign y9553 = ~n13182 ;
  assign y9554 = ~1'b0 ;
  assign y9555 = ~n15328 ;
  assign y9556 = n15333 ;
  assign y9557 = n15336 ;
  assign y9558 = n15337 ;
  assign y9559 = ~n15338 ;
  assign y9560 = n15339 ;
  assign y9561 = n15343 ;
  assign y9562 = ~n15347 ;
  assign y9563 = n15351 ;
  assign y9564 = ~n15355 ;
  assign y9565 = n15358 ;
  assign y9566 = ~1'b0 ;
  assign y9567 = ~1'b0 ;
  assign y9568 = n15359 ;
  assign y9569 = n15360 ;
  assign y9570 = n15361 ;
  assign y9571 = ~1'b0 ;
  assign y9572 = n15363 ;
  assign y9573 = ~1'b0 ;
  assign y9574 = ~n15366 ;
  assign y9575 = n15367 ;
  assign y9576 = ~1'b0 ;
  assign y9577 = ~n15369 ;
  assign y9578 = ~n15371 ;
  assign y9579 = n15375 ;
  assign y9580 = ~1'b0 ;
  assign y9581 = ~n15378 ;
  assign y9582 = ~n15379 ;
  assign y9583 = ~1'b0 ;
  assign y9584 = 1'b0 ;
  assign y9585 = ~n15382 ;
  assign y9586 = ~1'b0 ;
  assign y9587 = ~1'b0 ;
  assign y9588 = ~1'b0 ;
  assign y9589 = n15383 ;
  assign y9590 = ~n15384 ;
  assign y9591 = n15398 ;
  assign y9592 = ~1'b0 ;
  assign y9593 = n15400 ;
  assign y9594 = ~n15401 ;
  assign y9595 = ~n15404 ;
  assign y9596 = n15406 ;
  assign y9597 = 1'b0 ;
  assign y9598 = ~n2166 ;
  assign y9599 = n15408 ;
  assign y9600 = ~1'b0 ;
  assign y9601 = ~1'b0 ;
  assign y9602 = ~1'b0 ;
  assign y9603 = ~n15410 ;
  assign y9604 = n15412 ;
  assign y9605 = ~1'b0 ;
  assign y9606 = n3947 ;
  assign y9607 = ~n7453 ;
  assign y9608 = ~n7653 ;
  assign y9609 = n15414 ;
  assign y9610 = n2497 ;
  assign y9611 = ~n15415 ;
  assign y9612 = ~1'b0 ;
  assign y9613 = n15416 ;
  assign y9614 = ~n15418 ;
  assign y9615 = ~n15421 ;
  assign y9616 = ~1'b0 ;
  assign y9617 = 1'b0 ;
  assign y9618 = n15426 ;
  assign y9619 = ~1'b0 ;
  assign y9620 = ~1'b0 ;
  assign y9621 = ~1'b0 ;
  assign y9622 = n15427 ;
  assign y9623 = ~1'b0 ;
  assign y9624 = 1'b0 ;
  assign y9625 = ~n8509 ;
  assign y9626 = ~1'b0 ;
  assign y9627 = ~1'b0 ;
  assign y9628 = 1'b0 ;
  assign y9629 = ~n15429 ;
  assign y9630 = ~1'b0 ;
  assign y9631 = ~1'b0 ;
  assign y9632 = ~n15432 ;
  assign y9633 = ~1'b0 ;
  assign y9634 = ~1'b0 ;
  assign y9635 = ~1'b0 ;
  assign y9636 = ~n8398 ;
  assign y9637 = n15436 ;
  assign y9638 = ~1'b0 ;
  assign y9639 = n15441 ;
  assign y9640 = ~n15450 ;
  assign y9641 = ~n15454 ;
  assign y9642 = ~n15463 ;
  assign y9643 = ~1'b0 ;
  assign y9644 = n15465 ;
  assign y9645 = ~1'b0 ;
  assign y9646 = ~1'b0 ;
  assign y9647 = n15467 ;
  assign y9648 = n15468 ;
  assign y9649 = n15469 ;
  assign y9650 = 1'b0 ;
  assign y9651 = 1'b0 ;
  assign y9652 = ~n15471 ;
  assign y9653 = ~1'b0 ;
  assign y9654 = ~1'b0 ;
  assign y9655 = ~n15473 ;
  assign y9656 = ~1'b0 ;
  assign y9657 = ~n15474 ;
  assign y9658 = ~n15476 ;
  assign y9659 = n15478 ;
  assign y9660 = ~1'b0 ;
  assign y9661 = ~n15480 ;
  assign y9662 = n15482 ;
  assign y9663 = n15484 ;
  assign y9664 = n15486 ;
  assign y9665 = ~n15488 ;
  assign y9666 = 1'b0 ;
  assign y9667 = 1'b0 ;
  assign y9668 = ~n15489 ;
  assign y9669 = ~n15491 ;
  assign y9670 = ~1'b0 ;
  assign y9671 = n15494 ;
  assign y9672 = ~1'b0 ;
  assign y9673 = ~n15495 ;
  assign y9674 = ~1'b0 ;
  assign y9675 = n15500 ;
  assign y9676 = ~n15506 ;
  assign y9677 = ~n15512 ;
  assign y9678 = ~1'b0 ;
  assign y9679 = ~1'b0 ;
  assign y9680 = n15514 ;
  assign y9681 = ~n15516 ;
  assign y9682 = n15518 ;
  assign y9683 = ~1'b0 ;
  assign y9684 = ~n15522 ;
  assign y9685 = n15523 ;
  assign y9686 = ~1'b0 ;
  assign y9687 = ~n15525 ;
  assign y9688 = ~1'b0 ;
  assign y9689 = ~n15526 ;
  assign y9690 = ~n15529 ;
  assign y9691 = ~1'b0 ;
  assign y9692 = ~n15550 ;
  assign y9693 = ~1'b0 ;
  assign y9694 = ~1'b0 ;
  assign y9695 = n15551 ;
  assign y9696 = ~n15552 ;
  assign y9697 = ~1'b0 ;
  assign y9698 = ~n15553 ;
  assign y9699 = n1564 ;
  assign y9700 = ~1'b0 ;
  assign y9701 = ~1'b0 ;
  assign y9702 = n15555 ;
  assign y9703 = ~1'b0 ;
  assign y9704 = ~1'b0 ;
  assign y9705 = ~1'b0 ;
  assign y9706 = ~n3624 ;
  assign y9707 = n15556 ;
  assign y9708 = n15557 ;
  assign y9709 = n15559 ;
  assign y9710 = ~1'b0 ;
  assign y9711 = n15560 ;
  assign y9712 = ~1'b0 ;
  assign y9713 = ~n15564 ;
  assign y9714 = n15567 ;
  assign y9715 = ~1'b0 ;
  assign y9716 = ~n15568 ;
  assign y9717 = ~1'b0 ;
  assign y9718 = ~n1867 ;
  assign y9719 = n15571 ;
  assign y9720 = ~1'b0 ;
  assign y9721 = ~1'b0 ;
  assign y9722 = ~n12609 ;
  assign y9723 = 1'b0 ;
  assign y9724 = n15572 ;
  assign y9725 = n15574 ;
  assign y9726 = n15576 ;
  assign y9727 = ~n15578 ;
  assign y9728 = ~1'b0 ;
  assign y9729 = ~n15579 ;
  assign y9730 = ~1'b0 ;
  assign y9731 = ~1'b0 ;
  assign y9732 = n15580 ;
  assign y9733 = n15581 ;
  assign y9734 = 1'b0 ;
  assign y9735 = ~n15584 ;
  assign y9736 = ~n15585 ;
  assign y9737 = ~n15587 ;
  assign y9738 = n15588 ;
  assign y9739 = ~1'b0 ;
  assign y9740 = ~n15590 ;
  assign y9741 = n15592 ;
  assign y9742 = n15593 ;
  assign y9743 = n15594 ;
  assign y9744 = ~1'b0 ;
  assign y9745 = n15596 ;
  assign y9746 = ~n2425 ;
  assign y9747 = n8125 ;
  assign y9748 = ~n15598 ;
  assign y9749 = ~n15599 ;
  assign y9750 = n15602 ;
  assign y9751 = ~1'b0 ;
  assign y9752 = n6077 ;
  assign y9753 = ~n15603 ;
  assign y9754 = ~1'b0 ;
  assign y9755 = n15607 ;
  assign y9756 = ~1'b0 ;
  assign y9757 = ~n15612 ;
  assign y9758 = ~n15613 ;
  assign y9759 = ~1'b0 ;
  assign y9760 = n15617 ;
  assign y9761 = ~n15618 ;
  assign y9762 = n15621 ;
  assign y9763 = ~n15624 ;
  assign y9764 = ~1'b0 ;
  assign y9765 = n15626 ;
  assign y9766 = n15627 ;
  assign y9767 = 1'b0 ;
  assign y9768 = ~1'b0 ;
  assign y9769 = ~1'b0 ;
  assign y9770 = ~1'b0 ;
  assign y9771 = ~n15628 ;
  assign y9772 = n15630 ;
  assign y9773 = n652 ;
  assign y9774 = ~n15635 ;
  assign y9775 = ~1'b0 ;
  assign y9776 = n15637 ;
  assign y9777 = ~1'b0 ;
  assign y9778 = ~1'b0 ;
  assign y9779 = ~1'b0 ;
  assign y9780 = ~n15638 ;
  assign y9781 = n15641 ;
  assign y9782 = ~n15643 ;
  assign y9783 = n15647 ;
  assign y9784 = ~n2692 ;
  assign y9785 = ~n15648 ;
  assign y9786 = ~n15650 ;
  assign y9787 = n15651 ;
  assign y9788 = ~n15654 ;
  assign y9789 = ~1'b0 ;
  assign y9790 = ~n15407 ;
  assign y9791 = ~n15655 ;
  assign y9792 = ~1'b0 ;
  assign y9793 = ~n15658 ;
  assign y9794 = n15659 ;
  assign y9795 = n15661 ;
  assign y9796 = 1'b0 ;
  assign y9797 = ~n4444 ;
  assign y9798 = ~1'b0 ;
  assign y9799 = ~n15662 ;
  assign y9800 = ~n15664 ;
  assign y9801 = ~n15666 ;
  assign y9802 = ~1'b0 ;
  assign y9803 = ~1'b0 ;
  assign y9804 = 1'b0 ;
  assign y9805 = ~n4882 ;
  assign y9806 = ~1'b0 ;
  assign y9807 = 1'b0 ;
  assign y9808 = n526 ;
  assign y9809 = ~1'b0 ;
  assign y9810 = ~1'b0 ;
  assign y9811 = ~1'b0 ;
  assign y9812 = ~1'b0 ;
  assign y9813 = ~n15672 ;
  assign y9814 = ~1'b0 ;
  assign y9815 = ~n15675 ;
  assign y9816 = n15676 ;
  assign y9817 = ~1'b0 ;
  assign y9818 = ~n753 ;
  assign y9819 = ~1'b0 ;
  assign y9820 = ~1'b0 ;
  assign y9821 = 1'b0 ;
  assign y9822 = 1'b0 ;
  assign y9823 = ~1'b0 ;
  assign y9824 = ~n15677 ;
  assign y9825 = ~n15678 ;
  assign y9826 = ~1'b0 ;
  assign y9827 = ~n3359 ;
  assign y9828 = ~1'b0 ;
  assign y9829 = n15679 ;
  assign y9830 = ~1'b0 ;
  assign y9831 = n15680 ;
  assign y9832 = ~1'b0 ;
  assign y9833 = 1'b0 ;
  assign y9834 = n15684 ;
  assign y9835 = ~1'b0 ;
  assign y9836 = ~1'b0 ;
  assign y9837 = n15687 ;
  assign y9838 = ~n15689 ;
  assign y9839 = n15690 ;
  assign y9840 = ~1'b0 ;
  assign y9841 = 1'b0 ;
  assign y9842 = ~n15694 ;
  assign y9843 = ~1'b0 ;
  assign y9844 = n15695 ;
  assign y9845 = n5255 ;
  assign y9846 = ~n15697 ;
  assign y9847 = n15698 ;
  assign y9848 = ~n4377 ;
  assign y9849 = n15702 ;
  assign y9850 = ~n15705 ;
  assign y9851 = ~1'b0 ;
  assign y9852 = n15708 ;
  assign y9853 = ~n15710 ;
  assign y9854 = n15716 ;
  assign y9855 = ~1'b0 ;
  assign y9856 = n1324 ;
  assign y9857 = n15717 ;
  assign y9858 = n15719 ;
  assign y9859 = ~1'b0 ;
  assign y9860 = ~1'b0 ;
  assign y9861 = ~1'b0 ;
  assign y9862 = ~1'b0 ;
  assign y9863 = ~1'b0 ;
  assign y9864 = n15721 ;
  assign y9865 = ~n15722 ;
  assign y9866 = ~1'b0 ;
  assign y9867 = n15725 ;
  assign y9868 = ~1'b0 ;
  assign y9869 = ~n15727 ;
  assign y9870 = ~n15728 ;
  assign y9871 = n15729 ;
  assign y9872 = ~n15731 ;
  assign y9873 = ~1'b0 ;
  assign y9874 = n15732 ;
  assign y9875 = ~1'b0 ;
  assign y9876 = ~n15735 ;
  assign y9877 = ~n15742 ;
  assign y9878 = ~1'b0 ;
  assign y9879 = ~1'b0 ;
  assign y9880 = n15744 ;
  assign y9881 = n15746 ;
  assign y9882 = n8283 ;
  assign y9883 = ~n15747 ;
  assign y9884 = ~1'b0 ;
  assign y9885 = ~n15750 ;
  assign y9886 = n15753 ;
  assign y9887 = ~1'b0 ;
  assign y9888 = ~1'b0 ;
  assign y9889 = ~1'b0 ;
  assign y9890 = n15755 ;
  assign y9891 = ~1'b0 ;
  assign y9892 = ~1'b0 ;
  assign y9893 = ~n15756 ;
  assign y9894 = ~1'b0 ;
  assign y9895 = ~1'b0 ;
  assign y9896 = ~n15759 ;
  assign y9897 = n15762 ;
  assign y9898 = ~1'b0 ;
  assign y9899 = n15768 ;
  assign y9900 = ~1'b0 ;
  assign y9901 = ~1'b0 ;
  assign y9902 = n15769 ;
  assign y9903 = n15770 ;
  assign y9904 = 1'b0 ;
  assign y9905 = ~n15771 ;
  assign y9906 = n15772 ;
  assign y9907 = n15773 ;
  assign y9908 = n15775 ;
  assign y9909 = ~n15779 ;
  assign y9910 = n15780 ;
  assign y9911 = ~1'b0 ;
  assign y9912 = ~1'b0 ;
  assign y9913 = n15782 ;
  assign y9914 = n15783 ;
  assign y9915 = ~n15786 ;
  assign y9916 = ~1'b0 ;
  assign y9917 = n15788 ;
  assign y9918 = n15789 ;
  assign y9919 = n15790 ;
  assign y9920 = ~1'b0 ;
  assign y9921 = ~1'b0 ;
  assign y9922 = n15791 ;
  assign y9923 = ~1'b0 ;
  assign y9924 = ~n2115 ;
  assign y9925 = n15795 ;
  assign y9926 = n15799 ;
  assign y9927 = n7394 ;
  assign y9928 = n15801 ;
  assign y9929 = x112 ;
  assign y9930 = n15806 ;
  assign y9931 = ~1'b0 ;
  assign y9932 = ~1'b0 ;
  assign y9933 = ~1'b0 ;
  assign y9934 = ~1'b0 ;
  assign y9935 = ~1'b0 ;
  assign y9936 = ~n15807 ;
  assign y9937 = ~n15808 ;
  assign y9938 = n15810 ;
  assign y9939 = ~n15812 ;
  assign y9940 = n15814 ;
  assign y9941 = 1'b0 ;
  assign y9942 = n15820 ;
  assign y9943 = ~1'b0 ;
  assign y9944 = ~n10065 ;
  assign y9945 = n15823 ;
  assign y9946 = 1'b0 ;
  assign y9947 = ~n15824 ;
  assign y9948 = n15826 ;
  assign y9949 = n15828 ;
  assign y9950 = ~n9823 ;
  assign y9951 = ~n15832 ;
  assign y9952 = n15836 ;
  assign y9953 = n15844 ;
  assign y9954 = ~n15846 ;
  assign y9955 = ~n15848 ;
  assign y9956 = ~n15851 ;
  assign y9957 = ~1'b0 ;
  assign y9958 = ~1'b0 ;
  assign y9959 = n15852 ;
  assign y9960 = ~n15858 ;
  assign y9961 = n15859 ;
  assign y9962 = n15861 ;
  assign y9963 = ~1'b0 ;
  assign y9964 = 1'b0 ;
  assign y9965 = ~n15866 ;
  assign y9966 = n15869 ;
  assign y9967 = ~n15870 ;
  assign y9968 = ~1'b0 ;
  assign y9969 = n15872 ;
  assign y9970 = ~n15878 ;
  assign y9971 = ~1'b0 ;
  assign y9972 = ~1'b0 ;
  assign y9973 = ~n14368 ;
  assign y9974 = ~1'b0 ;
  assign y9975 = n15880 ;
  assign y9976 = ~n571 ;
  assign y9977 = n15882 ;
  assign y9978 = ~n5100 ;
  assign y9979 = n15883 ;
  assign y9980 = ~1'b0 ;
  assign y9981 = ~n15884 ;
  assign y9982 = ~1'b0 ;
  assign y9983 = ~1'b0 ;
  assign y9984 = n15886 ;
  assign y9985 = n15889 ;
  assign y9986 = ~n15892 ;
  assign y9987 = n15895 ;
  assign y9988 = ~n15897 ;
  assign y9989 = ~1'b0 ;
  assign y9990 = ~1'b0 ;
  assign y9991 = ~1'b0 ;
  assign y9992 = ~n15902 ;
  assign y9993 = 1'b0 ;
  assign y9994 = n15904 ;
  assign y9995 = ~n15906 ;
  assign y9996 = ~1'b0 ;
  assign y9997 = ~1'b0 ;
  assign y9998 = n415 ;
  assign y9999 = ~1'b0 ;
  assign y10000 = n15909 ;
  assign y10001 = ~n15912 ;
  assign y10002 = ~1'b0 ;
  assign y10003 = 1'b0 ;
  assign y10004 = ~1'b0 ;
  assign y10005 = 1'b0 ;
  assign y10006 = ~1'b0 ;
  assign y10007 = ~n15913 ;
  assign y10008 = ~n15916 ;
  assign y10009 = ~1'b0 ;
  assign y10010 = n15919 ;
  assign y10011 = ~n15921 ;
  assign y10012 = n15922 ;
  assign y10013 = n15923 ;
  assign y10014 = ~n15927 ;
  assign y10015 = n15931 ;
  assign y10016 = n15933 ;
  assign y10017 = ~n15935 ;
  assign y10018 = n15939 ;
  assign y10019 = ~n15944 ;
  assign y10020 = ~1'b0 ;
  assign y10021 = ~1'b0 ;
  assign y10022 = n15947 ;
  assign y10023 = ~n15949 ;
  assign y10024 = n8062 ;
  assign y10025 = ~n15950 ;
  assign y10026 = ~1'b0 ;
  assign y10027 = ~1'b0 ;
  assign y10028 = n15951 ;
  assign y10029 = ~1'b0 ;
  assign y10030 = ~n15953 ;
  assign y10031 = n2053 ;
  assign y10032 = n9904 ;
  assign y10033 = ~n15956 ;
  assign y10034 = n15959 ;
  assign y10035 = ~n6581 ;
  assign y10036 = n15960 ;
  assign y10037 = ~1'b0 ;
  assign y10038 = ~1'b0 ;
  assign y10039 = ~n15961 ;
  assign y10040 = ~n15964 ;
  assign y10041 = ~n2713 ;
  assign y10042 = 1'b0 ;
  assign y10043 = ~n15967 ;
  assign y10044 = n15969 ;
  assign y10045 = n354 ;
  assign y10046 = ~1'b0 ;
  assign y10047 = ~1'b0 ;
  assign y10048 = ~n15977 ;
  assign y10049 = n15982 ;
  assign y10050 = n15983 ;
  assign y10051 = ~n15984 ;
  assign y10052 = ~n15985 ;
  assign y10053 = n15989 ;
  assign y10054 = ~1'b0 ;
  assign y10055 = ~n986 ;
  assign y10056 = ~1'b0 ;
  assign y10057 = n15991 ;
  assign y10058 = ~n11663 ;
  assign y10059 = ~n15994 ;
  assign y10060 = ~n12324 ;
  assign y10061 = ~1'b0 ;
  assign y10062 = n15998 ;
  assign y10063 = ~1'b0 ;
  assign y10064 = ~1'b0 ;
  assign y10065 = ~n15999 ;
  assign y10066 = ~1'b0 ;
  assign y10067 = n16004 ;
  assign y10068 = n13270 ;
  assign y10069 = ~1'b0 ;
  assign y10070 = ~1'b0 ;
  assign y10071 = n16005 ;
  assign y10072 = n16007 ;
  assign y10073 = n16011 ;
  assign y10074 = n16012 ;
  assign y10075 = ~n16013 ;
  assign y10076 = ~1'b0 ;
  assign y10077 = ~n16015 ;
  assign y10078 = ~1'b0 ;
  assign y10079 = n16018 ;
  assign y10080 = ~n16022 ;
  assign y10081 = n8509 ;
  assign y10082 = ~1'b0 ;
  assign y10083 = ~1'b0 ;
  assign y10084 = n6933 ;
  assign y10085 = n16023 ;
  assign y10086 = n16024 ;
  assign y10087 = n16025 ;
  assign y10088 = ~1'b0 ;
  assign y10089 = n4882 ;
  assign y10090 = n16028 ;
  assign y10091 = ~n16029 ;
  assign y10092 = ~n2255 ;
  assign y10093 = ~1'b0 ;
  assign y10094 = ~1'b0 ;
  assign y10095 = n16030 ;
  assign y10096 = ~1'b0 ;
  assign y10097 = ~1'b0 ;
  assign y10098 = ~n16033 ;
  assign y10099 = n6217 ;
  assign y10100 = n1939 ;
  assign y10101 = n16034 ;
  assign y10102 = ~n16035 ;
  assign y10103 = ~n16036 ;
  assign y10104 = ~1'b0 ;
  assign y10105 = n375 ;
  assign y10106 = n16038 ;
  assign y10107 = n16042 ;
  assign y10108 = ~n16049 ;
  assign y10109 = ~1'b0 ;
  assign y10110 = ~n16052 ;
  assign y10111 = ~1'b0 ;
  assign y10112 = n16054 ;
  assign y10113 = 1'b0 ;
  assign y10114 = ~1'b0 ;
  assign y10115 = 1'b0 ;
  assign y10116 = n16055 ;
  assign y10117 = ~n16056 ;
  assign y10118 = ~1'b0 ;
  assign y10119 = ~n16058 ;
  assign y10120 = ~1'b0 ;
  assign y10121 = ~n4325 ;
  assign y10122 = ~n16063 ;
  assign y10123 = ~1'b0 ;
  assign y10124 = ~1'b0 ;
  assign y10125 = ~1'b0 ;
  assign y10126 = ~n16066 ;
  assign y10127 = n16067 ;
  assign y10128 = n16068 ;
  assign y10129 = ~n16070 ;
  assign y10130 = ~1'b0 ;
  assign y10131 = ~1'b0 ;
  assign y10132 = ~n16071 ;
  assign y10133 = ~n16073 ;
  assign y10134 = ~1'b0 ;
  assign y10135 = n16075 ;
  assign y10136 = n16078 ;
  assign y10137 = ~1'b0 ;
  assign y10138 = ~n16082 ;
  assign y10139 = ~n16083 ;
  assign y10140 = ~1'b0 ;
  assign y10141 = ~n16088 ;
  assign y10142 = ~n16090 ;
  assign y10143 = n13711 ;
  assign y10144 = ~1'b0 ;
  assign y10145 = 1'b0 ;
  assign y10146 = ~1'b0 ;
  assign y10147 = ~n16092 ;
  assign y10148 = ~n16095 ;
  assign y10149 = ~n16102 ;
  assign y10150 = ~1'b0 ;
  assign y10151 = ~1'b0 ;
  assign y10152 = ~1'b0 ;
  assign y10153 = ~n7735 ;
  assign y10154 = ~n16103 ;
  assign y10155 = ~1'b0 ;
  assign y10156 = ~1'b0 ;
  assign y10157 = ~1'b0 ;
  assign y10158 = n16104 ;
  assign y10159 = ~1'b0 ;
  assign y10160 = n11503 ;
  assign y10161 = ~1'b0 ;
  assign y10162 = ~1'b0 ;
  assign y10163 = n16106 ;
  assign y10164 = n16107 ;
  assign y10165 = ~n16110 ;
  assign y10166 = ~1'b0 ;
  assign y10167 = ~1'b0 ;
  assign y10168 = n16112 ;
  assign y10169 = n7668 ;
  assign y10170 = n16122 ;
  assign y10171 = ~n16125 ;
  assign y10172 = ~1'b0 ;
  assign y10173 = 1'b0 ;
  assign y10174 = n16126 ;
  assign y10175 = ~n16128 ;
  assign y10176 = n16129 ;
  assign y10177 = n16130 ;
  assign y10178 = ~n2561 ;
  assign y10179 = ~1'b0 ;
  assign y10180 = n16133 ;
  assign y10181 = n16134 ;
  assign y10182 = n1755 ;
  assign y10183 = n16138 ;
  assign y10184 = n16139 ;
  assign y10185 = ~1'b0 ;
  assign y10186 = ~1'b0 ;
  assign y10187 = ~n16140 ;
  assign y10188 = n4298 ;
  assign y10189 = 1'b0 ;
  assign y10190 = ~n1625 ;
  assign y10191 = n16144 ;
  assign y10192 = ~1'b0 ;
  assign y10193 = ~1'b0 ;
  assign y10194 = ~n16145 ;
  assign y10195 = n16148 ;
  assign y10196 = ~n16150 ;
  assign y10197 = ~n16151 ;
  assign y10198 = ~n16153 ;
  assign y10199 = n16155 ;
  assign y10200 = n16157 ;
  assign y10201 = ~n16158 ;
  assign y10202 = ~n16159 ;
  assign y10203 = ~1'b0 ;
  assign y10204 = ~1'b0 ;
  assign y10205 = ~n16163 ;
  assign y10206 = n5243 ;
  assign y10207 = ~n16166 ;
  assign y10208 = ~n16168 ;
  assign y10209 = ~n16170 ;
  assign y10210 = ~1'b0 ;
  assign y10211 = ~1'b0 ;
  assign y10212 = ~n16171 ;
  assign y10213 = ~1'b0 ;
  assign y10214 = ~n16172 ;
  assign y10215 = n16173 ;
  assign y10216 = ~1'b0 ;
  assign y10217 = ~1'b0 ;
  assign y10218 = ~1'b0 ;
  assign y10219 = ~n16176 ;
  assign y10220 = ~n16179 ;
  assign y10221 = ~n16180 ;
  assign y10222 = ~1'b0 ;
  assign y10223 = n16183 ;
  assign y10224 = n16185 ;
  assign y10225 = ~n16187 ;
  assign y10226 = n16188 ;
  assign y10227 = n16190 ;
  assign y10228 = ~1'b0 ;
  assign y10229 = n16191 ;
  assign y10230 = ~1'b0 ;
  assign y10231 = ~1'b0 ;
  assign y10232 = ~n983 ;
  assign y10233 = n16192 ;
  assign y10234 = n316 ;
  assign y10235 = n266 ;
  assign y10236 = ~n2427 ;
  assign y10237 = ~1'b0 ;
  assign y10238 = ~n8274 ;
  assign y10239 = n16193 ;
  assign y10240 = 1'b0 ;
  assign y10241 = ~n16194 ;
  assign y10242 = n16198 ;
  assign y10243 = n16204 ;
  assign y10244 = 1'b0 ;
  assign y10245 = ~n16205 ;
  assign y10246 = n12736 ;
  assign y10247 = n16207 ;
  assign y10248 = ~1'b0 ;
  assign y10249 = ~1'b0 ;
  assign y10250 = ~n16208 ;
  assign y10251 = n16211 ;
  assign y10252 = n16217 ;
  assign y10253 = n8462 ;
  assign y10254 = ~1'b0 ;
  assign y10255 = ~1'b0 ;
  assign y10256 = n2718 ;
  assign y10257 = n16218 ;
  assign y10258 = ~n16220 ;
  assign y10259 = ~1'b0 ;
  assign y10260 = ~n16221 ;
  assign y10261 = ~1'b0 ;
  assign y10262 = n16224 ;
  assign y10263 = n14399 ;
  assign y10264 = ~1'b0 ;
  assign y10265 = ~n16228 ;
  assign y10266 = n16229 ;
  assign y10267 = ~1'b0 ;
  assign y10268 = ~1'b0 ;
  assign y10269 = ~1'b0 ;
  assign y10270 = ~1'b0 ;
  assign y10271 = ~1'b0 ;
  assign y10272 = ~1'b0 ;
  assign y10273 = ~1'b0 ;
  assign y10274 = ~1'b0 ;
  assign y10275 = n3236 ;
  assign y10276 = ~1'b0 ;
  assign y10277 = ~1'b0 ;
  assign y10278 = ~n1724 ;
  assign y10279 = ~n16233 ;
  assign y10280 = ~n16234 ;
  assign y10281 = ~n16236 ;
  assign y10282 = ~n16237 ;
  assign y10283 = n16238 ;
  assign y10284 = n16240 ;
  assign y10285 = ~1'b0 ;
  assign y10286 = n16247 ;
  assign y10287 = n16248 ;
  assign y10288 = ~1'b0 ;
  assign y10289 = ~1'b0 ;
  assign y10290 = n16249 ;
  assign y10291 = ~1'b0 ;
  assign y10292 = ~n16250 ;
  assign y10293 = ~n16253 ;
  assign y10294 = n16254 ;
  assign y10295 = ~n13527 ;
  assign y10296 = ~1'b0 ;
  assign y10297 = n16256 ;
  assign y10298 = n16257 ;
  assign y10299 = ~1'b0 ;
  assign y10300 = ~n16259 ;
  assign y10301 = n14329 ;
  assign y10302 = n16261 ;
  assign y10303 = n3911 ;
  assign y10304 = ~1'b0 ;
  assign y10305 = n16265 ;
  assign y10306 = n16267 ;
  assign y10307 = ~n16269 ;
  assign y10308 = n16270 ;
  assign y10309 = ~n16272 ;
  assign y10310 = ~n16274 ;
  assign y10311 = ~n16275 ;
  assign y10312 = ~1'b0 ;
  assign y10313 = ~n16276 ;
  assign y10314 = ~1'b0 ;
  assign y10315 = ~1'b0 ;
  assign y10316 = ~n16280 ;
  assign y10317 = ~n16282 ;
  assign y10318 = n16284 ;
  assign y10319 = ~1'b0 ;
  assign y10320 = n16286 ;
  assign y10321 = 1'b0 ;
  assign y10322 = ~n16289 ;
  assign y10323 = n16290 ;
  assign y10324 = ~n16296 ;
  assign y10325 = ~1'b0 ;
  assign y10326 = ~1'b0 ;
  assign y10327 = n16299 ;
  assign y10328 = n16311 ;
  assign y10329 = ~n16314 ;
  assign y10330 = n16315 ;
  assign y10331 = ~n16318 ;
  assign y10332 = ~1'b0 ;
  assign y10333 = n16319 ;
  assign y10334 = ~1'b0 ;
  assign y10335 = n16323 ;
  assign y10336 = ~n16324 ;
  assign y10337 = n16326 ;
  assign y10338 = ~1'b0 ;
  assign y10339 = ~n7469 ;
  assign y10340 = ~n16327 ;
  assign y10341 = ~n16329 ;
  assign y10342 = ~1'b0 ;
  assign y10343 = n16331 ;
  assign y10344 = ~1'b0 ;
  assign y10345 = n16333 ;
  assign y10346 = ~1'b0 ;
  assign y10347 = ~1'b0 ;
  assign y10348 = n629 ;
  assign y10349 = ~1'b0 ;
  assign y10350 = ~n16334 ;
  assign y10351 = ~n16336 ;
  assign y10352 = ~1'b0 ;
  assign y10353 = n16337 ;
  assign y10354 = ~1'b0 ;
  assign y10355 = ~1'b0 ;
  assign y10356 = ~n16341 ;
  assign y10357 = ~1'b0 ;
  assign y10358 = ~1'b0 ;
  assign y10359 = ~n16344 ;
  assign y10360 = ~1'b0 ;
  assign y10361 = ~n16345 ;
  assign y10362 = ~1'b0 ;
  assign y10363 = ~n16346 ;
  assign y10364 = n16348 ;
  assign y10365 = ~n16350 ;
  assign y10366 = ~n16351 ;
  assign y10367 = ~1'b0 ;
  assign y10368 = n16354 ;
  assign y10369 = ~n16355 ;
  assign y10370 = ~n16357 ;
  assign y10371 = ~1'b0 ;
  assign y10372 = ~1'b0 ;
  assign y10373 = ~n16361 ;
  assign y10374 = n16362 ;
  assign y10375 = ~n16363 ;
  assign y10376 = 1'b0 ;
  assign y10377 = ~1'b0 ;
  assign y10378 = n16365 ;
  assign y10379 = ~1'b0 ;
  assign y10380 = ~n16367 ;
  assign y10381 = n16368 ;
  assign y10382 = ~x114 ;
  assign y10383 = n16373 ;
  assign y10384 = ~n16374 ;
  assign y10385 = ~1'b0 ;
  assign y10386 = n16378 ;
  assign y10387 = n16379 ;
  assign y10388 = ~1'b0 ;
  assign y10389 = n16389 ;
  assign y10390 = ~1'b0 ;
  assign y10391 = n16391 ;
  assign y10392 = ~n16392 ;
  assign y10393 = ~n16393 ;
  assign y10394 = ~1'b0 ;
  assign y10395 = ~1'b0 ;
  assign y10396 = n16396 ;
  assign y10397 = ~n16397 ;
  assign y10398 = ~1'b0 ;
  assign y10399 = 1'b0 ;
  assign y10400 = ~n16399 ;
  assign y10401 = ~n2530 ;
  assign y10402 = n16400 ;
  assign y10403 = ~1'b0 ;
  assign y10404 = ~n16404 ;
  assign y10405 = ~n16406 ;
  assign y10406 = n16410 ;
  assign y10407 = n16412 ;
  assign y10408 = n16413 ;
  assign y10409 = ~1'b0 ;
  assign y10410 = ~1'b0 ;
  assign y10411 = n16414 ;
  assign y10412 = ~n16417 ;
  assign y10413 = n6561 ;
  assign y10414 = ~n16420 ;
  assign y10415 = n1664 ;
  assign y10416 = ~1'b0 ;
  assign y10417 = n4098 ;
  assign y10418 = ~1'b0 ;
  assign y10419 = ~n16422 ;
  assign y10420 = ~n3664 ;
  assign y10421 = ~n16423 ;
  assign y10422 = ~1'b0 ;
  assign y10423 = n16424 ;
  assign y10424 = n16426 ;
  assign y10425 = n16427 ;
  assign y10426 = ~1'b0 ;
  assign y10427 = ~n8977 ;
  assign y10428 = ~n16431 ;
  assign y10429 = ~1'b0 ;
  assign y10430 = n7523 ;
  assign y10431 = ~n16432 ;
  assign y10432 = n16433 ;
  assign y10433 = n16436 ;
  assign y10434 = ~1'b0 ;
  assign y10435 = n5704 ;
  assign y10436 = ~n16437 ;
  assign y10437 = ~n16440 ;
  assign y10438 = ~n16441 ;
  assign y10439 = ~n16443 ;
  assign y10440 = n16445 ;
  assign y10441 = n16446 ;
  assign y10442 = n16447 ;
  assign y10443 = ~n16452 ;
  assign y10444 = n16455 ;
  assign y10445 = ~n11112 ;
  assign y10446 = ~n16462 ;
  assign y10447 = 1'b0 ;
  assign y10448 = ~n10526 ;
  assign y10449 = ~n16463 ;
  assign y10450 = ~1'b0 ;
  assign y10451 = n16464 ;
  assign y10452 = n16468 ;
  assign y10453 = ~n16471 ;
  assign y10454 = ~1'b0 ;
  assign y10455 = ~1'b0 ;
  assign y10456 = ~n16490 ;
  assign y10457 = ~n16491 ;
  assign y10458 = n16494 ;
  assign y10459 = ~1'b0 ;
  assign y10460 = n1176 ;
  assign y10461 = ~1'b0 ;
  assign y10462 = n16495 ;
  assign y10463 = ~1'b0 ;
  assign y10464 = ~n16496 ;
  assign y10465 = ~n16498 ;
  assign y10466 = n16500 ;
  assign y10467 = n16503 ;
  assign y10468 = n16504 ;
  assign y10469 = n12105 ;
  assign y10470 = ~1'b0 ;
  assign y10471 = ~1'b0 ;
  assign y10472 = ~1'b0 ;
  assign y10473 = ~n16506 ;
  assign y10474 = n16507 ;
  assign y10475 = ~n16510 ;
  assign y10476 = n16514 ;
  assign y10477 = n16516 ;
  assign y10478 = n16518 ;
  assign y10479 = ~n13882 ;
  assign y10480 = ~n16519 ;
  assign y10481 = ~n16520 ;
  assign y10482 = ~n16523 ;
  assign y10483 = ~n16524 ;
  assign y10484 = ~1'b0 ;
  assign y10485 = ~1'b0 ;
  assign y10486 = ~1'b0 ;
  assign y10487 = ~n16525 ;
  assign y10488 = ~n16530 ;
  assign y10489 = ~n16534 ;
  assign y10490 = ~1'b0 ;
  assign y10491 = 1'b0 ;
  assign y10492 = ~1'b0 ;
  assign y10493 = ~1'b0 ;
  assign y10494 = 1'b0 ;
  assign y10495 = n16535 ;
  assign y10496 = ~1'b0 ;
  assign y10497 = n16536 ;
  assign y10498 = ~n16540 ;
  assign y10499 = n1645 ;
  assign y10500 = ~n16544 ;
  assign y10501 = ~n16545 ;
  assign y10502 = n16546 ;
  assign y10503 = ~n16549 ;
  assign y10504 = ~n16552 ;
  assign y10505 = ~n16555 ;
  assign y10506 = ~n15769 ;
  assign y10507 = ~n16559 ;
  assign y10508 = n14134 ;
  assign y10509 = n16560 ;
  assign y10510 = ~1'b0 ;
  assign y10511 = ~1'b0 ;
  assign y10512 = ~n16561 ;
  assign y10513 = n16567 ;
  assign y10514 = ~n16575 ;
  assign y10515 = n16577 ;
  assign y10516 = 1'b0 ;
  assign y10517 = ~n16578 ;
  assign y10518 = ~n16580 ;
  assign y10519 = 1'b0 ;
  assign y10520 = ~1'b0 ;
  assign y10521 = ~n16581 ;
  assign y10522 = ~n16584 ;
  assign y10523 = 1'b0 ;
  assign y10524 = ~1'b0 ;
  assign y10525 = ~1'b0 ;
  assign y10526 = ~1'b0 ;
  assign y10527 = n16586 ;
  assign y10528 = ~1'b0 ;
  assign y10529 = ~1'b0 ;
  assign y10530 = n16590 ;
  assign y10531 = ~n16594 ;
  assign y10532 = ~n16595 ;
  assign y10533 = ~1'b0 ;
  assign y10534 = ~n6046 ;
  assign y10535 = n16599 ;
  assign y10536 = ~n16600 ;
  assign y10537 = ~n16601 ;
  assign y10538 = ~1'b0 ;
  assign y10539 = n16604 ;
  assign y10540 = n8738 ;
  assign y10541 = ~1'b0 ;
  assign y10542 = ~n16606 ;
  assign y10543 = n16608 ;
  assign y10544 = ~1'b0 ;
  assign y10545 = ~n16611 ;
  assign y10546 = n16613 ;
  assign y10547 = ~1'b0 ;
  assign y10548 = ~n16615 ;
  assign y10549 = ~1'b0 ;
  assign y10550 = ~n16618 ;
  assign y10551 = ~1'b0 ;
  assign y10552 = ~1'b0 ;
  assign y10553 = ~1'b0 ;
  assign y10554 = n16620 ;
  assign y10555 = n16625 ;
  assign y10556 = ~1'b0 ;
  assign y10557 = ~n16626 ;
  assign y10558 = n16629 ;
  assign y10559 = ~1'b0 ;
  assign y10560 = ~1'b0 ;
  assign y10561 = n10177 ;
  assign y10562 = ~1'b0 ;
  assign y10563 = ~n16632 ;
  assign y10564 = ~n16634 ;
  assign y10565 = ~1'b0 ;
  assign y10566 = ~n16636 ;
  assign y10567 = n16638 ;
  assign y10568 = ~1'b0 ;
  assign y10569 = ~1'b0 ;
  assign y10570 = ~n16639 ;
  assign y10571 = n16640 ;
  assign y10572 = n15947 ;
  assign y10573 = n16641 ;
  assign y10574 = n16642 ;
  assign y10575 = n16646 ;
  assign y10576 = ~n16648 ;
  assign y10577 = n16649 ;
  assign y10578 = ~1'b0 ;
  assign y10579 = ~1'b0 ;
  assign y10580 = ~1'b0 ;
  assign y10581 = ~n16651 ;
  assign y10582 = ~n6979 ;
  assign y10583 = n16652 ;
  assign y10584 = ~1'b0 ;
  assign y10585 = n16653 ;
  assign y10586 = ~1'b0 ;
  assign y10587 = ~1'b0 ;
  assign y10588 = ~1'b0 ;
  assign y10589 = n16655 ;
  assign y10590 = ~n4443 ;
  assign y10591 = n16656 ;
  assign y10592 = ~n16664 ;
  assign y10593 = ~n16667 ;
  assign y10594 = ~n16671 ;
  assign y10595 = ~1'b0 ;
  assign y10596 = ~n3083 ;
  assign y10597 = n16674 ;
  assign y10598 = n16677 ;
  assign y10599 = n16679 ;
  assign y10600 = ~1'b0 ;
  assign y10601 = ~n16681 ;
  assign y10602 = ~1'b0 ;
  assign y10603 = ~n16683 ;
  assign y10604 = ~n16684 ;
  assign y10605 = n16685 ;
  assign y10606 = ~1'b0 ;
  assign y10607 = ~n6396 ;
  assign y10608 = n16686 ;
  assign y10609 = ~n16687 ;
  assign y10610 = ~n16690 ;
  assign y10611 = n4878 ;
  assign y10612 = ~n16692 ;
  assign y10613 = 1'b0 ;
  assign y10614 = ~n16693 ;
  assign y10615 = ~1'b0 ;
  assign y10616 = ~1'b0 ;
  assign y10617 = ~1'b0 ;
  assign y10618 = ~n16694 ;
  assign y10619 = ~1'b0 ;
  assign y10620 = ~n16704 ;
  assign y10621 = n16705 ;
  assign y10622 = ~n8260 ;
  assign y10623 = ~1'b0 ;
  assign y10624 = n16709 ;
  assign y10625 = ~n16710 ;
  assign y10626 = ~1'b0 ;
  assign y10627 = ~n16712 ;
  assign y10628 = n16713 ;
  assign y10629 = ~1'b0 ;
  assign y10630 = ~1'b0 ;
  assign y10631 = n16715 ;
  assign y10632 = ~1'b0 ;
  assign y10633 = n16716 ;
  assign y10634 = n16718 ;
  assign y10635 = ~1'b0 ;
  assign y10636 = n16720 ;
  assign y10637 = n8927 ;
  assign y10638 = n16722 ;
  assign y10639 = n16723 ;
  assign y10640 = n16726 ;
  assign y10641 = ~n5727 ;
  assign y10642 = ~1'b0 ;
  assign y10643 = ~n16728 ;
  assign y10644 = ~1'b0 ;
  assign y10645 = ~1'b0 ;
  assign y10646 = ~n16729 ;
  assign y10647 = ~n4775 ;
  assign y10648 = ~1'b0 ;
  assign y10649 = n16732 ;
  assign y10650 = ~n16182 ;
  assign y10651 = ~n16733 ;
  assign y10652 = n16738 ;
  assign y10653 = ~n16739 ;
  assign y10654 = ~n16743 ;
  assign y10655 = n16745 ;
  assign y10656 = ~n16749 ;
  assign y10657 = n16753 ;
  assign y10658 = ~n16754 ;
  assign y10659 = n1002 ;
  assign y10660 = ~n16756 ;
  assign y10661 = ~n16758 ;
  assign y10662 = ~n16761 ;
  assign y10663 = ~n16762 ;
  assign y10664 = n16763 ;
  assign y10665 = n16764 ;
  assign y10666 = ~n6552 ;
  assign y10667 = ~1'b0 ;
  assign y10668 = ~1'b0 ;
  assign y10669 = n16765 ;
  assign y10670 = ~1'b0 ;
  assign y10671 = ~n16766 ;
  assign y10672 = ~n16769 ;
  assign y10673 = ~n16770 ;
  assign y10674 = n16773 ;
  assign y10675 = ~n16774 ;
  assign y10676 = ~n16775 ;
  assign y10677 = ~n16785 ;
  assign y10678 = ~n16786 ;
  assign y10679 = ~1'b0 ;
  assign y10680 = ~n16787 ;
  assign y10681 = ~n16788 ;
  assign y10682 = ~1'b0 ;
  assign y10683 = ~n16790 ;
  assign y10684 = n16791 ;
  assign y10685 = ~n16794 ;
  assign y10686 = ~n16795 ;
  assign y10687 = ~n12578 ;
  assign y10688 = n16798 ;
  assign y10689 = n16799 ;
  assign y10690 = n16800 ;
  assign y10691 = 1'b0 ;
  assign y10692 = ~n16802 ;
  assign y10693 = n16807 ;
  assign y10694 = ~1'b0 ;
  assign y10695 = ~1'b0 ;
  assign y10696 = ~n16809 ;
  assign y10697 = ~n16811 ;
  assign y10698 = ~n10142 ;
  assign y10699 = n16813 ;
  assign y10700 = ~1'b0 ;
  assign y10701 = ~n16814 ;
  assign y10702 = ~1'b0 ;
  assign y10703 = ~1'b0 ;
  assign y10704 = ~1'b0 ;
  assign y10705 = 1'b0 ;
  assign y10706 = n16815 ;
  assign y10707 = n16819 ;
  assign y10708 = ~n9801 ;
  assign y10709 = ~1'b0 ;
  assign y10710 = ~1'b0 ;
  assign y10711 = ~1'b0 ;
  assign y10712 = ~n16822 ;
  assign y10713 = ~1'b0 ;
  assign y10714 = ~n16824 ;
  assign y10715 = n12857 ;
  assign y10716 = ~n15697 ;
  assign y10717 = ~1'b0 ;
  assign y10718 = ~1'b0 ;
  assign y10719 = ~1'b0 ;
  assign y10720 = n16827 ;
  assign y10721 = n16830 ;
  assign y10722 = n16832 ;
  assign y10723 = 1'b0 ;
  assign y10724 = n16834 ;
  assign y10725 = ~1'b0 ;
  assign y10726 = 1'b0 ;
  assign y10727 = ~1'b0 ;
  assign y10728 = ~1'b0 ;
  assign y10729 = 1'b0 ;
  assign y10730 = n16835 ;
  assign y10731 = n3171 ;
  assign y10732 = ~1'b0 ;
  assign y10733 = n16836 ;
  assign y10734 = ~n16838 ;
  assign y10735 = ~n16840 ;
  assign y10736 = ~1'b0 ;
  assign y10737 = n16844 ;
  assign y10738 = ~1'b0 ;
  assign y10739 = n16849 ;
  assign y10740 = n16852 ;
  assign y10741 = ~1'b0 ;
  assign y10742 = 1'b0 ;
  assign y10743 = ~n16858 ;
  assign y10744 = ~n16859 ;
  assign y10745 = 1'b0 ;
  assign y10746 = ~1'b0 ;
  assign y10747 = n16861 ;
  assign y10748 = ~1'b0 ;
  assign y10749 = ~1'b0 ;
  assign y10750 = ~n16864 ;
  assign y10751 = n16865 ;
  assign y10752 = n16867 ;
  assign y10753 = ~n16870 ;
  assign y10754 = ~n16872 ;
  assign y10755 = ~1'b0 ;
  assign y10756 = ~1'b0 ;
  assign y10757 = ~n16873 ;
  assign y10758 = n16879 ;
  assign y10759 = n16881 ;
  assign y10760 = ~n16885 ;
  assign y10761 = ~1'b0 ;
  assign y10762 = ~n16886 ;
  assign y10763 = n16887 ;
  assign y10764 = ~1'b0 ;
  assign y10765 = ~n16889 ;
  assign y10766 = ~n16890 ;
  assign y10767 = ~n16892 ;
  assign y10768 = ~1'b0 ;
  assign y10769 = 1'b0 ;
  assign y10770 = n16893 ;
  assign y10771 = n16895 ;
  assign y10772 = n463 ;
  assign y10773 = n16896 ;
  assign y10774 = ~n16898 ;
  assign y10775 = n16899 ;
  assign y10776 = ~n16902 ;
  assign y10777 = n8260 ;
  assign y10778 = ~1'b0 ;
  assign y10779 = ~1'b0 ;
  assign y10780 = n16907 ;
  assign y10781 = n16908 ;
  assign y10782 = n16909 ;
  assign y10783 = n16910 ;
  assign y10784 = ~1'b0 ;
  assign y10785 = n16911 ;
  assign y10786 = n16918 ;
  assign y10787 = 1'b0 ;
  assign y10788 = ~1'b0 ;
  assign y10789 = ~1'b0 ;
  assign y10790 = ~1'b0 ;
  assign y10791 = n1952 ;
  assign y10792 = ~1'b0 ;
  assign y10793 = n16919 ;
  assign y10794 = ~1'b0 ;
  assign y10795 = ~1'b0 ;
  assign y10796 = ~n16921 ;
  assign y10797 = n16922 ;
  assign y10798 = ~n2773 ;
  assign y10799 = ~1'b0 ;
  assign y10800 = n16928 ;
  assign y10801 = ~n16929 ;
  assign y10802 = 1'b0 ;
  assign y10803 = n6398 ;
  assign y10804 = ~n16936 ;
  assign y10805 = ~n16938 ;
  assign y10806 = ~n16939 ;
  assign y10807 = ~1'b0 ;
  assign y10808 = ~1'b0 ;
  assign y10809 = 1'b0 ;
  assign y10810 = ~n16941 ;
  assign y10811 = ~1'b0 ;
  assign y10812 = n16942 ;
  assign y10813 = ~1'b0 ;
  assign y10814 = ~1'b0 ;
  assign y10815 = ~1'b0 ;
  assign y10816 = n16943 ;
  assign y10817 = ~1'b0 ;
  assign y10818 = ~n16948 ;
  assign y10819 = ~n16950 ;
  assign y10820 = ~1'b0 ;
  assign y10821 = ~1'b0 ;
  assign y10822 = ~1'b0 ;
  assign y10823 = 1'b0 ;
  assign y10824 = ~n16952 ;
  assign y10825 = n11532 ;
  assign y10826 = ~n16953 ;
  assign y10827 = ~n7184 ;
  assign y10828 = ~1'b0 ;
  assign y10829 = ~1'b0 ;
  assign y10830 = n16954 ;
  assign y10831 = ~n16956 ;
  assign y10832 = ~1'b0 ;
  assign y10833 = ~n16957 ;
  assign y10834 = ~n16961 ;
  assign y10835 = ~1'b0 ;
  assign y10836 = n16964 ;
  assign y10837 = ~1'b0 ;
  assign y10838 = ~1'b0 ;
  assign y10839 = ~n16967 ;
  assign y10840 = n14854 ;
  assign y10841 = ~n5870 ;
  assign y10842 = ~1'b0 ;
  assign y10843 = ~1'b0 ;
  assign y10844 = n4521 ;
  assign y10845 = n16969 ;
  assign y10846 = ~n7866 ;
  assign y10847 = ~n16970 ;
  assign y10848 = ~n16972 ;
  assign y10849 = n16974 ;
  assign y10850 = ~1'b0 ;
  assign y10851 = ~1'b0 ;
  assign y10852 = ~1'b0 ;
  assign y10853 = 1'b0 ;
  assign y10854 = n16976 ;
  assign y10855 = ~n16981 ;
  assign y10856 = n16984 ;
  assign y10857 = n16989 ;
  assign y10858 = ~1'b0 ;
  assign y10859 = n16999 ;
  assign y10860 = ~n17000 ;
  assign y10861 = ~n17005 ;
  assign y10862 = n17007 ;
  assign y10863 = ~1'b0 ;
  assign y10864 = ~1'b0 ;
  assign y10865 = ~n17011 ;
  assign y10866 = n17012 ;
  assign y10867 = ~1'b0 ;
  assign y10868 = n17020 ;
  assign y10869 = ~n17022 ;
  assign y10870 = ~n17026 ;
  assign y10871 = ~1'b0 ;
  assign y10872 = ~n17029 ;
  assign y10873 = ~1'b0 ;
  assign y10874 = n17030 ;
  assign y10875 = ~1'b0 ;
  assign y10876 = ~n17034 ;
  assign y10877 = ~1'b0 ;
  assign y10878 = ~n17038 ;
  assign y10879 = ~1'b0 ;
  assign y10880 = n17046 ;
  assign y10881 = ~n17049 ;
  assign y10882 = ~1'b0 ;
  assign y10883 = n17051 ;
  assign y10884 = ~n17056 ;
  assign y10885 = ~1'b0 ;
  assign y10886 = n17057 ;
  assign y10887 = ~n17059 ;
  assign y10888 = ~n17061 ;
  assign y10889 = ~n17062 ;
  assign y10890 = n17064 ;
  assign y10891 = n17067 ;
  assign y10892 = n17070 ;
  assign y10893 = ~n14788 ;
  assign y10894 = ~n17071 ;
  assign y10895 = ~1'b0 ;
  assign y10896 = ~1'b0 ;
  assign y10897 = n17072 ;
  assign y10898 = ~1'b0 ;
  assign y10899 = ~1'b0 ;
  assign y10900 = ~1'b0 ;
  assign y10901 = ~n17075 ;
  assign y10902 = ~n17081 ;
  assign y10903 = ~n17082 ;
  assign y10904 = 1'b0 ;
  assign y10905 = ~x127 ;
  assign y10906 = ~1'b0 ;
  assign y10907 = ~n17086 ;
  assign y10908 = ~n17091 ;
  assign y10909 = n17093 ;
  assign y10910 = ~n17094 ;
  assign y10911 = ~1'b0 ;
  assign y10912 = ~1'b0 ;
  assign y10913 = ~n17098 ;
  assign y10914 = 1'b0 ;
  assign y10915 = ~n17100 ;
  assign y10916 = ~n17102 ;
  assign y10917 = ~1'b0 ;
  assign y10918 = n17103 ;
  assign y10919 = ~n17104 ;
  assign y10920 = ~1'b0 ;
  assign y10921 = ~1'b0 ;
  assign y10922 = ~1'b0 ;
  assign y10923 = ~n17108 ;
  assign y10924 = n17109 ;
  assign y10925 = n17111 ;
  assign y10926 = n17113 ;
  assign y10927 = n17114 ;
  assign y10928 = n17116 ;
  assign y10929 = n1508 ;
  assign y10930 = n14038 ;
  assign y10931 = n17117 ;
  assign y10932 = ~n17128 ;
  assign y10933 = n17129 ;
  assign y10934 = n17133 ;
  assign y10935 = n17135 ;
  assign y10936 = n17138 ;
  assign y10937 = ~n17145 ;
  assign y10938 = ~1'b0 ;
  assign y10939 = n17147 ;
  assign y10940 = n17149 ;
  assign y10941 = ~1'b0 ;
  assign y10942 = n2149 ;
  assign y10943 = ~1'b0 ;
  assign y10944 = ~1'b0 ;
  assign y10945 = n17154 ;
  assign y10946 = ~n17155 ;
  assign y10947 = n17157 ;
  assign y10948 = ~1'b0 ;
  assign y10949 = ~1'b0 ;
  assign y10950 = ~1'b0 ;
  assign y10951 = ~1'b0 ;
  assign y10952 = ~n17158 ;
  assign y10953 = n17162 ;
  assign y10954 = ~n17164 ;
  assign y10955 = ~n4310 ;
  assign y10956 = ~n17197 ;
  assign y10957 = ~1'b0 ;
  assign y10958 = 1'b0 ;
  assign y10959 = 1'b0 ;
  assign y10960 = ~1'b0 ;
  assign y10961 = ~1'b0 ;
  assign y10962 = ~n13136 ;
  assign y10963 = ~1'b0 ;
  assign y10964 = ~n17199 ;
  assign y10965 = n17201 ;
  assign y10966 = n17203 ;
  assign y10967 = n17204 ;
  assign y10968 = ~1'b0 ;
  assign y10969 = ~n17206 ;
  assign y10970 = ~1'b0 ;
  assign y10971 = n14734 ;
  assign y10972 = ~n2773 ;
  assign y10973 = n17208 ;
  assign y10974 = ~1'b0 ;
  assign y10975 = n17209 ;
  assign y10976 = ~1'b0 ;
  assign y10977 = ~1'b0 ;
  assign y10978 = n15986 ;
  assign y10979 = n17211 ;
  assign y10980 = ~n17214 ;
  assign y10981 = ~1'b0 ;
  assign y10982 = ~1'b0 ;
  assign y10983 = n17216 ;
  assign y10984 = ~1'b0 ;
  assign y10985 = n17217 ;
  assign y10986 = n16612 ;
  assign y10987 = ~1'b0 ;
  assign y10988 = n17218 ;
  assign y10989 = ~n17220 ;
  assign y10990 = ~1'b0 ;
  assign y10991 = n17221 ;
  assign y10992 = n17223 ;
  assign y10993 = n17224 ;
  assign y10994 = 1'b0 ;
  assign y10995 = ~n17227 ;
  assign y10996 = ~n17228 ;
  assign y10997 = ~1'b0 ;
  assign y10998 = ~n17233 ;
  assign y10999 = 1'b0 ;
  assign y11000 = ~1'b0 ;
  assign y11001 = ~1'b0 ;
  assign y11002 = ~n17234 ;
  assign y11003 = n17235 ;
  assign y11004 = ~n17236 ;
  assign y11005 = ~n17240 ;
  assign y11006 = n17242 ;
  assign y11007 = n17243 ;
  assign y11008 = ~1'b0 ;
  assign y11009 = ~1'b0 ;
  assign y11010 = ~n2024 ;
  assign y11011 = ~1'b0 ;
  assign y11012 = ~n17244 ;
  assign y11013 = 1'b0 ;
  assign y11014 = ~n3322 ;
  assign y11015 = n9364 ;
  assign y11016 = ~1'b0 ;
  assign y11017 = ~n17247 ;
  assign y11018 = ~1'b0 ;
  assign y11019 = ~n17248 ;
  assign y11020 = n13694 ;
  assign y11021 = ~n17252 ;
  assign y11022 = ~n17256 ;
  assign y11023 = ~n17257 ;
  assign y11024 = ~1'b0 ;
  assign y11025 = ~n17260 ;
  assign y11026 = n17261 ;
  assign y11027 = ~1'b0 ;
  assign y11028 = ~1'b0 ;
  assign y11029 = ~n17263 ;
  assign y11030 = n17264 ;
  assign y11031 = n17265 ;
  assign y11032 = ~1'b0 ;
  assign y11033 = n17266 ;
  assign y11034 = ~n17267 ;
  assign y11035 = ~1'b0 ;
  assign y11036 = ~n6644 ;
  assign y11037 = n17276 ;
  assign y11038 = ~n17277 ;
  assign y11039 = ~n17280 ;
  assign y11040 = ~n17281 ;
  assign y11041 = ~1'b0 ;
  assign y11042 = n17282 ;
  assign y11043 = ~n3646 ;
  assign y11044 = ~1'b0 ;
  assign y11045 = n17289 ;
  assign y11046 = n17294 ;
  assign y11047 = ~n17296 ;
  assign y11048 = ~1'b0 ;
  assign y11049 = ~1'b0 ;
  assign y11050 = ~1'b0 ;
  assign y11051 = n17297 ;
  assign y11052 = n17301 ;
  assign y11053 = n967 ;
  assign y11054 = ~n17304 ;
  assign y11055 = ~1'b0 ;
  assign y11056 = ~1'b0 ;
  assign y11057 = ~n17305 ;
  assign y11058 = 1'b0 ;
  assign y11059 = ~n5458 ;
  assign y11060 = ~n17306 ;
  assign y11061 = n17308 ;
  assign y11062 = ~n6947 ;
  assign y11063 = ~n17311 ;
  assign y11064 = ~1'b0 ;
  assign y11065 = 1'b0 ;
  assign y11066 = n17314 ;
  assign y11067 = ~1'b0 ;
  assign y11068 = ~1'b0 ;
  assign y11069 = ~1'b0 ;
  assign y11070 = ~1'b0 ;
  assign y11071 = ~1'b0 ;
  assign y11072 = ~1'b0 ;
  assign y11073 = n17316 ;
  assign y11074 = 1'b0 ;
  assign y11075 = ~n1034 ;
  assign y11076 = ~n17318 ;
  assign y11077 = ~1'b0 ;
  assign y11078 = ~n17319 ;
  assign y11079 = ~n12518 ;
  assign y11080 = ~n17321 ;
  assign y11081 = ~n17322 ;
  assign y11082 = ~n17325 ;
  assign y11083 = ~1'b0 ;
  assign y11084 = ~1'b0 ;
  assign y11085 = n17331 ;
  assign y11086 = ~1'b0 ;
  assign y11087 = ~1'b0 ;
  assign y11088 = ~1'b0 ;
  assign y11089 = ~1'b0 ;
  assign y11090 = ~n17333 ;
  assign y11091 = n10186 ;
  assign y11092 = ~n17338 ;
  assign y11093 = ~n17340 ;
  assign y11094 = ~1'b0 ;
  assign y11095 = n17341 ;
  assign y11096 = n17343 ;
  assign y11097 = ~n12960 ;
  assign y11098 = ~n17344 ;
  assign y11099 = ~1'b0 ;
  assign y11100 = ~1'b0 ;
  assign y11101 = ~n17354 ;
  assign y11102 = ~1'b0 ;
  assign y11103 = ~n17355 ;
  assign y11104 = ~n17356 ;
  assign y11105 = ~1'b0 ;
  assign y11106 = n17357 ;
  assign y11107 = ~1'b0 ;
  assign y11108 = ~1'b0 ;
  assign y11109 = ~1'b0 ;
  assign y11110 = ~1'b0 ;
  assign y11111 = ~n17358 ;
  assign y11112 = n17362 ;
  assign y11113 = ~1'b0 ;
  assign y11114 = ~n17366 ;
  assign y11115 = ~n17375 ;
  assign y11116 = ~n17377 ;
  assign y11117 = n17379 ;
  assign y11118 = ~1'b0 ;
  assign y11119 = n17383 ;
  assign y11120 = n17384 ;
  assign y11121 = ~1'b0 ;
  assign y11122 = ~n17387 ;
  assign y11123 = ~n17389 ;
  assign y11124 = ~n17392 ;
  assign y11125 = ~1'b0 ;
  assign y11126 = n17394 ;
  assign y11127 = n17395 ;
  assign y11128 = n17400 ;
  assign y11129 = ~n17402 ;
  assign y11130 = ~n17405 ;
  assign y11131 = ~1'b0 ;
  assign y11132 = n17407 ;
  assign y11133 = n17410 ;
  assign y11134 = ~1'b0 ;
  assign y11135 = ~1'b0 ;
  assign y11136 = n17411 ;
  assign y11137 = ~1'b0 ;
  assign y11138 = n17416 ;
  assign y11139 = n17417 ;
  assign y11140 = n17419 ;
  assign y11141 = ~1'b0 ;
  assign y11142 = ~1'b0 ;
  assign y11143 = ~n8262 ;
  assign y11144 = ~1'b0 ;
  assign y11145 = ~n17421 ;
  assign y11146 = ~n17423 ;
  assign y11147 = ~n17425 ;
  assign y11148 = n17427 ;
  assign y11149 = n17429 ;
  assign y11150 = n17430 ;
  assign y11151 = ~1'b0 ;
  assign y11152 = n17431 ;
  assign y11153 = ~n17433 ;
  assign y11154 = n1216 ;
  assign y11155 = ~n17436 ;
  assign y11156 = ~n17439 ;
  assign y11157 = ~1'b0 ;
  assign y11158 = ~n17441 ;
  assign y11159 = n17446 ;
  assign y11160 = ~1'b0 ;
  assign y11161 = ~n17447 ;
  assign y11162 = ~n15309 ;
  assign y11163 = n17448 ;
  assign y11164 = n17449 ;
  assign y11165 = ~1'b0 ;
  assign y11166 = ~1'b0 ;
  assign y11167 = ~1'b0 ;
  assign y11168 = ~n17451 ;
  assign y11169 = ~n17453 ;
  assign y11170 = n17457 ;
  assign y11171 = ~1'b0 ;
  assign y11172 = ~n17458 ;
  assign y11173 = n17459 ;
  assign y11174 = ~1'b0 ;
  assign y11175 = ~n9713 ;
  assign y11176 = ~1'b0 ;
  assign y11177 = n17461 ;
  assign y11178 = ~1'b0 ;
  assign y11179 = n8705 ;
  assign y11180 = 1'b0 ;
  assign y11181 = n17464 ;
  assign y11182 = ~1'b0 ;
  assign y11183 = ~1'b0 ;
  assign y11184 = ~1'b0 ;
  assign y11185 = ~n17468 ;
  assign y11186 = n17469 ;
  assign y11187 = n17471 ;
  assign y11188 = n17475 ;
  assign y11189 = ~1'b0 ;
  assign y11190 = n17476 ;
  assign y11191 = ~1'b0 ;
  assign y11192 = ~n17481 ;
  assign y11193 = n17482 ;
  assign y11194 = ~1'b0 ;
  assign y11195 = ~1'b0 ;
  assign y11196 = ~n17484 ;
  assign y11197 = ~n17485 ;
  assign y11198 = ~1'b0 ;
  assign y11199 = ~n17487 ;
  assign y11200 = 1'b0 ;
  assign y11201 = ~1'b0 ;
  assign y11202 = n17488 ;
  assign y11203 = ~1'b0 ;
  assign y11204 = ~n17490 ;
  assign y11205 = 1'b0 ;
  assign y11206 = ~1'b0 ;
  assign y11207 = ~n17491 ;
  assign y11208 = ~1'b0 ;
  assign y11209 = ~n17495 ;
  assign y11210 = ~n17496 ;
  assign y11211 = ~1'b0 ;
  assign y11212 = n17498 ;
  assign y11213 = ~1'b0 ;
  assign y11214 = ~1'b0 ;
  assign y11215 = ~n17501 ;
  assign y11216 = ~1'b0 ;
  assign y11217 = ~n17503 ;
  assign y11218 = n4353 ;
  assign y11219 = n17505 ;
  assign y11220 = ~1'b0 ;
  assign y11221 = ~n17507 ;
  assign y11222 = ~1'b0 ;
  assign y11223 = n17509 ;
  assign y11224 = ~1'b0 ;
  assign y11225 = ~n17510 ;
  assign y11226 = n6463 ;
  assign y11227 = ~1'b0 ;
  assign y11228 = n17511 ;
  assign y11229 = ~1'b0 ;
  assign y11230 = ~1'b0 ;
  assign y11231 = ~1'b0 ;
  assign y11232 = n17512 ;
  assign y11233 = ~1'b0 ;
  assign y11234 = ~n17513 ;
  assign y11235 = ~n7852 ;
  assign y11236 = ~n17515 ;
  assign y11237 = n12198 ;
  assign y11238 = ~n17518 ;
  assign y11239 = ~1'b0 ;
  assign y11240 = n17520 ;
  assign y11241 = ~n17521 ;
  assign y11242 = n17524 ;
  assign y11243 = n17525 ;
  assign y11244 = n17531 ;
  assign y11245 = n17534 ;
  assign y11246 = n1554 ;
  assign y11247 = n17536 ;
  assign y11248 = ~1'b0 ;
  assign y11249 = ~1'b0 ;
  assign y11250 = n7001 ;
  assign y11251 = ~1'b0 ;
  assign y11252 = ~n17537 ;
  assign y11253 = n3391 ;
  assign y11254 = ~n17540 ;
  assign y11255 = ~n17545 ;
  assign y11256 = ~n17548 ;
  assign y11257 = n17550 ;
  assign y11258 = n14937 ;
  assign y11259 = n17551 ;
  assign y11260 = n9205 ;
  assign y11261 = ~n17553 ;
  assign y11262 = ~n17554 ;
  assign y11263 = ~n17556 ;
  assign y11264 = n17558 ;
  assign y11265 = ~1'b0 ;
  assign y11266 = n17560 ;
  assign y11267 = ~1'b0 ;
  assign y11268 = ~1'b0 ;
  assign y11269 = ~1'b0 ;
  assign y11270 = n17563 ;
  assign y11271 = ~1'b0 ;
  assign y11272 = ~1'b0 ;
  assign y11273 = ~n17565 ;
  assign y11274 = n17566 ;
  assign y11275 = ~n17567 ;
  assign y11276 = ~n17570 ;
  assign y11277 = n17572 ;
  assign y11278 = n863 ;
  assign y11279 = ~1'b0 ;
  assign y11280 = n17576 ;
  assign y11281 = ~1'b0 ;
  assign y11282 = ~1'b0 ;
  assign y11283 = ~n17581 ;
  assign y11284 = ~1'b0 ;
  assign y11285 = n17587 ;
  assign y11286 = ~n17593 ;
  assign y11287 = ~n6445 ;
  assign y11288 = ~1'b0 ;
  assign y11289 = ~n17597 ;
  assign y11290 = ~1'b0 ;
  assign y11291 = ~n17598 ;
  assign y11292 = 1'b0 ;
  assign y11293 = n7735 ;
  assign y11294 = ~n17604 ;
  assign y11295 = ~n17606 ;
  assign y11296 = n17607 ;
  assign y11297 = ~n17610 ;
  assign y11298 = n17612 ;
  assign y11299 = ~n17614 ;
  assign y11300 = n17621 ;
  assign y11301 = 1'b0 ;
  assign y11302 = ~1'b0 ;
  assign y11303 = 1'b0 ;
  assign y11304 = ~n17622 ;
  assign y11305 = n17627 ;
  assign y11306 = ~1'b0 ;
  assign y11307 = ~1'b0 ;
  assign y11308 = ~n17630 ;
  assign y11309 = n17632 ;
  assign y11310 = ~n17637 ;
  assign y11311 = ~1'b0 ;
  assign y11312 = ~1'b0 ;
  assign y11313 = ~n3632 ;
  assign y11314 = ~1'b0 ;
  assign y11315 = ~1'b0 ;
  assign y11316 = ~1'b0 ;
  assign y11317 = 1'b0 ;
  assign y11318 = n17641 ;
  assign y11319 = ~1'b0 ;
  assign y11320 = ~1'b0 ;
  assign y11321 = n17644 ;
  assign y11322 = n17645 ;
  assign y11323 = n17648 ;
  assign y11324 = n17649 ;
  assign y11325 = n17652 ;
  assign y11326 = n17653 ;
  assign y11327 = n17655 ;
  assign y11328 = n17656 ;
  assign y11329 = ~n9045 ;
  assign y11330 = ~1'b0 ;
  assign y11331 = ~1'b0 ;
  assign y11332 = n17664 ;
  assign y11333 = ~n17666 ;
  assign y11334 = n17668 ;
  assign y11335 = n17670 ;
  assign y11336 = ~n17671 ;
  assign y11337 = ~n17675 ;
  assign y11338 = ~n5245 ;
  assign y11339 = n17676 ;
  assign y11340 = ~1'b0 ;
  assign y11341 = n17677 ;
  assign y11342 = ~1'b0 ;
  assign y11343 = ~1'b0 ;
  assign y11344 = n17678 ;
  assign y11345 = ~n17682 ;
  assign y11346 = ~1'b0 ;
  assign y11347 = n17683 ;
  assign y11348 = ~n17685 ;
  assign y11349 = ~1'b0 ;
  assign y11350 = n17686 ;
  assign y11351 = n17691 ;
  assign y11352 = ~1'b0 ;
  assign y11353 = n17692 ;
  assign y11354 = ~1'b0 ;
  assign y11355 = ~n17694 ;
  assign y11356 = ~1'b0 ;
  assign y11357 = ~1'b0 ;
  assign y11358 = ~n17695 ;
  assign y11359 = n17699 ;
  assign y11360 = ~n17701 ;
  assign y11361 = 1'b0 ;
  assign y11362 = ~1'b0 ;
  assign y11363 = n17703 ;
  assign y11364 = ~1'b0 ;
  assign y11365 = ~1'b0 ;
  assign y11366 = ~1'b0 ;
  assign y11367 = ~n17704 ;
  assign y11368 = n17705 ;
  assign y11369 = n17708 ;
  assign y11370 = ~1'b0 ;
  assign y11371 = n17713 ;
  assign y11372 = n17375 ;
  assign y11373 = ~n17714 ;
  assign y11374 = ~n17716 ;
  assign y11375 = ~1'b0 ;
  assign y11376 = n17718 ;
  assign y11377 = n17719 ;
  assign y11378 = ~n17720 ;
  assign y11379 = ~1'b0 ;
  assign y11380 = ~1'b0 ;
  assign y11381 = ~n17723 ;
  assign y11382 = n17724 ;
  assign y11383 = ~1'b0 ;
  assign y11384 = n17727 ;
  assign y11385 = ~n17729 ;
  assign y11386 = ~n17732 ;
  assign y11387 = ~n17733 ;
  assign y11388 = 1'b0 ;
  assign y11389 = n14542 ;
  assign y11390 = n17734 ;
  assign y11391 = n17735 ;
  assign y11392 = 1'b0 ;
  assign y11393 = ~n17738 ;
  assign y11394 = 1'b0 ;
  assign y11395 = ~1'b0 ;
  assign y11396 = n17740 ;
  assign y11397 = ~n15390 ;
  assign y11398 = n17742 ;
  assign y11399 = n17745 ;
  assign y11400 = ~n17746 ;
  assign y11401 = n17747 ;
  assign y11402 = n17750 ;
  assign y11403 = n17751 ;
  assign y11404 = ~n17753 ;
  assign y11405 = ~1'b0 ;
  assign y11406 = ~n17754 ;
  assign y11407 = ~1'b0 ;
  assign y11408 = ~n17758 ;
  assign y11409 = n17759 ;
  assign y11410 = 1'b0 ;
  assign y11411 = 1'b0 ;
  assign y11412 = ~1'b0 ;
  assign y11413 = ~n17763 ;
  assign y11414 = ~n2154 ;
  assign y11415 = ~1'b0 ;
  assign y11416 = ~n17766 ;
  assign y11417 = n17767 ;
  assign y11418 = n13909 ;
  assign y11419 = ~1'b0 ;
  assign y11420 = ~1'b0 ;
  assign y11421 = 1'b0 ;
  assign y11422 = ~n17769 ;
  assign y11423 = ~1'b0 ;
  assign y11424 = ~1'b0 ;
  assign y11425 = ~n17770 ;
  assign y11426 = ~1'b0 ;
  assign y11427 = ~n17771 ;
  assign y11428 = ~1'b0 ;
  assign y11429 = ~1'b0 ;
  assign y11430 = ~1'b0 ;
  assign y11431 = ~n17773 ;
  assign y11432 = ~1'b0 ;
  assign y11433 = ~n17778 ;
  assign y11434 = n17779 ;
  assign y11435 = ~n17780 ;
  assign y11436 = ~n17784 ;
  assign y11437 = ~n17786 ;
  assign y11438 = ~n17788 ;
  assign y11439 = ~1'b0 ;
  assign y11440 = ~n17794 ;
  assign y11441 = n17799 ;
  assign y11442 = ~1'b0 ;
  assign y11443 = n17805 ;
  assign y11444 = ~n15643 ;
  assign y11445 = ~n2014 ;
  assign y11446 = n17806 ;
  assign y11447 = 1'b0 ;
  assign y11448 = ~1'b0 ;
  assign y11449 = 1'b0 ;
  assign y11450 = ~1'b0 ;
  assign y11451 = ~n17807 ;
  assign y11452 = ~n17809 ;
  assign y11453 = ~n17810 ;
  assign y11454 = ~n17814 ;
  assign y11455 = ~1'b0 ;
  assign y11456 = n17819 ;
  assign y11457 = n17820 ;
  assign y11458 = ~n17821 ;
  assign y11459 = ~1'b0 ;
  assign y11460 = ~n17822 ;
  assign y11461 = ~1'b0 ;
  assign y11462 = n17823 ;
  assign y11463 = n17826 ;
  assign y11464 = ~1'b0 ;
  assign y11465 = ~n17827 ;
  assign y11466 = n17828 ;
  assign y11467 = ~1'b0 ;
  assign y11468 = ~1'b0 ;
  assign y11469 = n17829 ;
  assign y11470 = ~n17831 ;
  assign y11471 = n17834 ;
  assign y11472 = n17836 ;
  assign y11473 = n17838 ;
  assign y11474 = ~1'b0 ;
  assign y11475 = ~n4001 ;
  assign y11476 = n17841 ;
  assign y11477 = ~n17843 ;
  assign y11478 = ~n17845 ;
  assign y11479 = ~n17846 ;
  assign y11480 = n17848 ;
  assign y11481 = n17850 ;
  assign y11482 = n17854 ;
  assign y11483 = ~1'b0 ;
  assign y11484 = ~1'b0 ;
  assign y11485 = ~n17858 ;
  assign y11486 = ~n17861 ;
  assign y11487 = ~1'b0 ;
  assign y11488 = ~n14489 ;
  assign y11489 = n17862 ;
  assign y11490 = ~n17865 ;
  assign y11491 = ~1'b0 ;
  assign y11492 = ~n17870 ;
  assign y11493 = n17871 ;
  assign y11494 = n17872 ;
  assign y11495 = ~1'b0 ;
  assign y11496 = ~n17873 ;
  assign y11497 = n2067 ;
  assign y11498 = ~1'b0 ;
  assign y11499 = ~n17874 ;
  assign y11500 = ~1'b0 ;
  assign y11501 = ~n17880 ;
  assign y11502 = ~1'b0 ;
  assign y11503 = ~n17881 ;
  assign y11504 = ~n4384 ;
  assign y11505 = n17882 ;
  assign y11506 = n17883 ;
  assign y11507 = ~1'b0 ;
  assign y11508 = ~1'b0 ;
  assign y11509 = ~1'b0 ;
  assign y11510 = ~1'b0 ;
  assign y11511 = ~n17885 ;
  assign y11512 = n17886 ;
  assign y11513 = n17888 ;
  assign y11514 = n17890 ;
  assign y11515 = ~1'b0 ;
  assign y11516 = 1'b0 ;
  assign y11517 = ~n17891 ;
  assign y11518 = ~1'b0 ;
  assign y11519 = ~n17894 ;
  assign y11520 = ~1'b0 ;
  assign y11521 = ~1'b0 ;
  assign y11522 = ~n17895 ;
  assign y11523 = ~n17897 ;
  assign y11524 = ~1'b0 ;
  assign y11525 = ~1'b0 ;
  assign y11526 = ~1'b0 ;
  assign y11527 = ~1'b0 ;
  assign y11528 = ~n17898 ;
  assign y11529 = ~1'b0 ;
  assign y11530 = n17458 ;
  assign y11531 = ~1'b0 ;
  assign y11532 = ~n2000 ;
  assign y11533 = ~n17907 ;
  assign y11534 = ~n17908 ;
  assign y11535 = n200 ;
  assign y11536 = ~n17914 ;
  assign y11537 = ~n4964 ;
  assign y11538 = n17916 ;
  assign y11539 = ~n17917 ;
  assign y11540 = ~1'b0 ;
  assign y11541 = ~1'b0 ;
  assign y11542 = ~1'b0 ;
  assign y11543 = ~1'b0 ;
  assign y11544 = ~n17920 ;
  assign y11545 = ~1'b0 ;
  assign y11546 = n3195 ;
  assign y11547 = ~n17923 ;
  assign y11548 = n17926 ;
  assign y11549 = ~n17951 ;
  assign y11550 = ~n17957 ;
  assign y11551 = n17958 ;
  assign y11552 = ~1'b0 ;
  assign y11553 = ~1'b0 ;
  assign y11554 = 1'b0 ;
  assign y11555 = n17959 ;
  assign y11556 = 1'b0 ;
  assign y11557 = ~1'b0 ;
  assign y11558 = ~1'b0 ;
  assign y11559 = ~n708 ;
  assign y11560 = ~n13866 ;
  assign y11561 = ~1'b0 ;
  assign y11562 = ~n17961 ;
  assign y11563 = ~n17963 ;
  assign y11564 = ~n17964 ;
  assign y11565 = ~n17966 ;
  assign y11566 = ~1'b0 ;
  assign y11567 = n17967 ;
  assign y11568 = n17968 ;
  assign y11569 = ~1'b0 ;
  assign y11570 = n17970 ;
  assign y11571 = ~n17971 ;
  assign y11572 = ~n17972 ;
  assign y11573 = ~n5168 ;
  assign y11574 = n17973 ;
  assign y11575 = n17974 ;
  assign y11576 = ~n17975 ;
  assign y11577 = n17977 ;
  assign y11578 = ~1'b0 ;
  assign y11579 = ~1'b0 ;
  assign y11580 = n17978 ;
  assign y11581 = ~1'b0 ;
  assign y11582 = n13507 ;
  assign y11583 = n17979 ;
  assign y11584 = n17980 ;
  assign y11585 = n17983 ;
  assign y11586 = ~1'b0 ;
  assign y11587 = ~1'b0 ;
  assign y11588 = ~n17986 ;
  assign y11589 = 1'b0 ;
  assign y11590 = 1'b0 ;
  assign y11591 = ~1'b0 ;
  assign y11592 = n17989 ;
  assign y11593 = n4265 ;
  assign y11594 = n8002 ;
  assign y11595 = ~1'b0 ;
  assign y11596 = ~n17991 ;
  assign y11597 = ~n14674 ;
  assign y11598 = ~1'b0 ;
  assign y11599 = ~n17992 ;
  assign y11600 = ~n7044 ;
  assign y11601 = ~1'b0 ;
  assign y11602 = ~n12484 ;
  assign y11603 = ~n17994 ;
  assign y11604 = ~1'b0 ;
  assign y11605 = ~n2542 ;
  assign y11606 = n17996 ;
  assign y11607 = ~1'b0 ;
  assign y11608 = n17998 ;
  assign y11609 = ~1'b0 ;
  assign y11610 = n18001 ;
  assign y11611 = ~1'b0 ;
  assign y11612 = n18002 ;
  assign y11613 = ~1'b0 ;
  assign y11614 = n18003 ;
  assign y11615 = ~1'b0 ;
  assign y11616 = ~1'b0 ;
  assign y11617 = n18005 ;
  assign y11618 = ~n18007 ;
  assign y11619 = n18008 ;
  assign y11620 = ~n18011 ;
  assign y11621 = ~1'b0 ;
  assign y11622 = ~1'b0 ;
  assign y11623 = ~n18017 ;
  assign y11624 = ~n18018 ;
  assign y11625 = ~n18019 ;
  assign y11626 = ~1'b0 ;
  assign y11627 = ~n18022 ;
  assign y11628 = n18024 ;
  assign y11629 = ~1'b0 ;
  assign y11630 = ~1'b0 ;
  assign y11631 = ~1'b0 ;
  assign y11632 = ~1'b0 ;
  assign y11633 = ~1'b0 ;
  assign y11634 = ~n5072 ;
  assign y11635 = n10968 ;
  assign y11636 = ~n18026 ;
  assign y11637 = n18027 ;
  assign y11638 = ~1'b0 ;
  assign y11639 = ~1'b0 ;
  assign y11640 = n2967 ;
  assign y11641 = ~1'b0 ;
  assign y11642 = ~1'b0 ;
  assign y11643 = n3898 ;
  assign y11644 = n18029 ;
  assign y11645 = ~n18030 ;
  assign y11646 = n18033 ;
  assign y11647 = n18034 ;
  assign y11648 = ~n18036 ;
  assign y11649 = n8665 ;
  assign y11650 = ~n18037 ;
  assign y11651 = ~1'b0 ;
  assign y11652 = ~1'b0 ;
  assign y11653 = ~n18039 ;
  assign y11654 = ~1'b0 ;
  assign y11655 = ~1'b0 ;
  assign y11656 = 1'b0 ;
  assign y11657 = n6824 ;
  assign y11658 = 1'b0 ;
  assign y11659 = n18040 ;
  assign y11660 = ~n4959 ;
  assign y11661 = ~n18041 ;
  assign y11662 = n18044 ;
  assign y11663 = 1'b0 ;
  assign y11664 = n18046 ;
  assign y11665 = ~1'b0 ;
  assign y11666 = n18047 ;
  assign y11667 = ~1'b0 ;
  assign y11668 = ~1'b0 ;
  assign y11669 = ~1'b0 ;
  assign y11670 = ~1'b0 ;
  assign y11671 = ~1'b0 ;
  assign y11672 = ~n18048 ;
  assign y11673 = ~n9635 ;
  assign y11674 = ~1'b0 ;
  assign y11675 = ~1'b0 ;
  assign y11676 = ~n18052 ;
  assign y11677 = n18053 ;
  assign y11678 = 1'b0 ;
  assign y11679 = ~n9991 ;
  assign y11680 = ~n18058 ;
  assign y11681 = ~1'b0 ;
  assign y11682 = ~1'b0 ;
  assign y11683 = ~n18060 ;
  assign y11684 = ~n18063 ;
  assign y11685 = ~n18066 ;
  assign y11686 = ~1'b0 ;
  assign y11687 = ~n18068 ;
  assign y11688 = ~1'b0 ;
  assign y11689 = ~1'b0 ;
  assign y11690 = ~1'b0 ;
  assign y11691 = ~1'b0 ;
  assign y11692 = ~1'b0 ;
  assign y11693 = n18069 ;
  assign y11694 = ~n18070 ;
  assign y11695 = ~n18071 ;
  assign y11696 = ~1'b0 ;
  assign y11697 = n18074 ;
  assign y11698 = 1'b0 ;
  assign y11699 = n2861 ;
  assign y11700 = 1'b0 ;
  assign y11701 = 1'b0 ;
  assign y11702 = ~n18078 ;
  assign y11703 = ~1'b0 ;
  assign y11704 = ~n18083 ;
  assign y11705 = ~n18085 ;
  assign y11706 = ~n18088 ;
  assign y11707 = ~n17722 ;
  assign y11708 = ~n18090 ;
  assign y11709 = ~1'b0 ;
  assign y11710 = n18091 ;
  assign y11711 = ~1'b0 ;
  assign y11712 = ~n18092 ;
  assign y11713 = n18097 ;
  assign y11714 = n994 ;
  assign y11715 = n18101 ;
  assign y11716 = n18102 ;
  assign y11717 = ~1'b0 ;
  assign y11718 = n18105 ;
  assign y11719 = n16834 ;
  assign y11720 = ~1'b0 ;
  assign y11721 = n18108 ;
  assign y11722 = ~n18109 ;
  assign y11723 = ~n18112 ;
  assign y11724 = n18113 ;
  assign y11725 = ~n18117 ;
  assign y11726 = ~n18119 ;
  assign y11727 = n18122 ;
  assign y11728 = ~1'b0 ;
  assign y11729 = ~1'b0 ;
  assign y11730 = ~n1070 ;
  assign y11731 = 1'b0 ;
  assign y11732 = ~n18123 ;
  assign y11733 = ~1'b0 ;
  assign y11734 = 1'b0 ;
  assign y11735 = ~n18126 ;
  assign y11736 = ~n18128 ;
  assign y11737 = ~n18134 ;
  assign y11738 = ~1'b0 ;
  assign y11739 = n18135 ;
  assign y11740 = n18137 ;
  assign y11741 = ~n18139 ;
  assign y11742 = ~n18143 ;
  assign y11743 = n18145 ;
  assign y11744 = ~n18146 ;
  assign y11745 = ~n18149 ;
  assign y11746 = n18153 ;
  assign y11747 = ~1'b0 ;
  assign y11748 = ~n18154 ;
  assign y11749 = ~1'b0 ;
  assign y11750 = ~n18156 ;
  assign y11751 = ~n18158 ;
  assign y11752 = ~n17523 ;
  assign y11753 = n18162 ;
  assign y11754 = n18164 ;
  assign y11755 = n18167 ;
  assign y11756 = n18173 ;
  assign y11757 = ~n18174 ;
  assign y11758 = ~1'b0 ;
  assign y11759 = ~1'b0 ;
  assign y11760 = ~n18178 ;
  assign y11761 = n18180 ;
  assign y11762 = n18184 ;
  assign y11763 = ~1'b0 ;
  assign y11764 = n18187 ;
  assign y11765 = n18191 ;
  assign y11766 = n18192 ;
  assign y11767 = n18193 ;
  assign y11768 = ~1'b0 ;
  assign y11769 = ~1'b0 ;
  assign y11770 = ~1'b0 ;
  assign y11771 = ~n5005 ;
  assign y11772 = ~n18194 ;
  assign y11773 = ~1'b0 ;
  assign y11774 = n18196 ;
  assign y11775 = 1'b0 ;
  assign y11776 = ~1'b0 ;
  assign y11777 = ~1'b0 ;
  assign y11778 = ~1'b0 ;
  assign y11779 = ~1'b0 ;
  assign y11780 = n18197 ;
  assign y11781 = n18203 ;
  assign y11782 = ~n18204 ;
  assign y11783 = n18205 ;
  assign y11784 = n2291 ;
  assign y11785 = n18208 ;
  assign y11786 = ~1'b0 ;
  assign y11787 = ~n18209 ;
  assign y11788 = ~1'b0 ;
  assign y11789 = ~1'b0 ;
  assign y11790 = ~1'b0 ;
  assign y11791 = ~n18210 ;
  assign y11792 = ~1'b0 ;
  assign y11793 = ~n18212 ;
  assign y11794 = ~n18219 ;
  assign y11795 = ~n18221 ;
  assign y11796 = ~1'b0 ;
  assign y11797 = 1'b0 ;
  assign y11798 = n18222 ;
  assign y11799 = ~n18224 ;
  assign y11800 = n18228 ;
  assign y11801 = n18230 ;
  assign y11802 = n18231 ;
  assign y11803 = ~n18232 ;
  assign y11804 = ~n18236 ;
  assign y11805 = ~n18238 ;
  assign y11806 = n18241 ;
  assign y11807 = ~1'b0 ;
  assign y11808 = ~n6274 ;
  assign y11809 = ~n5972 ;
  assign y11810 = ~n18244 ;
  assign y11811 = ~n18245 ;
  assign y11812 = n18246 ;
  assign y11813 = ~1'b0 ;
  assign y11814 = n18252 ;
  assign y11815 = ~n18258 ;
  assign y11816 = ~n18259 ;
  assign y11817 = ~1'b0 ;
  assign y11818 = ~1'b0 ;
  assign y11819 = ~1'b0 ;
  assign y11820 = n18260 ;
  assign y11821 = ~1'b0 ;
  assign y11822 = ~1'b0 ;
  assign y11823 = ~1'b0 ;
  assign y11824 = ~1'b0 ;
  assign y11825 = ~1'b0 ;
  assign y11826 = ~1'b0 ;
  assign y11827 = ~1'b0 ;
  assign y11828 = n18261 ;
  assign y11829 = 1'b0 ;
  assign y11830 = n18265 ;
  assign y11831 = ~n18268 ;
  assign y11832 = ~1'b0 ;
  assign y11833 = n18270 ;
  assign y11834 = ~n18272 ;
  assign y11835 = n18277 ;
  assign y11836 = n18280 ;
  assign y11837 = ~1'b0 ;
  assign y11838 = ~1'b0 ;
  assign y11839 = ~n18282 ;
  assign y11840 = ~1'b0 ;
  assign y11841 = n18285 ;
  assign y11842 = ~1'b0 ;
  assign y11843 = ~1'b0 ;
  assign y11844 = n18286 ;
  assign y11845 = ~1'b0 ;
  assign y11846 = n18290 ;
  assign y11847 = n18294 ;
  assign y11848 = n18295 ;
  assign y11849 = ~1'b0 ;
  assign y11850 = ~n18296 ;
  assign y11851 = n18299 ;
  assign y11852 = n18301 ;
  assign y11853 = ~1'b0 ;
  assign y11854 = ~n18304 ;
  assign y11855 = ~n707 ;
  assign y11856 = ~n18306 ;
  assign y11857 = ~n18310 ;
  assign y11858 = ~1'b0 ;
  assign y11859 = n12834 ;
  assign y11860 = ~n11110 ;
  assign y11861 = ~n6980 ;
  assign y11862 = n18313 ;
  assign y11863 = ~n18314 ;
  assign y11864 = ~1'b0 ;
  assign y11865 = n15904 ;
  assign y11866 = ~n5239 ;
  assign y11867 = ~n18317 ;
  assign y11868 = n18320 ;
  assign y11869 = n18327 ;
  assign y11870 = ~1'b0 ;
  assign y11871 = n18328 ;
  assign y11872 = n18329 ;
  assign y11873 = ~1'b0 ;
  assign y11874 = ~n2107 ;
  assign y11875 = n18332 ;
  assign y11876 = n18333 ;
  assign y11877 = n18334 ;
  assign y11878 = ~1'b0 ;
  assign y11879 = n18336 ;
  assign y11880 = ~1'b0 ;
  assign y11881 = n18339 ;
  assign y11882 = n3687 ;
  assign y11883 = 1'b0 ;
  assign y11884 = ~n18340 ;
  assign y11885 = ~n18342 ;
  assign y11886 = ~1'b0 ;
  assign y11887 = ~n18345 ;
  assign y11888 = ~n10445 ;
  assign y11889 = n18348 ;
  assign y11890 = ~1'b0 ;
  assign y11891 = ~n18349 ;
  assign y11892 = ~1'b0 ;
  assign y11893 = ~n16786 ;
  assign y11894 = ~n18353 ;
  assign y11895 = ~n2493 ;
  assign y11896 = ~1'b0 ;
  assign y11897 = ~n18357 ;
  assign y11898 = n18358 ;
  assign y11899 = n18360 ;
  assign y11900 = ~1'b0 ;
  assign y11901 = n18361 ;
  assign y11902 = ~n18364 ;
  assign y11903 = ~1'b0 ;
  assign y11904 = n18368 ;
  assign y11905 = ~1'b0 ;
  assign y11906 = ~1'b0 ;
  assign y11907 = n18369 ;
  assign y11908 = n9252 ;
  assign y11909 = ~n18376 ;
  assign y11910 = n18378 ;
  assign y11911 = ~1'b0 ;
  assign y11912 = ~n18380 ;
  assign y11913 = ~n18382 ;
  assign y11914 = ~1'b0 ;
  assign y11915 = ~1'b0 ;
  assign y11916 = 1'b0 ;
  assign y11917 = n3462 ;
  assign y11918 = ~n645 ;
  assign y11919 = ~n18383 ;
  assign y11920 = ~1'b0 ;
  assign y11921 = n18386 ;
  assign y11922 = ~1'b0 ;
  assign y11923 = ~n18390 ;
  assign y11924 = 1'b0 ;
  assign y11925 = 1'b0 ;
  assign y11926 = ~n18395 ;
  assign y11927 = ~n18397 ;
  assign y11928 = ~n18398 ;
  assign y11929 = n18401 ;
  assign y11930 = n18404 ;
  assign y11931 = n18406 ;
  assign y11932 = ~1'b0 ;
  assign y11933 = ~1'b0 ;
  assign y11934 = ~1'b0 ;
  assign y11935 = ~n18408 ;
  assign y11936 = ~n18410 ;
  assign y11937 = ~1'b0 ;
  assign y11938 = ~n18412 ;
  assign y11939 = n3862 ;
  assign y11940 = n18413 ;
  assign y11941 = ~1'b0 ;
  assign y11942 = ~n542 ;
  assign y11943 = ~n18415 ;
  assign y11944 = n1013 ;
  assign y11945 = ~1'b0 ;
  assign y11946 = ~n18421 ;
  assign y11947 = ~n14006 ;
  assign y11948 = n18425 ;
  assign y11949 = n18428 ;
  assign y11950 = ~1'b0 ;
  assign y11951 = ~1'b0 ;
  assign y11952 = ~1'b0 ;
  assign y11953 = ~n16081 ;
  assign y11954 = ~1'b0 ;
  assign y11955 = ~1'b0 ;
  assign y11956 = ~1'b0 ;
  assign y11957 = ~n18429 ;
  assign y11958 = n18433 ;
  assign y11959 = n18437 ;
  assign y11960 = n18438 ;
  assign y11961 = ~1'b0 ;
  assign y11962 = n11228 ;
  assign y11963 = ~1'b0 ;
  assign y11964 = n18441 ;
  assign y11965 = ~1'b0 ;
  assign y11966 = n18442 ;
  assign y11967 = ~1'b0 ;
  assign y11968 = ~n18443 ;
  assign y11969 = n18445 ;
  assign y11970 = 1'b0 ;
  assign y11971 = n18446 ;
  assign y11972 = ~1'b0 ;
  assign y11973 = ~n18448 ;
  assign y11974 = n18449 ;
  assign y11975 = ~n18452 ;
  assign y11976 = n18455 ;
  assign y11977 = ~n18457 ;
  assign y11978 = ~1'b0 ;
  assign y11979 = ~n18458 ;
  assign y11980 = n18460 ;
  assign y11981 = ~n18461 ;
  assign y11982 = ~x76 ;
  assign y11983 = ~n18463 ;
  assign y11984 = ~1'b0 ;
  assign y11985 = ~n18467 ;
  assign y11986 = ~1'b0 ;
  assign y11987 = ~1'b0 ;
  assign y11988 = ~n18469 ;
  assign y11989 = ~n18473 ;
  assign y11990 = n18475 ;
  assign y11991 = ~1'b0 ;
  assign y11992 = n18477 ;
  assign y11993 = ~1'b0 ;
  assign y11994 = ~n18480 ;
  assign y11995 = ~n18481 ;
  assign y11996 = ~n18483 ;
  assign y11997 = n18484 ;
  assign y11998 = n18485 ;
  assign y11999 = ~1'b0 ;
  assign y12000 = ~1'b0 ;
  assign y12001 = ~1'b0 ;
  assign y12002 = ~n18487 ;
  assign y12003 = ~n10018 ;
  assign y12004 = n18489 ;
  assign y12005 = ~n18490 ;
  assign y12006 = n18492 ;
  assign y12007 = ~n18493 ;
  assign y12008 = n18494 ;
  assign y12009 = n18496 ;
  assign y12010 = ~n18497 ;
  assign y12011 = ~1'b0 ;
  assign y12012 = ~n7348 ;
  assign y12013 = ~1'b0 ;
  assign y12014 = n18498 ;
  assign y12015 = n18504 ;
  assign y12016 = ~n18505 ;
  assign y12017 = ~1'b0 ;
  assign y12018 = ~1'b0 ;
  assign y12019 = n18506 ;
  assign y12020 = ~n18511 ;
  assign y12021 = ~1'b0 ;
  assign y12022 = ~n18514 ;
  assign y12023 = ~1'b0 ;
  assign y12024 = n18517 ;
  assign y12025 = n18518 ;
  assign y12026 = ~n18519 ;
  assign y12027 = ~1'b0 ;
  assign y12028 = ~n18520 ;
  assign y12029 = ~n6782 ;
  assign y12030 = n4602 ;
  assign y12031 = ~1'b0 ;
  assign y12032 = ~1'b0 ;
  assign y12033 = ~n5423 ;
  assign y12034 = ~n18522 ;
  assign y12035 = ~1'b0 ;
  assign y12036 = ~1'b0 ;
  assign y12037 = n18524 ;
  assign y12038 = ~n18525 ;
  assign y12039 = n18527 ;
  assign y12040 = ~n18528 ;
  assign y12041 = n18530 ;
  assign y12042 = n18533 ;
  assign y12043 = n18535 ;
  assign y12044 = ~n18537 ;
  assign y12045 = ~n18538 ;
  assign y12046 = ~1'b0 ;
  assign y12047 = ~1'b0 ;
  assign y12048 = ~n18540 ;
  assign y12049 = ~n18542 ;
  assign y12050 = ~n9506 ;
  assign y12051 = ~n18548 ;
  assign y12052 = ~n8302 ;
  assign y12053 = n18551 ;
  assign y12054 = n18552 ;
  assign y12055 = ~1'b0 ;
  assign y12056 = n15569 ;
  assign y12057 = n18554 ;
  assign y12058 = ~1'b0 ;
  assign y12059 = ~1'b0 ;
  assign y12060 = ~1'b0 ;
  assign y12061 = 1'b0 ;
  assign y12062 = n18555 ;
  assign y12063 = ~n18558 ;
  assign y12064 = ~n6495 ;
  assign y12065 = ~n18559 ;
  assign y12066 = ~n18560 ;
  assign y12067 = n18561 ;
  assign y12068 = ~n18562 ;
  assign y12069 = ~n18563 ;
  assign y12070 = ~1'b0 ;
  assign y12071 = ~n18564 ;
  assign y12072 = n11881 ;
  assign y12073 = ~n8221 ;
  assign y12074 = n8999 ;
  assign y12075 = ~1'b0 ;
  assign y12076 = ~1'b0 ;
  assign y12077 = n18566 ;
  assign y12078 = n18569 ;
  assign y12079 = ~1'b0 ;
  assign y12080 = n18576 ;
  assign y12081 = n18579 ;
  assign y12082 = ~n18581 ;
  assign y12083 = n18582 ;
  assign y12084 = n18589 ;
  assign y12085 = 1'b0 ;
  assign y12086 = ~1'b0 ;
  assign y12087 = ~1'b0 ;
  assign y12088 = n18590 ;
  assign y12089 = n7341 ;
  assign y12090 = n18592 ;
  assign y12091 = ~n13326 ;
  assign y12092 = ~1'b0 ;
  assign y12093 = n18594 ;
  assign y12094 = ~n7650 ;
  assign y12095 = ~1'b0 ;
  assign y12096 = ~x6 ;
  assign y12097 = ~n3904 ;
  assign y12098 = ~n18595 ;
  assign y12099 = ~1'b0 ;
  assign y12100 = ~1'b0 ;
  assign y12101 = ~n18596 ;
  assign y12102 = ~1'b0 ;
  assign y12103 = n18600 ;
  assign y12104 = n18605 ;
  assign y12105 = ~n18607 ;
  assign y12106 = ~1'b0 ;
  assign y12107 = ~1'b0 ;
  assign y12108 = ~x8 ;
  assign y12109 = ~1'b0 ;
  assign y12110 = ~1'b0 ;
  assign y12111 = n18609 ;
  assign y12112 = ~1'b0 ;
  assign y12113 = ~n18612 ;
  assign y12114 = ~n18613 ;
  assign y12115 = n18614 ;
  assign y12116 = ~n18617 ;
  assign y12117 = n18619 ;
  assign y12118 = ~1'b0 ;
  assign y12119 = ~1'b0 ;
  assign y12120 = n18621 ;
  assign y12121 = ~n18623 ;
  assign y12122 = ~1'b0 ;
  assign y12123 = ~n18624 ;
  assign y12124 = ~1'b0 ;
  assign y12125 = ~n18625 ;
  assign y12126 = ~n18626 ;
  assign y12127 = n18630 ;
  assign y12128 = ~1'b0 ;
  assign y12129 = n18633 ;
  assign y12130 = ~n18642 ;
  assign y12131 = n18643 ;
  assign y12132 = n18646 ;
  assign y12133 = ~1'b0 ;
  assign y12134 = n18648 ;
  assign y12135 = n18655 ;
  assign y12136 = n18656 ;
  assign y12137 = n18657 ;
  assign y12138 = ~n5234 ;
  assign y12139 = ~n18658 ;
  assign y12140 = ~n18660 ;
  assign y12141 = ~1'b0 ;
  assign y12142 = ~1'b0 ;
  assign y12143 = ~n18662 ;
  assign y12144 = ~1'b0 ;
  assign y12145 = ~1'b0 ;
  assign y12146 = n7139 ;
  assign y12147 = ~n18666 ;
  assign y12148 = ~1'b0 ;
  assign y12149 = ~1'b0 ;
  assign y12150 = ~1'b0 ;
  assign y12151 = 1'b0 ;
  assign y12152 = ~1'b0 ;
  assign y12153 = ~n12339 ;
  assign y12154 = n18667 ;
  assign y12155 = n18669 ;
  assign y12156 = ~1'b0 ;
  assign y12157 = ~1'b0 ;
  assign y12158 = ~1'b0 ;
  assign y12159 = ~1'b0 ;
  assign y12160 = ~n18671 ;
  assign y12161 = ~n18672 ;
  assign y12162 = ~n18674 ;
  assign y12163 = ~n18676 ;
  assign y12164 = ~n3644 ;
  assign y12165 = ~1'b0 ;
  assign y12166 = ~n18679 ;
  assign y12167 = n18688 ;
  assign y12168 = n18692 ;
  assign y12169 = 1'b0 ;
  assign y12170 = ~1'b0 ;
  assign y12171 = ~1'b0 ;
  assign y12172 = n1887 ;
  assign y12173 = ~n18693 ;
  assign y12174 = n18696 ;
  assign y12175 = ~1'b0 ;
  assign y12176 = ~1'b0 ;
  assign y12177 = ~n18698 ;
  assign y12178 = n18699 ;
  assign y12179 = ~n18700 ;
  assign y12180 = ~1'b0 ;
  assign y12181 = n18701 ;
  assign y12182 = ~n7659 ;
  assign y12183 = ~1'b0 ;
  assign y12184 = n18702 ;
  assign y12185 = ~1'b0 ;
  assign y12186 = ~1'b0 ;
  assign y12187 = ~n18704 ;
  assign y12188 = n18706 ;
  assign y12189 = n4312 ;
  assign y12190 = ~1'b0 ;
  assign y12191 = ~n12602 ;
  assign y12192 = ~n18708 ;
  assign y12193 = ~n11787 ;
  assign y12194 = ~1'b0 ;
  assign y12195 = n18709 ;
  assign y12196 = ~1'b0 ;
  assign y12197 = ~1'b0 ;
  assign y12198 = ~n18713 ;
  assign y12199 = ~n18714 ;
  assign y12200 = n18715 ;
  assign y12201 = n18719 ;
  assign y12202 = ~n18720 ;
  assign y12203 = ~1'b0 ;
  assign y12204 = ~1'b0 ;
  assign y12205 = n7242 ;
  assign y12206 = n18722 ;
  assign y12207 = n4805 ;
  assign y12208 = n18723 ;
  assign y12209 = ~n18725 ;
  assign y12210 = ~n18727 ;
  assign y12211 = ~1'b0 ;
  assign y12212 = 1'b0 ;
  assign y12213 = ~n2972 ;
  assign y12214 = ~1'b0 ;
  assign y12215 = ~1'b0 ;
  assign y12216 = ~n18731 ;
  assign y12217 = n8682 ;
  assign y12218 = ~n13914 ;
  assign y12219 = n18732 ;
  assign y12220 = ~1'b0 ;
  assign y12221 = n18736 ;
  assign y12222 = ~n8502 ;
  assign y12223 = n18741 ;
  assign y12224 = ~1'b0 ;
  assign y12225 = ~n18742 ;
  assign y12226 = ~1'b0 ;
  assign y12227 = ~1'b0 ;
  assign y12228 = ~n18744 ;
  assign y12229 = ~n18746 ;
  assign y12230 = n18747 ;
  assign y12231 = ~n18750 ;
  assign y12232 = n18752 ;
  assign y12233 = ~n18755 ;
  assign y12234 = ~n18758 ;
  assign y12235 = ~n18759 ;
  assign y12236 = ~1'b0 ;
  assign y12237 = n18762 ;
  assign y12238 = ~n18764 ;
  assign y12239 = n18766 ;
  assign y12240 = n18769 ;
  assign y12241 = n3230 ;
  assign y12242 = ~1'b0 ;
  assign y12243 = ~1'b0 ;
  assign y12244 = ~1'b0 ;
  assign y12245 = n18772 ;
  assign y12246 = ~1'b0 ;
  assign y12247 = ~n3120 ;
  assign y12248 = ~n18774 ;
  assign y12249 = ~n18775 ;
  assign y12250 = n18776 ;
  assign y12251 = ~n18778 ;
  assign y12252 = ~n18779 ;
  assign y12253 = ~n18782 ;
  assign y12254 = n11423 ;
  assign y12255 = ~1'b0 ;
  assign y12256 = 1'b0 ;
  assign y12257 = ~n18783 ;
  assign y12258 = ~1'b0 ;
  assign y12259 = n18785 ;
  assign y12260 = ~1'b0 ;
  assign y12261 = ~1'b0 ;
  assign y12262 = n18788 ;
  assign y12263 = ~n18789 ;
  assign y12264 = n18790 ;
  assign y12265 = ~n18791 ;
  assign y12266 = ~n18795 ;
  assign y12267 = n18796 ;
  assign y12268 = ~n18797 ;
  assign y12269 = n18798 ;
  assign y12270 = ~n18801 ;
  assign y12271 = ~n18803 ;
  assign y12272 = n16192 ;
  assign y12273 = n18805 ;
  assign y12274 = ~1'b0 ;
  assign y12275 = n14663 ;
  assign y12276 = ~1'b0 ;
  assign y12277 = ~1'b0 ;
  assign y12278 = ~1'b0 ;
  assign y12279 = n18808 ;
  assign y12280 = ~n18810 ;
  assign y12281 = ~1'b0 ;
  assign y12282 = ~n18812 ;
  assign y12283 = ~n18816 ;
  assign y12284 = ~1'b0 ;
  assign y12285 = n18819 ;
  assign y12286 = ~1'b0 ;
  assign y12287 = ~n18820 ;
  assign y12288 = n18821 ;
  assign y12289 = ~1'b0 ;
  assign y12290 = n18822 ;
  assign y12291 = ~1'b0 ;
  assign y12292 = ~n18826 ;
  assign y12293 = ~1'b0 ;
  assign y12294 = n18827 ;
  assign y12295 = ~n18829 ;
  assign y12296 = ~n18832 ;
  assign y12297 = ~n18834 ;
  assign y12298 = n18835 ;
  assign y12299 = ~n18838 ;
  assign y12300 = n18839 ;
  assign y12301 = n18841 ;
  assign y12302 = n18842 ;
  assign y12303 = ~n18845 ;
  assign y12304 = ~1'b0 ;
  assign y12305 = ~1'b0 ;
  assign y12306 = n18847 ;
  assign y12307 = ~n8723 ;
  assign y12308 = n18849 ;
  assign y12309 = n18853 ;
  assign y12310 = ~1'b0 ;
  assign y12311 = n18858 ;
  assign y12312 = ~n18861 ;
  assign y12313 = ~1'b0 ;
  assign y12314 = ~n18862 ;
  assign y12315 = n18863 ;
  assign y12316 = ~1'b0 ;
  assign y12317 = n18865 ;
  assign y12318 = n18866 ;
  assign y12319 = n17143 ;
  assign y12320 = ~n18867 ;
  assign y12321 = ~n18868 ;
  assign y12322 = ~n18870 ;
  assign y12323 = ~1'b0 ;
  assign y12324 = ~1'b0 ;
  assign y12325 = ~1'b0 ;
  assign y12326 = ~n18871 ;
  assign y12327 = ~1'b0 ;
  assign y12328 = ~n18873 ;
  assign y12329 = ~1'b0 ;
  assign y12330 = n18874 ;
  assign y12331 = ~n18877 ;
  assign y12332 = n18879 ;
  assign y12333 = ~n18883 ;
  assign y12334 = n18884 ;
  assign y12335 = n18885 ;
  assign y12336 = n18888 ;
  assign y12337 = n18890 ;
  assign y12338 = n18891 ;
  assign y12339 = n18892 ;
  assign y12340 = ~n18895 ;
  assign y12341 = ~n18898 ;
  assign y12342 = ~1'b0 ;
  assign y12343 = ~1'b0 ;
  assign y12344 = ~n18901 ;
  assign y12345 = ~1'b0 ;
  assign y12346 = n18904 ;
  assign y12347 = ~n6638 ;
  assign y12348 = ~1'b0 ;
  assign y12349 = ~n18906 ;
  assign y12350 = ~n2459 ;
  assign y12351 = n786 ;
  assign y12352 = n14882 ;
  assign y12353 = ~n11537 ;
  assign y12354 = ~1'b0 ;
  assign y12355 = ~1'b0 ;
  assign y12356 = n18908 ;
  assign y12357 = n18909 ;
  assign y12358 = 1'b0 ;
  assign y12359 = ~1'b0 ;
  assign y12360 = ~n18910 ;
  assign y12361 = ~1'b0 ;
  assign y12362 = n18912 ;
  assign y12363 = n6842 ;
  assign y12364 = ~n18915 ;
  assign y12365 = n18916 ;
  assign y12366 = ~1'b0 ;
  assign y12367 = ~1'b0 ;
  assign y12368 = ~n18917 ;
  assign y12369 = ~1'b0 ;
  assign y12370 = n18919 ;
  assign y12371 = ~n18921 ;
  assign y12372 = ~1'b0 ;
  assign y12373 = ~1'b0 ;
  assign y12374 = n18922 ;
  assign y12375 = ~n18926 ;
  assign y12376 = ~1'b0 ;
  assign y12377 = ~n18928 ;
  assign y12378 = ~n10410 ;
  assign y12379 = ~1'b0 ;
  assign y12380 = n18929 ;
  assign y12381 = ~1'b0 ;
  assign y12382 = ~1'b0 ;
  assign y12383 = n18931 ;
  assign y12384 = ~n18934 ;
  assign y12385 = ~n18941 ;
  assign y12386 = n18942 ;
  assign y12387 = n18944 ;
  assign y12388 = ~1'b0 ;
  assign y12389 = ~1'b0 ;
  assign y12390 = ~1'b0 ;
  assign y12391 = n18946 ;
  assign y12392 = ~1'b0 ;
  assign y12393 = ~n3890 ;
  assign y12394 = ~n18950 ;
  assign y12395 = n18952 ;
  assign y12396 = n18955 ;
  assign y12397 = ~1'b0 ;
  assign y12398 = ~1'b0 ;
  assign y12399 = ~n18956 ;
  assign y12400 = n18958 ;
  assign y12401 = n4306 ;
  assign y12402 = ~n18959 ;
  assign y12403 = n18962 ;
  assign y12404 = ~1'b0 ;
  assign y12405 = n18963 ;
  assign y12406 = ~1'b0 ;
  assign y12407 = ~n18965 ;
  assign y12408 = ~1'b0 ;
  assign y12409 = ~1'b0 ;
  assign y12410 = ~1'b0 ;
  assign y12411 = n18966 ;
  assign y12412 = ~1'b0 ;
  assign y12413 = ~n18967 ;
  assign y12414 = n18970 ;
  assign y12415 = n18971 ;
  assign y12416 = n18973 ;
  assign y12417 = ~n18975 ;
  assign y12418 = ~n18976 ;
  assign y12419 = ~n18977 ;
  assign y12420 = ~1'b0 ;
  assign y12421 = ~n18994 ;
  assign y12422 = ~n18996 ;
  assign y12423 = ~n18997 ;
  assign y12424 = ~n18998 ;
  assign y12425 = n19000 ;
  assign y12426 = ~n19001 ;
  assign y12427 = n7943 ;
  assign y12428 = ~1'b0 ;
  assign y12429 = ~1'b0 ;
  assign y12430 = n19019 ;
  assign y12431 = n19020 ;
  assign y12432 = n19021 ;
  assign y12433 = ~n717 ;
  assign y12434 = ~1'b0 ;
  assign y12435 = ~1'b0 ;
  assign y12436 = ~n19022 ;
  assign y12437 = ~1'b0 ;
  assign y12438 = ~1'b0 ;
  assign y12439 = ~1'b0 ;
  assign y12440 = n2343 ;
  assign y12441 = ~1'b0 ;
  assign y12442 = ~1'b0 ;
  assign y12443 = ~n19023 ;
  assign y12444 = ~n19031 ;
  assign y12445 = ~n19034 ;
  assign y12446 = n19035 ;
  assign y12447 = ~1'b0 ;
  assign y12448 = n2038 ;
  assign y12449 = n19041 ;
  assign y12450 = n19042 ;
  assign y12451 = n19044 ;
  assign y12452 = n19046 ;
  assign y12453 = n19047 ;
  assign y12454 = ~1'b0 ;
  assign y12455 = ~n1351 ;
  assign y12456 = ~n19048 ;
  assign y12457 = ~n19052 ;
  assign y12458 = ~1'b0 ;
  assign y12459 = n9839 ;
  assign y12460 = ~1'b0 ;
  assign y12461 = n19054 ;
  assign y12462 = n610 ;
  assign y12463 = ~n19055 ;
  assign y12464 = n19057 ;
  assign y12465 = ~n19059 ;
  assign y12466 = n19063 ;
  assign y12467 = ~n19067 ;
  assign y12468 = n19071 ;
  assign y12469 = ~n19072 ;
  assign y12470 = n19074 ;
  assign y12471 = ~1'b0 ;
  assign y12472 = n19076 ;
  assign y12473 = n19078 ;
  assign y12474 = ~n19079 ;
  assign y12475 = ~n19081 ;
  assign y12476 = ~n19083 ;
  assign y12477 = ~1'b0 ;
  assign y12478 = n19085 ;
  assign y12479 = n19087 ;
  assign y12480 = ~1'b0 ;
  assign y12481 = n1563 ;
  assign y12482 = ~1'b0 ;
  assign y12483 = 1'b0 ;
  assign y12484 = n19092 ;
  assign y12485 = n19093 ;
  assign y12486 = n19095 ;
  assign y12487 = ~1'b0 ;
  assign y12488 = n19097 ;
  assign y12489 = ~n19100 ;
  assign y12490 = ~1'b0 ;
  assign y12491 = n19102 ;
  assign y12492 = ~1'b0 ;
  assign y12493 = n19103 ;
  assign y12494 = n19105 ;
  assign y12495 = ~n19109 ;
  assign y12496 = ~1'b0 ;
  assign y12497 = ~1'b0 ;
  assign y12498 = ~n19110 ;
  assign y12499 = ~1'b0 ;
  assign y12500 = ~n19115 ;
  assign y12501 = ~n19119 ;
  assign y12502 = ~n19120 ;
  assign y12503 = 1'b0 ;
  assign y12504 = ~1'b0 ;
  assign y12505 = ~n19122 ;
  assign y12506 = ~1'b0 ;
  assign y12507 = ~n8504 ;
  assign y12508 = n19125 ;
  assign y12509 = ~n19129 ;
  assign y12510 = n19131 ;
  assign y12511 = ~n19133 ;
  assign y12512 = n19139 ;
  assign y12513 = ~n19141 ;
  assign y12514 = ~n7032 ;
  assign y12515 = ~1'b0 ;
  assign y12516 = ~n19142 ;
  assign y12517 = ~1'b0 ;
  assign y12518 = n19146 ;
  assign y12519 = ~1'b0 ;
  assign y12520 = 1'b0 ;
  assign y12521 = ~n19149 ;
  assign y12522 = ~1'b0 ;
  assign y12523 = n19150 ;
  assign y12524 = n19153 ;
  assign y12525 = ~1'b0 ;
  assign y12526 = ~n19154 ;
  assign y12527 = n19156 ;
  assign y12528 = ~n19158 ;
  assign y12529 = n19161 ;
  assign y12530 = ~n19163 ;
  assign y12531 = 1'b0 ;
  assign y12532 = n1387 ;
  assign y12533 = ~1'b0 ;
  assign y12534 = n19165 ;
  assign y12535 = ~n19166 ;
  assign y12536 = ~1'b0 ;
  assign y12537 = ~1'b0 ;
  assign y12538 = ~1'b0 ;
  assign y12539 = ~1'b0 ;
  assign y12540 = ~1'b0 ;
  assign y12541 = n3041 ;
  assign y12542 = ~1'b0 ;
  assign y12543 = n19167 ;
  assign y12544 = n19170 ;
  assign y12545 = ~n19173 ;
  assign y12546 = 1'b0 ;
  assign y12547 = ~n19174 ;
  assign y12548 = 1'b0 ;
  assign y12549 = ~n19177 ;
  assign y12550 = ~1'b0 ;
  assign y12551 = 1'b0 ;
  assign y12552 = n5374 ;
  assign y12553 = ~n19180 ;
  assign y12554 = ~n19181 ;
  assign y12555 = ~n19182 ;
  assign y12556 = ~n19185 ;
  assign y12557 = n19186 ;
  assign y12558 = n19189 ;
  assign y12559 = ~n19192 ;
  assign y12560 = n19193 ;
  assign y12561 = n4804 ;
  assign y12562 = ~n19199 ;
  assign y12563 = n19203 ;
  assign y12564 = ~1'b0 ;
  assign y12565 = ~n19205 ;
  assign y12566 = ~n19208 ;
  assign y12567 = ~n6539 ;
  assign y12568 = ~1'b0 ;
  assign y12569 = ~n19209 ;
  assign y12570 = n19210 ;
  assign y12571 = n19211 ;
  assign y12572 = n19213 ;
  assign y12573 = ~1'b0 ;
  assign y12574 = ~1'b0 ;
  assign y12575 = ~1'b0 ;
  assign y12576 = 1'b0 ;
  assign y12577 = ~n19219 ;
  assign y12578 = ~n19222 ;
  assign y12579 = n1628 ;
  assign y12580 = n19224 ;
  assign y12581 = ~1'b0 ;
  assign y12582 = ~1'b0 ;
  assign y12583 = ~n19226 ;
  assign y12584 = ~1'b0 ;
  assign y12585 = ~1'b0 ;
  assign y12586 = ~n17530 ;
  assign y12587 = ~1'b0 ;
  assign y12588 = 1'b0 ;
  assign y12589 = n19227 ;
  assign y12590 = ~1'b0 ;
  assign y12591 = ~n19230 ;
  assign y12592 = n14038 ;
  assign y12593 = ~1'b0 ;
  assign y12594 = n19234 ;
  assign y12595 = n19238 ;
  assign y12596 = 1'b0 ;
  assign y12597 = ~1'b0 ;
  assign y12598 = 1'b0 ;
  assign y12599 = ~n19242 ;
  assign y12600 = ~n19244 ;
  assign y12601 = ~n19246 ;
  assign y12602 = ~1'b0 ;
  assign y12603 = ~n19247 ;
  assign y12604 = ~1'b0 ;
  assign y12605 = ~n19250 ;
  assign y12606 = n2936 ;
  assign y12607 = ~1'b0 ;
  assign y12608 = ~n19251 ;
  assign y12609 = n19262 ;
  assign y12610 = 1'b0 ;
  assign y12611 = ~1'b0 ;
  assign y12612 = n19264 ;
  assign y12613 = n19265 ;
  assign y12614 = n19267 ;
  assign y12615 = ~n19269 ;
  assign y12616 = ~1'b0 ;
  assign y12617 = ~n19270 ;
  assign y12618 = ~n12101 ;
  assign y12619 = ~n19272 ;
  assign y12620 = ~1'b0 ;
  assign y12621 = ~1'b0 ;
  assign y12622 = ~n19276 ;
  assign y12623 = n19055 ;
  assign y12624 = ~1'b0 ;
  assign y12625 = ~1'b0 ;
  assign y12626 = n1610 ;
  assign y12627 = ~n19277 ;
  assign y12628 = n8015 ;
  assign y12629 = ~1'b0 ;
  assign y12630 = n19280 ;
  assign y12631 = n19282 ;
  assign y12632 = ~1'b0 ;
  assign y12633 = ~1'b0 ;
  assign y12634 = ~n19283 ;
  assign y12635 = ~n19284 ;
  assign y12636 = ~1'b0 ;
  assign y12637 = ~n19285 ;
  assign y12638 = ~n19293 ;
  assign y12639 = ~1'b0 ;
  assign y12640 = n19295 ;
  assign y12641 = ~n238 ;
  assign y12642 = n5235 ;
  assign y12643 = n6197 ;
  assign y12644 = ~1'b0 ;
  assign y12645 = ~n19298 ;
  assign y12646 = n19300 ;
  assign y12647 = 1'b0 ;
  assign y12648 = n1432 ;
  assign y12649 = n19302 ;
  assign y12650 = ~1'b0 ;
  assign y12651 = ~n5961 ;
  assign y12652 = n19303 ;
  assign y12653 = ~n19306 ;
  assign y12654 = n10612 ;
  assign y12655 = ~n8340 ;
  assign y12656 = n17271 ;
  assign y12657 = n19308 ;
  assign y12658 = ~1'b0 ;
  assign y12659 = n19309 ;
  assign y12660 = n19310 ;
  assign y12661 = n19312 ;
  assign y12662 = n19313 ;
  assign y12663 = ~n19314 ;
  assign y12664 = ~1'b0 ;
  assign y12665 = ~1'b0 ;
  assign y12666 = n19316 ;
  assign y12667 = ~1'b0 ;
  assign y12668 = n19317 ;
  assign y12669 = n13034 ;
  assign y12670 = n19318 ;
  assign y12671 = 1'b0 ;
  assign y12672 = n19321 ;
  assign y12673 = ~1'b0 ;
  assign y12674 = ~n19324 ;
  assign y12675 = ~n19327 ;
  assign y12676 = ~1'b0 ;
  assign y12677 = n19328 ;
  assign y12678 = ~1'b0 ;
  assign y12679 = n19329 ;
  assign y12680 = ~1'b0 ;
  assign y12681 = ~n19331 ;
  assign y12682 = ~n19333 ;
  assign y12683 = 1'b0 ;
  assign y12684 = ~n19335 ;
  assign y12685 = ~1'b0 ;
  assign y12686 = n19340 ;
  assign y12687 = ~n19343 ;
  assign y12688 = ~1'b0 ;
  assign y12689 = n19344 ;
  assign y12690 = 1'b0 ;
  assign y12691 = n19345 ;
  assign y12692 = ~1'b0 ;
  assign y12693 = ~n19347 ;
  assign y12694 = ~n19350 ;
  assign y12695 = ~n19354 ;
  assign y12696 = ~n19356 ;
  assign y12697 = n19357 ;
  assign y12698 = ~1'b0 ;
  assign y12699 = n19359 ;
  assign y12700 = ~1'b0 ;
  assign y12701 = ~1'b0 ;
  assign y12702 = ~n19363 ;
  assign y12703 = ~1'b0 ;
  assign y12704 = n19367 ;
  assign y12705 = ~1'b0 ;
  assign y12706 = ~1'b0 ;
  assign y12707 = ~n19369 ;
  assign y12708 = n19374 ;
  assign y12709 = n19380 ;
  assign y12710 = n19381 ;
  assign y12711 = ~1'b0 ;
  assign y12712 = ~n19384 ;
  assign y12713 = ~1'b0 ;
  assign y12714 = n19387 ;
  assign y12715 = ~n8982 ;
  assign y12716 = n19389 ;
  assign y12717 = ~1'b0 ;
  assign y12718 = ~1'b0 ;
  assign y12719 = ~n18098 ;
  assign y12720 = ~n19391 ;
  assign y12721 = ~n19392 ;
  assign y12722 = ~n19394 ;
  assign y12723 = ~n19395 ;
  assign y12724 = ~1'b0 ;
  assign y12725 = ~n19398 ;
  assign y12726 = ~1'b0 ;
  assign y12727 = ~1'b0 ;
  assign y12728 = ~1'b0 ;
  assign y12729 = ~n19402 ;
  assign y12730 = ~n19403 ;
  assign y12731 = ~n15456 ;
  assign y12732 = ~n19405 ;
  assign y12733 = n19406 ;
  assign y12734 = ~n19407 ;
  assign y12735 = ~n19409 ;
  assign y12736 = ~n12390 ;
  assign y12737 = ~1'b0 ;
  assign y12738 = n19410 ;
  assign y12739 = ~1'b0 ;
  assign y12740 = n19415 ;
  assign y12741 = 1'b0 ;
  assign y12742 = n19417 ;
  assign y12743 = n19418 ;
  assign y12744 = ~n19421 ;
  assign y12745 = ~n19422 ;
  assign y12746 = ~1'b0 ;
  assign y12747 = n19425 ;
  assign y12748 = ~1'b0 ;
  assign y12749 = n19427 ;
  assign y12750 = n12747 ;
  assign y12751 = ~n19428 ;
  assign y12752 = n19431 ;
  assign y12753 = ~1'b0 ;
  assign y12754 = ~1'b0 ;
  assign y12755 = ~1'b0 ;
  assign y12756 = ~n19434 ;
  assign y12757 = n19441 ;
  assign y12758 = n19442 ;
  assign y12759 = ~n10556 ;
  assign y12760 = ~n19445 ;
  assign y12761 = ~n19447 ;
  assign y12762 = ~1'b0 ;
  assign y12763 = ~1'b0 ;
  assign y12764 = ~1'b0 ;
  assign y12765 = ~n19451 ;
  assign y12766 = ~n19453 ;
  assign y12767 = ~n19455 ;
  assign y12768 = ~n19456 ;
  assign y12769 = ~n8888 ;
  assign y12770 = ~1'b0 ;
  assign y12771 = ~1'b0 ;
  assign y12772 = ~n2638 ;
  assign y12773 = ~1'b0 ;
  assign y12774 = ~n18866 ;
  assign y12775 = ~1'b0 ;
  assign y12776 = ~1'b0 ;
  assign y12777 = ~n586 ;
  assign y12778 = ~n2091 ;
  assign y12779 = ~1'b0 ;
  assign y12780 = ~1'b0 ;
  assign y12781 = ~n19457 ;
  assign y12782 = ~n19458 ;
  assign y12783 = n19460 ;
  assign y12784 = ~n19462 ;
  assign y12785 = ~1'b0 ;
  assign y12786 = ~n16996 ;
  assign y12787 = ~n19463 ;
  assign y12788 = n19464 ;
  assign y12789 = ~n19468 ;
  assign y12790 = n7206 ;
  assign y12791 = ~1'b0 ;
  assign y12792 = n19471 ;
  assign y12793 = ~1'b0 ;
  assign y12794 = ~n15581 ;
  assign y12795 = ~1'b0 ;
  assign y12796 = 1'b0 ;
  assign y12797 = n19472 ;
  assign y12798 = ~n19474 ;
  assign y12799 = n19475 ;
  assign y12800 = ~1'b0 ;
  assign y12801 = n19477 ;
  assign y12802 = n17794 ;
  assign y12803 = n240 ;
  assign y12804 = n19480 ;
  assign y12805 = 1'b0 ;
  assign y12806 = ~1'b0 ;
  assign y12807 = ~1'b0 ;
  assign y12808 = n19481 ;
  assign y12809 = ~1'b0 ;
  assign y12810 = ~n19482 ;
  assign y12811 = n19483 ;
  assign y12812 = n8232 ;
  assign y12813 = 1'b0 ;
  assign y12814 = ~n19484 ;
  assign y12815 = ~1'b0 ;
  assign y12816 = ~1'b0 ;
  assign y12817 = ~1'b0 ;
  assign y12818 = ~n19486 ;
  assign y12819 = ~n19488 ;
  assign y12820 = ~1'b0 ;
  assign y12821 = ~n19490 ;
  assign y12822 = ~n19492 ;
  assign y12823 = ~1'b0 ;
  assign y12824 = 1'b0 ;
  assign y12825 = n19495 ;
  assign y12826 = n19497 ;
  assign y12827 = ~1'b0 ;
  assign y12828 = ~n19499 ;
  assign y12829 = ~1'b0 ;
  assign y12830 = ~1'b0 ;
  assign y12831 = 1'b0 ;
  assign y12832 = ~1'b0 ;
  assign y12833 = ~1'b0 ;
  assign y12834 = ~1'b0 ;
  assign y12835 = ~n19505 ;
  assign y12836 = ~1'b0 ;
  assign y12837 = ~1'b0 ;
  assign y12838 = ~n15271 ;
  assign y12839 = n19510 ;
  assign y12840 = ~n19512 ;
  assign y12841 = ~1'b0 ;
  assign y12842 = n19517 ;
  assign y12843 = ~1'b0 ;
  assign y12844 = ~n19519 ;
  assign y12845 = ~n14807 ;
  assign y12846 = n19520 ;
  assign y12847 = 1'b0 ;
  assign y12848 = ~n3266 ;
  assign y12849 = ~1'b0 ;
  assign y12850 = 1'b0 ;
  assign y12851 = ~1'b0 ;
  assign y12852 = n19523 ;
  assign y12853 = n19524 ;
  assign y12854 = n19526 ;
  assign y12855 = ~1'b0 ;
  assign y12856 = n2396 ;
  assign y12857 = n19527 ;
  assign y12858 = ~n19529 ;
  assign y12859 = ~n19537 ;
  assign y12860 = ~n19538 ;
  assign y12861 = ~n19540 ;
  assign y12862 = ~n19542 ;
  assign y12863 = 1'b0 ;
  assign y12864 = n19548 ;
  assign y12865 = ~1'b0 ;
  assign y12866 = ~n19549 ;
  assign y12867 = n19551 ;
  assign y12868 = ~1'b0 ;
  assign y12869 = ~1'b0 ;
  assign y12870 = n19554 ;
  assign y12871 = ~1'b0 ;
  assign y12872 = ~n19556 ;
  assign y12873 = ~n19557 ;
  assign y12874 = ~1'b0 ;
  assign y12875 = n19558 ;
  assign y12876 = ~n19564 ;
  assign y12877 = ~1'b0 ;
  assign y12878 = 1'b0 ;
  assign y12879 = n19566 ;
  assign y12880 = n19569 ;
  assign y12881 = ~1'b0 ;
  assign y12882 = ~n19571 ;
  assign y12883 = 1'b0 ;
  assign y12884 = ~n645 ;
  assign y12885 = n19573 ;
  assign y12886 = ~n19578 ;
  assign y12887 = n6664 ;
  assign y12888 = ~n8406 ;
  assign y12889 = ~n19580 ;
  assign y12890 = ~1'b0 ;
  assign y12891 = ~1'b0 ;
  assign y12892 = ~1'b0 ;
  assign y12893 = ~1'b0 ;
  assign y12894 = ~n19583 ;
  assign y12895 = ~1'b0 ;
  assign y12896 = ~n19584 ;
  assign y12897 = ~1'b0 ;
  assign y12898 = 1'b0 ;
  assign y12899 = 1'b0 ;
  assign y12900 = ~1'b0 ;
  assign y12901 = n19587 ;
  assign y12902 = ~1'b0 ;
  assign y12903 = n19588 ;
  assign y12904 = ~1'b0 ;
  assign y12905 = ~1'b0 ;
  assign y12906 = n19590 ;
  assign y12907 = ~1'b0 ;
  assign y12908 = ~n19591 ;
  assign y12909 = ~1'b0 ;
  assign y12910 = n19594 ;
  assign y12911 = ~1'b0 ;
  assign y12912 = ~n19599 ;
  assign y12913 = ~1'b0 ;
  assign y12914 = n19600 ;
  assign y12915 = ~n19601 ;
  assign y12916 = n3012 ;
  assign y12917 = n19603 ;
  assign y12918 = 1'b0 ;
  assign y12919 = n19605 ;
  assign y12920 = ~n17533 ;
  assign y12921 = ~1'b0 ;
  assign y12922 = ~1'b0 ;
  assign y12923 = ~n15466 ;
  assign y12924 = ~n19606 ;
  assign y12925 = n19610 ;
  assign y12926 = ~1'b0 ;
  assign y12927 = n19611 ;
  assign y12928 = ~1'b0 ;
  assign y12929 = ~n12972 ;
  assign y12930 = ~1'b0 ;
  assign y12931 = ~1'b0 ;
  assign y12932 = ~n19613 ;
  assign y12933 = ~1'b0 ;
  assign y12934 = ~n19614 ;
  assign y12935 = ~1'b0 ;
  assign y12936 = ~1'b0 ;
  assign y12937 = ~n19618 ;
  assign y12938 = n19620 ;
  assign y12939 = ~n19622 ;
  assign y12940 = n19626 ;
  assign y12941 = ~n19627 ;
  assign y12942 = ~n19629 ;
  assign y12943 = n19631 ;
  assign y12944 = ~1'b0 ;
  assign y12945 = n19633 ;
  assign y12946 = n19635 ;
  assign y12947 = ~1'b0 ;
  assign y12948 = n19636 ;
  assign y12949 = n19638 ;
  assign y12950 = n1369 ;
  assign y12951 = ~n19640 ;
  assign y12952 = n6344 ;
  assign y12953 = n8390 ;
  assign y12954 = n19642 ;
  assign y12955 = n19643 ;
  assign y12956 = ~1'b0 ;
  assign y12957 = ~1'b0 ;
  assign y12958 = ~1'b0 ;
  assign y12959 = ~1'b0 ;
  assign y12960 = ~1'b0 ;
  assign y12961 = ~n19645 ;
  assign y12962 = ~n19647 ;
  assign y12963 = n19649 ;
  assign y12964 = ~n11423 ;
  assign y12965 = n19652 ;
  assign y12966 = n19653 ;
  assign y12967 = ~n19654 ;
  assign y12968 = ~n19656 ;
  assign y12969 = ~1'b0 ;
  assign y12970 = ~1'b0 ;
  assign y12971 = ~n19661 ;
  assign y12972 = ~n19662 ;
  assign y12973 = n19668 ;
  assign y12974 = ~1'b0 ;
  assign y12975 = ~1'b0 ;
  assign y12976 = ~n19670 ;
  assign y12977 = ~1'b0 ;
  assign y12978 = ~n19671 ;
  assign y12979 = ~1'b0 ;
  assign y12980 = ~n3934 ;
  assign y12981 = ~n19674 ;
  assign y12982 = n19676 ;
  assign y12983 = n19679 ;
  assign y12984 = ~1'b0 ;
  assign y12985 = ~1'b0 ;
  assign y12986 = ~1'b0 ;
  assign y12987 = ~1'b0 ;
  assign y12988 = n19680 ;
  assign y12989 = ~1'b0 ;
  assign y12990 = n19681 ;
  assign y12991 = ~n19684 ;
  assign y12992 = n19688 ;
  assign y12993 = n19690 ;
  assign y12994 = n19691 ;
  assign y12995 = ~1'b0 ;
  assign y12996 = ~1'b0 ;
  assign y12997 = ~1'b0 ;
  assign y12998 = ~1'b0 ;
  assign y12999 = ~1'b0 ;
  assign y13000 = ~n19692 ;
  assign y13001 = ~1'b0 ;
  assign y13002 = 1'b0 ;
  assign y13003 = ~1'b0 ;
  assign y13004 = ~1'b0 ;
  assign y13005 = ~1'b0 ;
  assign y13006 = ~1'b0 ;
  assign y13007 = n19693 ;
  assign y13008 = ~n19695 ;
  assign y13009 = ~1'b0 ;
  assign y13010 = n19696 ;
  assign y13011 = n19698 ;
  assign y13012 = ~1'b0 ;
  assign y13013 = ~n19702 ;
  assign y13014 = n19705 ;
  assign y13015 = ~1'b0 ;
  assign y13016 = 1'b0 ;
  assign y13017 = n19706 ;
  assign y13018 = ~n6821 ;
  assign y13019 = n19707 ;
  assign y13020 = ~1'b0 ;
  assign y13021 = ~n19709 ;
  assign y13022 = ~n19711 ;
  assign y13023 = ~n15244 ;
  assign y13024 = n19712 ;
  assign y13025 = ~1'b0 ;
  assign y13026 = n5374 ;
  assign y13027 = ~n19719 ;
  assign y13028 = n19723 ;
  assign y13029 = ~1'b0 ;
  assign y13030 = ~n19724 ;
  assign y13031 = ~1'b0 ;
  assign y13032 = n19725 ;
  assign y13033 = ~1'b0 ;
  assign y13034 = ~n19732 ;
  assign y13035 = ~n19734 ;
  assign y13036 = ~1'b0 ;
  assign y13037 = ~1'b0 ;
  assign y13038 = ~n19735 ;
  assign y13039 = ~1'b0 ;
  assign y13040 = ~n19736 ;
  assign y13041 = n14198 ;
  assign y13042 = ~1'b0 ;
  assign y13043 = ~1'b0 ;
  assign y13044 = n19740 ;
  assign y13045 = n19741 ;
  assign y13046 = ~n19742 ;
  assign y13047 = ~1'b0 ;
  assign y13048 = n19743 ;
  assign y13049 = ~1'b0 ;
  assign y13050 = ~n19745 ;
  assign y13051 = ~n19746 ;
  assign y13052 = ~1'b0 ;
  assign y13053 = n19749 ;
  assign y13054 = ~1'b0 ;
  assign y13055 = ~n19751 ;
  assign y13056 = ~1'b0 ;
  assign y13057 = ~1'b0 ;
  assign y13058 = ~n19752 ;
  assign y13059 = ~n19753 ;
  assign y13060 = ~1'b0 ;
  assign y13061 = ~1'b0 ;
  assign y13062 = ~1'b0 ;
  assign y13063 = 1'b0 ;
  assign y13064 = ~1'b0 ;
  assign y13065 = ~1'b0 ;
  assign y13066 = ~n19756 ;
  assign y13067 = ~1'b0 ;
  assign y13068 = n5208 ;
  assign y13069 = ~1'b0 ;
  assign y13070 = ~n19758 ;
  assign y13071 = ~1'b0 ;
  assign y13072 = n19759 ;
  assign y13073 = n19762 ;
  assign y13074 = ~n19764 ;
  assign y13075 = ~n6917 ;
  assign y13076 = ~n19765 ;
  assign y13077 = n19768 ;
  assign y13078 = ~1'b0 ;
  assign y13079 = ~n19770 ;
  assign y13080 = n19771 ;
  assign y13081 = n19774 ;
  assign y13082 = n10476 ;
  assign y13083 = ~1'b0 ;
  assign y13084 = ~1'b0 ;
  assign y13085 = n19778 ;
  assign y13086 = 1'b0 ;
  assign y13087 = ~n19779 ;
  assign y13088 = n19780 ;
  assign y13089 = ~n19781 ;
  assign y13090 = ~n19783 ;
  assign y13091 = ~n19784 ;
  assign y13092 = ~n19786 ;
  assign y13093 = ~n19788 ;
  assign y13094 = ~1'b0 ;
  assign y13095 = n19794 ;
  assign y13096 = n17846 ;
  assign y13097 = n19797 ;
  assign y13098 = n9459 ;
  assign y13099 = n19800 ;
  assign y13100 = ~1'b0 ;
  assign y13101 = ~1'b0 ;
  assign y13102 = ~n19803 ;
  assign y13103 = ~1'b0 ;
  assign y13104 = ~n19807 ;
  assign y13105 = ~1'b0 ;
  assign y13106 = n19808 ;
  assign y13107 = n19809 ;
  assign y13108 = ~n19810 ;
  assign y13109 = ~1'b0 ;
  assign y13110 = 1'b0 ;
  assign y13111 = ~n19814 ;
  assign y13112 = n19815 ;
  assign y13113 = n19818 ;
  assign y13114 = ~n19819 ;
  assign y13115 = ~n2862 ;
  assign y13116 = n19820 ;
  assign y13117 = n19821 ;
  assign y13118 = ~1'b0 ;
  assign y13119 = ~n19822 ;
  assign y13120 = n19824 ;
  assign y13121 = ~1'b0 ;
  assign y13122 = n19826 ;
  assign y13123 = ~n19828 ;
  assign y13124 = n19833 ;
  assign y13125 = ~1'b0 ;
  assign y13126 = ~n19834 ;
  assign y13127 = ~n19835 ;
  assign y13128 = n2831 ;
  assign y13129 = ~n19841 ;
  assign y13130 = ~1'b0 ;
  assign y13131 = ~1'b0 ;
  assign y13132 = ~n19846 ;
  assign y13133 = ~n19849 ;
  assign y13134 = n19854 ;
  assign y13135 = ~1'b0 ;
  assign y13136 = ~1'b0 ;
  assign y13137 = ~n19855 ;
  assign y13138 = ~1'b0 ;
  assign y13139 = ~1'b0 ;
  assign y13140 = 1'b0 ;
  assign y13141 = n19856 ;
  assign y13142 = n19858 ;
  assign y13143 = ~n19861 ;
  assign y13144 = n19863 ;
  assign y13145 = ~n19865 ;
  assign y13146 = n19868 ;
  assign y13147 = n19870 ;
  assign y13148 = ~n19873 ;
  assign y13149 = ~1'b0 ;
  assign y13150 = ~n19875 ;
  assign y13151 = 1'b0 ;
  assign y13152 = ~n13866 ;
  assign y13153 = n19877 ;
  assign y13154 = n19879 ;
  assign y13155 = ~1'b0 ;
  assign y13156 = n19885 ;
  assign y13157 = n19886 ;
  assign y13158 = n19889 ;
  assign y13159 = ~1'b0 ;
  assign y13160 = n1228 ;
  assign y13161 = ~1'b0 ;
  assign y13162 = n19891 ;
  assign y13163 = 1'b0 ;
  assign y13164 = ~1'b0 ;
  assign y13165 = ~n19894 ;
  assign y13166 = ~n19895 ;
  assign y13167 = ~x48 ;
  assign y13168 = ~1'b0 ;
  assign y13169 = ~n19898 ;
  assign y13170 = n19899 ;
  assign y13171 = n19900 ;
  assign y13172 = ~n19903 ;
  assign y13173 = n19904 ;
  assign y13174 = ~n2951 ;
  assign y13175 = ~n19906 ;
  assign y13176 = ~1'b0 ;
  assign y13177 = ~1'b0 ;
  assign y13178 = ~n19909 ;
  assign y13179 = ~1'b0 ;
  assign y13180 = n19915 ;
  assign y13181 = n16091 ;
  assign y13182 = n19916 ;
  assign y13183 = n5582 ;
  assign y13184 = ~1'b0 ;
  assign y13185 = ~n19917 ;
  assign y13186 = ~1'b0 ;
  assign y13187 = ~n19918 ;
  assign y13188 = ~1'b0 ;
  assign y13189 = n19919 ;
  assign y13190 = n4906 ;
  assign y13191 = ~n19920 ;
  assign y13192 = n19922 ;
  assign y13193 = ~n19923 ;
  assign y13194 = n19926 ;
  assign y13195 = n19928 ;
  assign y13196 = n3855 ;
  assign y13197 = ~n19930 ;
  assign y13198 = ~1'b0 ;
  assign y13199 = ~n11634 ;
  assign y13200 = ~n19931 ;
  assign y13201 = ~1'b0 ;
  assign y13202 = ~n19935 ;
  assign y13203 = ~1'b0 ;
  assign y13204 = n19938 ;
  assign y13205 = ~n19939 ;
  assign y13206 = n19942 ;
  assign y13207 = ~1'b0 ;
  assign y13208 = ~n19943 ;
  assign y13209 = ~1'b0 ;
  assign y13210 = ~n19945 ;
  assign y13211 = ~1'b0 ;
  assign y13212 = 1'b0 ;
  assign y13213 = ~n19948 ;
  assign y13214 = ~1'b0 ;
  assign y13215 = ~n19949 ;
  assign y13216 = ~n19955 ;
  assign y13217 = n4206 ;
  assign y13218 = ~n19959 ;
  assign y13219 = n19962 ;
  assign y13220 = n19964 ;
  assign y13221 = n16144 ;
  assign y13222 = ~n19966 ;
  assign y13223 = ~1'b0 ;
  assign y13224 = n19968 ;
  assign y13225 = n19970 ;
  assign y13226 = ~1'b0 ;
  assign y13227 = ~n19974 ;
  assign y13228 = n19975 ;
  assign y13229 = ~n19977 ;
  assign y13230 = ~n19983 ;
  assign y13231 = ~n19985 ;
  assign y13232 = ~n19986 ;
  assign y13233 = ~1'b0 ;
  assign y13234 = n19989 ;
  assign y13235 = n19990 ;
  assign y13236 = ~n19992 ;
  assign y13237 = ~n6205 ;
  assign y13238 = n19993 ;
  assign y13239 = ~1'b0 ;
  assign y13240 = ~n19995 ;
  assign y13241 = n19997 ;
  assign y13242 = ~1'b0 ;
  assign y13243 = n20000 ;
  assign y13244 = n20002 ;
  assign y13245 = n20004 ;
  assign y13246 = n20005 ;
  assign y13247 = ~1'b0 ;
  assign y13248 = ~n20007 ;
  assign y13249 = ~n20009 ;
  assign y13250 = n20010 ;
  assign y13251 = ~n20015 ;
  assign y13252 = n20016 ;
  assign y13253 = ~1'b0 ;
  assign y13254 = ~n20019 ;
  assign y13255 = ~1'b0 ;
  assign y13256 = n4941 ;
  assign y13257 = ~n20024 ;
  assign y13258 = ~1'b0 ;
  assign y13259 = ~1'b0 ;
  assign y13260 = n20025 ;
  assign y13261 = n20027 ;
  assign y13262 = ~n20029 ;
  assign y13263 = 1'b0 ;
  assign y13264 = n20030 ;
  assign y13265 = n20033 ;
  assign y13266 = n20034 ;
  assign y13267 = ~1'b0 ;
  assign y13268 = n20035 ;
  assign y13269 = n20037 ;
  assign y13270 = n20039 ;
  assign y13271 = ~n20040 ;
  assign y13272 = ~1'b0 ;
  assign y13273 = n20042 ;
  assign y13274 = n20045 ;
  assign y13275 = ~1'b0 ;
  assign y13276 = ~n2089 ;
  assign y13277 = ~1'b0 ;
  assign y13278 = ~1'b0 ;
  assign y13279 = ~1'b0 ;
  assign y13280 = ~1'b0 ;
  assign y13281 = n20048 ;
  assign y13282 = n20050 ;
  assign y13283 = n20051 ;
  assign y13284 = ~n20053 ;
  assign y13285 = ~n20057 ;
  assign y13286 = ~1'b0 ;
  assign y13287 = ~n20062 ;
  assign y13288 = ~1'b0 ;
  assign y13289 = n19131 ;
  assign y13290 = ~1'b0 ;
  assign y13291 = n20063 ;
  assign y13292 = ~n20064 ;
  assign y13293 = n20066 ;
  assign y13294 = ~1'b0 ;
  assign y13295 = ~n20068 ;
  assign y13296 = n20071 ;
  assign y13297 = ~n20076 ;
  assign y13298 = n13226 ;
  assign y13299 = n20078 ;
  assign y13300 = ~n20079 ;
  assign y13301 = ~n5475 ;
  assign y13302 = n9271 ;
  assign y13303 = ~n8269 ;
  assign y13304 = ~n20081 ;
  assign y13305 = ~n20085 ;
  assign y13306 = ~1'b0 ;
  assign y13307 = ~n20088 ;
  assign y13308 = n20090 ;
  assign y13309 = n6322 ;
  assign y13310 = n20094 ;
  assign y13311 = n20095 ;
  assign y13312 = 1'b0 ;
  assign y13313 = ~n20096 ;
  assign y13314 = n20097 ;
  assign y13315 = ~1'b0 ;
  assign y13316 = ~n20098 ;
  assign y13317 = n20099 ;
  assign y13318 = ~n7634 ;
  assign y13319 = ~1'b0 ;
  assign y13320 = ~1'b0 ;
  assign y13321 = n20103 ;
  assign y13322 = ~n20104 ;
  assign y13323 = n20106 ;
  assign y13324 = ~n20107 ;
  assign y13325 = n20109 ;
  assign y13326 = n20110 ;
  assign y13327 = n20117 ;
  assign y13328 = ~1'b0 ;
  assign y13329 = n20118 ;
  assign y13330 = n20120 ;
  assign y13331 = ~1'b0 ;
  assign y13332 = ~n20123 ;
  assign y13333 = ~n20124 ;
  assign y13334 = n20125 ;
  assign y13335 = n20126 ;
  assign y13336 = ~n13330 ;
  assign y13337 = ~1'b0 ;
  assign y13338 = n18111 ;
  assign y13339 = ~1'b0 ;
  assign y13340 = ~n20132 ;
  assign y13341 = ~n20134 ;
  assign y13342 = n20142 ;
  assign y13343 = ~1'b0 ;
  assign y13344 = ~1'b0 ;
  assign y13345 = ~1'b0 ;
  assign y13346 = n20143 ;
  assign y13347 = 1'b0 ;
  assign y13348 = ~1'b0 ;
  assign y13349 = ~1'b0 ;
  assign y13350 = ~n20144 ;
  assign y13351 = n20145 ;
  assign y13352 = ~n20148 ;
  assign y13353 = n12091 ;
  assign y13354 = ~n20152 ;
  assign y13355 = n9931 ;
  assign y13356 = n828 ;
  assign y13357 = ~1'b0 ;
  assign y13358 = ~n20155 ;
  assign y13359 = ~n19112 ;
  assign y13360 = ~1'b0 ;
  assign y13361 = ~1'b0 ;
  assign y13362 = ~1'b0 ;
  assign y13363 = ~n4314 ;
  assign y13364 = ~n20159 ;
  assign y13365 = n20160 ;
  assign y13366 = ~1'b0 ;
  assign y13367 = n20161 ;
  assign y13368 = ~n20169 ;
  assign y13369 = ~n20170 ;
  assign y13370 = ~1'b0 ;
  assign y13371 = ~1'b0 ;
  assign y13372 = n20172 ;
  assign y13373 = ~n20173 ;
  assign y13374 = ~1'b0 ;
  assign y13375 = n20175 ;
  assign y13376 = n20177 ;
  assign y13377 = ~1'b0 ;
  assign y13378 = n20178 ;
  assign y13379 = ~1'b0 ;
  assign y13380 = n3987 ;
  assign y13381 = n20180 ;
  assign y13382 = ~1'b0 ;
  assign y13383 = n20182 ;
  assign y13384 = ~n19311 ;
  assign y13385 = ~n20183 ;
  assign y13386 = n20184 ;
  assign y13387 = ~n20187 ;
  assign y13388 = n20192 ;
  assign y13389 = ~1'b0 ;
  assign y13390 = ~1'b0 ;
  assign y13391 = ~1'b0 ;
  assign y13392 = n20194 ;
  assign y13393 = ~1'b0 ;
  assign y13394 = ~1'b0 ;
  assign y13395 = n20196 ;
  assign y13396 = ~1'b0 ;
  assign y13397 = ~1'b0 ;
  assign y13398 = 1'b0 ;
  assign y13399 = ~1'b0 ;
  assign y13400 = 1'b0 ;
  assign y13401 = n20197 ;
  assign y13402 = ~1'b0 ;
  assign y13403 = ~n2804 ;
  assign y13404 = ~n3651 ;
  assign y13405 = n745 ;
  assign y13406 = n20198 ;
  assign y13407 = ~n20199 ;
  assign y13408 = n20202 ;
  assign y13409 = ~n20203 ;
  assign y13410 = n20204 ;
  assign y13411 = n20206 ;
  assign y13412 = 1'b0 ;
  assign y13413 = n20207 ;
  assign y13414 = ~n20208 ;
  assign y13415 = ~n20209 ;
  assign y13416 = ~n20210 ;
  assign y13417 = n4974 ;
  assign y13418 = n8673 ;
  assign y13419 = 1'b0 ;
  assign y13420 = ~n20211 ;
  assign y13421 = n20212 ;
  assign y13422 = ~n20217 ;
  assign y13423 = ~n20218 ;
  assign y13424 = ~x59 ;
  assign y13425 = ~n20219 ;
  assign y13426 = n20221 ;
  assign y13427 = ~n20222 ;
  assign y13428 = ~n20226 ;
  assign y13429 = ~n20227 ;
  assign y13430 = 1'b0 ;
  assign y13431 = n20229 ;
  assign y13432 = n20230 ;
  assign y13433 = n20235 ;
  assign y13434 = ~1'b0 ;
  assign y13435 = n20237 ;
  assign y13436 = ~1'b0 ;
  assign y13437 = ~n20240 ;
  assign y13438 = ~1'b0 ;
  assign y13439 = ~n20243 ;
  assign y13440 = ~1'b0 ;
  assign y13441 = ~n20245 ;
  assign y13442 = n20247 ;
  assign y13443 = ~1'b0 ;
  assign y13444 = ~n20251 ;
  assign y13445 = 1'b0 ;
  assign y13446 = n20253 ;
  assign y13447 = ~1'b0 ;
  assign y13448 = ~1'b0 ;
  assign y13449 = ~1'b0 ;
  assign y13450 = n20254 ;
  assign y13451 = n20255 ;
  assign y13452 = ~1'b0 ;
  assign y13453 = n20258 ;
  assign y13454 = ~1'b0 ;
  assign y13455 = n20259 ;
  assign y13456 = ~n7814 ;
  assign y13457 = n20263 ;
  assign y13458 = ~1'b0 ;
  assign y13459 = n20268 ;
  assign y13460 = ~1'b0 ;
  assign y13461 = n20273 ;
  assign y13462 = n20274 ;
  assign y13463 = n20276 ;
  assign y13464 = ~1'b0 ;
  assign y13465 = ~1'b0 ;
  assign y13466 = ~1'b0 ;
  assign y13467 = n20278 ;
  assign y13468 = ~n20279 ;
  assign y13469 = n20280 ;
  assign y13470 = ~n20281 ;
  assign y13471 = n20284 ;
  assign y13472 = ~n20288 ;
  assign y13473 = n20290 ;
  assign y13474 = ~n20293 ;
  assign y13475 = ~n20294 ;
  assign y13476 = n20295 ;
  assign y13477 = ~n20299 ;
  assign y13478 = n20301 ;
  assign y13479 = ~n20302 ;
  assign y13480 = n20307 ;
  assign y13481 = ~n20308 ;
  assign y13482 = n20309 ;
  assign y13483 = ~n20311 ;
  assign y13484 = ~n20313 ;
  assign y13485 = ~n20315 ;
  assign y13486 = ~n20317 ;
  assign y13487 = ~1'b0 ;
  assign y13488 = ~n1623 ;
  assign y13489 = ~1'b0 ;
  assign y13490 = n20318 ;
  assign y13491 = ~n20320 ;
  assign y13492 = ~1'b0 ;
  assign y13493 = ~n2091 ;
  assign y13494 = n20324 ;
  assign y13495 = n20325 ;
  assign y13496 = n20330 ;
  assign y13497 = ~n20335 ;
  assign y13498 = n20336 ;
  assign y13499 = n20338 ;
  assign y13500 = ~n20340 ;
  assign y13501 = n20342 ;
  assign y13502 = ~n20344 ;
  assign y13503 = ~1'b0 ;
  assign y13504 = ~1'b0 ;
  assign y13505 = ~1'b0 ;
  assign y13506 = ~n20346 ;
  assign y13507 = n8292 ;
  assign y13508 = ~n20349 ;
  assign y13509 = ~n20353 ;
  assign y13510 = ~n8067 ;
  assign y13511 = ~n5309 ;
  assign y13512 = ~1'b0 ;
  assign y13513 = ~n20354 ;
  assign y13514 = ~1'b0 ;
  assign y13515 = n20355 ;
  assign y13516 = ~n20356 ;
  assign y13517 = ~1'b0 ;
  assign y13518 = n20359 ;
  assign y13519 = n20364 ;
  assign y13520 = n20367 ;
  assign y13521 = 1'b0 ;
  assign y13522 = ~1'b0 ;
  assign y13523 = 1'b0 ;
  assign y13524 = ~1'b0 ;
  assign y13525 = n20370 ;
  assign y13526 = n9089 ;
  assign y13527 = ~n1999 ;
  assign y13528 = ~n20372 ;
  assign y13529 = n20376 ;
  assign y13530 = ~1'b0 ;
  assign y13531 = n20378 ;
  assign y13532 = ~n20380 ;
  assign y13533 = ~1'b0 ;
  assign y13534 = ~n20382 ;
  assign y13535 = n20384 ;
  assign y13536 = ~1'b0 ;
  assign y13537 = ~1'b0 ;
  assign y13538 = ~1'b0 ;
  assign y13539 = n20385 ;
  assign y13540 = ~1'b0 ;
  assign y13541 = n9625 ;
  assign y13542 = n20389 ;
  assign y13543 = n20390 ;
  assign y13544 = n20414 ;
  assign y13545 = ~1'b0 ;
  assign y13546 = ~1'b0 ;
  assign y13547 = n20417 ;
  assign y13548 = ~1'b0 ;
  assign y13549 = ~1'b0 ;
  assign y13550 = ~n20418 ;
  assign y13551 = ~n20419 ;
  assign y13552 = ~1'b0 ;
  assign y13553 = ~n20424 ;
  assign y13554 = ~1'b0 ;
  assign y13555 = ~n20429 ;
  assign y13556 = ~1'b0 ;
  assign y13557 = ~1'b0 ;
  assign y13558 = ~n20431 ;
  assign y13559 = n20432 ;
  assign y13560 = ~1'b0 ;
  assign y13561 = ~1'b0 ;
  assign y13562 = n20435 ;
  assign y13563 = n20437 ;
  assign y13564 = ~1'b0 ;
  assign y13565 = n20439 ;
  assign y13566 = ~n20443 ;
  assign y13567 = n20446 ;
  assign y13568 = n20449 ;
  assign y13569 = n20450 ;
  assign y13570 = ~n20451 ;
  assign y13571 = ~1'b0 ;
  assign y13572 = ~1'b0 ;
  assign y13573 = ~n20452 ;
  assign y13574 = n20456 ;
  assign y13575 = ~n20458 ;
  assign y13576 = ~1'b0 ;
  assign y13577 = ~1'b0 ;
  assign y13578 = ~1'b0 ;
  assign y13579 = ~n20460 ;
  assign y13580 = n20462 ;
  assign y13581 = n20463 ;
  assign y13582 = ~1'b0 ;
  assign y13583 = n20468 ;
  assign y13584 = ~n20472 ;
  assign y13585 = n20474 ;
  assign y13586 = n20475 ;
  assign y13587 = n10619 ;
  assign y13588 = ~1'b0 ;
  assign y13589 = ~n20477 ;
  assign y13590 = ~1'b0 ;
  assign y13591 = n20480 ;
  assign y13592 = n20482 ;
  assign y13593 = ~n20484 ;
  assign y13594 = ~1'b0 ;
  assign y13595 = ~1'b0 ;
  assign y13596 = ~n20488 ;
  assign y13597 = ~n20490 ;
  assign y13598 = ~1'b0 ;
  assign y13599 = ~n20492 ;
  assign y13600 = ~1'b0 ;
  assign y13601 = ~n20493 ;
  assign y13602 = n20495 ;
  assign y13603 = ~1'b0 ;
  assign y13604 = n20499 ;
  assign y13605 = ~1'b0 ;
  assign y13606 = n20500 ;
  assign y13607 = ~1'b0 ;
  assign y13608 = n20501 ;
  assign y13609 = n20503 ;
  assign y13610 = ~1'b0 ;
  assign y13611 = ~n6226 ;
  assign y13612 = 1'b0 ;
  assign y13613 = n20504 ;
  assign y13614 = n20507 ;
  assign y13615 = n20509 ;
  assign y13616 = ~1'b0 ;
  assign y13617 = ~n17097 ;
  assign y13618 = ~1'b0 ;
  assign y13619 = ~1'b0 ;
  assign y13620 = n20512 ;
  assign y13621 = ~1'b0 ;
  assign y13622 = n20514 ;
  assign y13623 = ~1'b0 ;
  assign y13624 = n20515 ;
  assign y13625 = n20517 ;
  assign y13626 = ~1'b0 ;
  assign y13627 = ~1'b0 ;
  assign y13628 = n6835 ;
  assign y13629 = ~n20519 ;
  assign y13630 = n20520 ;
  assign y13631 = ~1'b0 ;
  assign y13632 = n20522 ;
  assign y13633 = ~n904 ;
  assign y13634 = ~n4800 ;
  assign y13635 = ~n20523 ;
  assign y13636 = ~1'b0 ;
  assign y13637 = ~n4033 ;
  assign y13638 = 1'b0 ;
  assign y13639 = n20525 ;
  assign y13640 = 1'b0 ;
  assign y13641 = n20532 ;
  assign y13642 = n20534 ;
  assign y13643 = ~1'b0 ;
  assign y13644 = n20535 ;
  assign y13645 = ~n20536 ;
  assign y13646 = ~n20542 ;
  assign y13647 = ~n20544 ;
  assign y13648 = ~n20546 ;
  assign y13649 = 1'b0 ;
  assign y13650 = n20548 ;
  assign y13651 = ~1'b0 ;
  assign y13652 = n12378 ;
  assign y13653 = ~n20551 ;
  assign y13654 = ~n20552 ;
  assign y13655 = ~n20553 ;
  assign y13656 = n20554 ;
  assign y13657 = ~1'b0 ;
  assign y13658 = ~1'b0 ;
  assign y13659 = n20558 ;
  assign y13660 = ~n5708 ;
  assign y13661 = ~n20563 ;
  assign y13662 = ~1'b0 ;
  assign y13663 = ~1'b0 ;
  assign y13664 = n20566 ;
  assign y13665 = ~n20567 ;
  assign y13666 = ~n1536 ;
  assign y13667 = ~n20569 ;
  assign y13668 = 1'b0 ;
  assign y13669 = ~n20573 ;
  assign y13670 = ~n20575 ;
  assign y13671 = ~n20578 ;
  assign y13672 = ~1'b0 ;
  assign y13673 = ~n20580 ;
  assign y13674 = n20582 ;
  assign y13675 = ~n20583 ;
  assign y13676 = ~n13930 ;
  assign y13677 = n20584 ;
  assign y13678 = n20586 ;
  assign y13679 = n20592 ;
  assign y13680 = ~n20596 ;
  assign y13681 = ~1'b0 ;
  assign y13682 = ~1'b0 ;
  assign y13683 = ~n20598 ;
  assign y13684 = ~1'b0 ;
  assign y13685 = ~1'b0 ;
  assign y13686 = n20599 ;
  assign y13687 = ~n20602 ;
  assign y13688 = 1'b0 ;
  assign y13689 = ~1'b0 ;
  assign y13690 = ~n20603 ;
  assign y13691 = ~n20604 ;
  assign y13692 = n1162 ;
  assign y13693 = ~1'b0 ;
  assign y13694 = ~n20608 ;
  assign y13695 = n20609 ;
  assign y13696 = ~n20610 ;
  assign y13697 = ~n20611 ;
  assign y13698 = ~n20616 ;
  assign y13699 = ~1'b0 ;
  assign y13700 = n20618 ;
  assign y13701 = ~n20620 ;
  assign y13702 = n20624 ;
  assign y13703 = ~1'b0 ;
  assign y13704 = ~1'b0 ;
  assign y13705 = ~1'b0 ;
  assign y13706 = ~1'b0 ;
  assign y13707 = ~1'b0 ;
  assign y13708 = 1'b0 ;
  assign y13709 = ~n20628 ;
  assign y13710 = ~1'b0 ;
  assign y13711 = n20629 ;
  assign y13712 = n20630 ;
  assign y13713 = ~n20635 ;
  assign y13714 = ~1'b0 ;
  assign y13715 = ~1'b0 ;
  assign y13716 = ~n20637 ;
  assign y13717 = ~1'b0 ;
  assign y13718 = ~1'b0 ;
  assign y13719 = n20641 ;
  assign y13720 = ~n20643 ;
  assign y13721 = ~n20645 ;
  assign y13722 = ~1'b0 ;
  assign y13723 = n20647 ;
  assign y13724 = ~n20650 ;
  assign y13725 = n3998 ;
  assign y13726 = n20652 ;
  assign y13727 = ~1'b0 ;
  assign y13728 = n20654 ;
  assign y13729 = ~1'b0 ;
  assign y13730 = ~n20655 ;
  assign y13731 = ~n2722 ;
  assign y13732 = ~n20660 ;
  assign y13733 = n20664 ;
  assign y13734 = n2733 ;
  assign y13735 = 1'b0 ;
  assign y13736 = ~1'b0 ;
  assign y13737 = ~n20665 ;
  assign y13738 = 1'b0 ;
  assign y13739 = ~1'b0 ;
  assign y13740 = ~1'b0 ;
  assign y13741 = ~n11927 ;
  assign y13742 = n20667 ;
  assign y13743 = n20668 ;
  assign y13744 = ~1'b0 ;
  assign y13745 = ~n20669 ;
  assign y13746 = n20672 ;
  assign y13747 = n20673 ;
  assign y13748 = n20674 ;
  assign y13749 = ~n20675 ;
  assign y13750 = ~1'b0 ;
  assign y13751 = ~1'b0 ;
  assign y13752 = ~1'b0 ;
  assign y13753 = ~1'b0 ;
  assign y13754 = ~1'b0 ;
  assign y13755 = ~n20677 ;
  assign y13756 = ~n20681 ;
  assign y13757 = n1277 ;
  assign y13758 = ~1'b0 ;
  assign y13759 = n20682 ;
  assign y13760 = ~n20683 ;
  assign y13761 = n20685 ;
  assign y13762 = n20690 ;
  assign y13763 = ~n20693 ;
  assign y13764 = ~n20696 ;
  assign y13765 = n20700 ;
  assign y13766 = n17534 ;
  assign y13767 = ~1'b0 ;
  assign y13768 = 1'b0 ;
  assign y13769 = ~n20701 ;
  assign y13770 = ~1'b0 ;
  assign y13771 = ~n20705 ;
  assign y13772 = ~1'b0 ;
  assign y13773 = n20706 ;
  assign y13774 = ~1'b0 ;
  assign y13775 = ~n20707 ;
  assign y13776 = ~1'b0 ;
  assign y13777 = n20713 ;
  assign y13778 = ~n20714 ;
  assign y13779 = ~1'b0 ;
  assign y13780 = ~1'b0 ;
  assign y13781 = ~n20716 ;
  assign y13782 = ~n20717 ;
  assign y13783 = ~1'b0 ;
  assign y13784 = ~n20719 ;
  assign y13785 = n18325 ;
  assign y13786 = ~1'b0 ;
  assign y13787 = ~n20721 ;
  assign y13788 = ~1'b0 ;
  assign y13789 = ~n20724 ;
  assign y13790 = n20725 ;
  assign y13791 = ~1'b0 ;
  assign y13792 = n20728 ;
  assign y13793 = ~n20729 ;
  assign y13794 = n20733 ;
  assign y13795 = ~1'b0 ;
  assign y13796 = n20734 ;
  assign y13797 = ~1'b0 ;
  assign y13798 = n1069 ;
  assign y13799 = ~1'b0 ;
  assign y13800 = n20737 ;
  assign y13801 = n20742 ;
  assign y13802 = n15478 ;
  assign y13803 = ~n20743 ;
  assign y13804 = n20746 ;
  assign y13805 = n20747 ;
  assign y13806 = ~1'b0 ;
  assign y13807 = n20748 ;
  assign y13808 = ~n20750 ;
  assign y13809 = n20752 ;
  assign y13810 = ~1'b0 ;
  assign y13811 = ~n20753 ;
  assign y13812 = n20756 ;
  assign y13813 = ~1'b0 ;
  assign y13814 = n20758 ;
  assign y13815 = n12482 ;
  assign y13816 = ~1'b0 ;
  assign y13817 = n20759 ;
  assign y13818 = ~n20760 ;
  assign y13819 = ~1'b0 ;
  assign y13820 = ~n20763 ;
  assign y13821 = ~1'b0 ;
  assign y13822 = ~n20765 ;
  assign y13823 = ~n20766 ;
  assign y13824 = n20767 ;
  assign y13825 = 1'b0 ;
  assign y13826 = ~n20768 ;
  assign y13827 = ~n20770 ;
  assign y13828 = n20772 ;
  assign y13829 = n20773 ;
  assign y13830 = n20775 ;
  assign y13831 = ~n20776 ;
  assign y13832 = ~1'b0 ;
  assign y13833 = ~n20779 ;
  assign y13834 = ~n20782 ;
  assign y13835 = n20783 ;
  assign y13836 = ~1'b0 ;
  assign y13837 = n20785 ;
  assign y13838 = n20788 ;
  assign y13839 = n20789 ;
  assign y13840 = n20791 ;
  assign y13841 = ~1'b0 ;
  assign y13842 = ~n20792 ;
  assign y13843 = n20794 ;
  assign y13844 = ~1'b0 ;
  assign y13845 = n11659 ;
  assign y13846 = ~1'b0 ;
  assign y13847 = ~n20795 ;
  assign y13848 = ~1'b0 ;
  assign y13849 = ~n2227 ;
  assign y13850 = ~1'b0 ;
  assign y13851 = ~1'b0 ;
  assign y13852 = ~n20797 ;
  assign y13853 = n20800 ;
  assign y13854 = ~1'b0 ;
  assign y13855 = n20803 ;
  assign y13856 = n20804 ;
  assign y13857 = ~n4859 ;
  assign y13858 = ~n20808 ;
  assign y13859 = ~1'b0 ;
  assign y13860 = ~1'b0 ;
  assign y13861 = ~1'b0 ;
  assign y13862 = ~n20812 ;
  assign y13863 = ~n20813 ;
  assign y13864 = ~1'b0 ;
  assign y13865 = ~n20822 ;
  assign y13866 = ~1'b0 ;
  assign y13867 = ~1'b0 ;
  assign y13868 = ~1'b0 ;
  assign y13869 = ~1'b0 ;
  assign y13870 = ~n20827 ;
  assign y13871 = n1782 ;
  assign y13872 = ~n20829 ;
  assign y13873 = ~1'b0 ;
  assign y13874 = ~n20832 ;
  assign y13875 = ~n20833 ;
  assign y13876 = ~1'b0 ;
  assign y13877 = ~n20836 ;
  assign y13878 = ~1'b0 ;
  assign y13879 = ~1'b0 ;
  assign y13880 = ~1'b0 ;
  assign y13881 = ~1'b0 ;
  assign y13882 = n5768 ;
  assign y13883 = 1'b0 ;
  assign y13884 = ~1'b0 ;
  assign y13885 = ~1'b0 ;
  assign y13886 = n20837 ;
  assign y13887 = n6147 ;
  assign y13888 = ~n20838 ;
  assign y13889 = ~n20839 ;
  assign y13890 = n20840 ;
  assign y13891 = ~n20844 ;
  assign y13892 = n20846 ;
  assign y13893 = ~1'b0 ;
  assign y13894 = n8342 ;
  assign y13895 = ~1'b0 ;
  assign y13896 = ~n20849 ;
  assign y13897 = n20850 ;
  assign y13898 = n20852 ;
  assign y13899 = n20854 ;
  assign y13900 = ~n20856 ;
  assign y13901 = n20860 ;
  assign y13902 = 1'b0 ;
  assign y13903 = n20862 ;
  assign y13904 = ~1'b0 ;
  assign y13905 = ~1'b0 ;
  assign y13906 = n20867 ;
  assign y13907 = n20872 ;
  assign y13908 = ~n20873 ;
  assign y13909 = ~1'b0 ;
  assign y13910 = ~n20878 ;
  assign y13911 = ~n20879 ;
  assign y13912 = n20880 ;
  assign y13913 = ~1'b0 ;
  assign y13914 = ~1'b0 ;
  assign y13915 = n20884 ;
  assign y13916 = n20887 ;
  assign y13917 = ~1'b0 ;
  assign y13918 = x66 ;
  assign y13919 = n7631 ;
  assign y13920 = ~1'b0 ;
  assign y13921 = ~1'b0 ;
  assign y13922 = ~1'b0 ;
  assign y13923 = ~1'b0 ;
  assign y13924 = ~n20890 ;
  assign y13925 = n20891 ;
  assign y13926 = ~1'b0 ;
  assign y13927 = ~n20894 ;
  assign y13928 = ~1'b0 ;
  assign y13929 = n18653 ;
  assign y13930 = ~n20895 ;
  assign y13931 = ~1'b0 ;
  assign y13932 = ~n20897 ;
  assign y13933 = ~1'b0 ;
  assign y13934 = ~n20898 ;
  assign y13935 = 1'b0 ;
  assign y13936 = n20899 ;
  assign y13937 = ~n20900 ;
  assign y13938 = n20904 ;
  assign y13939 = ~1'b0 ;
  assign y13940 = n20906 ;
  assign y13941 = n20908 ;
  assign y13942 = ~n20909 ;
  assign y13943 = 1'b0 ;
  assign y13944 = ~n3622 ;
  assign y13945 = ~n20915 ;
  assign y13946 = ~n20917 ;
  assign y13947 = ~1'b0 ;
  assign y13948 = ~1'b0 ;
  assign y13949 = n20920 ;
  assign y13950 = n20922 ;
  assign y13951 = ~n20924 ;
  assign y13952 = ~1'b0 ;
  assign y13953 = ~1'b0 ;
  assign y13954 = ~n20926 ;
  assign y13955 = ~1'b0 ;
  assign y13956 = ~n20927 ;
  assign y13957 = ~1'b0 ;
  assign y13958 = ~n20931 ;
  assign y13959 = ~n20933 ;
  assign y13960 = n20938 ;
  assign y13961 = ~1'b0 ;
  assign y13962 = ~n20944 ;
  assign y13963 = n20950 ;
  assign y13964 = ~n20952 ;
  assign y13965 = n20953 ;
  assign y13966 = ~n20958 ;
  assign y13967 = ~n20959 ;
  assign y13968 = ~n20962 ;
  assign y13969 = ~n18060 ;
  assign y13970 = ~n20965 ;
  assign y13971 = ~n20966 ;
  assign y13972 = ~1'b0 ;
  assign y13973 = n20967 ;
  assign y13974 = ~1'b0 ;
  assign y13975 = n11859 ;
  assign y13976 = n20975 ;
  assign y13977 = ~n20976 ;
  assign y13978 = ~1'b0 ;
  assign y13979 = n20979 ;
  assign y13980 = ~1'b0 ;
  assign y13981 = ~n20980 ;
  assign y13982 = ~n20982 ;
  assign y13983 = ~1'b0 ;
  assign y13984 = ~n20985 ;
  assign y13985 = ~1'b0 ;
  assign y13986 = ~n9928 ;
  assign y13987 = ~n20987 ;
  assign y13988 = n20990 ;
  assign y13989 = n20992 ;
  assign y13990 = ~1'b0 ;
  assign y13991 = ~1'b0 ;
  assign y13992 = ~n20994 ;
  assign y13993 = 1'b0 ;
  assign y13994 = ~1'b0 ;
  assign y13995 = ~n20995 ;
  assign y13996 = ~1'b0 ;
  assign y13997 = ~1'b0 ;
  assign y13998 = ~1'b0 ;
  assign y13999 = ~1'b0 ;
  assign y14000 = n20996 ;
  assign y14001 = ~1'b0 ;
  assign y14002 = n20998 ;
  assign y14003 = n21000 ;
  assign y14004 = ~1'b0 ;
  assign y14005 = ~1'b0 ;
  assign y14006 = ~n21002 ;
  assign y14007 = ~1'b0 ;
  assign y14008 = ~n21003 ;
  assign y14009 = n21004 ;
  assign y14010 = ~1'b0 ;
  assign y14011 = n21005 ;
  assign y14012 = ~n21010 ;
  assign y14013 = ~n21012 ;
  assign y14014 = ~n21013 ;
  assign y14015 = x103 ;
  assign y14016 = ~1'b0 ;
  assign y14017 = ~n21016 ;
  assign y14018 = ~1'b0 ;
  assign y14019 = n15340 ;
  assign y14020 = ~1'b0 ;
  assign y14021 = ~n21017 ;
  assign y14022 = n21019 ;
  assign y14023 = ~1'b0 ;
  assign y14024 = ~n21021 ;
  assign y14025 = ~1'b0 ;
  assign y14026 = ~1'b0 ;
  assign y14027 = ~1'b0 ;
  assign y14028 = ~n19773 ;
  assign y14029 = ~1'b0 ;
  assign y14030 = n21023 ;
  assign y14031 = n21024 ;
  assign y14032 = ~1'b0 ;
  assign y14033 = ~1'b0 ;
  assign y14034 = n21027 ;
  assign y14035 = ~n21028 ;
  assign y14036 = n21030 ;
  assign y14037 = n21031 ;
  assign y14038 = ~1'b0 ;
  assign y14039 = ~n21032 ;
  assign y14040 = ~1'b0 ;
  assign y14041 = ~n4366 ;
  assign y14042 = ~1'b0 ;
  assign y14043 = ~n21033 ;
  assign y14044 = n21034 ;
  assign y14045 = ~n21035 ;
  assign y14046 = n20875 ;
  assign y14047 = ~1'b0 ;
  assign y14048 = ~n21037 ;
  assign y14049 = ~1'b0 ;
  assign y14050 = ~n21039 ;
  assign y14051 = ~1'b0 ;
  assign y14052 = n1566 ;
  assign y14053 = ~1'b0 ;
  assign y14054 = ~n21044 ;
  assign y14055 = 1'b0 ;
  assign y14056 = n21045 ;
  assign y14057 = ~1'b0 ;
  assign y14058 = 1'b0 ;
  assign y14059 = n10095 ;
  assign y14060 = ~n10235 ;
  assign y14061 = n21046 ;
  assign y14062 = ~1'b0 ;
  assign y14063 = ~1'b0 ;
  assign y14064 = ~1'b0 ;
  assign y14065 = n21048 ;
  assign y14066 = ~n20292 ;
  assign y14067 = ~n21050 ;
  assign y14068 = ~1'b0 ;
  assign y14069 = ~1'b0 ;
  assign y14070 = ~n9544 ;
  assign y14071 = ~n21051 ;
  assign y14072 = ~n21015 ;
  assign y14073 = n21052 ;
  assign y14074 = n21054 ;
  assign y14075 = ~1'b0 ;
  assign y14076 = n21057 ;
  assign y14077 = 1'b0 ;
  assign y14078 = ~n7383 ;
  assign y14079 = ~1'b0 ;
  assign y14080 = ~n21061 ;
  assign y14081 = ~n21063 ;
  assign y14082 = 1'b0 ;
  assign y14083 = ~n21066 ;
  assign y14084 = ~1'b0 ;
  assign y14085 = ~1'b0 ;
  assign y14086 = n21067 ;
  assign y14087 = ~n21069 ;
  assign y14088 = ~1'b0 ;
  assign y14089 = ~1'b0 ;
  assign y14090 = ~1'b0 ;
  assign y14091 = n21071 ;
  assign y14092 = n21073 ;
  assign y14093 = ~n1935 ;
  assign y14094 = ~n21075 ;
  assign y14095 = ~n21076 ;
  assign y14096 = 1'b0 ;
  assign y14097 = ~1'b0 ;
  assign y14098 = ~1'b0 ;
  assign y14099 = ~1'b0 ;
  assign y14100 = ~1'b0 ;
  assign y14101 = ~n9787 ;
  assign y14102 = ~1'b0 ;
  assign y14103 = ~n21080 ;
  assign y14104 = ~1'b0 ;
  assign y14105 = ~1'b0 ;
  assign y14106 = n21081 ;
  assign y14107 = ~n21082 ;
  assign y14108 = n21085 ;
  assign y14109 = ~1'b0 ;
  assign y14110 = ~1'b0 ;
  assign y14111 = ~1'b0 ;
  assign y14112 = n21086 ;
  assign y14113 = ~n21089 ;
  assign y14114 = ~n21091 ;
  assign y14115 = ~1'b0 ;
  assign y14116 = n12514 ;
  assign y14117 = ~1'b0 ;
  assign y14118 = n21092 ;
  assign y14119 = ~1'b0 ;
  assign y14120 = ~1'b0 ;
  assign y14121 = ~1'b0 ;
  assign y14122 = n21096 ;
  assign y14123 = ~1'b0 ;
  assign y14124 = n21097 ;
  assign y14125 = n21102 ;
  assign y14126 = ~1'b0 ;
  assign y14127 = n21105 ;
  assign y14128 = n11623 ;
  assign y14129 = n21106 ;
  assign y14130 = ~1'b0 ;
  assign y14131 = n21107 ;
  assign y14132 = ~n16224 ;
  assign y14133 = n21108 ;
  assign y14134 = n21109 ;
  assign y14135 = n21110 ;
  assign y14136 = n21113 ;
  assign y14137 = ~1'b0 ;
  assign y14138 = n21114 ;
  assign y14139 = ~1'b0 ;
  assign y14140 = n19624 ;
  assign y14141 = n21117 ;
  assign y14142 = ~1'b0 ;
  assign y14143 = ~1'b0 ;
  assign y14144 = ~n1103 ;
  assign y14145 = ~n5603 ;
  assign y14146 = ~1'b0 ;
  assign y14147 = ~n21118 ;
  assign y14148 = n21121 ;
  assign y14149 = n21124 ;
  assign y14150 = n21128 ;
  assign y14151 = ~n21130 ;
  assign y14152 = ~1'b0 ;
  assign y14153 = n21131 ;
  assign y14154 = ~n21133 ;
  assign y14155 = n15292 ;
  assign y14156 = ~n21138 ;
  assign y14157 = n21139 ;
  assign y14158 = ~n17755 ;
  assign y14159 = n21140 ;
  assign y14160 = ~n21141 ;
  assign y14161 = n8619 ;
  assign y14162 = ~n21142 ;
  assign y14163 = n21145 ;
  assign y14164 = ~1'b0 ;
  assign y14165 = n4847 ;
  assign y14166 = ~n21147 ;
  assign y14167 = ~n21148 ;
  assign y14168 = n21149 ;
  assign y14169 = ~n13969 ;
  assign y14170 = ~n21154 ;
  assign y14171 = n21157 ;
  assign y14172 = ~1'b0 ;
  assign y14173 = ~n11563 ;
  assign y14174 = ~n21158 ;
  assign y14175 = ~n21161 ;
  assign y14176 = n4901 ;
  assign y14177 = ~n21163 ;
  assign y14178 = ~n21169 ;
  assign y14179 = ~n21172 ;
  assign y14180 = ~1'b0 ;
  assign y14181 = ~1'b0 ;
  assign y14182 = ~n21174 ;
  assign y14183 = n21175 ;
  assign y14184 = 1'b0 ;
  assign y14185 = n623 ;
  assign y14186 = n21176 ;
  assign y14187 = ~1'b0 ;
  assign y14188 = 1'b0 ;
  assign y14189 = ~n21178 ;
  assign y14190 = ~1'b0 ;
  assign y14191 = ~n21180 ;
  assign y14192 = n21186 ;
  assign y14193 = ~n21191 ;
  assign y14194 = ~1'b0 ;
  assign y14195 = ~1'b0 ;
  assign y14196 = n1635 ;
  assign y14197 = n21192 ;
  assign y14198 = n21194 ;
  assign y14199 = ~1'b0 ;
  assign y14200 = n21197 ;
  assign y14201 = n21198 ;
  assign y14202 = ~n21200 ;
  assign y14203 = ~1'b0 ;
  assign y14204 = n21202 ;
  assign y14205 = ~1'b0 ;
  assign y14206 = ~1'b0 ;
  assign y14207 = ~1'b0 ;
  assign y14208 = ~1'b0 ;
  assign y14209 = ~n15908 ;
  assign y14210 = ~1'b0 ;
  assign y14211 = ~n21204 ;
  assign y14212 = n19856 ;
  assign y14213 = ~1'b0 ;
  assign y14214 = ~1'b0 ;
  assign y14215 = ~n8831 ;
  assign y14216 = ~1'b0 ;
  assign y14217 = x50 ;
  assign y14218 = n21205 ;
  assign y14219 = n21208 ;
  assign y14220 = ~1'b0 ;
  assign y14221 = ~n21210 ;
  assign y14222 = ~n21214 ;
  assign y14223 = n21216 ;
  assign y14224 = n21218 ;
  assign y14225 = n21220 ;
  assign y14226 = ~n21223 ;
  assign y14227 = ~1'b0 ;
  assign y14228 = n15181 ;
  assign y14229 = ~1'b0 ;
  assign y14230 = n21225 ;
  assign y14231 = ~1'b0 ;
  assign y14232 = n21227 ;
  assign y14233 = ~n21228 ;
  assign y14234 = ~n21229 ;
  assign y14235 = ~n21230 ;
  assign y14236 = ~n21233 ;
  assign y14237 = 1'b0 ;
  assign y14238 = ~1'b0 ;
  assign y14239 = n21234 ;
  assign y14240 = ~n21235 ;
  assign y14241 = ~1'b0 ;
  assign y14242 = ~1'b0 ;
  assign y14243 = ~n4394 ;
  assign y14244 = n21237 ;
  assign y14245 = n21238 ;
  assign y14246 = ~n21239 ;
  assign y14247 = ~n21240 ;
  assign y14248 = n10816 ;
  assign y14249 = ~n21241 ;
  assign y14250 = ~1'b0 ;
  assign y14251 = ~n21246 ;
  assign y14252 = ~1'b0 ;
  assign y14253 = ~n21247 ;
  assign y14254 = n21251 ;
  assign y14255 = n21253 ;
  assign y14256 = n21254 ;
  assign y14257 = n21256 ;
  assign y14258 = n21257 ;
  assign y14259 = ~1'b0 ;
  assign y14260 = ~1'b0 ;
  assign y14261 = n21259 ;
  assign y14262 = ~n21260 ;
  assign y14263 = ~n21261 ;
  assign y14264 = ~x16 ;
  assign y14265 = n21265 ;
  assign y14266 = ~1'b0 ;
  assign y14267 = ~1'b0 ;
  assign y14268 = ~1'b0 ;
  assign y14269 = ~n21267 ;
  assign y14270 = ~1'b0 ;
  assign y14271 = ~1'b0 ;
  assign y14272 = ~1'b0 ;
  assign y14273 = n21268 ;
  assign y14274 = ~n17311 ;
  assign y14275 = n21269 ;
  assign y14276 = ~1'b0 ;
  assign y14277 = n21272 ;
  assign y14278 = ~n19582 ;
  assign y14279 = n21274 ;
  assign y14280 = ~n21277 ;
  assign y14281 = ~n21279 ;
  assign y14282 = ~1'b0 ;
  assign y14283 = n21282 ;
  assign y14284 = ~n21283 ;
  assign y14285 = ~n21286 ;
  assign y14286 = n21288 ;
  assign y14287 = 1'b0 ;
  assign y14288 = ~n21289 ;
  assign y14289 = n21290 ;
  assign y14290 = n21291 ;
  assign y14291 = ~1'b0 ;
  assign y14292 = ~1'b0 ;
  assign y14293 = n21292 ;
  assign y14294 = n21295 ;
  assign y14295 = n21296 ;
  assign y14296 = ~n21297 ;
  assign y14297 = n5861 ;
  assign y14298 = n21301 ;
  assign y14299 = ~1'b0 ;
  assign y14300 = ~1'b0 ;
  assign y14301 = ~n21302 ;
  assign y14302 = ~n21303 ;
  assign y14303 = ~1'b0 ;
  assign y14304 = ~n21308 ;
  assign y14305 = ~n21310 ;
  assign y14306 = ~n21312 ;
  assign y14307 = ~1'b0 ;
  assign y14308 = n21314 ;
  assign y14309 = ~1'b0 ;
  assign y14310 = ~n21319 ;
  assign y14311 = n21321 ;
  assign y14312 = n21323 ;
  assign y14313 = ~1'b0 ;
  assign y14314 = ~1'b0 ;
  assign y14315 = ~1'b0 ;
  assign y14316 = ~n21324 ;
  assign y14317 = n21326 ;
  assign y14318 = n21327 ;
  assign y14319 = n21330 ;
  assign y14320 = n21331 ;
  assign y14321 = ~n15752 ;
  assign y14322 = n21332 ;
  assign y14323 = n21334 ;
  assign y14324 = ~1'b0 ;
  assign y14325 = n21335 ;
  assign y14326 = n21337 ;
  assign y14327 = n21338 ;
  assign y14328 = ~n21344 ;
  assign y14329 = n21347 ;
  assign y14330 = n21348 ;
  assign y14331 = ~1'b0 ;
  assign y14332 = ~1'b0 ;
  assign y14333 = ~1'b0 ;
  assign y14334 = ~1'b0 ;
  assign y14335 = ~1'b0 ;
  assign y14336 = ~n9778 ;
  assign y14337 = ~n21349 ;
  assign y14338 = ~n21352 ;
  assign y14339 = ~1'b0 ;
  assign y14340 = ~1'b0 ;
  assign y14341 = ~n6648 ;
  assign y14342 = ~n21353 ;
  assign y14343 = ~n21355 ;
  assign y14344 = n21357 ;
  assign y14345 = ~1'b0 ;
  assign y14346 = ~n21359 ;
  assign y14347 = 1'b0 ;
  assign y14348 = ~n21360 ;
  assign y14349 = ~n21362 ;
  assign y14350 = ~n21367 ;
  assign y14351 = ~1'b0 ;
  assign y14352 = ~n21369 ;
  assign y14353 = n21370 ;
  assign y14354 = n21372 ;
  assign y14355 = ~n21378 ;
  assign y14356 = ~n21383 ;
  assign y14357 = ~1'b0 ;
  assign y14358 = ~1'b0 ;
  assign y14359 = ~1'b0 ;
  assign y14360 = ~n21385 ;
  assign y14361 = ~1'b0 ;
  assign y14362 = ~1'b0 ;
  assign y14363 = ~n21386 ;
  assign y14364 = ~1'b0 ;
  assign y14365 = n21387 ;
  assign y14366 = ~n21391 ;
  assign y14367 = n21392 ;
  assign y14368 = ~1'b0 ;
  assign y14369 = n21394 ;
  assign y14370 = ~1'b0 ;
  assign y14371 = ~n21399 ;
  assign y14372 = 1'b0 ;
  assign y14373 = ~n877 ;
  assign y14374 = ~n21402 ;
  assign y14375 = ~1'b0 ;
  assign y14376 = n16041 ;
  assign y14377 = n21403 ;
  assign y14378 = n21406 ;
  assign y14379 = n15127 ;
  assign y14380 = ~1'b0 ;
  assign y14381 = ~n21407 ;
  assign y14382 = n21410 ;
  assign y14383 = ~n21411 ;
  assign y14384 = n20183 ;
  assign y14385 = ~1'b0 ;
  assign y14386 = n21414 ;
  assign y14387 = n21416 ;
  assign y14388 = ~1'b0 ;
  assign y14389 = ~1'b0 ;
  assign y14390 = ~n15937 ;
  assign y14391 = ~n21419 ;
  assign y14392 = ~1'b0 ;
  assign y14393 = ~1'b0 ;
  assign y14394 = ~n21422 ;
  assign y14395 = ~n21424 ;
  assign y14396 = n21425 ;
  assign y14397 = n21426 ;
  assign y14398 = ~n21427 ;
  assign y14399 = ~n21430 ;
  assign y14400 = 1'b0 ;
  assign y14401 = 1'b0 ;
  assign y14402 = 1'b0 ;
  assign y14403 = ~n185 ;
  assign y14404 = ~1'b0 ;
  assign y14405 = ~1'b0 ;
  assign y14406 = n21432 ;
  assign y14407 = ~n21433 ;
  assign y14408 = ~1'b0 ;
  assign y14409 = ~1'b0 ;
  assign y14410 = ~n17393 ;
  assign y14411 = ~1'b0 ;
  assign y14412 = ~1'b0 ;
  assign y14413 = ~n21434 ;
  assign y14414 = ~1'b0 ;
  assign y14415 = ~n21436 ;
  assign y14416 = ~1'b0 ;
  assign y14417 = ~1'b0 ;
endmodule
