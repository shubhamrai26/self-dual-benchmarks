module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 ;
  assign n129 = ( x70 & ~x93 ) | ( x70 & x110 ) | ( ~x93 & x110 ) ;
  assign n130 = x17 & x125 ;
  assign n131 = ~x107 & n130 ;
  assign n132 = x75 ^ x3 ^ 1'b0 ;
  assign n133 = x93 & n132 ;
  assign n134 = ( x15 & ~x18 ) | ( x15 & x40 ) | ( ~x18 & x40 ) ;
  assign n136 = x9 & x91 ;
  assign n137 = n136 ^ x102 ^ 1'b0 ;
  assign n135 = x18 & x86 ;
  assign n138 = n137 ^ n135 ^ 1'b0 ;
  assign n139 = ( ~x83 & x112 ) | ( ~x83 & n129 ) | ( x112 & n129 ) ;
  assign n140 = x81 & x105 ;
  assign n141 = ~x67 & n140 ;
  assign n142 = x95 ^ x49 ^ 1'b0 ;
  assign n143 = x1 & n142 ;
  assign n144 = ( ~x65 & x109 ) | ( ~x65 & n143 ) | ( x109 & n143 ) ;
  assign n145 = x67 & ~x77 ;
  assign n146 = x57 & x104 ;
  assign n147 = ~x123 & n146 ;
  assign n148 = x108 ^ x68 ^ x60 ;
  assign n149 = x22 & ~n148 ;
  assign n150 = ~x56 & n149 ;
  assign n151 = x33 & x92 ;
  assign n152 = n151 ^ x11 ^ 1'b0 ;
  assign n153 = x17 & x111 ;
  assign n154 = n152 & n153 ;
  assign n155 = x33 & x65 ;
  assign n156 = n155 ^ x28 ^ 1'b0 ;
  assign n157 = n156 ^ n138 ^ x34 ;
  assign n158 = x65 & x79 ;
  assign n159 = n158 ^ x8 ^ 1'b0 ;
  assign n160 = x31 & x40 ;
  assign n161 = n160 ^ n154 ^ 1'b0 ;
  assign n162 = n134 ^ x21 ^ 1'b0 ;
  assign n163 = x109 & n162 ;
  assign n164 = x47 & x95 ;
  assign n165 = ~x38 & n164 ;
  assign n166 = ( ~x86 & x112 ) | ( ~x86 & n165 ) | ( x112 & n165 ) ;
  assign n167 = ~x4 & x59 ;
  assign n172 = x80 & x92 ;
  assign n168 = x84 & x106 ;
  assign n169 = ~x2 & n168 ;
  assign n170 = x46 & ~n169 ;
  assign n171 = ~x64 & n170 ;
  assign n173 = n172 ^ n171 ^ 1'b0 ;
  assign n174 = n167 | n173 ;
  assign n175 = x123 ^ x90 ^ 1'b0 ;
  assign n176 = x61 & ~n175 ;
  assign n177 = n156 & n176 ;
  assign n178 = x19 ^ x17 ^ 1'b0 ;
  assign n179 = x4 & n178 ;
  assign n180 = x96 ^ x54 ^ x41 ;
  assign n181 = x76 & ~n180 ;
  assign n182 = ~n179 & n181 ;
  assign n183 = x5 & x31 ;
  assign n184 = n183 ^ x64 ^ 1'b0 ;
  assign n185 = x49 & x91 ;
  assign n186 = n185 ^ x103 ^ 1'b0 ;
  assign n187 = x7 & x56 ;
  assign n188 = n186 & n187 ;
  assign n189 = n166 ^ x17 ^ 1'b0 ;
  assign n190 = x111 & ~n189 ;
  assign n191 = n143 ^ x123 ^ 1'b0 ;
  assign n192 = ~n175 & n191 ;
  assign n193 = x88 & n192 ;
  assign n194 = ~x116 & n193 ;
  assign n195 = x45 & ~x53 ;
  assign n196 = x63 & x96 ;
  assign n197 = x82 ^ x81 ^ 1'b0 ;
  assign n198 = x33 & n197 ;
  assign n199 = x117 ^ x14 ^ 1'b0 ;
  assign n200 = n198 & n199 ;
  assign n201 = x38 & n200 ;
  assign n202 = ~x89 & n201 ;
  assign n203 = n138 ^ x113 ^ x53 ;
  assign n204 = x39 ^ x32 ^ x28 ;
  assign n205 = ( x12 & n203 ) | ( x12 & ~n204 ) | ( n203 & ~n204 ) ;
  assign n207 = x93 & x99 ;
  assign n208 = n131 & n207 ;
  assign n209 = x78 & n208 ;
  assign n206 = x66 & n198 ;
  assign n210 = n209 ^ n206 ^ 1'b0 ;
  assign n212 = x49 ^ x34 ^ 1'b0 ;
  assign n213 = x65 & n212 ;
  assign n214 = n133 & n213 ;
  assign n215 = n214 ^ x80 ^ 1'b0 ;
  assign n216 = n215 ^ x91 ^ 1'b0 ;
  assign n217 = x47 & ~n216 ;
  assign n211 = x8 & x35 ;
  assign n218 = n217 ^ n211 ^ 1'b0 ;
  assign n219 = n182 ^ x52 ^ 1'b0 ;
  assign n220 = n147 | n219 ;
  assign n221 = x26 & x125 ;
  assign n222 = n221 ^ x2 ^ 1'b0 ;
  assign n223 = n222 ^ x16 ^ 1'b0 ;
  assign n224 = n156 | n223 ;
  assign n225 = ~x121 & n179 ;
  assign n226 = n159 ^ x39 ^ 1'b0 ;
  assign n227 = x37 & ~n226 ;
  assign n228 = n133 ^ x14 ^ 1'b0 ;
  assign n229 = x65 & n228 ;
  assign n230 = x96 ^ x88 ^ 1'b0 ;
  assign n231 = n229 & n230 ;
  assign n232 = ( x56 & x105 ) | ( x56 & ~x111 ) | ( x105 & ~x111 ) ;
  assign n233 = x77 ^ x71 ^ 1'b0 ;
  assign n234 = ~n180 & n233 ;
  assign n235 = n232 & n234 ;
  assign n236 = n235 ^ n200 ^ 1'b0 ;
  assign n237 = x45 & x66 ;
  assign n238 = ~x2 & n237 ;
  assign n239 = x1 & x33 ;
  assign n240 = n179 ^ x55 ^ 1'b0 ;
  assign n241 = ( x22 & n188 ) | ( x22 & n240 ) | ( n188 & n240 ) ;
  assign n242 = x126 & n241 ;
  assign n243 = ~n239 & n242 ;
  assign n244 = n243 ^ n196 ^ x25 ;
  assign n245 = n244 ^ x86 ^ 1'b0 ;
  assign n246 = n213 & n245 ;
  assign n248 = x113 ^ x16 ^ 1'b0 ;
  assign n249 = x115 & n248 ;
  assign n247 = ~n141 & n234 ;
  assign n250 = n249 ^ n247 ^ 1'b0 ;
  assign n251 = x72 & x82 ;
  assign n252 = ~n240 & n251 ;
  assign n253 = x0 & x25 ;
  assign n254 = ~x15 & n253 ;
  assign n255 = n229 | n254 ;
  assign n256 = x61 & ~x66 ;
  assign n257 = n167 ^ x94 ^ 1'b0 ;
  assign n258 = n171 ^ n138 ^ x34 ;
  assign n259 = x106 & x122 ;
  assign n260 = ~n258 & n259 ;
  assign n261 = n205 ^ x34 ^ 1'b0 ;
  assign n268 = x83 ^ x17 ^ 1'b0 ;
  assign n269 = n239 & n268 ;
  assign n271 = x89 & ~n148 ;
  assign n272 = ~x121 & n271 ;
  assign n270 = x91 & n234 ;
  assign n273 = n272 ^ n270 ^ 1'b0 ;
  assign n274 = n269 & n273 ;
  assign n275 = n274 ^ x11 ^ 1'b0 ;
  assign n264 = x67 & x106 ;
  assign n265 = n264 ^ n131 ^ 1'b0 ;
  assign n262 = ~x34 & x38 ;
  assign n263 = ~n186 & n262 ;
  assign n266 = n265 ^ n263 ^ 1'b0 ;
  assign n267 = n266 ^ x71 ^ x57 ;
  assign n276 = n275 ^ n267 ^ x31 ;
  assign n277 = ( x6 & x49 ) | ( x6 & n182 ) | ( x49 & n182 ) ;
  assign n278 = x113 ^ x64 ^ x53 ;
  assign n279 = n278 ^ n157 ^ 1'b0 ;
  assign n280 = ~n222 & n279 ;
  assign n281 = ~x7 & n280 ;
  assign n282 = n195 & ~n220 ;
  assign n283 = n281 & n282 ;
  assign n284 = ~n150 & n231 ;
  assign n285 = n284 ^ x117 ^ 1'b0 ;
  assign n286 = x102 & n217 ;
  assign n287 = n286 ^ x31 ^ 1'b0 ;
  assign n288 = ~x58 & x60 ;
  assign n289 = x6 & x12 ;
  assign n290 = n289 ^ x47 ^ 1'b0 ;
  assign n291 = n137 | n141 ;
  assign n292 = n291 ^ x91 ^ 1'b0 ;
  assign n293 = n290 & n292 ;
  assign n294 = n250 ^ x24 ^ 1'b0 ;
  assign n295 = x78 & x107 ;
  assign n296 = n295 ^ x52 ^ 1'b0 ;
  assign n297 = x96 & ~n296 ;
  assign n298 = x60 & x96 ;
  assign n299 = ~x79 & n298 ;
  assign n300 = n255 & ~n299 ;
  assign n301 = ~x121 & n300 ;
  assign n302 = x10 & n204 ;
  assign n303 = x65 ^ x62 ^ x51 ;
  assign n304 = n302 | n303 ;
  assign n305 = n266 & ~n304 ;
  assign n306 = x57 & ~n305 ;
  assign n307 = ~x16 & n306 ;
  assign n308 = x8 & n179 ;
  assign n309 = n308 ^ x39 ^ 1'b0 ;
  assign n310 = n229 & ~n309 ;
  assign n311 = n310 ^ n243 ^ 1'b0 ;
  assign n312 = x26 & n311 ;
  assign n313 = ~x50 & n312 ;
  assign n314 = x77 ^ x72 ^ 1'b0 ;
  assign n315 = x26 & n314 ;
  assign n316 = ~n147 & n315 ;
  assign n317 = ~x60 & n316 ;
  assign n318 = n137 ^ x87 ^ 1'b0 ;
  assign n319 = n318 ^ n275 ^ x79 ;
  assign n320 = n319 ^ x52 ^ 1'b0 ;
  assign n321 = ~n317 & n320 ;
  assign n322 = x27 & n133 ;
  assign n323 = n322 ^ n303 ^ 1'b0 ;
  assign n324 = n323 ^ n141 ^ x49 ;
  assign n325 = ~n203 & n324 ;
  assign n326 = n325 ^ n258 ^ 1'b0 ;
  assign n329 = x91 & n279 ;
  assign n330 = ~x65 & n329 ;
  assign n327 = ( x27 & x29 ) | ( x27 & ~n323 ) | ( x29 & ~n323 ) ;
  assign n328 = n192 & n327 ;
  assign n331 = n330 ^ n328 ^ 1'b0 ;
  assign n332 = n262 ^ n177 ^ x125 ;
  assign n333 = n332 ^ x104 ^ 1'b0 ;
  assign n334 = x55 & n333 ;
  assign n335 = ( ~x115 & x124 ) | ( ~x115 & n154 ) | ( x124 & n154 ) ;
  assign n336 = n335 ^ x44 ^ 1'b0 ;
  assign n337 = n150 | n278 ;
  assign n338 = n215 & ~n337 ;
  assign n339 = ( x73 & n283 ) | ( x73 & ~n338 ) | ( n283 & ~n338 ) ;
  assign n340 = x103 & ~n186 ;
  assign n341 = x116 ^ x12 ^ 1'b0 ;
  assign n342 = n279 & n341 ;
  assign n343 = n340 & n342 ;
  assign n344 = ~x24 & n343 ;
  assign n345 = x121 ^ x100 ^ 1'b0 ;
  assign n346 = x48 & x99 ;
  assign n347 = n346 ^ x123 ^ 1'b0 ;
  assign n348 = n208 | n347 ;
  assign n349 = n348 ^ x85 ^ 1'b0 ;
  assign n350 = x57 & n349 ;
  assign n351 = ~x51 & n350 ;
  assign n352 = x14 & ~n186 ;
  assign n353 = n352 ^ n129 ^ 1'b0 ;
  assign n354 = n190 & ~n236 ;
  assign n355 = n335 & n354 ;
  assign n356 = n355 ^ n210 ^ 1'b0 ;
  assign n357 = n353 | n356 ;
  assign n358 = ( x58 & n159 ) | ( x58 & n357 ) | ( n159 & n357 ) ;
  assign n359 = n177 | n277 ;
  assign n360 = x74 & n319 ;
  assign n361 = n224 & n360 ;
  assign n362 = x92 ^ x84 ^ 1'b0 ;
  assign n363 = x105 & n362 ;
  assign n364 = ~n196 & n239 ;
  assign n365 = n172 ^ x87 ^ 1'b0 ;
  assign n366 = x72 & n365 ;
  assign n367 = ~n364 & n366 ;
  assign n368 = ~n359 & n367 ;
  assign n369 = n281 ^ n180 ^ x115 ;
  assign n370 = n315 ^ n213 ^ 1'b0 ;
  assign n371 = x49 & n370 ;
  assign n372 = x67 & x122 ;
  assign n373 = ~n231 & n372 ;
  assign n374 = n373 ^ n326 ^ 1'b0 ;
  assign n375 = x125 ^ x23 ^ 1'b0 ;
  assign n376 = n234 & n375 ;
  assign n377 = n182 & n376 ;
  assign n378 = n377 ^ n363 ^ 1'b0 ;
  assign n379 = x0 & n378 ;
  assign n380 = x89 & ~n299 ;
  assign n381 = n208 & n380 ;
  assign n382 = n287 ^ x39 ^ 1'b0 ;
  assign n383 = n238 | n382 ;
  assign n384 = n383 ^ n163 ^ 1'b0 ;
  assign n385 = ~n351 & n384 ;
  assign n386 = n381 & n385 ;
  assign n387 = n205 ^ x56 ^ x19 ;
  assign n388 = ( x105 & ~n225 ) | ( x105 & n387 ) | ( ~n225 & n387 ) ;
  assign n390 = n232 ^ x18 ^ 1'b0 ;
  assign n391 = x26 & n390 ;
  assign n389 = n236 ^ n209 ^ x39 ;
  assign n392 = n391 ^ n389 ^ 1'b0 ;
  assign n393 = x18 & ~x63 ;
  assign n396 = n303 ^ x38 ^ 1'b0 ;
  assign n397 = x115 & ~n396 ;
  assign n394 = x104 & ~n224 ;
  assign n395 = n394 ^ n134 ^ 1'b0 ;
  assign n398 = n397 ^ n395 ^ x65 ;
  assign n399 = x65 | n148 ;
  assign n400 = n399 ^ n299 ^ 1'b0 ;
  assign n401 = x103 | n400 ;
  assign n402 = n364 ^ x109 ^ 1'b0 ;
  assign n403 = ~n401 & n402 ;
  assign n404 = ~n166 & n302 ;
  assign n406 = x108 ^ x86 ^ 1'b0 ;
  assign n405 = n184 | n381 ;
  assign n407 = n406 ^ n405 ^ 1'b0 ;
  assign n408 = x53 & x54 ;
  assign n409 = n194 & n408 ;
  assign n410 = x43 & n138 ;
  assign n411 = ~x29 & n410 ;
  assign n412 = ( x105 & ~n231 ) | ( x105 & n256 ) | ( ~n231 & n256 ) ;
  assign n413 = n411 | n412 ;
  assign n414 = n409 & ~n413 ;
  assign n415 = x8 & ~x25 ;
  assign n416 = x124 & n179 ;
  assign n417 = n416 ^ n205 ^ 1'b0 ;
  assign n418 = x61 & x112 ;
  assign n419 = n418 ^ n138 ^ 1'b0 ;
  assign n420 = n419 ^ x5 ^ 1'b0 ;
  assign n421 = n147 | n420 ;
  assign n422 = x119 & ~n381 ;
  assign n423 = ~x26 & n422 ;
  assign n424 = n166 | n423 ;
  assign n425 = x50 | n424 ;
  assign n426 = n261 ^ x92 ^ 1'b0 ;
  assign n427 = x80 & n426 ;
  assign n428 = ( x94 & n225 ) | ( x94 & ~n427 ) | ( n225 & ~n427 ) ;
  assign n435 = ( x0 & x8 ) | ( x0 & ~x29 ) | ( x8 & ~x29 ) ;
  assign n436 = n215 ^ x65 ^ 1'b0 ;
  assign n437 = n435 & n436 ;
  assign n429 = n347 ^ x116 ^ 1'b0 ;
  assign n430 = x103 & ~n429 ;
  assign n431 = n430 ^ x115 ^ x50 ;
  assign n432 = x31 & ~n165 ;
  assign n433 = ~n273 & n432 ;
  assign n434 = n431 | n433 ;
  assign n438 = n437 ^ n434 ^ 1'b0 ;
  assign n439 = x120 & ~n171 ;
  assign n440 = n439 ^ x32 ^ 1'b0 ;
  assign n441 = n362 ^ x56 ^ 1'b0 ;
  assign n442 = x121 & ~n441 ;
  assign n443 = n331 & n442 ;
  assign n444 = n440 & n443 ;
  assign n445 = n204 ^ x24 ^ 1'b0 ;
  assign n446 = x88 | n287 ;
  assign n447 = ~n377 & n446 ;
  assign n448 = ~n129 & n447 ;
  assign n449 = n400 ^ x115 ^ 1'b0 ;
  assign n450 = n330 | n449 ;
  assign n451 = n156 | n450 ;
  assign n452 = n451 ^ n252 ^ 1'b0 ;
  assign n453 = n433 ^ n276 ^ 1'b0 ;
  assign n454 = n453 ^ n311 ^ 1'b0 ;
  assign n455 = n452 | n454 ;
  assign n456 = n137 & n276 ;
  assign n457 = n381 ^ n258 ^ 1'b0 ;
  assign n458 = x34 & ~n457 ;
  assign n459 = ~n154 & n283 ;
  assign n460 = n393 ^ n144 ^ 1'b0 ;
  assign n461 = n459 | n460 ;
  assign n462 = ( x64 & ~x72 ) | ( x64 & x77 ) | ( ~x72 & x77 ) ;
  assign n463 = n260 ^ n227 ^ 1'b0 ;
  assign n464 = n462 | n463 ;
  assign n465 = x64 & ~n381 ;
  assign n466 = n464 & n465 ;
  assign n467 = x17 & ~n420 ;
  assign n468 = n466 & n467 ;
  assign n469 = x29 & x78 ;
  assign n470 = n241 & n469 ;
  assign n471 = n470 ^ n208 ^ 1'b0 ;
  assign n472 = ~x74 & n471 ;
  assign n474 = x68 ^ x38 ^ 1'b0 ;
  assign n475 = x67 & n474 ;
  assign n473 = ~n147 & n196 ;
  assign n476 = n475 ^ n473 ^ 1'b0 ;
  assign n477 = ~x117 & n198 ;
  assign n478 = x115 | n477 ;
  assign n479 = ( ~n278 & n427 ) | ( ~n278 & n478 ) | ( n427 & n478 ) ;
  assign n480 = n145 ^ x65 ^ 1'b0 ;
  assign n481 = n480 ^ n208 ^ x97 ;
  assign n482 = n326 | n409 ;
  assign n483 = n482 ^ n387 ^ 1'b0 ;
  assign n484 = n243 ^ n171 ^ 1'b0 ;
  assign n485 = n484 ^ n260 ^ 1'b0 ;
  assign n486 = ~n387 & n485 ;
  assign n487 = ( n171 & n236 ) | ( n171 & n438 ) | ( n236 & n438 ) ;
  assign n488 = n213 ^ x81 ^ 1'b0 ;
  assign n489 = ( x90 & n134 ) | ( x90 & n488 ) | ( n134 & n488 ) ;
  assign n490 = x52 & x65 ;
  assign n491 = n161 & n490 ;
  assign n492 = x41 & ~n362 ;
  assign n493 = n492 ^ n309 ^ 1'b0 ;
  assign n494 = ~n491 & n493 ;
  assign n495 = n373 ^ x70 ^ 1'b0 ;
  assign n496 = n234 & ~n495 ;
  assign n497 = x25 & x120 ;
  assign n498 = n497 ^ n277 ^ 1'b0 ;
  assign n499 = n498 ^ n347 ^ n200 ;
  assign n500 = ~n186 & n499 ;
  assign n501 = n500 ^ n336 ^ 1'b0 ;
  assign n502 = n336 ^ n252 ^ 1'b0 ;
  assign n503 = x40 & ~n502 ;
  assign n504 = x57 & ~n503 ;
  assign n505 = n446 & ~n452 ;
  assign n506 = n505 ^ x91 ^ 1'b0 ;
  assign n507 = x61 & ~n395 ;
  assign n508 = x108 & ~n145 ;
  assign n509 = n508 ^ n267 ^ 1'b0 ;
  assign n510 = x81 ^ x44 ^ 1'b0 ;
  assign n511 = x6 & n510 ;
  assign n512 = n511 ^ n180 ^ 1'b0 ;
  assign n513 = n509 | n512 ;
  assign n514 = n409 ^ x109 ^ 1'b0 ;
  assign n515 = x110 & ~n514 ;
  assign n516 = n192 & n515 ;
  assign n517 = n513 & n516 ;
  assign n518 = ( x117 & n507 ) | ( x117 & n517 ) | ( n507 & n517 ) ;
  assign n519 = ( n244 & n435 ) | ( n244 & ~n518 ) | ( n435 & ~n518 ) ;
  assign n520 = x35 & ~n252 ;
  assign n521 = ~n349 & n520 ;
  assign n522 = n150 | n521 ;
  assign n523 = x30 | n522 ;
  assign n524 = ~n335 & n523 ;
  assign n525 = n524 ^ n513 ^ 1'b0 ;
  assign n526 = n444 ^ n401 ^ 1'b0 ;
  assign n527 = n525 & n526 ;
  assign n528 = x41 & ~n141 ;
  assign n529 = n528 ^ x75 ^ 1'b0 ;
  assign n530 = n529 ^ n141 ^ 1'b0 ;
  assign n531 = n366 & ~n530 ;
  assign n532 = x63 & n327 ;
  assign n533 = ~n234 & n532 ;
  assign n534 = x115 & n148 ;
  assign n535 = n190 & ~n309 ;
  assign n536 = ~x97 & n535 ;
  assign n537 = x20 ^ x14 ^ 1'b0 ;
  assign n538 = ~n536 & n537 ;
  assign n539 = n475 ^ x95 ^ 1'b0 ;
  assign n540 = n404 ^ n377 ^ n254 ;
  assign n541 = n281 | n330 ;
  assign n542 = x3 & ~x114 ;
  assign n543 = n315 ^ n220 ^ x34 ;
  assign n544 = n511 & n543 ;
  assign n545 = ~x62 & n544 ;
  assign n546 = x110 ^ x22 ^ 1'b0 ;
  assign n547 = ~n256 & n546 ;
  assign n548 = n547 ^ n507 ^ 1'b0 ;
  assign n549 = n156 ^ x14 ^ 1'b0 ;
  assign n550 = ~n260 & n511 ;
  assign n551 = ~n549 & n550 ;
  assign n552 = x78 ^ x48 ^ 1'b0 ;
  assign n553 = ~n152 & n552 ;
  assign n554 = ~n166 & n553 ;
  assign n555 = n309 & n554 ;
  assign n556 = ( x11 & n290 ) | ( x11 & ~n301 ) | ( n290 & ~n301 ) ;
  assign n557 = n555 | n556 ;
  assign n558 = n430 ^ n261 ^ 1'b0 ;
  assign n559 = x117 & n558 ;
  assign n560 = ( x61 & x71 ) | ( x61 & n165 ) | ( x71 & n165 ) ;
  assign n561 = x21 & x109 ;
  assign n562 = n561 ^ n488 ^ 1'b0 ;
  assign n563 = n244 & n562 ;
  assign n564 = n560 & n563 ;
  assign n565 = n564 ^ x10 ^ 1'b0 ;
  assign n566 = n565 ^ n364 ^ 1'b0 ;
  assign n567 = x18 & n566 ;
  assign n568 = n567 ^ n478 ^ 1'b0 ;
  assign n569 = n559 & ~n568 ;
  assign n570 = ~n456 & n569 ;
  assign n571 = n570 ^ n401 ^ 1'b0 ;
  assign n572 = x63 & x103 ;
  assign n573 = ~n240 & n572 ;
  assign n574 = x93 ^ x32 ^ 1'b0 ;
  assign n575 = ~n415 & n574 ;
  assign n576 = x112 & n575 ;
  assign n577 = n573 & n576 ;
  assign n578 = ( x118 & n509 ) | ( x118 & ~n539 ) | ( n509 & ~n539 ) ;
  assign n579 = n411 ^ x82 ^ 1'b0 ;
  assign n580 = x114 & ~n579 ;
  assign n581 = n500 ^ n353 ^ x101 ;
  assign n582 = n581 ^ n249 ^ 1'b0 ;
  assign n583 = ~n521 & n582 ;
  assign n584 = n275 ^ x39 ^ 1'b0 ;
  assign n585 = n553 & ~n584 ;
  assign n586 = ( x1 & n131 ) | ( x1 & n165 ) | ( n131 & n165 ) ;
  assign n587 = x91 & n452 ;
  assign n588 = ( n227 & n586 ) | ( n227 & n587 ) | ( n586 & n587 ) ;
  assign n589 = n588 ^ n389 ^ x6 ;
  assign n590 = n459 ^ x89 ^ 1'b0 ;
  assign n591 = n589 & ~n590 ;
  assign n592 = x99 & n402 ;
  assign n593 = ~x38 & n592 ;
  assign n594 = x88 & ~n417 ;
  assign n595 = ~x72 & n594 ;
  assign n596 = n595 ^ n236 ^ 1'b0 ;
  assign n597 = x68 & n596 ;
  assign n603 = x45 ^ x18 ^ 1'b0 ;
  assign n604 = ~n177 & n603 ;
  assign n598 = ~x69 & n179 ;
  assign n599 = n198 & n397 ;
  assign n600 = n599 ^ x10 ^ 1'b0 ;
  assign n601 = ( x0 & n180 ) | ( x0 & n600 ) | ( n180 & n600 ) ;
  assign n602 = n598 & ~n601 ;
  assign n605 = n604 ^ n602 ^ 1'b0 ;
  assign n611 = n301 ^ x86 ^ 1'b0 ;
  assign n606 = x14 & x16 ;
  assign n607 = ~x97 & n606 ;
  assign n608 = n344 ^ n232 ^ 1'b0 ;
  assign n609 = n607 | n608 ;
  assign n610 = n455 | n609 ;
  assign n612 = n611 ^ n610 ^ 1'b0 ;
  assign n613 = n574 ^ x46 ^ 1'b0 ;
  assign n614 = n613 ^ x116 ^ 1'b0 ;
  assign n615 = n614 ^ n585 ^ 1'b0 ;
  assign n616 = n152 ^ x79 ^ 1'b0 ;
  assign n617 = x45 & ~n377 ;
  assign n618 = ~n265 & n617 ;
  assign n619 = n186 | n450 ;
  assign n620 = n340 | n619 ;
  assign n621 = n620 ^ n188 ^ n154 ;
  assign n622 = ~n618 & n621 ;
  assign n623 = ~n560 & n622 ;
  assign n624 = x25 & ~n466 ;
  assign n625 = n355 & n624 ;
  assign n626 = x123 & ~n625 ;
  assign n627 = n626 ^ n414 ^ 1'b0 ;
  assign n628 = n244 ^ x61 ^ 1'b0 ;
  assign n629 = n147 & ~n377 ;
  assign n630 = n629 ^ n445 ^ 1'b0 ;
  assign n631 = n244 & n340 ;
  assign n632 = n631 ^ n283 ^ 1'b0 ;
  assign n633 = n330 & n366 ;
  assign n634 = n633 ^ n548 ^ n484 ;
  assign n635 = n456 ^ n376 ^ 1'b0 ;
  assign n636 = n327 & ~n635 ;
  assign n637 = n309 ^ n262 ^ 1'b0 ;
  assign n638 = x67 & ~n266 ;
  assign n639 = ~x53 & n638 ;
  assign n640 = n342 & ~n639 ;
  assign n641 = ( n402 & n637 ) | ( n402 & ~n640 ) | ( n637 & ~n640 ) ;
  assign n642 = ~n236 & n412 ;
  assign n647 = n490 ^ n278 ^ 1'b0 ;
  assign n648 = x102 & n647 ;
  assign n644 = n305 ^ x38 ^ 1'b0 ;
  assign n645 = n265 & ~n644 ;
  assign n643 = n493 ^ n296 ^ 1'b0 ;
  assign n646 = n645 ^ n643 ^ x3 ;
  assign n649 = n648 ^ n646 ^ n369 ;
  assign n651 = n389 | n489 ;
  assign n650 = n139 & ~n299 ;
  assign n652 = n651 ^ n650 ^ 1'b0 ;
  assign n653 = x77 | n278 ;
  assign n654 = n652 & ~n653 ;
  assign n655 = ~x99 & n654 ;
  assign n656 = n209 | n655 ;
  assign n657 = n374 ^ n293 ^ n275 ;
  assign n658 = n657 ^ n625 ^ n395 ;
  assign n659 = ~n545 & n658 ;
  assign n660 = n659 ^ n321 ^ 1'b0 ;
  assign n661 = ~n299 & n324 ;
  assign n662 = n661 ^ n415 ^ n218 ;
  assign n663 = n612 ^ x26 ^ 1'b0 ;
  assign n664 = n446 & n663 ;
  assign n665 = ~n335 & n643 ;
  assign n666 = ( ~x74 & n415 ) | ( ~x74 & n665 ) | ( n415 & n665 ) ;
  assign n667 = n666 ^ x106 ^ 1'b0 ;
  assign n668 = ~n278 & n288 ;
  assign n669 = n668 ^ n466 ^ 1'b0 ;
  assign n670 = ~n533 & n669 ;
  assign n671 = n670 ^ n433 ^ 1'b0 ;
  assign n672 = ( x37 & ~n359 ) | ( x37 & n518 ) | ( ~n359 & n518 ) ;
  assign n673 = x103 ^ x92 ^ 1'b0 ;
  assign n674 = n673 ^ n349 ^ x62 ;
  assign n675 = n129 ^ x93 ^ 1'b0 ;
  assign n676 = n234 & n307 ;
  assign n677 = x67 & n676 ;
  assign n678 = ~n607 & n651 ;
  assign n679 = n315 ^ n186 ^ 1'b0 ;
  assign n680 = n523 ^ n283 ^ n250 ;
  assign n681 = x46 ^ x20 ^ 1'b0 ;
  assign n682 = n681 ^ n359 ^ n194 ;
  assign n683 = n682 ^ n169 ^ 1'b0 ;
  assign n684 = x15 & ~n182 ;
  assign n685 = ~x23 & n684 ;
  assign n686 = n257 & ~n685 ;
  assign n687 = ~x33 & n686 ;
  assign n688 = ~n395 & n442 ;
  assign n689 = x33 & ~n293 ;
  assign n690 = ~n688 & n689 ;
  assign n691 = n605 ^ n487 ^ 1'b0 ;
  assign n692 = ~n690 & n691 ;
  assign n693 = x62 & ~n548 ;
  assign n694 = n693 ^ x12 ^ 1'b0 ;
  assign n695 = n402 ^ n217 ^ 1'b0 ;
  assign n696 = n695 ^ x38 ^ 1'b0 ;
  assign n697 = ~n694 & n696 ;
  assign n698 = x18 & ~n662 ;
  assign n699 = ~x35 & n698 ;
  assign n700 = n200 & ~n699 ;
  assign n701 = n700 ^ x10 ^ 1'b0 ;
  assign n702 = n229 ^ x84 ^ 1'b0 ;
  assign n703 = x31 & n279 ;
  assign n704 = ~n702 & n703 ;
  assign n705 = x37 & x50 ;
  assign n706 = n705 ^ n695 ^ 1'b0 ;
  assign n707 = n706 ^ n573 ^ 1'b0 ;
  assign n708 = ~n704 & n707 ;
  assign n709 = ( ~x77 & n208 ) | ( ~x77 & n273 ) | ( n208 & n273 ) ;
  assign n710 = ~n252 & n709 ;
  assign n712 = x79 & x120 ;
  assign n713 = n712 ^ n195 ^ 1'b0 ;
  assign n711 = n240 & n342 ;
  assign n714 = n713 ^ n711 ^ 1'b0 ;
  assign n715 = n479 ^ x20 ^ 1'b0 ;
  assign n716 = ~n499 & n715 ;
  assign n717 = x6 & n716 ;
  assign n718 = n452 & n717 ;
  assign n719 = n147 & n384 ;
  assign n720 = ~n186 & n719 ;
  assign n721 = n720 ^ x4 ^ 1'b0 ;
  assign n722 = n721 ^ n152 ^ 1'b0 ;
  assign n723 = ( ~n265 & n471 ) | ( ~n265 & n639 ) | ( n471 & n639 ) ;
  assign n724 = n723 ^ n653 ^ 1'b0 ;
  assign n725 = n374 & n724 ;
  assign n726 = x77 & ~n374 ;
  assign n729 = ( ~x47 & x97 ) | ( ~x47 & n137 ) | ( x97 & n137 ) ;
  assign n727 = x97 & n340 ;
  assign n728 = n727 ^ x72 ^ 1'b0 ;
  assign n730 = n729 ^ n728 ^ n156 ;
  assign n731 = x66 & ~n536 ;
  assign n732 = n731 ^ n379 ^ 1'b0 ;
  assign n733 = n397 & ~n511 ;
  assign n734 = n406 ^ n351 ^ 1'b0 ;
  assign n735 = n733 & ~n734 ;
  assign n736 = n735 ^ n166 ^ 1'b0 ;
  assign n737 = n169 | n736 ;
  assign n738 = n607 ^ n580 ^ x62 ;
  assign n739 = n509 | n681 ;
  assign n740 = n442 | n739 ;
  assign n741 = ~n487 & n740 ;
  assign n742 = ( ~x86 & n163 ) | ( ~x86 & n645 ) | ( n163 & n645 ) ;
  assign n743 = x26 & ~n490 ;
  assign n744 = n743 ^ n656 ^ 1'b0 ;
  assign n745 = n509 | n744 ;
  assign n746 = n701 ^ x62 ^ 1'b0 ;
  assign n747 = x69 & n267 ;
  assign n748 = x51 & ~n633 ;
  assign n749 = n748 ^ n642 ^ 1'b0 ;
  assign n750 = n749 ^ n144 ^ 1'b0 ;
  assign n751 = n477 | n750 ;
  assign n753 = x51 & ~x74 ;
  assign n752 = n379 & n695 ;
  assign n754 = n753 ^ n752 ^ 1'b0 ;
  assign n756 = n137 ^ x52 ^ 1'b0 ;
  assign n755 = n260 ^ x48 ^ 1'b0 ;
  assign n757 = n756 ^ n755 ^ 1'b0 ;
  assign n758 = ~n729 & n757 ;
  assign n759 = ~n613 & n620 ;
  assign n760 = n759 ^ n533 ^ 1'b0 ;
  assign n761 = n145 | n760 ;
  assign n762 = n761 ^ x55 ^ 1'b0 ;
  assign n763 = x41 ^ x16 ^ 1'b0 ;
  assign n764 = n763 ^ n345 ^ 1'b0 ;
  assign n765 = x6 | n764 ;
  assign n766 = ( ~n519 & n742 ) | ( ~n519 & n765 ) | ( n742 & n765 ) ;
  assign n767 = x102 & ~n607 ;
  assign n768 = n297 & ~n767 ;
  assign n769 = x97 & ~n392 ;
  assign n770 = ~n261 & n519 ;
  assign n771 = x17 | n749 ;
  assign n772 = n462 ^ x80 ^ 1'b0 ;
  assign n773 = x125 & ~n772 ;
  assign n774 = ( x95 & n484 ) | ( x95 & ~n773 ) | ( n484 & ~n773 ) ;
  assign n775 = n632 ^ n401 ^ 1'b0 ;
  assign n776 = n774 | n775 ;
  assign n777 = n776 ^ n718 ^ 1'b0 ;
  assign n778 = n234 & n452 ;
  assign n779 = ~n406 & n778 ;
  assign n780 = n440 | n472 ;
  assign n781 = n780 ^ x69 ^ 1'b0 ;
  assign n782 = n395 ^ n334 ^ x122 ;
  assign n783 = n345 ^ x73 ^ 1'b0 ;
  assign n784 = n782 & ~n783 ;
  assign n785 = n382 | n587 ;
  assign n786 = x110 | n785 ;
  assign n787 = ( n215 & n784 ) | ( n215 & n786 ) | ( n784 & n786 ) ;
  assign n788 = n144 & n787 ;
  assign n789 = n563 & ~n788 ;
  assign n794 = n231 ^ x37 ^ 1'b0 ;
  assign n795 = ( x127 & ~n134 ) | ( x127 & n794 ) | ( ~n134 & n794 ) ;
  assign n790 = n147 | n574 ;
  assign n791 = n790 ^ x71 ^ 1'b0 ;
  assign n792 = ~n477 & n791 ;
  assign n793 = n569 & n792 ;
  assign n796 = n795 ^ n793 ^ 1'b0 ;
  assign n797 = n713 ^ n636 ^ 1'b0 ;
  assign n798 = n129 ^ x50 ^ 1'b0 ;
  assign n799 = x29 & n798 ;
  assign n800 = n417 | n677 ;
  assign n801 = x35 | n800 ;
  assign n802 = ~n799 & n801 ;
  assign n803 = x40 & n165 ;
  assign n804 = x109 & ~n803 ;
  assign n805 = n275 & n804 ;
  assign n806 = ( ~x56 & n667 ) | ( ~x56 & n805 ) | ( n667 & n805 ) ;
  assign n807 = n702 & ~n806 ;
  assign n808 = n807 ^ n208 ^ 1'b0 ;
  assign n809 = n806 ^ n481 ^ 1'b0 ;
  assign n810 = x51 & n620 ;
  assign n811 = n261 ^ x123 ^ x54 ;
  assign n812 = x93 & n213 ;
  assign n813 = n266 & n812 ;
  assign n814 = n609 ^ x37 ^ 1'b0 ;
  assign n815 = ( n427 & n813 ) | ( n427 & ~n814 ) | ( n813 & ~n814 ) ;
  assign n816 = n210 | n541 ;
  assign n819 = n353 | n682 ;
  assign n820 = n819 ^ n347 ^ 1'b0 ;
  assign n817 = x74 | n509 ;
  assign n818 = n742 & n817 ;
  assign n821 = n820 ^ n818 ^ 1'b0 ;
  assign n822 = x127 & n208 ;
  assign n823 = x80 & ~n585 ;
  assign n824 = ( n630 & n740 ) | ( n630 & ~n823 ) | ( n740 & ~n823 ) ;
  assign n825 = n824 ^ x28 ^ 1'b0 ;
  assign n826 = n362 | n613 ;
  assign n827 = ( n363 & ~n398 ) | ( n363 & n826 ) | ( ~n398 & n826 ) ;
  assign n828 = n501 & n827 ;
  assign n829 = n828 ^ n334 ^ 1'b0 ;
  assign n832 = n477 ^ x34 ^ 1'b0 ;
  assign n833 = x38 & ~n209 ;
  assign n834 = x52 & n833 ;
  assign n835 = ~x91 & n834 ;
  assign n836 = ( n445 & ~n832 ) | ( n445 & n835 ) | ( ~n832 & n835 ) ;
  assign n830 = ~n154 & n674 ;
  assign n831 = n287 & n830 ;
  assign n837 = n836 ^ n831 ^ 1'b0 ;
  assign n838 = ~n829 & n837 ;
  assign n839 = n747 ^ n549 ^ 1'b0 ;
  assign n840 = ~n338 & n839 ;
  assign n841 = n267 ^ x106 ^ 1'b0 ;
  assign n842 = ( n675 & n730 ) | ( n675 & n754 ) | ( n730 & n754 ) ;
  assign n843 = n317 & ~n389 ;
  assign n844 = x118 & n371 ;
  assign n845 = x66 & n243 ;
  assign n846 = n845 ^ n709 ^ 1'b0 ;
  assign n847 = ~n487 & n846 ;
  assign n848 = n239 & ~n362 ;
  assign n849 = n848 ^ x25 ^ 1'b0 ;
  assign n850 = x102 & ~n849 ;
  assign n851 = ~n227 & n850 ;
  assign n852 = n851 ^ n639 ^ 1'b0 ;
  assign n853 = n730 ^ n134 ^ 1'b0 ;
  assign n854 = n733 ^ x1 ^ 1'b0 ;
  assign n855 = n542 ^ n265 ^ 1'b0 ;
  assign n856 = n855 ^ x25 ^ 1'b0 ;
  assign n857 = ( n648 & ~n854 ) | ( n648 & n856 ) | ( ~n854 & n856 ) ;
  assign n858 = n553 ^ n412 ^ 1'b0 ;
  assign n859 = n244 ^ n215 ^ n131 ;
  assign n860 = n859 ^ n491 ^ 1'b0 ;
  assign n861 = ( n137 & n620 ) | ( n137 & n687 ) | ( n620 & n687 ) ;
  assign n862 = n200 & ~n533 ;
  assign n863 = ~x43 & n862 ;
  assign n864 = n332 ^ n200 ^ 1'b0 ;
  assign n865 = ~n452 & n864 ;
  assign n866 = n607 | n865 ;
  assign n867 = n863 | n866 ;
  assign n868 = n327 ^ n283 ^ n148 ;
  assign n869 = ( x6 & ~n553 ) | ( x6 & n868 ) | ( ~n553 & n868 ) ;
  assign n870 = n167 | n869 ;
  assign n871 = n409 & ~n870 ;
  assign n873 = n849 ^ n574 ^ 1'b0 ;
  assign n874 = ~n147 & n873 ;
  assign n872 = n634 & n762 ;
  assign n875 = n874 ^ n872 ^ 1'b0 ;
  assign n876 = ( x10 & n486 ) | ( x10 & ~n556 ) | ( n486 & ~n556 ) ;
  assign n877 = x44 & ~n281 ;
  assign n878 = n877 ^ x6 ^ 1'b0 ;
  assign n880 = x34 & n129 ;
  assign n881 = ~x109 & n880 ;
  assign n879 = n403 & n448 ;
  assign n882 = n881 ^ n879 ^ n357 ;
  assign n883 = ( ~x14 & x111 ) | ( ~x14 & n144 ) | ( x111 & n144 ) ;
  assign n884 = n883 ^ n577 ^ 1'b0 ;
  assign n885 = n677 ^ n469 ^ 1'b0 ;
  assign n886 = ~n137 & n496 ;
  assign n887 = n224 | n886 ;
  assign n888 = n702 | n887 ;
  assign n889 = n531 & n888 ;
  assign n890 = ~x119 & n889 ;
  assign n891 = ~n355 & n397 ;
  assign n892 = ~n769 & n891 ;
  assign n893 = x29 & n735 ;
  assign n894 = ~x109 & n893 ;
  assign n895 = x79 & x94 ;
  assign n896 = n895 ^ n515 ^ 1'b0 ;
  assign n897 = n896 ^ n172 ^ 1'b0 ;
  assign n898 = n709 | n813 ;
  assign n899 = n446 & ~n481 ;
  assign n900 = n899 ^ n849 ^ 1'b0 ;
  assign n901 = ( x106 & n196 ) | ( x106 & n357 ) | ( n196 & n357 ) ;
  assign n902 = n901 ^ n377 ^ 1'b0 ;
  assign n903 = ~n900 & n902 ;
  assign n904 = n403 & n409 ;
  assign n905 = ~n903 & n904 ;
  assign n906 = n905 ^ n152 ^ 1'b0 ;
  assign n907 = n898 | n906 ;
  assign n908 = n213 & ~n395 ;
  assign n909 = ~x75 & n908 ;
  assign n910 = n909 ^ n719 ^ 1'b0 ;
  assign n911 = n402 & ~n910 ;
  assign n912 = n567 & n902 ;
  assign n913 = n912 ^ n258 ^ 1'b0 ;
  assign n914 = n809 ^ x69 ^ 1'b0 ;
  assign n915 = ~n381 & n914 ;
  assign n916 = ~n157 & n915 ;
  assign n917 = x29 & n569 ;
  assign n918 = n917 ^ x96 ^ 1'b0 ;
  assign n919 = n527 & n771 ;
  assign n920 = n919 ^ x34 ^ 1'b0 ;
  assign n921 = n657 | n920 ;
  assign n922 = n918 & ~n921 ;
  assign n923 = ~n147 & n866 ;
  assign n924 = n511 ^ n273 ^ 1'b0 ;
  assign n925 = x110 & n924 ;
  assign n926 = n925 ^ n897 ^ x105 ;
  assign n927 = x65 & ~n305 ;
  assign n928 = x103 ^ x47 ^ 1'b0 ;
  assign n929 = n928 ^ n462 ^ 1'b0 ;
  assign n930 = n927 & ~n929 ;
  assign n931 = n581 ^ n541 ^ 1'b0 ;
  assign n932 = n782 ^ n427 ^ 1'b0 ;
  assign n933 = x24 & n932 ;
  assign n934 = n931 & n933 ;
  assign n935 = n257 & ~n934 ;
  assign n936 = n234 & ~n478 ;
  assign n937 = n936 ^ n604 ^ 1'b0 ;
  assign n938 = n774 ^ x74 ^ 1'b0 ;
  assign n939 = n194 | n938 ;
  assign n940 = n515 ^ n401 ^ 1'b0 ;
  assign n941 = n682 | n940 ;
  assign n942 = n941 ^ n250 ^ 1'b0 ;
  assign n943 = n540 ^ n359 ^ 1'b0 ;
  assign n944 = n585 & ~n943 ;
  assign n945 = ~x58 & n944 ;
  assign n946 = n546 & ~n751 ;
  assign n947 = ~n435 & n946 ;
  assign n948 = n431 ^ n387 ^ 1'b0 ;
  assign n949 = ~n630 & n948 ;
  assign n950 = n184 & n949 ;
  assign n951 = n950 ^ n213 ^ 1'b0 ;
  assign n952 = n556 & ~n614 ;
  assign n953 = n529 ^ n166 ^ 1'b0 ;
  assign n954 = x55 & ~n277 ;
  assign n955 = n262 ^ x13 ^ 1'b0 ;
  assign n956 = x68 & n955 ;
  assign n957 = n133 & n956 ;
  assign n958 = ~n753 & n957 ;
  assign n959 = ( ~n445 & n549 ) | ( ~n445 & n958 ) | ( n549 & n958 ) ;
  assign n960 = n959 ^ n634 ^ 1'b0 ;
  assign n961 = n954 & ~n960 ;
  assign n962 = ~n953 & n961 ;
  assign n963 = x30 & x91 ;
  assign n964 = ~n882 & n963 ;
  assign n965 = n687 ^ n680 ^ 1'b0 ;
  assign n966 = n179 & n462 ;
  assign n967 = n639 & n966 ;
  assign n968 = n575 ^ n412 ^ 1'b0 ;
  assign n969 = n205 & ~n968 ;
  assign n970 = n234 & n969 ;
  assign n971 = n970 ^ n435 ^ 1'b0 ;
  assign n972 = n967 | n971 ;
  assign n973 = n777 & ~n972 ;
  assign n974 = n165 | n499 ;
  assign n975 = n974 ^ n719 ^ 1'b0 ;
  assign n976 = ~x58 & n163 ;
  assign n977 = ( ~n444 & n466 ) | ( ~n444 & n976 ) | ( n466 & n976 ) ;
  assign n978 = n977 ^ n765 ^ 1'b0 ;
  assign n979 = x29 & ~n978 ;
  assign n980 = ~x24 & n979 ;
  assign n981 = n690 ^ x114 ^ 1'b0 ;
  assign n982 = ~n980 & n981 ;
  assign n983 = n913 ^ n768 ^ 1'b0 ;
  assign n984 = n682 ^ x20 ^ 1'b0 ;
  assign n985 = n613 & ~n984 ;
  assign n986 = n985 ^ n888 ^ n204 ;
  assign n991 = x6 & ~n338 ;
  assign n992 = ~x31 & n991 ;
  assign n993 = ~n480 & n992 ;
  assign n987 = n303 ^ x82 ^ 1'b0 ;
  assign n988 = n384 ^ n194 ^ 1'b0 ;
  assign n989 = ( ~n257 & n987 ) | ( ~n257 & n988 ) | ( n987 & n988 ) ;
  assign n990 = ~n533 & n989 ;
  assign n994 = n993 ^ n990 ^ 1'b0 ;
  assign n995 = n994 ^ n330 ^ 1'b0 ;
  assign n996 = n628 ^ n525 ^ 1'b0 ;
  assign n997 = n240 & n996 ;
  assign n998 = n377 & ~n607 ;
  assign n999 = n863 ^ n143 ^ 1'b0 ;
  assign n1000 = x65 & ~n721 ;
  assign n1001 = n1000 ^ n759 ^ 1'b0 ;
  assign n1002 = n409 | n1001 ;
  assign n1003 = x30 | n1002 ;
  assign n1007 = x20 & n139 ;
  assign n1008 = ~n560 & n1007 ;
  assign n1004 = n309 ^ n157 ^ 1'b0 ;
  assign n1005 = n881 | n1004 ;
  assign n1006 = n911 & ~n1005 ;
  assign n1009 = n1008 ^ n1006 ^ 1'b0 ;
  assign n1010 = ~n521 & n1009 ;
  assign n1011 = n218 & n1010 ;
  assign n1012 = x23 & ~n303 ;
  assign n1013 = n1012 ^ n747 ^ n327 ;
  assign n1014 = x120 & ~n682 ;
  assign n1015 = ~x36 & n1014 ;
  assign n1016 = x23 & x69 ;
  assign n1017 = ~n791 & n1016 ;
  assign n1018 = n1017 ^ n327 ^ 1'b0 ;
  assign n1019 = n1015 | n1018 ;
  assign n1020 = n695 & ~n751 ;
  assign n1021 = n344 & n1020 ;
  assign n1022 = n217 & ~n1021 ;
  assign n1023 = ~n144 & n1022 ;
  assign n1024 = n1023 ^ x74 ^ 1'b0 ;
  assign n1025 = n885 ^ n435 ^ 1'b0 ;
  assign n1026 = ~n662 & n1025 ;
  assign n1027 = x65 & ~n166 ;
  assign n1028 = n1027 ^ n586 ^ x80 ;
  assign n1029 = n1028 ^ x54 ^ 1'b0 ;
  assign n1030 = n498 | n1029 ;
  assign n1031 = n342 & ~n1030 ;
  assign n1032 = n412 ^ n305 ^ 1'b0 ;
  assign n1033 = ~n477 & n1032 ;
  assign n1034 = ~n685 & n1033 ;
  assign n1035 = n1034 ^ n349 ^ 1'b0 ;
  assign n1036 = n255 & ~n484 ;
  assign n1037 = n468 & n1036 ;
  assign n1038 = ( ~n680 & n1035 ) | ( ~n680 & n1037 ) | ( n1035 & n1037 ) ;
  assign n1039 = n1015 ^ n753 ^ 1'b0 ;
  assign n1040 = ~x33 & n468 ;
  assign n1041 = n1039 ^ n460 ^ 1'b0 ;
  assign n1042 = n152 | n1041 ;
  assign n1043 = n675 ^ n539 ^ 1'b0 ;
  assign n1044 = n1027 | n1043 ;
  assign n1045 = n393 & n1044 ;
  assign n1046 = n933 ^ n358 ^ x42 ;
  assign n1047 = n583 ^ n296 ^ 1'b0 ;
  assign n1048 = n565 ^ x34 ^ 1'b0 ;
  assign n1049 = x116 & ~n1048 ;
  assign n1050 = n279 & ~n296 ;
  assign n1051 = n1050 ^ x52 ^ 1'b0 ;
  assign n1052 = n1049 & n1051 ;
  assign n1053 = ( ~x62 & n1015 ) | ( ~x62 & n1052 ) | ( n1015 & n1052 ) ;
  assign n1054 = n737 ^ x57 ^ 1'b0 ;
  assign n1055 = x6 & ~n448 ;
  assign n1056 = ~n133 & n1055 ;
  assign n1057 = n1056 ^ n607 ^ x107 ;
  assign n1058 = n665 ^ n601 ^ 1'b0 ;
  assign n1059 = n745 ^ n137 ^ 1'b0 ;
  assign n1060 = ~n452 & n1059 ;
  assign n1061 = n1060 ^ n238 ^ 1'b0 ;
  assign n1062 = n1054 & ~n1061 ;
  assign n1063 = n258 & ~n1037 ;
  assign n1064 = ~n332 & n1063 ;
  assign n1065 = ( ~n366 & n548 ) | ( ~n366 & n925 ) | ( n548 & n925 ) ;
  assign n1066 = n292 & ~n794 ;
  assign n1067 = n262 & n1066 ;
  assign n1068 = n281 | n292 ;
  assign n1069 = n448 | n952 ;
  assign n1070 = n1069 ^ n1015 ^ 1'b0 ;
  assign n1071 = ( x113 & n869 ) | ( x113 & ~n913 ) | ( n869 & ~n913 ) ;
  assign n1072 = n285 | n701 ;
  assign n1073 = n503 | n1072 ;
  assign n1077 = x21 | n177 ;
  assign n1074 = n279 ^ n244 ^ 1'b0 ;
  assign n1075 = n1074 ^ x111 ^ 1'b0 ;
  assign n1076 = n622 & ~n1075 ;
  assign n1078 = n1077 ^ n1076 ^ 1'b0 ;
  assign n1079 = ( x54 & n1008 ) | ( x54 & ~n1078 ) | ( n1008 & ~n1078 ) ;
  assign n1080 = n1073 & ~n1079 ;
  assign n1081 = ~n491 & n1080 ;
  assign n1082 = ~n362 & n833 ;
  assign n1083 = n335 & n1082 ;
  assign n1084 = n1076 & ~n1083 ;
  assign n1085 = n1084 ^ n840 ^ 1'b0 ;
  assign n1086 = n730 | n1085 ;
  assign n1087 = n1086 ^ n391 ^ 1'b0 ;
  assign n1088 = n930 & n1087 ;
  assign n1091 = n258 ^ x81 ^ 1'b0 ;
  assign n1092 = n585 & n1091 ;
  assign n1093 = n1092 ^ x72 ^ 1'b0 ;
  assign n1094 = n1093 ^ n855 ^ n687 ;
  assign n1089 = n411 ^ n395 ^ n265 ;
  assign n1090 = n371 & ~n1089 ;
  assign n1095 = n1094 ^ n1090 ^ 1'b0 ;
  assign n1096 = n1095 ^ n500 ^ n220 ;
  assign n1097 = x97 ^ x50 ^ 1'b0 ;
  assign n1098 = x54 ^ x53 ^ 1'b0 ;
  assign n1099 = x70 & n1098 ;
  assign n1100 = n1099 ^ n471 ^ 1'b0 ;
  assign n1101 = n1097 | n1100 ;
  assign n1102 = n1101 ^ n954 ^ 1'b0 ;
  assign n1103 = n305 & n767 ;
  assign n1104 = n1102 & ~n1103 ;
  assign n1105 = n236 & n1104 ;
  assign n1106 = x116 & x122 ;
  assign n1107 = ~x30 & n1106 ;
  assign n1108 = n612 & ~n1107 ;
  assign n1109 = n1108 ^ n621 ^ 1'b0 ;
  assign n1110 = x107 & ~n250 ;
  assign n1111 = n431 & n1110 ;
  assign n1112 = n244 & ~n278 ;
  assign n1113 = x105 ^ x101 ^ x33 ;
  assign n1114 = n1112 | n1113 ;
  assign n1115 = n305 & n611 ;
  assign n1116 = n1114 & ~n1115 ;
  assign n1117 = n1116 ^ n401 ^ 1'b0 ;
  assign n1118 = ( n583 & n960 ) | ( n583 & ~n994 ) | ( n960 & ~n994 ) ;
  assign n1119 = n607 ^ n541 ^ n344 ;
  assign n1120 = n1119 ^ n967 ^ x14 ;
  assign n1121 = n148 & ~n1027 ;
  assign n1122 = x52 & ~n1121 ;
  assign n1123 = ~n702 & n1122 ;
  assign n1124 = n472 & ~n478 ;
  assign n1125 = n1066 & ~n1124 ;
  assign n1126 = n409 & n1125 ;
  assign n1127 = n1123 | n1126 ;
  assign n1128 = n639 & ~n1127 ;
  assign n1129 = n215 | n1128 ;
  assign n1130 = n656 ^ n613 ^ 1'b0 ;
  assign n1131 = n543 ^ n533 ^ 1'b0 ;
  assign n1132 = n1130 & ~n1131 ;
  assign n1133 = n344 ^ x2 ^ 1'b0 ;
  assign n1134 = n1133 ^ x121 ^ 1'b0 ;
  assign n1135 = ( n255 & ~n266 ) | ( n255 & n1134 ) | ( ~n266 & n1134 ) ;
  assign n1136 = x65 & n975 ;
  assign n1137 = n1136 ^ n1078 ^ 1'b0 ;
  assign n1138 = n453 | n1001 ;
  assign n1139 = n674 ^ n575 ^ 1'b0 ;
  assign n1140 = x21 & n1139 ;
  assign n1142 = n529 ^ n150 ^ 1'b0 ;
  assign n1141 = n327 & ~n414 ;
  assign n1143 = n1142 ^ n1141 ^ 1'b0 ;
  assign n1144 = n1143 ^ x70 ^ 1'b0 ;
  assign n1145 = n262 & ~n1144 ;
  assign n1148 = x41 & n581 ;
  assign n1149 = n1148 ^ n384 ^ 1'b0 ;
  assign n1146 = x43 & ~n344 ;
  assign n1147 = n573 & n1146 ;
  assign n1150 = n1149 ^ n1147 ^ 1'b0 ;
  assign n1154 = ( x126 & ~n131 ) | ( x126 & n729 ) | ( ~n131 & n729 ) ;
  assign n1151 = x76 & ~n290 ;
  assign n1152 = ~n315 & n1151 ;
  assign n1153 = n364 | n1152 ;
  assign n1155 = n1154 ^ n1153 ^ 1'b0 ;
  assign n1156 = x73 & n1155 ;
  assign n1157 = n760 & n1156 ;
  assign n1158 = x117 ^ x22 ^ 1'b0 ;
  assign n1159 = ~n203 & n1158 ;
  assign n1161 = x25 & n249 ;
  assign n1162 = ~n265 & n1161 ;
  assign n1160 = x111 & n827 ;
  assign n1163 = n1162 ^ n1160 ^ 1'b0 ;
  assign n1164 = ( n534 & n1159 ) | ( n534 & ~n1163 ) | ( n1159 & ~n1163 ) ;
  assign n1165 = ~x68 & x80 ;
  assign n1166 = n1165 ^ n368 ^ 1'b0 ;
  assign n1167 = x42 & ~n573 ;
  assign n1168 = n1167 ^ n1035 ^ n138 ;
  assign n1169 = n1168 ^ n989 ^ n879 ;
  assign n1170 = ( ~n777 & n781 ) | ( ~n777 & n881 ) | ( n781 & n881 ) ;
  assign n1171 = x125 & n1170 ;
  assign n1172 = n1171 ^ n290 ^ 1'b0 ;
  assign n1173 = n1083 ^ n466 ^ 1'b0 ;
  assign n1174 = n195 & n1173 ;
  assign n1175 = n1174 ^ n1057 ^ n860 ;
  assign n1176 = n481 ^ n302 ^ 1'b0 ;
  assign n1177 = n177 & ~n1176 ;
  assign n1178 = n1177 ^ n548 ^ 1'b0 ;
  assign n1179 = n345 | n1178 ;
  assign n1180 = n483 | n675 ;
  assign n1181 = ~n381 & n885 ;
  assign n1182 = n1181 ^ n364 ^ 1'b0 ;
  assign n1183 = n952 ^ n632 ^ 1'b0 ;
  assign n1184 = ~n386 & n507 ;
  assign n1185 = n1184 ^ n918 ^ 1'b0 ;
  assign n1186 = n256 | n1185 ;
  assign n1187 = n557 ^ n437 ^ 1'b0 ;
  assign n1188 = n486 & n1187 ;
  assign n1189 = ~n1186 & n1188 ;
  assign n1190 = ~x37 & n279 ;
  assign n1191 = x121 & n900 ;
  assign n1192 = n1191 ^ n1067 ^ x113 ;
  assign n1193 = n1192 ^ n1121 ^ n573 ;
  assign n1194 = n517 | n855 ;
  assign n1195 = x75 | n1194 ;
  assign n1196 = x10 & x58 ;
  assign n1197 = ~n801 & n1196 ;
  assign n1198 = n827 ^ x27 ^ 1'b0 ;
  assign n1199 = n1197 | n1198 ;
  assign n1200 = ( n167 & n246 ) | ( n167 & n437 ) | ( n246 & n437 ) ;
  assign n1201 = ~n716 & n1200 ;
  assign n1202 = n1089 ^ n855 ^ 1'b0 ;
  assign n1203 = n1202 ^ n813 ^ 1'b0 ;
  assign n1204 = ~n1201 & n1203 ;
  assign n1205 = n1204 ^ n236 ^ 1'b0 ;
  assign n1206 = n1205 ^ n562 ^ n327 ;
  assign n1207 = n741 & n860 ;
  assign n1208 = n1207 ^ n709 ^ 1'b0 ;
  assign n1209 = ( n262 & n730 ) | ( n262 & n1017 ) | ( n730 & n1017 ) ;
  assign n1210 = ~n420 & n1209 ;
  assign n1211 = n959 & n1210 ;
  assign n1212 = ( ~n200 & n362 ) | ( ~n200 & n421 ) | ( n362 & n421 ) ;
  assign n1213 = n1212 ^ n673 ^ x121 ;
  assign n1214 = ~n421 & n738 ;
  assign n1215 = n1214 ^ n923 ^ 1'b0 ;
  assign n1216 = n988 ^ n721 ^ 1'b0 ;
  assign n1217 = n983 & ~n1216 ;
  assign n1218 = ~n995 & n1217 ;
  assign n1219 = n154 & n1218 ;
  assign n1220 = n144 & n695 ;
  assign n1221 = n1220 ^ x65 ^ 1'b0 ;
  assign n1222 = n1221 ^ n831 ^ 1'b0 ;
  assign n1223 = n977 | n1167 ;
  assign n1224 = n557 ^ x72 ^ 1'b0 ;
  assign n1227 = n419 | n881 ;
  assign n1228 = x109 | n1227 ;
  assign n1226 = x107 & ~n618 ;
  assign n1229 = n1228 ^ n1226 ^ 1'b0 ;
  assign n1225 = x111 ^ x74 ^ 1'b0 ;
  assign n1230 = n1229 ^ n1225 ^ 1'b0 ;
  assign n1231 = n1176 & n1230 ;
  assign n1232 = n633 | n763 ;
  assign n1233 = ( n692 & n978 ) | ( n692 & n1232 ) | ( n978 & n1232 ) ;
  assign n1234 = n614 ^ n258 ^ 1'b0 ;
  assign n1235 = x34 & n1234 ;
  assign n1236 = n246 & n905 ;
  assign n1237 = ~n797 & n1236 ;
  assign n1238 = n1056 ^ x0 ^ 1'b0 ;
  assign n1239 = n261 & ~n1238 ;
  assign n1240 = ~x43 & n523 ;
  assign n1241 = n945 & n1240 ;
  assign n1242 = n1239 & n1241 ;
  assign n1243 = ~x12 & n133 ;
  assign n1244 = n1243 ^ n1117 ^ 1'b0 ;
  assign n1245 = n437 ^ x58 ^ 1'b0 ;
  assign n1246 = n1245 ^ n763 ^ 1'b0 ;
  assign n1247 = n1015 | n1246 ;
  assign n1248 = ~x127 & n621 ;
  assign n1249 = n489 ^ n290 ^ 1'b0 ;
  assign n1250 = n692 & ~n1249 ;
  assign n1251 = n1248 & n1250 ;
  assign n1252 = n770 ^ x75 ^ 1'b0 ;
  assign n1253 = n1252 ^ n718 ^ 1'b0 ;
  assign n1254 = n1251 & ~n1253 ;
  assign n1257 = n803 ^ n690 ^ 1'b0 ;
  assign n1255 = x101 & ~n388 ;
  assign n1256 = n1255 ^ n896 ^ 1'b0 ;
  assign n1258 = n1257 ^ n1256 ^ n562 ;
  assign n1259 = n746 & ~n1237 ;
  assign n1260 = n773 & n1052 ;
  assign n1261 = n732 & n1260 ;
  assign n1262 = n1083 ^ n357 ^ 1'b0 ;
  assign n1263 = ~n894 & n1262 ;
  assign n1264 = n1263 ^ n622 ^ 1'b0 ;
  assign n1265 = n660 ^ n420 ^ 1'b0 ;
  assign n1266 = x55 & n1265 ;
  assign n1267 = x89 & ~n718 ;
  assign n1268 = n415 & n1267 ;
  assign n1269 = n269 & ~n1268 ;
  assign n1270 = n1143 & n1269 ;
  assign n1271 = n437 & ~n1270 ;
  assign n1272 = n620 & n1088 ;
  assign n1273 = ~x103 & n1272 ;
  assign n1274 = x77 & n1204 ;
  assign n1275 = n455 & n1274 ;
  assign n1276 = n1275 ^ x102 ^ 1'b0 ;
  assign n1278 = n174 | n709 ;
  assign n1279 = n307 & ~n1278 ;
  assign n1277 = n359 ^ n275 ^ n157 ;
  assign n1280 = n1279 ^ n1277 ^ 1'b0 ;
  assign n1281 = n420 | n1280 ;
  assign n1282 = n227 & ~n1281 ;
  assign n1283 = n301 & n1282 ;
  assign n1284 = n472 | n1283 ;
  assign n1285 = n1284 ^ x84 ^ 1'b0 ;
  assign n1288 = n202 | n499 ;
  assign n1289 = n661 | n1288 ;
  assign n1286 = ~n254 & n546 ;
  assign n1287 = n1286 ^ n649 ^ 1'b0 ;
  assign n1290 = n1289 ^ n1287 ^ 1'b0 ;
  assign n1291 = n569 & ~n1290 ;
  assign n1292 = n323 & n1291 ;
  assign n1293 = ~n1285 & n1292 ;
  assign n1294 = n844 & ~n1293 ;
  assign n1295 = ~n1182 & n1294 ;
  assign n1296 = n628 & ~n883 ;
  assign n1301 = n567 ^ n400 ^ n386 ;
  assign n1299 = x75 & ~n154 ;
  assign n1300 = n1299 ^ x54 ^ 1'b0 ;
  assign n1302 = n1301 ^ n1300 ^ 1'b0 ;
  assign n1303 = ~n726 & n1302 ;
  assign n1297 = n393 & n543 ;
  assign n1298 = n1297 ^ n860 ^ 1'b0 ;
  assign n1304 = n1303 ^ n1298 ^ n677 ;
  assign n1305 = n258 & n515 ;
  assign n1306 = n760 & n1305 ;
  assign n1307 = n878 ^ n393 ^ 1'b0 ;
  assign n1308 = n1142 & n1307 ;
  assign n1309 = n827 ^ n673 ^ 1'b0 ;
  assign n1310 = n1309 ^ n894 ^ 1'b0 ;
  assign n1311 = n1308 & n1310 ;
  assign n1312 = n161 ^ x61 ^ 1'b0 ;
  assign n1313 = ~n643 & n1312 ;
  assign n1314 = n847 & n1313 ;
  assign n1315 = n1314 ^ n195 ^ 1'b0 ;
  assign n1316 = n1005 ^ n192 ^ 1'b0 ;
  assign n1317 = n565 | n1316 ;
  assign n1318 = n150 | n1317 ;
  assign n1319 = n1318 ^ n897 ^ 1'b0 ;
  assign n1320 = ~n1124 & n1319 ;
  assign n1321 = ~x108 & n1320 ;
  assign n1322 = n1257 ^ x90 ^ 1'b0 ;
  assign n1323 = n620 & n1289 ;
  assign n1324 = ~n446 & n1323 ;
  assign n1325 = n1324 ^ n934 ^ 1'b0 ;
  assign n1326 = n336 & ~n950 ;
  assign n1327 = ~n1325 & n1326 ;
  assign n1328 = n1067 & ~n1327 ;
  assign n1329 = ~n1322 & n1328 ;
  assign n1330 = n1277 ^ n747 ^ n382 ;
  assign n1331 = n133 & n371 ;
  assign n1332 = ~x83 & x112 ;
  assign n1333 = ~n1331 & n1332 ;
  assign n1335 = x19 & ~n1083 ;
  assign n1336 = ~x47 & n1335 ;
  assign n1334 = n476 & ~n863 ;
  assign n1337 = n1336 ^ n1334 ^ 1'b0 ;
  assign n1338 = n1337 ^ n922 ^ 1'b0 ;
  assign n1339 = n1338 ^ n379 ^ 1'b0 ;
  assign n1340 = n1133 & n1339 ;
  assign n1341 = n831 ^ n791 ^ 1'b0 ;
  assign n1342 = n621 ^ n215 ^ 1'b0 ;
  assign n1343 = x13 & ~n412 ;
  assign n1344 = x79 ^ x6 ^ 1'b0 ;
  assign n1345 = n1343 & n1344 ;
  assign n1346 = ~x80 & n1345 ;
  assign n1347 = x39 & ~n272 ;
  assign n1348 = n1346 & n1347 ;
  assign n1349 = n478 | n1348 ;
  assign n1350 = n562 | n1349 ;
  assign n1351 = n1342 & ~n1350 ;
  assign n1352 = ~n174 & n1343 ;
  assign n1353 = n995 & n1352 ;
  assign n1354 = n640 ^ n393 ^ n389 ;
  assign n1355 = ( x38 & n472 ) | ( x38 & n1354 ) | ( n472 & n1354 ) ;
  assign n1356 = n1066 & n1355 ;
  assign n1357 = n1356 ^ n215 ^ 1'b0 ;
  assign n1358 = n1357 ^ n589 ^ 1'b0 ;
  assign n1359 = ~n1353 & n1358 ;
  assign n1360 = n1107 ^ n190 ^ 1'b0 ;
  assign n1361 = x36 & ~n1360 ;
  assign n1362 = n937 ^ n701 ^ 1'b0 ;
  assign n1363 = n1361 & ~n1362 ;
  assign n1364 = x109 & n435 ;
  assign n1365 = n1364 ^ n275 ^ 1'b0 ;
  assign n1366 = n496 & ~n1105 ;
  assign n1367 = n1366 ^ n814 ^ 1'b0 ;
  assign n1368 = n1174 ^ n297 ^ 1'b0 ;
  assign n1369 = ~n836 & n1368 ;
  assign n1370 = ( n231 & n751 ) | ( n231 & n1369 ) | ( n751 & n1369 ) ;
  assign n1371 = n763 ^ n272 ^ 1'b0 ;
  assign n1372 = n278 | n1371 ;
  assign n1373 = n1092 & ~n1372 ;
  assign n1374 = n1011 & n1373 ;
  assign n1375 = n381 | n960 ;
  assign n1376 = x60 | n1375 ;
  assign n1377 = n1376 ^ n1115 ^ 1'b0 ;
  assign n1378 = ( ~n417 & n459 ) | ( ~n417 & n1289 ) | ( n459 & n1289 ) ;
  assign n1379 = n349 & ~n863 ;
  assign n1380 = n779 & n1379 ;
  assign n1385 = x112 ^ x97 ^ 1'b0 ;
  assign n1381 = n196 & ~n1035 ;
  assign n1382 = n1381 ^ n620 ^ 1'b0 ;
  assign n1383 = n1044 & ~n1382 ;
  assign n1384 = n1067 & ~n1383 ;
  assign n1386 = n1385 ^ n1384 ^ 1'b0 ;
  assign n1387 = n1291 ^ n649 ^ 1'b0 ;
  assign n1388 = ~n415 & n1387 ;
  assign n1389 = n288 & n1388 ;
  assign n1390 = ~x83 & n1389 ;
  assign n1391 = n1191 & n1390 ;
  assign n1392 = n430 ^ x52 ^ 1'b0 ;
  assign n1393 = n1027 ^ n888 ^ n745 ;
  assign n1394 = n210 & n671 ;
  assign n1395 = n476 ^ x126 ^ 1'b0 ;
  assign n1396 = n580 | n1395 ;
  assign n1397 = x100 & n753 ;
  assign n1398 = n1397 ^ n336 ^ 1'b0 ;
  assign n1399 = ( x8 & x96 ) | ( x8 & ~x110 ) | ( x96 & ~x110 ) ;
  assign n1400 = ~n542 & n1399 ;
  assign n1401 = n1400 ^ n494 ^ 1'b0 ;
  assign n1402 = n440 | n460 ;
  assign n1403 = n813 ^ n180 ^ 1'b0 ;
  assign n1404 = ~n1402 & n1403 ;
  assign n1405 = n175 & n1404 ;
  assign n1406 = n728 & ~n1324 ;
  assign n1407 = n660 | n1406 ;
  assign n1408 = n766 & ~n1407 ;
  assign n1409 = n671 & ~n1408 ;
  assign n1410 = ~x71 & n1409 ;
  assign n1411 = n1410 ^ n1120 ^ 1'b0 ;
  assign n1412 = n484 ^ n477 ^ 1'b0 ;
  assign n1413 = x28 & ~n978 ;
  assign n1414 = n680 & n1413 ;
  assign n1415 = n753 & ~n1414 ;
  assign n1416 = n976 & n1415 ;
  assign n1417 = x1 & n138 ;
  assign n1418 = n1417 ^ n523 ^ 1'b0 ;
  assign n1419 = ( n1167 & n1281 ) | ( n1167 & n1418 ) | ( n1281 & n1418 ) ;
  assign n1420 = n545 | n1419 ;
  assign n1421 = n1330 & n1420 ;
  assign n1424 = x127 & n803 ;
  assign n1425 = ( ~n143 & n419 ) | ( ~n143 & n1424 ) | ( n419 & n1424 ) ;
  assign n1423 = x42 & n589 ;
  assign n1426 = n1425 ^ n1423 ^ 1'b0 ;
  assign n1427 = n1426 ^ x98 ^ 1'b0 ;
  assign n1428 = n1229 ^ n278 ^ 1'b0 ;
  assign n1429 = n1427 & n1428 ;
  assign n1422 = ( ~x38 & n491 ) | ( ~x38 & n1204 ) | ( n491 & n1204 ) ;
  assign n1430 = n1429 ^ n1422 ^ 1'b0 ;
  assign n1431 = ~n1211 & n1430 ;
  assign n1432 = n147 | n499 ;
  assign n1433 = n902 ^ n200 ^ 1'b0 ;
  assign n1434 = n1078 & n1433 ;
  assign n1435 = n324 & n1434 ;
  assign n1436 = n1398 ^ x85 ^ 1'b0 ;
  assign n1437 = n740 & ~n1436 ;
  assign n1439 = n753 ^ n400 ^ 1'b0 ;
  assign n1438 = n521 ^ x57 ^ 1'b0 ;
  assign n1440 = n1439 ^ n1438 ^ 1'b0 ;
  assign n1441 = x15 ^ x3 ^ 1'b0 ;
  assign n1442 = ~n1097 & n1441 ;
  assign n1443 = n171 | n243 ;
  assign n1444 = x22 | n1443 ;
  assign n1445 = ~n1089 & n1444 ;
  assign n1446 = ~n1442 & n1445 ;
  assign n1447 = n1331 ^ n479 ^ 1'b0 ;
  assign n1448 = n1446 | n1447 ;
  assign n1449 = n1448 ^ n169 ^ 1'b0 ;
  assign n1450 = ~n1083 & n1449 ;
  assign n1451 = x63 & n1450 ;
  assign n1452 = ~n1188 & n1451 ;
  assign n1453 = n279 & n778 ;
  assign n1454 = n1453 ^ n1088 ^ 1'b0 ;
  assign n1455 = ( n404 & ~n605 ) | ( n404 & n1454 ) | ( ~n605 & n1454 ) ;
  assign n1460 = n227 ^ x104 ^ 1'b0 ;
  assign n1461 = x12 & n1460 ;
  assign n1462 = n713 ^ n428 ^ 1'b0 ;
  assign n1463 = n1461 & ~n1462 ;
  assign n1464 = ( x90 & n548 ) | ( x90 & n1463 ) | ( n548 & n1463 ) ;
  assign n1456 = n539 ^ n182 ^ 1'b0 ;
  assign n1457 = ~n147 & n1456 ;
  assign n1458 = n1457 ^ n695 ^ n324 ;
  assign n1459 = ~n252 & n1458 ;
  assign n1465 = n1464 ^ n1459 ^ 1'b0 ;
  assign n1466 = x98 & n430 ;
  assign n1467 = ~n359 & n1466 ;
  assign n1468 = n293 | n1467 ;
  assign n1469 = n1008 & ~n1468 ;
  assign n1470 = n843 ^ x99 ^ 1'b0 ;
  assign n1471 = ~x31 & n882 ;
  assign n1472 = n645 ^ n198 ^ 1'b0 ;
  assign n1473 = ~n881 & n1472 ;
  assign n1474 = ~n709 & n1473 ;
  assign n1475 = n1474 ^ n1174 ^ 1'b0 ;
  assign n1476 = n612 & n1475 ;
  assign n1485 = n225 ^ x21 ^ x3 ;
  assign n1479 = n208 & ~n252 ;
  assign n1480 = n756 | n1479 ;
  assign n1481 = n138 | n1480 ;
  assign n1482 = n1481 ^ n706 ^ 1'b0 ;
  assign n1483 = n728 | n1482 ;
  assign n1477 = n1049 & n1424 ;
  assign n1478 = ~x1 & n1477 ;
  assign n1484 = n1483 ^ n1478 ^ x48 ;
  assign n1486 = n1485 ^ n1484 ^ 1'b0 ;
  assign n1487 = ~n992 & n1486 ;
  assign n1488 = x16 & ~x33 ;
  assign n1489 = n133 & ~n1488 ;
  assign n1490 = n1488 | n1489 ;
  assign n1491 = n721 & n1490 ;
  assign n1492 = n1421 ^ n260 ^ 1'b0 ;
  assign n1493 = ~n131 & n1492 ;
  assign n1494 = x6 & ~n150 ;
  assign n1495 = n1494 ^ n621 ^ 1'b0 ;
  assign n1496 = n1495 ^ n479 ^ 1'b0 ;
  assign n1497 = n433 | n1496 ;
  assign n1498 = ~n1137 & n1497 ;
  assign n1499 = x121 & ~n1097 ;
  assign n1500 = n1499 ^ n205 ^ 1'b0 ;
  assign n1501 = n565 | n1500 ;
  assign n1502 = n1498 & ~n1501 ;
  assign n1503 = ~n637 & n1424 ;
  assign n1504 = ~n186 & n827 ;
  assign n1505 = ~x58 & n1504 ;
  assign n1506 = n676 & ~n1505 ;
  assign n1507 = n1506 ^ n805 ^ 1'b0 ;
  assign n1508 = n843 & n1464 ;
  assign n1509 = ~x90 & n1508 ;
  assign n1510 = x118 & n200 ;
  assign n1511 = n1510 ^ n740 ^ 1'b0 ;
  assign n1512 = ( x50 & ~x81 ) | ( x50 & n598 ) | ( ~x81 & n598 ) ;
  assign n1513 = n1439 & n1512 ;
  assign n1514 = ~x90 & n1513 ;
  assign n1515 = n144 & n721 ;
  assign n1516 = x55 & n1230 ;
  assign n1517 = ~n832 & n1516 ;
  assign n1518 = n400 & ~n710 ;
  assign n1519 = n801 & ~n1243 ;
  assign n1520 = ~n138 & n1519 ;
  assign n1521 = n147 & ~n1520 ;
  assign n1522 = n1521 ^ n1489 ^ 1'b0 ;
  assign n1523 = n973 & ~n1522 ;
  assign n1524 = ~x70 & n161 ;
  assign n1525 = n222 ^ n200 ^ 1'b0 ;
  assign n1526 = n243 | n1525 ;
  assign n1527 = n1526 ^ n688 ^ 1'b0 ;
  assign n1528 = n1527 ^ n371 ^ 1'b0 ;
  assign n1529 = n911 & ~n1528 ;
  assign n1530 = n1529 ^ x75 ^ 1'b0 ;
  assign n1531 = n687 | n1530 ;
  assign n1532 = n1344 ^ n1092 ^ 1'b0 ;
  assign n1533 = ~n208 & n557 ;
  assign n1534 = ~n1532 & n1533 ;
  assign n1535 = ~n374 & n479 ;
  assign n1536 = x72 & n1535 ;
  assign n1537 = n190 & ~n546 ;
  assign n1538 = n823 | n1537 ;
  assign n1539 = n157 & n486 ;
  assign n1540 = n1538 & n1539 ;
  assign n1541 = x7 | n194 ;
  assign n1542 = ~n978 & n1432 ;
  assign n1543 = ~n1541 & n1542 ;
  assign n1548 = n871 ^ x18 ^ 1'b0 ;
  assign n1549 = n363 | n1548 ;
  assign n1544 = n695 & n1424 ;
  assign n1545 = ~n1325 & n1544 ;
  assign n1546 = n1243 ^ x20 ^ 1'b0 ;
  assign n1547 = n1545 | n1546 ;
  assign n1550 = n1549 ^ n1547 ^ 1'b0 ;
  assign n1551 = x78 & ~n760 ;
  assign n1552 = n302 & n1551 ;
  assign n1555 = n1149 ^ n947 ^ n414 ;
  assign n1553 = ( n148 & ~n246 ) | ( n148 & n620 ) | ( ~n246 & n620 ) ;
  assign n1554 = x34 & ~n1553 ;
  assign n1556 = n1555 ^ n1554 ^ 1'b0 ;
  assign n1557 = x16 & n292 ;
  assign n1558 = n1557 ^ n815 ^ 1'b0 ;
  assign n1559 = n781 & n1558 ;
  assign n1560 = ~n1507 & n1559 ;
  assign n1561 = n989 ^ n756 ^ 1'b0 ;
  assign n1562 = n716 & ~n1561 ;
  assign n1563 = n1562 ^ n976 ^ n475 ;
  assign n1564 = n672 ^ x80 ^ 1'b0 ;
  assign n1565 = n161 & n1564 ;
  assign n1566 = ( x74 & n694 ) | ( x74 & ~n1565 ) | ( n694 & ~n1565 ) ;
  assign n1567 = n1021 ^ n909 ^ n156 ;
  assign n1568 = n1300 ^ x47 ^ 1'b0 ;
  assign n1569 = n1567 & ~n1568 ;
  assign n1570 = ~n462 & n1064 ;
  assign n1571 = n1570 ^ n157 ^ 1'b0 ;
  assign n1572 = n632 & n1571 ;
  assign n1573 = n334 & ~n1107 ;
  assign n1574 = ~n827 & n1573 ;
  assign n1575 = x75 & n381 ;
  assign n1577 = n1361 ^ n632 ^ 1'b0 ;
  assign n1578 = ~n344 & n1577 ;
  assign n1576 = n249 & n587 ;
  assign n1579 = n1578 ^ n1576 ^ 1'b0 ;
  assign n1580 = n1575 & ~n1579 ;
  assign n1581 = n1574 & n1580 ;
  assign n1582 = n976 ^ n257 ^ 1'b0 ;
  assign n1583 = n1581 & ~n1582 ;
  assign n1584 = n527 ^ n180 ^ 1'b0 ;
  assign n1585 = n683 | n1584 ;
  assign n1586 = n475 | n805 ;
  assign n1587 = n1586 ^ n826 ^ n319 ;
  assign n1588 = ( n769 & ~n1291 ) | ( n769 & n1587 ) | ( ~n1291 & n1587 ) ;
  assign n1589 = n1588 ^ n630 ^ 1'b0 ;
  assign n1590 = ~n1585 & n1589 ;
  assign n1591 = n498 | n849 ;
  assign n1592 = n1591 ^ n1488 ^ 1'b0 ;
  assign n1593 = n1592 ^ n1497 ^ 1'b0 ;
  assign n1594 = n1324 | n1593 ;
  assign n1595 = n1165 ^ n477 ^ 1'b0 ;
  assign n1596 = n294 & ~n1595 ;
  assign n1597 = n1596 ^ x16 ^ 1'b0 ;
  assign n1598 = n476 | n1083 ;
  assign n1599 = n1598 ^ n311 ^ 1'b0 ;
  assign n1600 = n1132 & n1594 ;
  assign n1601 = ( n702 & n1003 ) | ( n702 & ~n1241 ) | ( n1003 & ~n1241 ) ;
  assign n1602 = n1601 ^ n1365 ^ 1'b0 ;
  assign n1603 = ~n452 & n1264 ;
  assign n1604 = x4 & x103 ;
  assign n1605 = n1604 ^ x34 ^ 1'b0 ;
  assign n1606 = n1060 | n1605 ;
  assign n1607 = n1606 ^ n1579 ^ 1'b0 ;
  assign n1608 = n1313 & ~n1607 ;
  assign n1609 = ~n710 & n1319 ;
  assign n1610 = x121 & n1609 ;
  assign n1611 = ~x26 & n1610 ;
  assign n1612 = n1611 ^ n1086 ^ 1'b0 ;
  assign n1614 = ( n652 & ~n730 ) | ( n652 & n1457 ) | ( ~n730 & n1457 ) ;
  assign n1613 = ~n534 & n695 ;
  assign n1615 = n1614 ^ n1613 ^ 1'b0 ;
  assign n1616 = n1615 ^ n330 ^ 1'b0 ;
  assign n1617 = ~n489 & n722 ;
  assign n1618 = n911 ^ n266 ^ 1'b0 ;
  assign n1619 = n1617 | n1618 ;
  assign n1621 = ( n649 & ~n833 ) | ( n649 & n915 ) | ( ~n833 & n915 ) ;
  assign n1620 = n1221 ^ n639 ^ 1'b0 ;
  assign n1622 = n1621 ^ n1620 ^ 1'b0 ;
  assign n1623 = n1619 | n1622 ;
  assign n1624 = n1056 ^ n994 ^ 1'b0 ;
  assign n1625 = n456 & n1624 ;
  assign n1626 = x1 & n1489 ;
  assign n1627 = n290 & n1626 ;
  assign n1628 = n595 | n1627 ;
  assign n1629 = n1628 ^ n373 ^ 1'b0 ;
  assign n1630 = x20 & n543 ;
  assign n1631 = ~x97 & n1630 ;
  assign n1632 = n1631 ^ n1518 ^ 1'b0 ;
  assign n1633 = n252 & ~n994 ;
  assign n1634 = x89 | n704 ;
  assign n1635 = x106 | n1027 ;
  assign n1636 = n1256 & ~n1635 ;
  assign n1637 = n204 & n1636 ;
  assign n1638 = ( n549 & n1372 ) | ( n549 & ~n1637 ) | ( n1372 & ~n1637 ) ;
  assign n1639 = ( ~x64 & n165 ) | ( ~x64 & n1638 ) | ( n165 & n1638 ) ;
  assign n1640 = n1639 ^ n1467 ^ 1'b0 ;
  assign n1641 = ~n1634 & n1640 ;
  assign n1642 = n1641 ^ n721 ^ n543 ;
  assign n1643 = n491 & ~n726 ;
  assign n1644 = n719 & n1256 ;
  assign n1645 = ~n1643 & n1644 ;
  assign n1646 = x66 | n531 ;
  assign n1647 = n1642 & n1646 ;
  assign n1648 = ~n499 & n1277 ;
  assign n1649 = n1648 ^ n591 ^ 1'b0 ;
  assign n1650 = n1649 ^ x44 ^ 1'b0 ;
  assign n1651 = x45 & ~n1650 ;
  assign n1652 = n175 & ~n1651 ;
  assign n1653 = x72 & ~n625 ;
  assign n1654 = n1653 ^ n1109 ^ 1'b0 ;
  assign n1655 = x13 & n1439 ;
  assign n1656 = n1655 ^ x81 ^ 1'b0 ;
  assign n1657 = n1510 & n1656 ;
  assign n1658 = ( n200 & ~n376 ) | ( n200 & n1243 ) | ( ~n376 & n1243 ) ;
  assign n1659 = n615 | n1496 ;
  assign n1660 = n1658 | n1659 ;
  assign n1661 = n423 & ~n1660 ;
  assign n1662 = ( n374 & ~n879 ) | ( n374 & n1661 ) | ( ~n879 & n1661 ) ;
  assign n1663 = n1632 | n1662 ;
  assign n1664 = n1663 ^ n556 ^ 1'b0 ;
  assign n1665 = n143 & ~n324 ;
  assign n1666 = n1367 & n1665 ;
  assign n1667 = n1558 ^ n823 ^ 1'b0 ;
  assign n1668 = n1553 | n1667 ;
  assign n1669 = n198 & ~n577 ;
  assign n1670 = n836 & n1669 ;
  assign n1671 = n1089 ^ n147 ^ 1'b0 ;
  assign n1672 = n1670 | n1671 ;
  assign n1673 = n232 ^ x125 ^ 1'b0 ;
  assign n1674 = ~n1672 & n1673 ;
  assign n1675 = x108 ^ x31 ^ 1'b0 ;
  assign n1676 = n902 & n1675 ;
  assign n1678 = n826 & ~n859 ;
  assign n1679 = n1678 ^ n129 ^ 1'b0 ;
  assign n1680 = n541 | n1679 ;
  assign n1677 = n294 & n1183 ;
  assign n1681 = n1680 ^ n1677 ^ 1'b0 ;
  assign n1682 = n593 ^ n254 ^ 1'b0 ;
  assign n1683 = n1256 & ~n1682 ;
  assign n1684 = ~n935 & n1683 ;
  assign n1685 = n148 & n1684 ;
  assign n1686 = n1685 ^ n486 ^ n353 ;
  assign n1687 = ~x58 & n491 ;
  assign n1688 = n667 | n892 ;
  assign n1689 = ( n1382 & ~n1687 ) | ( n1382 & n1688 ) | ( ~n1687 & n1688 ) ;
  assign n1691 = n791 ^ x119 ^ 1'b0 ;
  assign n1692 = n1691 ^ n941 ^ x60 ;
  assign n1690 = x102 & n244 ;
  assign n1693 = n1692 ^ n1690 ^ 1'b0 ;
  assign n1694 = x110 & ~n903 ;
  assign n1695 = ~n1558 & n1694 ;
  assign n1696 = x102 ^ x27 ^ 1'b0 ;
  assign n1697 = n632 & n1696 ;
  assign n1698 = x101 & n1697 ;
  assign n1699 = n560 & n1241 ;
  assign n1700 = ~n1698 & n1699 ;
  assign n1707 = x73 & ~n1229 ;
  assign n1708 = n859 & n1707 ;
  assign n1709 = n1708 ^ n781 ^ 1'b0 ;
  assign n1710 = n1638 & ~n1709 ;
  assign n1701 = n679 ^ x42 ^ 1'b0 ;
  assign n1702 = n521 | n1035 ;
  assign n1703 = n1701 & ~n1702 ;
  assign n1704 = n139 & ~n1703 ;
  assign n1705 = n1704 ^ n379 ^ 1'b0 ;
  assign n1706 = x21 & ~n1705 ;
  assign n1711 = n1710 ^ n1706 ^ 1'b0 ;
  assign n1712 = n549 ^ n139 ^ 1'b0 ;
  assign n1713 = n273 & n1712 ;
  assign n1714 = ~n163 & n1713 ;
  assign n1715 = n1179 ^ n709 ^ 1'b0 ;
  assign n1716 = ~n1714 & n1715 ;
  assign n1717 = n653 ^ x46 ^ 1'b0 ;
  assign n1718 = n283 | n1717 ;
  assign n1719 = n157 & ~n1718 ;
  assign n1720 = n1313 ^ n1250 ^ 1'b0 ;
  assign n1721 = x21 & ~n1627 ;
  assign n1722 = n1721 ^ x17 ^ 1'b0 ;
  assign n1723 = n437 & n479 ;
  assign n1724 = n820 | n1329 ;
  assign n1725 = n1724 ^ n180 ^ 1'b0 ;
  assign n1726 = n323 | n1013 ;
  assign n1727 = n1726 ^ n699 ^ 1'b0 ;
  assign n1728 = n531 & ~n1727 ;
  assign n1731 = n1047 ^ n775 ^ 1'b0 ;
  assign n1732 = n154 | n1731 ;
  assign n1729 = ~x105 & n632 ;
  assign n1730 = n987 & ~n1729 ;
  assign n1733 = n1732 ^ n1730 ^ 1'b0 ;
  assign n1734 = n1596 ^ n616 ^ 1'b0 ;
  assign n1735 = n1354 & n1734 ;
  assign n1736 = n993 ^ x5 ^ 1'b0 ;
  assign n1737 = n195 & n1736 ;
  assign n1738 = ( n976 & n1735 ) | ( n976 & n1737 ) | ( n1735 & n1737 ) ;
  assign n1739 = n1733 & n1738 ;
  assign n1740 = n789 & n1739 ;
  assign n1741 = n1467 ^ n871 ^ 1'b0 ;
  assign n1742 = n1100 ^ n472 ^ 1'b0 ;
  assign n1743 = n1742 ^ x44 ^ 1'b0 ;
  assign n1744 = ~n303 & n781 ;
  assign n1745 = n1744 ^ n1448 ^ 1'b0 ;
  assign n1746 = n1074 ^ n738 ^ 1'b0 ;
  assign n1747 = n1745 & ~n1746 ;
  assign n1748 = ~n1681 & n1687 ;
  assign n1749 = n826 ^ n601 ^ 1'b0 ;
  assign n1750 = n713 | n1749 ;
  assign n1751 = n881 & ~n1750 ;
  assign n1752 = ~n959 & n1751 ;
  assign n1753 = n1205 & n1752 ;
  assign n1754 = n478 ^ n445 ^ x95 ;
  assign n1755 = ( n518 & n1753 ) | ( n518 & n1754 ) | ( n1753 & n1754 ) ;
  assign n1756 = ~n1021 & n1166 ;
  assign n1757 = x80 & ~n673 ;
  assign n1758 = n1757 ^ n293 ^ x79 ;
  assign n1759 = n930 & ~n1758 ;
  assign n1760 = x82 & n1062 ;
  assign n1761 = n1760 ^ n794 ^ 1'b0 ;
  assign n1762 = x28 & x59 ;
  assign n1763 = n202 & n1762 ;
  assign n1764 = n1763 ^ n1324 ^ 1'b0 ;
  assign n1765 = ~n1761 & n1764 ;
  assign n1766 = n1240 ^ n718 ^ x46 ;
  assign n1767 = n1766 ^ n855 ^ 1'b0 ;
  assign n1768 = ~n845 & n1133 ;
  assign n1769 = n529 & n1768 ;
  assign n1770 = n505 | n1769 ;
  assign n1771 = n768 | n1770 ;
  assign n1772 = x48 & ~n1771 ;
  assign n1773 = x15 & x82 ;
  assign n1774 = x103 & n1773 ;
  assign n1775 = n1535 ^ x70 ^ 1'b0 ;
  assign n1776 = n753 & ~n1775 ;
  assign n1777 = ~n283 & n1776 ;
  assign n1778 = ~n1774 & n1777 ;
  assign n1779 = n708 | n779 ;
  assign n1780 = ~n1778 & n1779 ;
  assign n1781 = x27 & n175 ;
  assign n1782 = ~n879 & n1781 ;
  assign n1783 = n1546 | n1782 ;
  assign n1784 = n1410 & ~n1783 ;
  assign n1785 = n504 | n1661 ;
  assign n1786 = ~n605 & n1785 ;
  assign n1787 = x99 & ~n262 ;
  assign n1788 = n1221 & n1787 ;
  assign n1789 = n1788 ^ n1293 ^ 1'b0 ;
  assign n1790 = n1786 & ~n1789 ;
  assign n1791 = ~n404 & n1300 ;
  assign n1792 = n740 & ~n1791 ;
  assign n1793 = n1183 & ~n1558 ;
  assign n1794 = ~n1792 & n1793 ;
  assign n1795 = n180 & n753 ;
  assign n1796 = ~x5 & n1795 ;
  assign n1797 = n1155 ^ n530 ^ x5 ;
  assign n1798 = n1693 | n1797 ;
  assign n1799 = n1796 & ~n1798 ;
  assign n1800 = n569 ^ n527 ^ 1'b0 ;
  assign n1801 = ~n541 & n1800 ;
  assign n1802 = n1801 ^ n1336 ^ 1'b0 ;
  assign n1803 = n1361 & ~n1802 ;
  assign n1804 = n1097 ^ n787 ^ n236 ;
  assign n1805 = ( n1155 & ~n1313 ) | ( n1155 & n1484 ) | ( ~n1313 & n1484 ) ;
  assign n1806 = x23 & n1291 ;
  assign n1807 = n1806 ^ n1183 ^ 1'b0 ;
  assign n1808 = n391 & ~n713 ;
  assign n1809 = n431 & n1808 ;
  assign n1810 = n1809 ^ n1426 ^ 1'b0 ;
  assign n1811 = n758 & n1094 ;
  assign n1812 = n1811 ^ x61 ^ 1'b0 ;
  assign n1813 = n1273 ^ n323 ^ 1'b0 ;
  assign n1814 = ( n431 & ~n468 ) | ( n431 & n733 ) | ( ~n468 & n733 ) ;
  assign n1815 = n935 ^ n791 ^ 1'b0 ;
  assign n1816 = n1814 & ~n1815 ;
  assign n1817 = n1103 | n1816 ;
  assign n1818 = n288 & n645 ;
  assign n1819 = ~x34 & n1818 ;
  assign n1820 = n531 ^ n371 ^ 1'b0 ;
  assign n1821 = ~n595 & n1820 ;
  assign n1822 = ~n1040 & n1821 ;
  assign n1823 = n1027 & n1822 ;
  assign n1824 = n1823 ^ n184 ^ 1'b0 ;
  assign n1825 = n567 ^ n133 ^ 1'b0 ;
  assign n1826 = n1735 & ~n1825 ;
  assign n1827 = ~n1692 & n1826 ;
  assign n1828 = n301 | n1827 ;
  assign n1829 = n620 ^ n353 ^ 1'b0 ;
  assign n1830 = n488 | n1829 ;
  assign n1831 = n1830 ^ n1496 ^ x94 ;
  assign n1832 = n1819 & n1831 ;
  assign n1833 = n305 ^ x11 ^ 1'b0 ;
  assign n1834 = x43 & ~n1833 ;
  assign n1835 = n1834 ^ n401 ^ 1'b0 ;
  assign n1836 = ~n892 & n1056 ;
  assign n1837 = n213 & ~n272 ;
  assign n1838 = ~n1713 & n1837 ;
  assign n1839 = n542 | n1838 ;
  assign n1840 = n484 & ~n1839 ;
  assign n1841 = x109 & ~n1840 ;
  assign n1842 = n382 & n1841 ;
  assign n1843 = n1842 ^ n477 ^ 1'b0 ;
  assign n1844 = n1836 & n1843 ;
  assign n1845 = x58 & n694 ;
  assign n1846 = n1735 & ~n1845 ;
  assign n1847 = n1846 ^ n1164 ^ 1'b0 ;
  assign n1848 = n1847 ^ n704 ^ 1'b0 ;
  assign n1849 = n468 & ~n1848 ;
  assign n1850 = n607 ^ n444 ^ 1'b0 ;
  assign n1851 = n440 | n1850 ;
  assign n1852 = n1527 ^ x40 ^ 1'b0 ;
  assign n1853 = n1348 | n1852 ;
  assign n1854 = n658 & n1853 ;
  assign n1855 = n1321 ^ n238 ^ 1'b0 ;
  assign n1856 = ~n1040 & n1855 ;
  assign n1857 = n1856 ^ n1263 ^ 1'b0 ;
  assign n1858 = ~n1854 & n1857 ;
  assign n1859 = ~n886 & n1713 ;
  assign n1860 = n1859 ^ n1856 ^ 1'b0 ;
  assign n1861 = n1510 ^ n147 ^ 1'b0 ;
  assign n1862 = x69 & ~n1467 ;
  assign n1863 = n1723 ^ n1040 ^ 1'b0 ;
  assign n1864 = n868 | n1767 ;
  assign n1865 = n1037 & ~n1864 ;
  assign n1866 = n732 ^ n499 ^ 1'b0 ;
  assign n1867 = ~n290 & n1866 ;
  assign n1868 = ( n468 & ~n527 ) | ( n468 & n1867 ) | ( ~n527 & n1867 ) ;
  assign n1869 = x63 ^ x6 ^ 1'b0 ;
  assign n1870 = n581 & n667 ;
  assign n1871 = n1870 ^ n147 ^ 1'b0 ;
  assign n1872 = n1869 & n1871 ;
  assign n1873 = n1872 ^ n1740 ^ 1'b0 ;
  assign n1874 = ~n1868 & n1873 ;
  assign n1875 = x18 & n1033 ;
  assign n1876 = ~n1450 & n1875 ;
  assign n1877 = ( n1044 & n1467 ) | ( n1044 & ~n1689 ) | ( n1467 & ~n1689 ) ;
  assign n1878 = n574 ^ n209 ^ 1'b0 ;
  assign n1879 = n1878 ^ n1301 ^ 1'b0 ;
  assign n1880 = n842 & ~n1879 ;
  assign n1881 = ( x43 & n256 ) | ( x43 & n546 ) | ( n256 & n546 ) ;
  assign n1882 = n704 | n1881 ;
  assign n1883 = n556 & n876 ;
  assign n1884 = n1883 ^ n640 ^ 1'b0 ;
  assign n1885 = n679 ^ n317 ^ 1'b0 ;
  assign n1886 = ~n1884 & n1885 ;
  assign n1887 = x57 & n1331 ;
  assign n1888 = n1887 ^ n651 ^ 1'b0 ;
  assign n1889 = n381 | n1118 ;
  assign n1890 = ( n1353 & n1888 ) | ( n1353 & n1889 ) | ( n1888 & n1889 ) ;
  assign n1891 = n742 & n1890 ;
  assign n1892 = ~n222 & n1221 ;
  assign n1893 = n1353 & ~n1416 ;
  assign n1894 = n1892 & ~n1893 ;
  assign n1895 = n1435 & n1894 ;
  assign n1896 = n730 ^ n182 ^ 1'b0 ;
  assign n1897 = n1012 & ~n1896 ;
  assign n1898 = n1897 ^ n1473 ^ 1'b0 ;
  assign n1899 = n1898 ^ n1845 ^ n1019 ;
  assign n1900 = n1092 & ~n1585 ;
  assign n1901 = n1900 ^ n184 ^ 1'b0 ;
  assign n1902 = n788 ^ n147 ^ 1'b0 ;
  assign n1903 = x12 & n1902 ;
  assign n1904 = n1903 ^ n791 ^ n507 ;
  assign n1905 = n1901 & ~n1904 ;
  assign n1906 = n1899 & n1905 ;
  assign n1907 = n983 | n1346 ;
  assign n1908 = n190 & n1092 ;
  assign n1909 = ( ~n1772 & n1907 ) | ( ~n1772 & n1908 ) | ( n1907 & n1908 ) ;
  assign n1910 = n694 ^ x50 ^ 1'b0 ;
  assign n1911 = n1910 ^ n630 ^ 1'b0 ;
  assign n1912 = ~n855 & n1432 ;
  assign n1913 = ( n688 & ~n795 ) | ( n688 & n1301 ) | ( ~n795 & n1301 ) ;
  assign n1914 = x70 & n1471 ;
  assign n1915 = n797 & n1914 ;
  assign n1916 = n1915 ^ n1776 ^ 1'b0 ;
  assign n1917 = n293 | n925 ;
  assign n1918 = n774 | n1408 ;
  assign n1919 = n1918 ^ n788 ^ 1'b0 ;
  assign n1920 = n1263 & n1919 ;
  assign n1921 = x24 & ~n442 ;
  assign n1922 = n1921 ^ n1276 ^ 1'b0 ;
  assign n1923 = ~n252 & n791 ;
  assign n1924 = ~n163 & n1923 ;
  assign n1925 = ( n200 & ~n671 ) | ( n200 & n1924 ) | ( ~n671 & n1924 ) ;
  assign n1926 = ( n480 & ~n1632 ) | ( n480 & n1925 ) | ( ~n1632 & n1925 ) ;
  assign n1927 = n1252 | n1926 ;
  assign n1928 = x31 & ~n243 ;
  assign n1929 = ~n427 & n1928 ;
  assign n1930 = n1279 ^ n369 ^ 1'b0 ;
  assign n1931 = ~n464 & n1930 ;
  assign n1932 = n1931 ^ n1096 ^ 1'b0 ;
  assign n1933 = n1932 ^ n1076 ^ 1'b0 ;
  assign n1934 = x97 & n1933 ;
  assign n1935 = n1929 & n1934 ;
  assign n1936 = n706 ^ x67 ^ x24 ;
  assign n1937 = n428 & n675 ;
  assign n1938 = n371 & n1077 ;
  assign n1939 = n1938 ^ n303 ^ 1'b0 ;
  assign n1940 = n210 & n393 ;
  assign n1941 = n1301 & n1940 ;
  assign n1942 = n1590 & ~n1941 ;
  assign n1943 = ~n1939 & n1942 ;
  assign n1948 = n993 & ~n1576 ;
  assign n1944 = n147 & ~n1149 ;
  assign n1945 = n1944 ^ n760 ^ 1'b0 ;
  assign n1946 = n597 & n1945 ;
  assign n1947 = n1013 & n1946 ;
  assign n1949 = n1948 ^ n1947 ^ 1'b0 ;
  assign n1950 = n1471 | n1949 ;
  assign n1951 = n995 ^ n293 ^ 1'b0 ;
  assign n1952 = ~n1756 & n1951 ;
  assign n1953 = n1952 ^ n297 ^ 1'b0 ;
  assign n1954 = n134 & ~n1616 ;
  assign n1955 = n1582 & n1954 ;
  assign n1958 = n1881 ^ n287 ^ 1'b0 ;
  assign n1959 = n147 & ~n1958 ;
  assign n1956 = x111 & ~n500 ;
  assign n1957 = n1956 ^ n1073 ^ 1'b0 ;
  assign n1960 = n1959 ^ n1957 ^ 1'b0 ;
  assign n1961 = n1058 & n1960 ;
  assign n1962 = n1961 ^ n398 ^ 1'b0 ;
  assign n1963 = n781 & n904 ;
  assign n1964 = n1962 & ~n1963 ;
  assign n1965 = n1964 ^ n808 ^ 1'b0 ;
  assign n1966 = n817 ^ n389 ^ 1'b0 ;
  assign n1967 = n1204 & ~n1295 ;
  assign n1968 = n1473 ^ n419 ^ 1'b0 ;
  assign n1969 = n1350 & ~n1968 ;
  assign n1970 = n1325 & ~n1969 ;
  assign n1971 = n224 & n1049 ;
  assign n1972 = n1567 ^ n988 ^ 1'b0 ;
  assign n1976 = n1051 ^ n453 ^ 1'b0 ;
  assign n1977 = x12 & n1976 ;
  assign n1973 = n392 ^ n236 ^ x61 ;
  assign n1974 = n817 & n1973 ;
  assign n1975 = n1974 ^ n487 ^ 1'b0 ;
  assign n1978 = n1977 ^ n1975 ^ 1'b0 ;
  assign n1979 = n1495 ^ x127 ^ 1'b0 ;
  assign n1980 = n1979 ^ n1909 ^ 1'b0 ;
  assign n1981 = ~n1019 & n1980 ;
  assign n1982 = n1981 ^ n1888 ^ 1'b0 ;
  assign n1983 = x30 & ~n808 ;
  assign n1984 = n194 | n387 ;
  assign n1985 = n1984 ^ n1614 ^ 1'b0 ;
  assign n1986 = ~n1681 & n1985 ;
  assign n1987 = ~n1983 & n1986 ;
  assign n1988 = n1840 & ~n1987 ;
  assign n1990 = n369 ^ n166 ^ 1'b0 ;
  assign n1989 = x88 & n661 ;
  assign n1991 = n1990 ^ n1989 ^ 1'b0 ;
  assign n1992 = n674 ^ n655 ^ 1'b0 ;
  assign n1993 = ~n685 & n1992 ;
  assign n1994 = n1993 ^ n1713 ^ 1'b0 ;
  assign n1995 = n808 & n1994 ;
  assign n1996 = n1867 ^ n1664 ^ 1'b0 ;
  assign n1997 = ~n319 & n1524 ;
  assign n1998 = n1997 ^ n1133 ^ 1'b0 ;
  assign n1999 = n1689 | n1998 ;
  assign n2000 = n632 ^ n462 ^ 1'b0 ;
  assign n2001 = n2000 ^ n1495 ^ 1'b0 ;
  assign n2002 = n2001 ^ x15 ^ 1'b0 ;
  assign n2003 = n956 & n2002 ;
  assign n2004 = x56 & n1200 ;
  assign n2005 = ~n709 & n2004 ;
  assign n2006 = n330 | n1124 ;
  assign n2007 = n2006 ^ n541 ^ 1'b0 ;
  assign n2008 = n1932 & n2007 ;
  assign n2009 = n1057 | n2008 ;
  assign n2010 = n943 ^ x43 ^ 1'b0 ;
  assign n2011 = n1147 | n2010 ;
  assign n2012 = n293 | n2011 ;
  assign n2013 = n730 | n1797 ;
  assign n2014 = x34 | n145 ;
  assign n2015 = ~n307 & n2014 ;
  assign n2016 = n2013 & n2015 ;
  assign n2018 = n1250 ^ n567 ^ 1'b0 ;
  assign n2019 = n2018 ^ n1111 ^ 1'b0 ;
  assign n2020 = n1674 & n2019 ;
  assign n2017 = x44 & n1165 ;
  assign n2021 = n2020 ^ n2017 ^ 1'b0 ;
  assign n2022 = n315 & ~n710 ;
  assign n2025 = x47 & n1204 ;
  assign n2026 = ~n232 & n2025 ;
  assign n2023 = n277 & ~n1143 ;
  assign n2024 = n2023 ^ n1879 ^ 1'b0 ;
  assign n2027 = n2026 ^ n2024 ^ 1'b0 ;
  assign n2028 = n926 & n1217 ;
  assign n2029 = x15 & n2028 ;
  assign n2030 = n1493 ^ n1429 ^ x110 ;
  assign n2031 = ~n363 & n863 ;
  assign n2032 = n1510 & n2031 ;
  assign n2033 = n2032 ^ n175 ^ 1'b0 ;
  assign n2034 = n620 ^ x79 ^ 1'b0 ;
  assign n2035 = n1491 & n2034 ;
  assign n2036 = ~n1757 & n2035 ;
  assign n2037 = n332 & n1450 ;
  assign n2038 = ~x69 & n2037 ;
  assign n2039 = n2038 ^ n1333 ^ 1'b0 ;
  assign n2041 = n277 & ~n1661 ;
  assign n2042 = n2041 ^ n1192 ^ 1'b0 ;
  assign n2040 = n1365 & n1873 ;
  assign n2043 = n2042 ^ n2040 ^ 1'b0 ;
  assign n2044 = n2043 ^ n1180 ^ 1'b0 ;
  assign n2045 = n1117 | n1518 ;
  assign n2046 = n2045 ^ x50 ^ 1'b0 ;
  assign n2050 = n1670 ^ n729 ^ n503 ;
  assign n2047 = n144 & ~n1074 ;
  assign n2048 = n2047 ^ x0 ^ 1'b0 ;
  assign n2049 = ~n749 & n2048 ;
  assign n2051 = n2050 ^ n2049 ^ n943 ;
  assign n2052 = n1662 ^ n1095 ^ 1'b0 ;
  assign n2053 = n578 & ~n2052 ;
  assign n2054 = n2053 ^ n842 ^ n246 ;
  assign n2056 = ~n305 & n1424 ;
  assign n2057 = n2056 ^ n1081 ^ 1'b0 ;
  assign n2058 = n1654 & n2057 ;
  assign n2059 = n1535 & n2058 ;
  assign n2055 = n637 ^ x98 ^ 1'b0 ;
  assign n2060 = n2059 ^ n2055 ^ x99 ;
  assign n2061 = x26 & n1646 ;
  assign n2062 = n2061 ^ x20 ^ 1'b0 ;
  assign n2063 = n915 & n1102 ;
  assign n2064 = ~n1385 & n2063 ;
  assign n2065 = n1693 | n2064 ;
  assign n2066 = n952 & ~n2065 ;
  assign n2067 = n1017 ^ n637 ^ 1'b0 ;
  assign n2068 = n920 | n1791 ;
  assign n2069 = n838 & n901 ;
  assign n2070 = ~n229 & n2069 ;
  assign n2071 = n969 ^ x35 ^ 1'b0 ;
  assign n2072 = ~n1587 & n2071 ;
  assign n2073 = ~n809 & n2072 ;
  assign n2074 = n1165 & n1279 ;
  assign n2075 = n1078 & n2074 ;
  assign n2076 = ( x37 & x99 ) | ( x37 & n2075 ) | ( x99 & n2075 ) ;
  assign n2077 = ~n1152 & n1881 ;
  assign n2078 = ~n435 & n2077 ;
  assign n2079 = n2078 ^ x112 ^ 1'b0 ;
  assign n2080 = n2076 & ~n2079 ;
  assign n2081 = n225 & ~n490 ;
  assign n2082 = n357 & n2081 ;
  assign n2083 = n678 & ~n2082 ;
  assign n2084 = n1186 & n2083 ;
  assign n2085 = ~n2080 & n2084 ;
  assign n2086 = n723 & ~n1309 ;
  assign n2087 = ( n287 & n645 ) | ( n287 & n685 ) | ( n645 & n685 ) ;
  assign n2088 = n960 | n2087 ;
  assign n2089 = n832 ^ x18 ^ 1'b0 ;
  assign n2090 = n246 & n2089 ;
  assign n2091 = n2090 ^ n875 ^ n397 ;
  assign n2092 = n1563 & n2091 ;
  assign n2093 = ~n1614 & n2092 ;
  assign n2094 = n1300 ^ n1027 ^ 1'b0 ;
  assign n2095 = n988 & n2094 ;
  assign n2096 = n1553 ^ n1329 ^ 1'b0 ;
  assign n2097 = n777 | n1860 ;
  assign n2098 = n1688 | n2097 ;
  assign n2100 = ~n440 & n1541 ;
  assign n2101 = n2100 ^ n384 ^ 1'b0 ;
  assign n2099 = n722 & ~n802 ;
  assign n2102 = n2101 ^ n2099 ^ 1'b0 ;
  assign n2103 = ~n913 & n2102 ;
  assign n2104 = ~n444 & n2055 ;
  assign n2105 = ~n2103 & n2104 ;
  assign n2106 = ~n204 & n1077 ;
  assign n2107 = n2106 ^ n1830 ^ 1'b0 ;
  assign n2108 = n667 & n1552 ;
  assign n2109 = n504 ^ x18 ^ 1'b0 ;
  assign n2110 = n2109 ^ n2048 ^ 1'b0 ;
  assign n2111 = n1541 & n2110 ;
  assign n2112 = n1321 ^ n788 ^ 1'b0 ;
  assign n2113 = n556 & ~n2112 ;
  assign n2114 = n1382 | n2113 ;
  assign n2115 = n1461 | n2114 ;
  assign n2116 = n2115 ^ n1746 ^ n1199 ;
  assign n2117 = n1033 ^ n489 ^ 1'b0 ;
  assign n2118 = n879 & n2117 ;
  assign n2119 = n2118 ^ n729 ^ 1'b0 ;
  assign n2120 = n1884 ^ n985 ^ 1'b0 ;
  assign n2126 = ( x27 & n279 ) | ( x27 & ~n1457 ) | ( n279 & ~n1457 ) ;
  assign n2127 = n861 | n2126 ;
  assign n2124 = ( x44 & n393 ) | ( x44 & ~n768 ) | ( n393 & ~n768 ) ;
  assign n2125 = ~n254 & n2124 ;
  assign n2121 = n1266 ^ x3 ^ 1'b0 ;
  assign n2122 = n1121 & ~n1553 ;
  assign n2123 = ~n2121 & n2122 ;
  assign n2128 = n2127 ^ n2125 ^ n2123 ;
  assign n2129 = n1809 ^ n1562 ^ 1'b0 ;
  assign n2130 = n1538 | n2129 ;
  assign n2131 = n2130 ^ n459 ^ 1'b0 ;
  assign n2132 = n1772 ^ n1627 ^ 1'b0 ;
  assign n2133 = n2131 & n2132 ;
  assign n2134 = ~n2024 & n2133 ;
  assign n2135 = n1529 ^ n489 ^ 1'b0 ;
  assign n2143 = x36 & n336 ;
  assign n2136 = ( n349 & n519 ) | ( n349 & n836 ) | ( n519 & n836 ) ;
  assign n2137 = n565 ^ n553 ^ 1'b0 ;
  assign n2138 = n2137 ^ n1939 ^ n1838 ;
  assign n2139 = n2138 ^ n815 ^ 1'b0 ;
  assign n2140 = n2136 & n2139 ;
  assign n2141 = n2140 ^ n927 ^ 1'b0 ;
  assign n2142 = n632 & n2141 ;
  assign n2144 = n2143 ^ n2142 ^ 1'b0 ;
  assign n2145 = n345 ^ n303 ^ 1'b0 ;
  assign n2146 = n645 & n2145 ;
  assign n2147 = n1507 ^ n464 ^ 1'b0 ;
  assign n2148 = n746 | n2147 ;
  assign n2149 = n1574 | n2148 ;
  assign n2150 = n2149 ^ n1971 ^ 1'b0 ;
  assign n2151 = n475 & ~n604 ;
  assign n2152 = n1558 & ~n2151 ;
  assign n2153 = n2152 ^ n571 ^ 1'b0 ;
  assign n2155 = n445 & n874 ;
  assign n2156 = n1248 & n2155 ;
  assign n2157 = n2156 ^ x89 ^ 1'b0 ;
  assign n2158 = n1078 & ~n2157 ;
  assign n2159 = n737 | n2158 ;
  assign n2154 = n756 ^ n321 ^ 1'b0 ;
  assign n2160 = n2159 ^ n2154 ^ 1'b0 ;
  assign n2161 = ~n609 & n2140 ;
  assign n2162 = n2161 ^ n1313 ^ 1'b0 ;
  assign n2163 = n959 ^ n756 ^ 1'b0 ;
  assign n2164 = ~n2162 & n2163 ;
  assign n2165 = n975 ^ n366 ^ 1'b0 ;
  assign n2166 = n2164 & n2165 ;
  assign n2167 = n2166 ^ n1933 ^ 1'b0 ;
  assign n2176 = n988 & n1342 ;
  assign n2177 = n649 & n2176 ;
  assign n2178 = n2177 ^ n883 ^ 1'b0 ;
  assign n2168 = ( x118 & ~n411 ) | ( x118 & n601 ) | ( ~n411 & n601 ) ;
  assign n2169 = n985 & n2168 ;
  assign n2170 = ~n1565 & n2169 ;
  assign n2171 = n397 | n1522 ;
  assign n2172 = n1344 ^ n525 ^ 1'b0 ;
  assign n2173 = n2172 ^ n1264 ^ 1'b0 ;
  assign n2174 = n2171 & ~n2173 ;
  assign n2175 = ~n2170 & n2174 ;
  assign n2179 = n2178 ^ n2175 ^ 1'b0 ;
  assign n2180 = x54 & n1273 ;
  assign n2181 = n1697 ^ n240 ^ 1'b0 ;
  assign n2182 = ~n1659 & n2181 ;
  assign n2183 = n143 & ~n2098 ;
  assign n2184 = ~n442 & n1076 ;
  assign n2185 = n478 & n2184 ;
  assign n2186 = ~n387 & n714 ;
  assign n2187 = n2186 ^ x125 ^ 1'b0 ;
  assign n2188 = n2187 ^ n1003 ^ 1'b0 ;
  assign n2189 = ( n1270 & n1916 ) | ( n1270 & ~n2188 ) | ( n1916 & ~n2188 ) ;
  assign n2191 = n2102 ^ n1809 ^ n1567 ;
  assign n2190 = n534 | n1452 ;
  assign n2192 = n2191 ^ n2190 ^ 1'b0 ;
  assign n2193 = n1566 ^ n392 ^ 1'b0 ;
  assign n2194 = n615 | n2193 ;
  assign n2195 = n2194 ^ n1761 ^ 1'b0 ;
  assign n2196 = n1001 ^ n342 ^ 1'b0 ;
  assign n2197 = ~n1398 & n2196 ;
  assign n2198 = ~n1353 & n2156 ;
  assign n2199 = n2006 ^ n796 ^ 1'b0 ;
  assign n2200 = ~n209 & n2199 ;
  assign n2201 = ( n2127 & n2198 ) | ( n2127 & ~n2200 ) | ( n2198 & ~n2200 ) ;
  assign n2202 = x33 & ~n1396 ;
  assign n2203 = n2202 ^ n1233 ^ 1'b0 ;
  assign n2204 = ( n1750 & n1769 ) | ( n1750 & ~n2203 ) | ( n1769 & ~n2203 ) ;
  assign n2205 = n755 | n2204 ;
  assign n2206 = n2205 ^ n681 ^ 1'b0 ;
  assign n2209 = n427 ^ x29 ^ 1'b0 ;
  assign n2210 = ~n831 & n2209 ;
  assign n2207 = n147 | n1484 ;
  assign n2208 = ~n1605 & n2207 ;
  assign n2211 = n2210 ^ n2208 ^ 1'b0 ;
  assign n2212 = n2024 ^ x116 ^ 1'b0 ;
  assign n2213 = n2211 | n2212 ;
  assign n2214 = ( ~x82 & n1889 ) | ( ~x82 & n2118 ) | ( n1889 & n2118 ) ;
  assign n2215 = ( n605 & n1842 ) | ( n605 & n2214 ) | ( n1842 & n2214 ) ;
  assign n2216 = ~n1639 & n1713 ;
  assign n2217 = n2216 ^ n1092 ^ 1'b0 ;
  assign n2218 = n2217 ^ n1510 ^ 1'b0 ;
  assign n2219 = n1427 ^ n335 ^ 1'b0 ;
  assign n2220 = n675 & ~n2219 ;
  assign n2221 = n2220 ^ x37 ^ 1'b0 ;
  assign n2222 = n1703 ^ x93 ^ x31 ;
  assign n2223 = ( n229 & ~n500 ) | ( n229 & n2222 ) | ( ~n500 & n2222 ) ;
  assign n2224 = x78 & n685 ;
  assign n2225 = n1823 | n2224 ;
  assign n2226 = n2223 | n2225 ;
  assign n2227 = n1612 ^ n175 ^ 1'b0 ;
  assign n2228 = n400 ^ x94 ^ 1'b0 ;
  assign n2229 = ~x89 & n2228 ;
  assign n2230 = n2227 & n2229 ;
  assign n2231 = ~n2226 & n2230 ;
  assign n2232 = n148 | n741 ;
  assign n2233 = ~n729 & n1686 ;
  assign n2234 = n2233 ^ n1920 ^ n1015 ;
  assign n2235 = n500 ^ n323 ^ 1'b0 ;
  assign n2236 = n2235 ^ n459 ^ 1'b0 ;
  assign n2237 = n1124 & n2236 ;
  assign n2238 = n1701 ^ n954 ^ 1'b0 ;
  assign n2239 = n505 & ~n2059 ;
  assign n2240 = n2238 & n2239 ;
  assign n2242 = n664 ^ x119 ^ 1'b0 ;
  assign n2243 = x1 | n2242 ;
  assign n2244 = n1529 ^ n215 ^ 1'b0 ;
  assign n2245 = n2243 & ~n2244 ;
  assign n2246 = n2245 ^ n1057 ^ 1'b0 ;
  assign n2247 = n423 | n2246 ;
  assign n2248 = x77 | n2247 ;
  assign n2241 = n208 | n431 ;
  assign n2249 = n2248 ^ n2241 ^ 1'b0 ;
  assign n2250 = n721 | n735 ;
  assign n2251 = ~n1703 & n2250 ;
  assign n2252 = n2251 ^ x65 ^ 1'b0 ;
  assign n2253 = n382 | n2252 ;
  assign n2254 = n2253 ^ n411 ^ 1'b0 ;
  assign n2255 = n2254 ^ n1372 ^ 1'b0 ;
  assign n2256 = n252 | n2170 ;
  assign n2257 = n218 & ~n2256 ;
  assign n2258 = x102 | n154 ;
  assign n2259 = n2258 ^ n234 ^ 1'b0 ;
  assign n2260 = x11 & n2090 ;
  assign n2261 = n2260 ^ n433 ^ 1'b0 ;
  assign n2262 = ~x94 & n2261 ;
  assign n2263 = n273 & ~n2262 ;
  assign n2264 = n2263 ^ n646 ^ 1'b0 ;
  assign n2265 = n987 & ~n2264 ;
  assign n2266 = n2085 & n2265 ;
  assign n2267 = n555 | n1574 ;
  assign n2268 = n858 ^ n669 ^ 1'b0 ;
  assign n2269 = n2268 ^ n1089 ^ 1'b0 ;
  assign n2270 = n1118 & n2269 ;
  assign n2271 = ( n1096 & ~n1361 ) | ( n1096 & n2270 ) | ( ~n1361 & n2270 ) ;
  assign n2272 = n246 & ~n625 ;
  assign n2273 = n2271 & n2272 ;
  assign n2274 = ~n2095 & n2273 ;
  assign n2275 = ( ~n795 & n808 ) | ( ~n795 & n1523 ) | ( n808 & n1523 ) ;
  assign n2276 = ~n448 & n2217 ;
  assign n2277 = x2 & ~n2276 ;
  assign n2278 = ~n1691 & n2277 ;
  assign n2279 = n364 | n1021 ;
  assign n2280 = n1230 | n2279 ;
  assign n2281 = n897 ^ n277 ^ 1'b0 ;
  assign n2282 = n1190 & ~n2281 ;
  assign n2283 = ~n2280 & n2282 ;
  assign n2284 = n2283 ^ n1119 ^ 1'b0 ;
  assign n2285 = n2278 | n2284 ;
  assign n2286 = x101 | n950 ;
  assign n2287 = n2286 ^ n745 ^ 1'b0 ;
  assign n2288 = n595 & ~n922 ;
  assign n2289 = n1738 ^ n601 ^ 1'b0 ;
  assign n2290 = n1198 | n1416 ;
  assign n2291 = n332 & ~n2290 ;
  assign n2292 = ~n1643 & n2291 ;
  assign n2293 = n2292 ^ n1429 ^ 1'b0 ;
  assign n2295 = ~x12 & n827 ;
  assign n2296 = n134 & ~n2295 ;
  assign n2297 = n718 & n2296 ;
  assign n2298 = n1732 & ~n2297 ;
  assign n2299 = n1115 | n2298 ;
  assign n2294 = n143 & n1250 ;
  assign n2300 = n2299 ^ n2294 ^ 1'b0 ;
  assign n2301 = n1365 & n1606 ;
  assign n2302 = n2301 ^ n1348 ^ 1'b0 ;
  assign n2303 = n559 ^ x121 ^ 1'b0 ;
  assign n2304 = x60 & n1143 ;
  assign n2305 = n1448 & n2304 ;
  assign n2306 = n2305 ^ n803 ^ n740 ;
  assign n2307 = x12 & ~n666 ;
  assign n2308 = n2170 | n2307 ;
  assign n2309 = n1190 ^ n723 ^ 1'b0 ;
  assign n2310 = n1811 | n2309 ;
  assign n2312 = n366 & ~n460 ;
  assign n2311 = n729 | n1581 ;
  assign n2313 = n2312 ^ n2311 ^ 1'b0 ;
  assign n2314 = x62 & ~n2313 ;
  assign n2315 = ~n2227 & n2314 ;
  assign n2316 = n759 & n787 ;
  assign n2317 = n2316 ^ n1617 ^ 1'b0 ;
  assign n2318 = ( n2105 & ~n2307 ) | ( n2105 & n2317 ) | ( ~n2307 & n2317 ) ;
  assign n2321 = n589 ^ n267 ^ 1'b0 ;
  assign n2320 = ~n656 & n801 ;
  assign n2322 = n2321 ^ n2320 ^ 1'b0 ;
  assign n2319 = n1213 ^ n669 ^ 1'b0 ;
  assign n2323 = n2322 ^ n2319 ^ n2005 ;
  assign n2324 = n540 ^ n269 ^ 1'b0 ;
  assign n2325 = n1649 | n2324 ;
  assign n2326 = n1202 & ~n2325 ;
  assign n2327 = n1511 & n2326 ;
  assign n2328 = n1773 ^ n1264 ^ x95 ;
  assign n2329 = n2003 & ~n2328 ;
  assign n2330 = n1583 & n2329 ;
  assign n2331 = ( ~n701 & n1167 ) | ( ~n701 & n2330 ) | ( n1167 & n2330 ) ;
  assign n2332 = n556 ^ n279 ^ 1'b0 ;
  assign n2333 = n1257 ^ x93 ^ 1'b0 ;
  assign n2334 = n896 & ~n2333 ;
  assign n2335 = n784 & n2146 ;
  assign n2336 = n2335 ^ x69 ^ 1'b0 ;
  assign n2337 = n2336 ^ n2164 ^ n1081 ;
  assign n2338 = n427 & ~n1276 ;
  assign n2339 = ( n507 & ~n768 ) | ( n507 & n1301 ) | ( ~n768 & n1301 ) ;
  assign n2340 = n1535 ^ n833 ^ 1'b0 ;
  assign n2341 = ~x126 & n1209 ;
  assign n2342 = x74 | n2341 ;
  assign n2343 = n2340 & n2342 ;
  assign n2344 = n2343 ^ n611 ^ 1'b0 ;
  assign n2345 = n2271 ^ n1405 ^ 1'b0 ;
  assign n2346 = ~n444 & n2345 ;
  assign n2347 = n1625 ^ n243 ^ 1'b0 ;
  assign n2348 = n2346 & ~n2347 ;
  assign n2349 = ~n362 & n716 ;
  assign n2350 = n2349 ^ n916 ^ 1'b0 ;
  assign n2351 = n911 & n2350 ;
  assign n2352 = x106 & ~n421 ;
  assign n2353 = ~n2351 & n2352 ;
  assign n2354 = ( n177 & n1204 ) | ( n177 & n1588 ) | ( n1204 & n1588 ) ;
  assign n2355 = n2354 ^ n1450 ^ 1'b0 ;
  assign n2356 = ~n1510 & n2355 ;
  assign n2357 = n171 | n620 ;
  assign n2358 = n679 | n2011 ;
  assign n2359 = n2358 ^ n366 ^ 1'b0 ;
  assign n2360 = n137 ^ x114 ^ x87 ;
  assign n2361 = n1567 & n2360 ;
  assign n2362 = n2361 ^ n2031 ^ 1'b0 ;
  assign n2363 = n1211 & n1748 ;
  assign n2364 = n941 | n1285 ;
  assign n2368 = ~n161 & n1973 ;
  assign n2369 = n1183 & ~n1825 ;
  assign n2370 = ~n2368 & n2369 ;
  assign n2365 = ~n373 & n2049 ;
  assign n2366 = n1797 | n2365 ;
  assign n2367 = n1809 | n2366 ;
  assign n2371 = n2370 ^ n2367 ^ 1'b0 ;
  assign n2372 = n683 & ~n1982 ;
  assign n2373 = n1697 ^ n1552 ^ 1'b0 ;
  assign n2374 = n1396 ^ n685 ^ 1'b0 ;
  assign n2375 = ~n952 & n2136 ;
  assign n2376 = n1605 & n2375 ;
  assign n2377 = n1771 ^ n704 ^ 1'b0 ;
  assign n2378 = ~n2376 & n2377 ;
  assign n2379 = n2378 ^ x37 ^ 1'b0 ;
  assign n2380 = ~n2264 & n2379 ;
  assign n2381 = n1058 ^ n1003 ^ 1'b0 ;
  assign n2382 = n661 & ~n1599 ;
  assign n2383 = n890 ^ x125 ^ 1'b0 ;
  assign n2384 = n311 & ~n2383 ;
  assign n2385 = x11 & n2384 ;
  assign n2386 = n2385 ^ n538 ^ 1'b0 ;
  assign n2387 = n1503 | n2386 ;
  assign n2388 = x59 & n2116 ;
  assign n2389 = n2196 ^ n679 ^ 1'b0 ;
  assign n2390 = x70 & ~n299 ;
  assign n2391 = n1357 & n2390 ;
  assign n2392 = ~x78 & n172 ;
  assign n2393 = ~n1515 & n1698 ;
  assign n2394 = n1661 & n2393 ;
  assign n2395 = n2200 | n2394 ;
  assign n2396 = n799 & ~n1641 ;
  assign n2397 = n1229 & n2396 ;
  assign n2398 = n1635 ^ n1634 ^ 1'b0 ;
  assign n2399 = x22 & ~n878 ;
  assign n2400 = ~n361 & n1155 ;
  assign n2401 = ~x74 & n2400 ;
  assign n2403 = n1496 ^ n1124 ^ 1'b0 ;
  assign n2402 = ( ~x72 & n505 ) | ( ~x72 & n1510 ) | ( n505 & n1510 ) ;
  assign n2404 = n2403 ^ n2402 ^ 1'b0 ;
  assign n2405 = n885 & n2404 ;
  assign n2406 = n2405 ^ n1021 ^ 1'b0 ;
  assign n2407 = n2401 | n2406 ;
  assign n2409 = n1099 ^ n1015 ^ x14 ;
  assign n2408 = n986 & ~n1085 ;
  assign n2410 = n2409 ^ n2408 ^ 1'b0 ;
  assign n2411 = n1722 | n2410 ;
  assign n2412 = n2407 & ~n2411 ;
  assign n2413 = n2121 ^ n1155 ^ n868 ;
  assign n2414 = ~n355 & n1869 ;
  assign n2415 = n719 ^ n250 ^ 1'b0 ;
  assign n2416 = n327 & ~n2415 ;
  assign n2417 = n2416 ^ n1550 ^ 1'b0 ;
  assign n2418 = n2417 ^ x122 ^ 1'b0 ;
  assign n2419 = n898 ^ n770 ^ n438 ;
  assign n2420 = n652 & ~n2419 ;
  assign n2421 = ~n808 & n2420 ;
  assign n2422 = n2421 ^ n377 ^ 1'b0 ;
  assign n2423 = ~n755 & n2422 ;
  assign n2424 = ~n2418 & n2423 ;
  assign n2425 = n900 & n1507 ;
  assign n2426 = n357 & ~n1588 ;
  assign n2427 = n2426 ^ n943 ^ 1'b0 ;
  assign n2428 = n1740 ^ n1154 ^ n651 ;
  assign n2429 = n172 | n1963 ;
  assign n2430 = x16 & n163 ;
  assign n2431 = n2430 ^ n407 ^ 1'b0 ;
  assign n2434 = ( x31 & n392 ) | ( x31 & n1549 ) | ( n392 & n1549 ) ;
  assign n2435 = n665 & n2434 ;
  assign n2432 = n208 | n1695 ;
  assign n2433 = n1638 | n2432 ;
  assign n2436 = n2435 ^ n2433 ^ 1'b0 ;
  assign n2437 = ~n600 & n1184 ;
  assign n2438 = n2437 ^ n685 ^ 1'b0 ;
  assign n2440 = n2146 ^ n139 ^ 1'b0 ;
  assign n2439 = n134 & n1003 ;
  assign n2441 = n2440 ^ n2439 ^ 1'b0 ;
  assign n2447 = n260 | n1761 ;
  assign n2442 = n675 | n913 ;
  assign n2443 = x4 & n1228 ;
  assign n2444 = n2443 ^ n1123 ^ 1'b0 ;
  assign n2445 = ( x21 & n2048 ) | ( x21 & n2444 ) | ( n2048 & n2444 ) ;
  assign n2446 = ~n2442 & n2445 ;
  assign n2448 = n2447 ^ n2446 ^ 1'b0 ;
  assign n2449 = n1281 ^ n1129 ^ 1'b0 ;
  assign n2450 = n437 & ~n1120 ;
  assign n2451 = ~n1401 & n1816 ;
  assign n2452 = n824 & ~n1705 ;
  assign n2453 = n753 & ~n1527 ;
  assign n2454 = n2453 ^ n1444 ^ 1'b0 ;
  assign n2455 = n499 | n2454 ;
  assign n2456 = n1854 & ~n2455 ;
  assign n2457 = n674 & ~n1270 ;
  assign n2458 = n517 & n2457 ;
  assign n2460 = n1085 ^ n829 ^ n673 ;
  assign n2459 = n174 | n283 ;
  assign n2461 = n2460 ^ n2459 ^ 1'b0 ;
  assign n2462 = n2458 | n2461 ;
  assign n2463 = x78 & n1977 ;
  assign n2464 = n2463 ^ n450 ^ n244 ;
  assign n2465 = n353 ^ n338 ^ 1'b0 ;
  assign n2466 = n133 & n2465 ;
  assign n2467 = x66 & n2466 ;
  assign n2468 = n2467 ^ n683 ^ 1'b0 ;
  assign n2469 = n1562 & ~n2044 ;
  assign n2470 = n2469 ^ n580 ^ 1'b0 ;
  assign n2471 = n2076 ^ x59 ^ 1'b0 ;
  assign n2472 = n499 ^ n148 ^ 1'b0 ;
  assign n2473 = n2471 & n2472 ;
  assign n2474 = n1008 | n1941 ;
  assign n2475 = n2474 ^ n937 ^ 1'b0 ;
  assign n2476 = ( n2470 & ~n2473 ) | ( n2470 & n2475 ) | ( ~n2473 & n2475 ) ;
  assign n2477 = n218 & n953 ;
  assign n2478 = ~n387 & n2207 ;
  assign n2479 = n2478 ^ n738 ^ 1'b0 ;
  assign n2480 = n1753 ^ n444 ^ 1'b0 ;
  assign n2481 = n496 & n2480 ;
  assign n2482 = ~n243 & n905 ;
  assign n2483 = ~x24 & n791 ;
  assign n2484 = ( x57 & ~n844 ) | ( x57 & n1801 ) | ( ~n844 & n1801 ) ;
  assign n2485 = ~n444 & n2484 ;
  assign n2486 = n174 & n2485 ;
  assign n2487 = n2486 ^ n2156 ^ n1341 ;
  assign n2488 = n805 ^ n657 ^ 1'b0 ;
  assign n2489 = ~n1103 & n2488 ;
  assign n2492 = n1881 ^ x120 ^ 1'b0 ;
  assign n2490 = n471 & n1089 ;
  assign n2491 = n1903 & ~n2490 ;
  assign n2493 = n2492 ^ n2491 ^ 1'b0 ;
  assign n2494 = n2489 & ~n2493 ;
  assign n2495 = n1962 ^ n1251 ^ 1'b0 ;
  assign n2496 = ~n400 & n2495 ;
  assign n2497 = n1687 ^ n934 ^ 1'b0 ;
  assign n2498 = n2497 ^ n725 ^ 1'b0 ;
  assign n2499 = x84 & ~n2498 ;
  assign n2500 = ~n175 & n2499 ;
  assign n2501 = n2500 ^ n1164 ^ 1'b0 ;
  assign n2502 = x77 | n1332 ;
  assign n2503 = ( ~n1023 & n1256 ) | ( ~n1023 & n2502 ) | ( n1256 & n2502 ) ;
  assign n2504 = ( n978 & n2501 ) | ( n978 & n2503 ) | ( n2501 & n2503 ) ;
  assign n2505 = n509 | n1531 ;
  assign n2506 = n2505 ^ n971 ^ 1'b0 ;
  assign n2507 = n817 & n2131 ;
  assign n2508 = n2506 & n2507 ;
  assign n2509 = n509 ^ n398 ^ 1'b0 ;
  assign n2510 = ~n2508 & n2509 ;
  assign n2511 = n2021 ^ n943 ^ 1'b0 ;
  assign n2512 = ~n1211 & n2511 ;
  assign n2513 = n1118 & n2475 ;
  assign n2514 = n2513 ^ n1038 ^ 1'b0 ;
  assign n2515 = n1882 & n2514 ;
  assign n2516 = n1754 ^ n660 ^ 1'b0 ;
  assign n2517 = ~n1947 & n2132 ;
  assign n2518 = n1135 & n2106 ;
  assign n2519 = n2131 & n2518 ;
  assign n2520 = ~n1871 & n2519 ;
  assign n2521 = n1892 ^ n1123 ^ 1'b0 ;
  assign n2522 = n1053 ^ x55 ^ 1'b0 ;
  assign n2523 = n382 | n2522 ;
  assign n2524 = n1204 ^ n856 ^ 1'b0 ;
  assign n2525 = n2523 | n2524 ;
  assign n2526 = n1661 ^ n309 ^ 1'b0 ;
  assign n2527 = n277 & n2526 ;
  assign n2528 = n2527 ^ n357 ^ 1'b0 ;
  assign n2529 = n144 & ~n2528 ;
  assign n2530 = ~n2087 & n2529 ;
  assign n2531 = n481 ^ n137 ^ x31 ;
  assign n2532 = n2531 ^ n586 ^ 1'b0 ;
  assign n2533 = n294 & n2532 ;
  assign n2534 = n2533 ^ n1142 ^ 1'b0 ;
  assign n2535 = ~n529 & n2534 ;
  assign n2536 = n511 & ~n2535 ;
  assign n2537 = n2536 ^ n655 ^ 1'b0 ;
  assign n2538 = n2373 ^ x10 ^ 1'b0 ;
  assign n2539 = n2003 & n2538 ;
  assign n2540 = n2539 ^ n1413 ^ n1008 ;
  assign n2551 = n484 | n498 ;
  assign n2541 = n1901 ^ n1243 ^ 1'b0 ;
  assign n2542 = n236 | n2541 ;
  assign n2543 = n722 & ~n777 ;
  assign n2544 = n1656 ^ n163 ^ 1'b0 ;
  assign n2545 = x8 & ~n2544 ;
  assign n2546 = n2341 | n2545 ;
  assign n2547 = n2543 & n2546 ;
  assign n2548 = n2547 ^ n1251 ^ 1'b0 ;
  assign n2549 = n2542 | n2548 ;
  assign n2550 = n420 & ~n2549 ;
  assign n2552 = n2551 ^ n2550 ^ 1'b0 ;
  assign n2553 = n371 & n2552 ;
  assign n2554 = ~n137 & n1805 ;
  assign n2555 = n1520 ^ x69 ^ 1'b0 ;
  assign n2556 = n476 | n2555 ;
  assign n2557 = ( ~n1586 & n1835 ) | ( ~n1586 & n2556 ) | ( n1835 & n2556 ) ;
  assign n2558 = n347 ^ x64 ^ 1'b0 ;
  assign n2559 = ( n1679 & n2409 ) | ( n1679 & n2558 ) | ( n2409 & n2558 ) ;
  assign n2560 = ~n1495 & n2398 ;
  assign n2561 = n1787 ^ n1088 ^ 1'b0 ;
  assign n2562 = ( n277 & ~n317 ) | ( n277 & n373 ) | ( ~n317 & n373 ) ;
  assign n2563 = ( n1682 & n2083 ) | ( n1682 & ~n2562 ) | ( n2083 & ~n2562 ) ;
  assign n2564 = n1209 ^ n1123 ^ 1'b0 ;
  assign n2565 = n653 ^ n571 ^ 1'b0 ;
  assign n2566 = x19 & ~n2565 ;
  assign n2567 = n2176 & ~n2566 ;
  assign n2568 = n1895 ^ n1005 ^ 1'b0 ;
  assign n2569 = n2567 | n2568 ;
  assign n2570 = n815 | n1955 ;
  assign n2571 = n2570 ^ n1722 ^ 1'b0 ;
  assign n2572 = x38 & ~n358 ;
  assign n2573 = n1013 & n2572 ;
  assign n2574 = n1810 ^ n826 ^ 1'b0 ;
  assign n2575 = n2573 | n2574 ;
  assign n2576 = n2525 | n2575 ;
  assign n2577 = n741 & ~n2576 ;
  assign n2578 = n1165 & ~n1270 ;
  assign n2579 = ~n810 & n2578 ;
  assign n2580 = n1567 & ~n2579 ;
  assign n2581 = ~n2372 & n2580 ;
  assign n2582 = n2305 ^ n395 ^ 1'b0 ;
  assign n2583 = ~n374 & n1319 ;
  assign n2584 = n2136 ^ n1520 ^ 1'b0 ;
  assign n2585 = n738 & ~n2584 ;
  assign n2586 = n2583 & n2585 ;
  assign n2587 = n2586 ^ n1163 ^ 1'b0 ;
  assign n2588 = n1406 ^ n355 ^ 1'b0 ;
  assign n2589 = n1102 & n2588 ;
  assign n2590 = ~n174 & n865 ;
  assign n2591 = ~n2589 & n2590 ;
  assign n2592 = n1567 ^ n509 ^ 1'b0 ;
  assign n2593 = n2591 | n2592 ;
  assign n2594 = n1926 | n1935 ;
  assign n2595 = n324 & ~n2594 ;
  assign n2596 = n141 | n2595 ;
  assign n2597 = n2558 ^ n1639 ^ 1'b0 ;
  assign n2598 = ~n710 & n900 ;
  assign n2599 = n2598 ^ n339 ^ 1'b0 ;
  assign n2600 = n2148 | n2599 ;
  assign n2601 = n2600 ^ n1939 ^ 1'b0 ;
  assign n2602 = n1102 ^ n695 ^ x24 ;
  assign n2603 = n2387 ^ n678 ^ 1'b0 ;
  assign n2604 = ( ~n475 & n1631 ) | ( ~n475 & n1871 ) | ( n1631 & n1871 ) ;
  assign n2605 = n925 ^ n886 ^ n787 ;
  assign n2606 = ~n1395 & n2464 ;
  assign n2607 = ~n2605 & n2606 ;
  assign n2608 = n2210 ^ n1046 ^ 1'b0 ;
  assign n2609 = n2608 ^ n2394 ^ 1'b0 ;
  assign n2610 = ~n1587 & n2609 ;
  assign n2611 = ( n232 & ~n1198 ) | ( n232 & n2531 ) | ( ~n1198 & n2531 ) ;
  assign n2612 = ( ~n265 & n469 ) | ( ~n265 & n2611 ) | ( n469 & n2611 ) ;
  assign n2613 = n1586 ^ n1163 ^ 1'b0 ;
  assign n2614 = n437 & n730 ;
  assign n2615 = n856 & n2614 ;
  assign n2616 = n1997 | n2615 ;
  assign n2617 = n2613 | n2616 ;
  assign n2618 = ( ~n377 & n857 ) | ( ~n377 & n2075 ) | ( n857 & n2075 ) ;
  assign n2619 = ~n2617 & n2618 ;
  assign n2620 = n1266 & ~n2619 ;
  assign n2621 = ~n1641 & n2620 ;
  assign n2622 = ~x61 & n2125 ;
  assign n2623 = n1396 ^ n680 ^ 1'b0 ;
  assign n2624 = x47 & n2623 ;
  assign n2625 = n1880 ^ n428 ^ 1'b0 ;
  assign n2626 = n1728 & ~n2625 ;
  assign n2627 = n784 ^ x61 ^ 1'b0 ;
  assign n2632 = x83 & n213 ;
  assign n2628 = n169 & ~n1402 ;
  assign n2629 = n2409 | n2628 ;
  assign n2630 = x17 & ~n2629 ;
  assign n2631 = n2200 & n2630 ;
  assign n2633 = n2632 ^ n2631 ^ 1'b0 ;
  assign n2634 = n2451 ^ n1263 ^ 1'b0 ;
  assign n2635 = n297 ^ x51 ^ 1'b0 ;
  assign n2636 = n928 & ~n2635 ;
  assign n2637 = n1814 ^ n1380 ^ 1'b0 ;
  assign n2638 = n2637 ^ n2388 ^ 1'b0 ;
  assign n2639 = n1163 ^ x65 ^ 1'b0 ;
  assign n2640 = n2639 ^ n1635 ^ x40 ;
  assign n2644 = n569 | n945 ;
  assign n2641 = n1168 & n1257 ;
  assign n2642 = ~n1009 & n2641 ;
  assign n2643 = n1315 | n2642 ;
  assign n2645 = n2644 ^ n2643 ^ 1'b0 ;
  assign n2646 = n1374 | n2645 ;
  assign n2647 = n2306 & ~n2646 ;
  assign n2648 = n2502 ^ n1311 ^ n646 ;
  assign n2649 = n1485 | n2328 ;
  assign n2650 = x77 | n2649 ;
  assign n2651 = ~n854 & n2650 ;
  assign n2652 = ~n2648 & n2651 ;
  assign n2653 = n1017 ^ x87 ^ 1'b0 ;
  assign n2654 = n1235 & ~n2653 ;
  assign n2655 = n1100 ^ x78 ^ 1'b0 ;
  assign n2657 = n498 | n1484 ;
  assign n2658 = n2499 | n2657 ;
  assign n2659 = n2242 ^ n287 ^ 1'b0 ;
  assign n2660 = n2658 & n2659 ;
  assign n2656 = n425 | n1030 ;
  assign n2661 = n2660 ^ n2656 ^ 1'b0 ;
  assign n2662 = n344 | n2661 ;
  assign n2663 = n2189 ^ n1654 ^ 1'b0 ;
  assign n2664 = n1856 & ~n2663 ;
  assign n2665 = n2662 & n2664 ;
  assign n2666 = n636 & n640 ;
  assign n2667 = n499 & n2666 ;
  assign n2668 = n2667 ^ n2492 ^ n1147 ;
  assign n2669 = n2668 ^ n1511 ^ 1'b0 ;
  assign n2670 = ~n1190 & n2669 ;
  assign n2671 = n2670 ^ n1133 ^ 1'b0 ;
  assign n2672 = n1204 ^ n735 ^ 1'b0 ;
  assign n2673 = n741 & n2672 ;
  assign n2674 = n1763 | n2673 ;
  assign n2675 = n2071 & n2674 ;
  assign n2676 = n2675 ^ n2431 ^ 1'b0 ;
  assign n2677 = ( n487 & ~n756 ) | ( n487 & n1102 ) | ( ~n756 & n1102 ) ;
  assign n2678 = ( n775 & n2371 ) | ( n775 & n2677 ) | ( n2371 & n2677 ) ;
  assign n2679 = n2262 ^ n489 ^ n435 ;
  assign n2680 = ~n1089 & n2679 ;
  assign n2681 = n2315 | n2515 ;
  assign n2682 = ~n694 & n2499 ;
  assign n2683 = n2682 ^ n317 ^ 1'b0 ;
  assign n2684 = ( ~n531 & n560 ) | ( ~n531 & n2683 ) | ( n560 & n2683 ) ;
  assign n2685 = n2684 ^ n898 ^ 1'b0 ;
  assign n2686 = n2685 ^ n2452 ^ n1354 ;
  assign n2687 = n2013 ^ n1420 ^ 1'b0 ;
  assign n2688 = n2611 ^ n791 ^ 1'b0 ;
  assign n2689 = n2514 | n2688 ;
  assign n2690 = n766 | n2326 ;
  assign n2691 = n622 | n2690 ;
  assign n2692 = n1081 ^ n745 ^ 1'b0 ;
  assign n2693 = n1755 ^ n787 ^ 1'b0 ;
  assign n2694 = n1279 & ~n2442 ;
  assign n2695 = n811 | n2694 ;
  assign n2696 = n2693 | n2695 ;
  assign n2697 = ~n1612 & n1679 ;
  assign n2698 = n1322 & ~n2697 ;
  assign n2699 = n2698 ^ n1534 ^ 1'b0 ;
  assign n2707 = n672 & ~n1028 ;
  assign n2708 = n2707 ^ x7 ^ 1'b0 ;
  assign n2709 = n2708 ^ n814 ^ 1'b0 ;
  assign n2706 = n521 | n1083 ;
  assign n2710 = n2709 ^ n2706 ^ 1'b0 ;
  assign n2700 = n1390 ^ x32 ^ 1'b0 ;
  assign n2701 = n713 | n2700 ;
  assign n2702 = ( n1344 & ~n1535 ) | ( n1344 & n2701 ) | ( ~n1535 & n2701 ) ;
  assign n2703 = n929 & n2702 ;
  assign n2704 = ~n2517 & n2703 ;
  assign n2705 = n2704 ^ n598 ^ 1'b0 ;
  assign n2711 = n2710 ^ n2705 ^ 1'b0 ;
  assign n2712 = n2699 & ~n2711 ;
  assign n2713 = n652 & n2673 ;
  assign n2714 = n2713 ^ n1985 ^ 1'b0 ;
  assign n2715 = n2714 ^ n1981 ^ n1229 ;
  assign n2716 = n1844 & n2462 ;
  assign n2717 = n2716 ^ n1275 ^ 1'b0 ;
  assign n2718 = n810 ^ n797 ^ 1'b0 ;
  assign n2719 = n419 | n2718 ;
  assign n2720 = n2719 ^ x17 ^ 1'b0 ;
  assign n2721 = n2720 ^ n1085 ^ 1'b0 ;
  assign n2722 = n163 & ~n2721 ;
  assign n2723 = ~n664 & n1745 ;
  assign n2724 = n2723 ^ x104 ^ 1'b0 ;
  assign n2725 = n227 & ~n431 ;
  assign n2726 = n1222 & n2725 ;
  assign n2727 = ~n1879 & n2589 ;
  assign n2728 = n1811 & n2727 ;
  assign n2729 = n782 & n2307 ;
  assign n2730 = n2729 ^ n2392 ^ 1'b0 ;
  assign n2731 = x53 & n180 ;
  assign n2732 = x8 & n2731 ;
  assign n2733 = n2732 ^ x53 ^ 1'b0 ;
  assign n2734 = n2733 ^ n2515 ^ 1'b0 ;
  assign n2735 = n1174 & ~n2734 ;
  assign n2736 = n1078 & ~n2431 ;
  assign n2737 = n2736 ^ n1647 ^ 1'b0 ;
  assign n2738 = n1957 ^ n133 ^ 1'b0 ;
  assign n2739 = ( n615 & n786 ) | ( n615 & n925 ) | ( n786 & n925 ) ;
  assign n2740 = n340 & n2739 ;
  assign n2741 = n2740 ^ n2200 ^ 1'b0 ;
  assign n2742 = n1529 & n2741 ;
  assign n2743 = n615 & n1754 ;
  assign n2744 = n186 | n1666 ;
  assign n2745 = x72 | n2744 ;
  assign n2746 = ( n442 & n459 ) | ( n442 & ~n1587 ) | ( n459 & ~n1587 ) ;
  assign n2747 = n331 & n2746 ;
  assign n2748 = n2747 ^ n760 ^ 1'b0 ;
  assign n2749 = n2748 ^ n139 ^ 1'b0 ;
  assign n2750 = ~n182 & n2749 ;
  assign n2751 = n1193 ^ n425 ^ 1'b0 ;
  assign n2752 = n2751 ^ n1713 ^ 1'b0 ;
  assign n2757 = n1044 ^ n588 ^ 1'b0 ;
  assign n2758 = n1253 & n2757 ;
  assign n2759 = n2758 ^ n1303 ^ 1'b0 ;
  assign n2753 = ~n305 & n1473 ;
  assign n2754 = n2753 ^ n747 ^ 1'b0 ;
  assign n2755 = x23 & ~n2754 ;
  assign n2756 = n283 & n2755 ;
  assign n2760 = n2759 ^ n2756 ^ n1271 ;
  assign n2761 = n2760 ^ n2054 ^ 1'b0 ;
  assign n2762 = ~n194 & n2761 ;
  assign n2763 = n1483 & n2762 ;
  assign n2767 = ~n344 & n833 ;
  assign n2768 = ~n261 & n2767 ;
  assign n2764 = n1971 & ~n2170 ;
  assign n2765 = ~n1121 & n2764 ;
  assign n2766 = n1805 | n2765 ;
  assign n2769 = n2768 ^ n2766 ^ 1'b0 ;
  assign n2773 = x98 & n833 ;
  assign n2774 = ~n334 & n2773 ;
  assign n2770 = n1119 ^ n767 ^ 1'b0 ;
  assign n2771 = ~n254 & n2770 ;
  assign n2772 = n2771 ^ n1620 ^ 1'b0 ;
  assign n2775 = n2774 ^ n2772 ^ 1'b0 ;
  assign n2776 = ~n1039 & n2775 ;
  assign n2777 = n1960 ^ n1582 ^ n1327 ;
  assign n2778 = n238 | n658 ;
  assign n2779 = n2778 ^ n487 ^ 1'b0 ;
  assign n2780 = ( n1245 & n2629 ) | ( n1245 & ~n2779 ) | ( n2629 & ~n2779 ) ;
  assign n2781 = n277 & n324 ;
  assign n2782 = ~x118 & n2781 ;
  assign n2783 = n1563 ^ n863 ^ 1'b0 ;
  assign n2784 = n2782 & ~n2783 ;
  assign n2785 = ~n832 & n2784 ;
  assign n2787 = n867 & n2499 ;
  assign n2786 = x97 & n446 ;
  assign n2788 = n2787 ^ n2786 ^ 1'b0 ;
  assign n2789 = n2788 ^ n1343 ^ 1'b0 ;
  assign n2790 = n134 & ~n2789 ;
  assign n2791 = x44 & ~n2454 ;
  assign n2792 = ~n937 & n2791 ;
  assign n2793 = n369 & ~n1273 ;
  assign n2794 = n2793 ^ n1587 ^ 1'b0 ;
  assign n2795 = ~n2337 & n2414 ;
  assign n2796 = n2795 ^ n381 ^ 1'b0 ;
  assign n2797 = ( n1331 & n1543 ) | ( n1331 & n2796 ) | ( n1543 & n2796 ) ;
  assign n2798 = n2421 ^ n1479 ^ 1'b0 ;
  assign n2799 = n2127 & n2798 ;
  assign n2800 = n1943 & n2799 ;
  assign n2801 = x7 ^ x6 ^ 1'b0 ;
  assign n2802 = n1287 | n2801 ;
  assign n2803 = n407 ^ n222 ^ 1'b0 ;
  assign n2804 = n2802 | n2803 ;
  assign n2805 = n2090 ^ n1910 ^ 1'b0 ;
  assign n2806 = ~n1152 & n1844 ;
  assign n2807 = n2708 ^ n2308 ^ n2275 ;
  assign n2808 = n651 | n973 ;
  assign n2809 = n1556 & ~n2808 ;
  assign n2810 = n2809 ^ n2542 ^ 1'b0 ;
  assign n2811 = n2805 & ~n2810 ;
  assign n2812 = ~n2530 & n2811 ;
  assign n2813 = n2127 ^ n1058 ^ 1'b0 ;
  assign n2814 = n2776 ^ n1761 ^ 1'b0 ;
  assign n2818 = ~n167 & n1538 ;
  assign n2819 = n695 | n2818 ;
  assign n2820 = n138 ^ x56 ^ 1'b0 ;
  assign n2821 = ~n2819 & n2820 ;
  assign n2815 = n1100 ^ n523 ^ 1'b0 ;
  assign n2816 = n1649 | n2815 ;
  assign n2817 = n1258 | n2816 ;
  assign n2822 = n2821 ^ n2817 ^ 1'b0 ;
  assign n2823 = n1729 ^ n238 ^ x66 ;
  assign n2824 = n2468 ^ n1129 ^ 1'b0 ;
  assign n2831 = n364 | n681 ;
  assign n2832 = n344 | n2831 ;
  assign n2829 = n726 & ~n1627 ;
  assign n2830 = n2401 & n2829 ;
  assign n2825 = n239 & ~n1138 ;
  assign n2826 = ~n1858 & n2825 ;
  assign n2827 = n2826 ^ n1128 ^ 1'b0 ;
  assign n2828 = ( x32 & n616 ) | ( x32 & n2827 ) | ( n616 & n2827 ) ;
  assign n2833 = n2832 ^ n2830 ^ n2828 ;
  assign n2834 = ~n163 & n2833 ;
  assign n2837 = n1256 ^ n133 ^ 1'b0 ;
  assign n2835 = n1473 ^ n243 ^ 1'b0 ;
  assign n2836 = n1922 & n2835 ;
  assign n2838 = n2837 ^ n2836 ^ 1'b0 ;
  assign n2839 = ~n139 & n340 ;
  assign n2840 = n2839 ^ x8 ^ 1'b0 ;
  assign n2841 = ~n651 & n1973 ;
  assign n2842 = n1658 & n2841 ;
  assign n2843 = n922 ^ n726 ^ 1'b0 ;
  assign n2844 = ~n2842 & n2843 ;
  assign n2845 = n2844 ^ n1741 ^ 1'b0 ;
  assign n2846 = n2845 ^ n1902 ^ n927 ;
  assign n2847 = n1396 ^ x38 ^ 1'b0 ;
  assign n2848 = ~n2168 & n2200 ;
  assign n2849 = n1515 & n2848 ;
  assign n2850 = n817 & n2492 ;
  assign n2851 = n2850 ^ n1346 ^ 1'b0 ;
  assign n2852 = ~n1810 & n2851 ;
  assign n2853 = ~x92 & n2852 ;
  assign n2854 = n2853 ^ n2548 ^ 1'b0 ;
  assign n2855 = n1180 ^ n902 ^ 1'b0 ;
  assign n2856 = n292 & n1485 ;
  assign n2857 = n2038 ^ n1723 ^ 1'b0 ;
  assign n2858 = n1609 & ~n2857 ;
  assign n2859 = ( ~n575 & n2856 ) | ( ~n575 & n2858 ) | ( n2856 & n2858 ) ;
  assign n2860 = ~n330 & n1077 ;
  assign n2861 = n2860 ^ n266 ^ 1'b0 ;
  assign n2862 = ( n338 & n1361 ) | ( n338 & n2861 ) | ( n1361 & n2861 ) ;
  assign n2863 = n875 ^ n760 ^ n279 ;
  assign n2864 = ~n498 & n1073 ;
  assign n2865 = n2366 & n2864 ;
  assign n2866 = n2865 ^ n1241 ^ 1'b0 ;
  assign n2867 = ~n1336 & n1969 ;
  assign n2868 = n1079 & n2867 ;
  assign n2869 = x6 & ~n362 ;
  assign n2870 = n2170 & ~n2188 ;
  assign n2871 = n161 & ~n2870 ;
  assign n2872 = n2871 ^ n2540 ^ 1'b0 ;
  assign n2873 = ~n1111 & n1359 ;
  assign n2874 = n2873 ^ n382 ^ 1'b0 ;
  assign n2875 = ~n513 & n1427 ;
  assign n2876 = n1204 ^ n740 ^ 1'b0 ;
  assign n2877 = n800 ^ x19 ^ 1'b0 ;
  assign n2878 = n2877 ^ n2426 ^ n1523 ;
  assign n2879 = n838 & n1962 ;
  assign n2880 = n2879 ^ n723 ^ 1'b0 ;
  assign n2881 = n1743 & n2880 ;
  assign n2882 = n2881 ^ n1510 ^ 1'b0 ;
  assign n2883 = n425 ^ n157 ^ 1'b0 ;
  assign n2884 = n737 ^ n499 ^ 1'b0 ;
  assign n2885 = ( x94 & n1647 ) | ( x94 & n2884 ) | ( n1647 & n2884 ) ;
  assign n2886 = n1529 ^ x31 ^ 1'b0 ;
  assign n2888 = n1496 ^ n147 ^ 1'b0 ;
  assign n2889 = n1361 & ~n2888 ;
  assign n2887 = n754 | n2224 ;
  assign n2890 = n2889 ^ n2887 ^ 1'b0 ;
  assign n2894 = n1243 ^ n421 ^ 1'b0 ;
  assign n2895 = n2894 ^ n569 ^ 1'b0 ;
  assign n2896 = ~n1129 & n2895 ;
  assign n2891 = x17 & x126 ;
  assign n2892 = n2891 ^ n639 ^ 1'b0 ;
  assign n2893 = ~n1939 & n2892 ;
  assign n2897 = n2896 ^ n2893 ^ 1'b0 ;
  assign n2898 = n2330 & ~n2897 ;
  assign n2899 = n2295 ^ n1176 ^ 1'b0 ;
  assign n2901 = n1317 ^ n458 ^ 1'b0 ;
  assign n2902 = ~n1105 & n2901 ;
  assign n2903 = n2902 ^ n1778 ^ 1'b0 ;
  assign n2904 = n666 & n2903 ;
  assign n2900 = n1121 ^ n679 ^ n540 ;
  assign n2905 = n2904 ^ n2900 ^ 1'b0 ;
  assign n2906 = n2899 | n2905 ;
  assign n2908 = ~n382 & n414 ;
  assign n2907 = n445 & n507 ;
  assign n2909 = n2908 ^ n2907 ^ 1'b0 ;
  assign n2910 = n2909 ^ n290 ^ 1'b0 ;
  assign n2911 = n2910 ^ n1167 ^ 1'b0 ;
  assign n2912 = n2607 | n2911 ;
  assign n2913 = n2599 ^ n1047 ^ n860 ;
  assign n2914 = n2913 ^ n1242 ^ 1'b0 ;
  assign n2915 = ~n338 & n2087 ;
  assign n2916 = n2686 ^ n2596 ^ n1009 ;
  assign n2917 = ( n369 & ~n468 ) | ( n369 & n1097 ) | ( ~n468 & n1097 ) ;
  assign n2918 = n392 & ~n2917 ;
  assign n2919 = n2918 ^ n1585 ^ 1'b0 ;
  assign n2920 = n2919 ^ n1877 ^ n1067 ;
  assign n2921 = n509 & n2031 ;
  assign n2922 = n2605 ^ n1605 ^ n791 ;
  assign n2923 = n1045 & n2922 ;
  assign n2924 = n774 & n2923 ;
  assign n2925 = ( n1750 & n2921 ) | ( n1750 & n2924 ) | ( n2921 & n2924 ) ;
  assign n2926 = n336 & ~n358 ;
  assign n2927 = n2926 ^ n194 ^ 1'b0 ;
  assign n2928 = n2927 ^ n1825 ^ 1'b0 ;
  assign n2930 = n505 & n1382 ;
  assign n2929 = ~x75 & n2758 ;
  assign n2931 = n2930 ^ n2929 ^ 1'b0 ;
  assign n2932 = n1659 & n2931 ;
  assign n2933 = n714 ^ n232 ^ 1'b0 ;
  assign n2934 = x68 & ~n777 ;
  assign n2935 = ~n2933 & n2934 ;
  assign n2936 = n2816 & ~n2935 ;
  assign n2937 = n445 ^ n157 ^ n144 ;
  assign n2938 = n290 | n1510 ;
  assign n2939 = n2938 ^ n2771 ^ 1'b0 ;
  assign n2940 = ~n2937 & n2939 ;
  assign n2941 = ~n855 & n1180 ;
  assign n2942 = ~n2940 & n2941 ;
  assign n2943 = n315 ^ n141 ^ 1'b0 ;
  assign n2944 = n1404 & ~n2943 ;
  assign n2945 = n1386 & n2944 ;
  assign n2946 = n1287 ^ x110 ^ 1'b0 ;
  assign n2947 = n2687 ^ n157 ^ 1'b0 ;
  assign n2948 = n2048 ^ n637 ^ 1'b0 ;
  assign n2949 = n2101 ^ n1871 ^ n1642 ;
  assign n2950 = n2949 ^ n1534 ^ 1'b0 ;
  assign n2951 = n565 | n2950 ;
  assign n2952 = x48 & n2951 ;
  assign n2953 = n143 & n2048 ;
  assign n2954 = ~n1566 & n2953 ;
  assign n2955 = n2954 ^ n1103 ^ 1'b0 ;
  assign n2956 = n2229 ^ n1990 ^ 1'b0 ;
  assign n2957 = n2090 ^ n959 ^ 1'b0 ;
  assign n2958 = ( n523 & n1553 ) | ( n523 & ~n2378 ) | ( n1553 & ~n2378 ) ;
  assign n2959 = n1637 ^ n1315 ^ 1'b0 ;
  assign n2960 = n2286 ^ n401 ^ 1'b0 ;
  assign n2966 = ~n236 & n791 ;
  assign n2967 = n941 & n2966 ;
  assign n2968 = n2967 ^ n1086 ^ 1'b0 ;
  assign n2969 = n1124 | n2968 ;
  assign n2962 = n809 & ~n976 ;
  assign n2963 = n2962 ^ n1263 ^ 1'b0 ;
  assign n2961 = n1666 ^ n1081 ^ 1'b0 ;
  assign n2964 = n2963 ^ n2961 ^ 1'b0 ;
  assign n2965 = x39 & ~n2964 ;
  assign n2970 = n2969 ^ n2965 ^ 1'b0 ;
  assign n2971 = n430 & ~n2005 ;
  assign n2972 = n1109 & n2971 ;
  assign n2973 = x14 & ~n2972 ;
  assign n2974 = n2088 | n2193 ;
  assign n2975 = n148 | n859 ;
  assign n2976 = n2975 ^ n2333 ^ 1'b0 ;
  assign n2977 = n951 & n2746 ;
  assign n2978 = n254 & n2977 ;
  assign n2979 = n2978 ^ n506 ^ n442 ;
  assign n2981 = n1177 & ~n1588 ;
  assign n2982 = ~n1361 & n2981 ;
  assign n2980 = n2963 ^ n2272 ^ n1232 ;
  assign n2983 = n2982 ^ n2980 ^ 1'b0 ;
  assign n2984 = n2583 & ~n2983 ;
  assign n2985 = ~n1140 & n2423 ;
  assign n2988 = ~n1425 & n2756 ;
  assign n2989 = n1697 & ~n2988 ;
  assign n2986 = n802 | n2566 ;
  assign n2987 = n2986 ^ n1244 ^ 1'b0 ;
  assign n2990 = n2989 ^ n2987 ^ n1567 ;
  assign n2992 = n1013 | n2083 ;
  assign n2993 = n2992 ^ n726 ^ 1'b0 ;
  assign n2991 = n1197 ^ n425 ^ 1'b0 ;
  assign n2994 = n2993 ^ n2991 ^ n2701 ;
  assign n2995 = n855 ^ n186 ^ 1'b0 ;
  assign n2996 = n2589 & n2995 ;
  assign n2997 = n527 & n1354 ;
  assign n2998 = n2997 ^ n841 ^ 1'b0 ;
  assign n2999 = n2996 & n2998 ;
  assign n3000 = n2999 ^ n1049 ^ 1'b0 ;
  assign n3001 = n3000 ^ n1147 ^ x47 ;
  assign n3002 = x19 & ~n1634 ;
  assign n3003 = n3002 ^ n2300 ^ 1'b0 ;
  assign n3004 = n1281 ^ n722 ^ 1'b0 ;
  assign n3005 = ~n1056 & n1361 ;
  assign n3006 = n679 & n3005 ;
  assign n3007 = n3006 ^ n2931 ^ 1'b0 ;
  assign n3008 = n1374 & n3007 ;
  assign n3009 = n2039 ^ n1668 ^ n277 ;
  assign n3010 = n1670 ^ x126 ^ 1'b0 ;
  assign n3011 = x6 | n3010 ;
  assign n3012 = n3011 ^ n2059 ^ 1'b0 ;
  assign n3013 = ~n2937 & n3012 ;
  assign n3014 = n1738 ^ n511 ^ 1'b0 ;
  assign n3015 = n1118 & n3014 ;
  assign n3016 = n3015 ^ n186 ^ 1'b0 ;
  assign n3017 = ( n886 & ~n1429 ) | ( n886 & n3016 ) | ( ~n1429 & n3016 ) ;
  assign n3018 = n1484 ^ n194 ^ 1'b0 ;
  assign n3019 = n1184 & n3018 ;
  assign n3020 = n420 & n3019 ;
  assign n3021 = n499 ^ x118 ^ 1'b0 ;
  assign n3022 = n1222 ^ n875 ^ 1'b0 ;
  assign n3023 = n1133 ^ n682 ^ 1'b0 ;
  assign n3026 = x55 & n827 ;
  assign n3027 = ~n2286 & n3026 ;
  assign n3024 = n1914 ^ n1276 ^ 1'b0 ;
  assign n3025 = n1422 & ~n3024 ;
  assign n3028 = n3027 ^ n3025 ^ 1'b0 ;
  assign n3029 = n1632 | n3028 ;
  assign n3031 = n224 | n2708 ;
  assign n3032 = n588 & ~n3031 ;
  assign n3030 = n1771 & n2118 ;
  assign n3033 = n3032 ^ n3030 ^ 1'b0 ;
  assign n3034 = n1450 & n1816 ;
  assign n3035 = n2642 & n3034 ;
  assign n3036 = n2165 ^ n987 ^ 1'b0 ;
  assign n3037 = ~n3035 & n3036 ;
  assign n3038 = n1565 ^ n888 ^ 1'b0 ;
  assign n3039 = n2629 & n3038 ;
  assign n3040 = n3037 & n3039 ;
  assign n3041 = n3040 ^ n505 ^ 1'b0 ;
  assign n3042 = n1723 & n2083 ;
  assign n3043 = n2756 & n3042 ;
  assign n3044 = n2603 & ~n3043 ;
  assign n3045 = n3044 ^ x34 ^ 1'b0 ;
  assign n3046 = n679 ^ n427 ^ 1'b0 ;
  assign n3047 = n794 & ~n2462 ;
  assign n3048 = n2006 ^ n240 ^ 1'b0 ;
  assign n3049 = ( n2113 & ~n2697 ) | ( n2113 & n3048 ) | ( ~n2697 & n3048 ) ;
  assign n3050 = ~n2823 & n3049 ;
  assign n3051 = n1309 & n3050 ;
  assign n3053 = n1046 | n1675 ;
  assign n3054 = n1298 | n3053 ;
  assign n3052 = x14 & ~n1074 ;
  assign n3055 = n3054 ^ n3052 ^ 1'b0 ;
  assign n3056 = n2123 & n2288 ;
  assign n3057 = n836 | n3056 ;
  assign n3058 = n2102 | n3057 ;
  assign n3059 = ( n469 & n733 ) | ( n469 & ~n1221 ) | ( n733 & ~n1221 ) ;
  assign n3060 = n3059 ^ n1327 ^ 1'b0 ;
  assign n3061 = n855 | n3060 ;
  assign n3062 = ( n305 & n1399 ) | ( n305 & n2363 ) | ( n1399 & n2363 ) ;
  assign n3063 = n2441 & ~n2678 ;
  assign n3064 = n2634 & n3063 ;
  assign n3065 = n3064 ^ n2105 ^ 1'b0 ;
  assign n3066 = ~n1461 & n1511 ;
  assign n3067 = n1811 ^ n1250 ^ 1'b0 ;
  assign n3068 = n2553 ^ n1457 ^ 1'b0 ;
  assign n3069 = n915 & n2153 ;
  assign n3070 = n913 & n1710 ;
  assign n3071 = n2118 & n3070 ;
  assign n3072 = n1230 ^ n1094 ^ 1'b0 ;
  assign n3073 = ( n150 & n1193 ) | ( n150 & ~n3072 ) | ( n1193 & ~n3072 ) ;
  assign n3074 = n675 & ~n2346 ;
  assign n3075 = n3074 ^ n1176 ^ n660 ;
  assign n3076 = n2648 ^ n959 ^ 1'b0 ;
  assign n3077 = ~n1013 & n2613 ;
  assign n3078 = n3077 ^ n195 ^ 1'b0 ;
  assign n3079 = n2816 | n3078 ;
  assign n3080 = n1507 | n3079 ;
  assign n3081 = n1904 ^ n1794 ^ 1'b0 ;
  assign n3082 = n1672 ^ n1301 ^ x19 ;
  assign n3083 = n3082 ^ n442 ^ 1'b0 ;
  assign n3084 = n3083 ^ n2948 ^ 1'b0 ;
  assign n3085 = n1426 ^ n521 ^ 1'b0 ;
  assign n3086 = n975 & ~n3085 ;
  assign n3087 = ~n1129 & n2908 ;
  assign n3088 = n1195 & n3087 ;
  assign n3089 = n2596 & n3088 ;
  assign n3090 = n1264 & n1810 ;
  assign n3091 = n3090 ^ n1253 ^ 1'b0 ;
  assign n3092 = n1889 ^ n1495 ^ x30 ;
  assign n3093 = n2376 | n2683 ;
  assign n3094 = n1849 ^ n1212 ^ 1'b0 ;
  assign n3095 = n3093 | n3094 ;
  assign n3096 = ~n967 & n1737 ;
  assign n3097 = ~n1621 & n3096 ;
  assign n3098 = n1247 & ~n3097 ;
  assign n3099 = n1315 & n3098 ;
  assign n3100 = n930 & n1615 ;
  assign n3101 = n1204 ^ x71 ^ 1'b0 ;
  assign n3102 = n3101 ^ n754 ^ 1'b0 ;
  assign n3103 = n939 | n1514 ;
  assign n3104 = n3103 ^ n330 ^ 1'b0 ;
  assign n3105 = n612 | n3104 ;
  assign n3106 = n175 & n1361 ;
  assign n3107 = n1300 ^ n1056 ^ 1'b0 ;
  assign n3108 = n2428 ^ n695 ^ 1'b0 ;
  assign n3109 = n3107 | n3108 ;
  assign n3110 = n2131 ^ n1175 ^ 1'b0 ;
  assign n3113 = n1270 & n1774 ;
  assign n3111 = n1502 & n1575 ;
  assign n3112 = n1778 & ~n3111 ;
  assign n3114 = n3113 ^ n3112 ^ 1'b0 ;
  assign n3115 = n3110 | n3114 ;
  assign n3116 = n1689 ^ n1390 ^ n762 ;
  assign n3117 = x95 & ~n2283 ;
  assign n3118 = n1374 & n3117 ;
  assign n3119 = n208 | n3118 ;
  assign n3120 = n2390 & ~n3119 ;
  assign n3121 = n3120 ^ n1132 ^ 1'b0 ;
  assign n3122 = n2575 ^ n2101 ^ 1'b0 ;
  assign n3123 = n2647 ^ n1619 ^ 1'b0 ;
  assign n3124 = ~n326 & n3123 ;
  assign n3129 = n421 | n1406 ;
  assign n3130 = n1701 & ~n3129 ;
  assign n3125 = n1473 & ~n2486 ;
  assign n3126 = n3125 ^ n735 ^ 1'b0 ;
  assign n3127 = n3126 ^ n2710 ^ 1'b0 ;
  assign n3128 = n2673 & n3127 ;
  assign n3131 = n3130 ^ n3128 ^ n1163 ;
  assign n3132 = n382 ^ x6 ^ 1'b0 ;
  assign n3133 = n3131 & n3132 ;
  assign n3134 = n1408 | n1863 ;
  assign n3135 = n3134 ^ n1189 ^ 1'b0 ;
  assign n3136 = ~n488 & n1074 ;
  assign n3137 = x48 & ~n1497 ;
  assign n3138 = n577 & n3137 ;
  assign n3139 = ( n2575 & ~n3136 ) | ( n2575 & n3138 ) | ( ~n3136 & n3138 ) ;
  assign n3140 = n621 & ~n1592 ;
  assign n3141 = ~n1028 & n2280 ;
  assign n3142 = ~n714 & n3141 ;
  assign n3143 = n3142 ^ n605 ^ 1'b0 ;
  assign n3144 = n925 & ~n1150 ;
  assign n3145 = n2101 & n3144 ;
  assign n3146 = n3145 ^ n2908 ^ 1'b0 ;
  assign n3147 = n3146 ^ n1332 ^ x18 ;
  assign n3148 = n1186 & ~n1485 ;
  assign n3149 = n2880 ^ n1810 ^ 1'b0 ;
  assign n3150 = n878 & ~n3149 ;
  assign n3151 = ~n565 & n3150 ;
  assign n3152 = n3148 & n3151 ;
  assign n3153 = ~n3147 & n3152 ;
  assign n3154 = n2632 ^ n2224 ^ 1'b0 ;
  assign n3155 = ~n555 & n2433 ;
  assign n3156 = n1367 & n3155 ;
  assign n3157 = n683 | n1661 ;
  assign n3158 = x115 | n3157 ;
  assign n3159 = x3 & ~n760 ;
  assign n3160 = ~n2988 & n3159 ;
  assign n3161 = n3158 & n3160 ;
  assign n3162 = n3161 ^ n208 ^ 1'b0 ;
  assign n3163 = n133 & n2477 ;
  assign n3164 = n3163 ^ n1965 ^ 1'b0 ;
  assign n3165 = n1073 ^ n869 ^ 1'b0 ;
  assign n3167 = ~x108 & n695 ;
  assign n3166 = x28 & ~n2673 ;
  assign n3168 = n3167 ^ n3166 ^ 1'b0 ;
  assign n3169 = ~n1011 & n3168 ;
  assign n3170 = n883 & ~n1537 ;
  assign n3171 = ( n675 & n1026 ) | ( n675 & n3170 ) | ( n1026 & n3170 ) ;
  assign n3172 = ~n503 & n3171 ;
  assign n3173 = n1703 ^ x82 ^ 1'b0 ;
  assign n3174 = n1562 & ~n3173 ;
  assign n3175 = n3172 & n3174 ;
  assign n3176 = n262 & n2022 ;
  assign n3177 = n3176 ^ x72 ^ 1'b0 ;
  assign n3180 = n2227 ^ n1261 ^ n849 ;
  assign n3178 = x23 & ~n1804 ;
  assign n3179 = n3178 ^ n878 ^ 1'b0 ;
  assign n3181 = n3180 ^ n3179 ^ 1'b0 ;
  assign n3182 = x34 & ~n3181 ;
  assign n3183 = n3182 ^ n1979 ^ 1'b0 ;
  assign n3184 = n648 & n2200 ;
  assign n3185 = n3184 ^ n1927 ^ 1'b0 ;
  assign n3186 = ~n427 & n1183 ;
  assign n3187 = n143 & ~n710 ;
  assign n3188 = n1520 & n3187 ;
  assign n3189 = n301 ^ x83 ^ 1'b0 ;
  assign n3190 = ( n349 & ~n655 ) | ( n349 & n1588 ) | ( ~n655 & n1588 ) ;
  assign n3191 = n3190 ^ n1541 ^ 1'b0 ;
  assign n3192 = ~n2853 & n3191 ;
  assign n3193 = ( ~n2434 & n3189 ) | ( ~n2434 & n3192 ) | ( n3189 & n3192 ) ;
  assign n3194 = ~x38 & n2477 ;
  assign n3195 = n3194 ^ n2103 ^ 1'b0 ;
  assign n3196 = n2006 ^ n988 ^ 1'b0 ;
  assign n3197 = ~n395 & n3196 ;
  assign n3198 = ~n792 & n3197 ;
  assign n3199 = n3198 ^ n2931 ^ 1'b0 ;
  assign n3200 = n1860 | n3199 ;
  assign n3201 = n1927 & ~n2162 ;
  assign n3202 = ~n1735 & n3201 ;
  assign n3203 = n3202 ^ n1309 ^ 1'b0 ;
  assign n3204 = n175 & n1439 ;
  assign n3205 = n2883 & n3204 ;
  assign n3206 = n555 | n585 ;
  assign n3207 = n3206 ^ n1510 ^ 1'b0 ;
  assign n3209 = n2340 ^ n621 ^ 1'b0 ;
  assign n3208 = n327 & n2126 ;
  assign n3210 = n3209 ^ n3208 ^ 1'b0 ;
  assign n3211 = n1691 & n3210 ;
  assign n3212 = n999 & n3211 ;
  assign n3213 = n3212 ^ n1572 ^ 1'b0 ;
  assign n3214 = n802 | n3213 ;
  assign n3215 = x119 | n2337 ;
  assign n3216 = n335 ^ n243 ^ 1'b0 ;
  assign n3217 = n1424 & n3216 ;
  assign n3218 = ~n1924 & n3217 ;
  assign n3219 = n3218 ^ n1296 ^ 1'b0 ;
  assign n3220 = n1985 ^ n591 ^ 1'b0 ;
  assign n3221 = n2903 & n3220 ;
  assign n3222 = ( n958 & n3219 ) | ( n958 & ~n3221 ) | ( n3219 & ~n3221 ) ;
  assign n3223 = n1038 | n3222 ;
  assign n3224 = n649 | n3223 ;
  assign n3225 = n1027 ^ n557 ^ n459 ;
  assign n3226 = n3225 ^ n1682 ^ 1'b0 ;
  assign n3227 = n2292 | n3226 ;
  assign n3228 = ~n231 & n911 ;
  assign n3229 = n3228 ^ n3087 ^ 1'b0 ;
  assign n3230 = n2150 & n3229 ;
  assign n3231 = n2489 ^ n276 ^ 1'b0 ;
  assign n3232 = n1769 ^ n956 ^ 1'b0 ;
  assign n3233 = n935 | n3232 ;
  assign n3234 = n3233 ^ n1279 ^ 1'b0 ;
  assign n3235 = ~n643 & n744 ;
  assign n3236 = n1212 & n3235 ;
  assign n3237 = n460 & n2414 ;
  assign n3238 = n254 | n1773 ;
  assign n3239 = ~n836 & n3238 ;
  assign n3240 = ( ~n2945 & n3237 ) | ( ~n2945 & n3239 ) | ( n3237 & n3239 ) ;
  assign n3241 = n174 ^ x75 ^ 1'b0 ;
  assign n3242 = ~n3010 & n3241 ;
  assign n3243 = n3242 ^ n2930 ^ 1'b0 ;
  assign n3247 = n234 & ~n719 ;
  assign n3248 = ( n147 & ~n277 ) | ( n147 & n3247 ) | ( ~n277 & n3247 ) ;
  assign n3244 = n973 | n1325 ;
  assign n3245 = n1575 | n3244 ;
  assign n3246 = n3212 & n3245 ;
  assign n3249 = n3248 ^ n3246 ^ 1'b0 ;
  assign n3256 = n867 & n1174 ;
  assign n3257 = n894 & n3256 ;
  assign n3258 = n1361 & ~n3257 ;
  assign n3259 = n3258 ^ x65 ^ 1'b0 ;
  assign n3260 = n3259 ^ n1877 ^ 1'b0 ;
  assign n3261 = ~n2948 & n3260 ;
  assign n3250 = n1473 & n2543 ;
  assign n3251 = n3250 ^ n505 ^ 1'b0 ;
  assign n3252 = ~n694 & n1912 ;
  assign n3253 = n3251 & n3252 ;
  assign n3254 = n2628 | n3253 ;
  assign n3255 = n3254 ^ n2953 ^ 1'b0 ;
  assign n3262 = n3261 ^ n3255 ^ n204 ;
  assign n3263 = ~n180 & n2806 ;
  assign n3264 = ~n1012 & n3263 ;
  assign n3270 = x6 | n498 ;
  assign n3271 = n741 & n3270 ;
  assign n3272 = n3271 ^ n241 ^ 1'b0 ;
  assign n3265 = n1524 & ~n2130 ;
  assign n3266 = n3265 ^ n469 ^ 1'b0 ;
  assign n3267 = n1074 | n2275 ;
  assign n3268 = n3266 & ~n3267 ;
  assign n3269 = n1890 & ~n3268 ;
  assign n3273 = n3272 ^ n3269 ^ n1471 ;
  assign n3274 = n627 & ~n2779 ;
  assign n3275 = n1046 & n1562 ;
  assign n3276 = n3275 ^ x26 ^ 1'b0 ;
  assign n3277 = n2211 | n3276 ;
  assign n3278 = n1594 & ~n3277 ;
  assign n3279 = n3278 ^ n2543 ^ 1'b0 ;
  assign n3280 = n2898 ^ n1497 ^ 1'b0 ;
  assign n3281 = n1095 ^ n604 ^ 1'b0 ;
  assign n3282 = n3280 & n3281 ;
  assign n3283 = n1189 ^ n796 ^ 1'b0 ;
  assign n3284 = n1129 | n1588 ;
  assign n3285 = n3284 ^ n462 ^ 1'b0 ;
  assign n3286 = n3283 | n3285 ;
  assign n3287 = n2551 & n2715 ;
  assign n3288 = n3287 ^ x47 ^ 1'b0 ;
  assign n3289 = n688 & ~n714 ;
  assign n3290 = n662 & ~n3289 ;
  assign n3291 = n3290 ^ n857 ^ 1'b0 ;
  assign n3292 = x26 & ~n3291 ;
  assign n3293 = n875 | n2856 ;
  assign n3294 = n2416 | n3293 ;
  assign n3295 = n3294 ^ n139 ^ 1'b0 ;
  assign n3297 = ~n433 & n1481 ;
  assign n3296 = n297 & n2413 ;
  assign n3298 = n3297 ^ n3296 ^ 1'b0 ;
  assign n3299 = n1621 & n1966 ;
  assign n3300 = n2188 & n3299 ;
  assign n3301 = n886 | n2525 ;
  assign n3302 = n3301 ^ n2948 ^ 1'b0 ;
  assign n3303 = n2144 | n2745 ;
  assign n3305 = n542 ^ x98 ^ 1'b0 ;
  assign n3306 = ~n456 & n3305 ;
  assign n3307 = n1750 ^ n154 ^ 1'b0 ;
  assign n3308 = n3306 & n3307 ;
  assign n3304 = n1605 ^ n857 ^ 1'b0 ;
  assign n3309 = n3308 ^ n3304 ^ 1'b0 ;
  assign n3310 = n1790 & ~n3309 ;
  assign n3311 = n190 & n3166 ;
  assign n3313 = n1190 & n1503 ;
  assign n3312 = ~n1117 & n1433 ;
  assign n3314 = n3313 ^ n3312 ^ 1'b0 ;
  assign n3315 = n538 & n1132 ;
  assign n3316 = n3315 ^ n389 ^ 1'b0 ;
  assign n3317 = n3316 ^ n2197 ^ 1'b0 ;
  assign n3318 = ~n1039 & n3317 ;
  assign n3319 = n1121 ^ n922 ^ 1'b0 ;
  assign n3321 = ~n545 & n2787 ;
  assign n3320 = ( ~n400 & n464 ) | ( ~n400 & n614 ) | ( n464 & n614 ) ;
  assign n3322 = n3321 ^ n3320 ^ 1'b0 ;
  assign n3323 = n3322 ^ n1812 ^ 1'b0 ;
  assign n3324 = n3323 ^ n3162 ^ 1'b0 ;
  assign n3325 = n260 | n2701 ;
  assign n3326 = n3325 ^ n3320 ^ 1'b0 ;
  assign n3327 = n3145 ^ n1102 ^ 1'b0 ;
  assign n3328 = n3327 ^ n2759 ^ n1674 ;
  assign n3330 = n2658 ^ x58 ^ 1'b0 ;
  assign n3329 = n2255 & n2913 ;
  assign n3331 = n3330 ^ n3329 ^ 1'b0 ;
  assign n3332 = n593 | n1825 ;
  assign n3333 = n3332 ^ n929 ^ 1'b0 ;
  assign n3334 = n2953 & n3333 ;
  assign n3335 = n1523 | n2832 ;
  assign n3338 = ~x48 & x62 ;
  assign n3336 = n297 & n1293 ;
  assign n3337 = n1411 & ~n3336 ;
  assign n3339 = n3338 ^ n3337 ^ 1'b0 ;
  assign n3340 = ~n1515 & n1757 ;
  assign n3341 = n2681 & ~n3032 ;
  assign n3342 = n3341 ^ n2073 ^ 1'b0 ;
  assign n3343 = n1670 ^ n138 ^ 1'b0 ;
  assign n3344 = n1414 & ~n3343 ;
  assign n3345 = n411 ^ x38 ^ 1'b0 ;
  assign n3346 = n588 | n3345 ;
  assign n3347 = ~n875 & n2091 ;
  assign n3348 = n1085 & n3347 ;
  assign n3349 = n3346 | n3348 ;
  assign n3350 = n3344 | n3349 ;
  assign n3356 = x106 & ~n878 ;
  assign n3351 = n1670 | n1828 ;
  assign n3352 = n2083 | n3351 ;
  assign n3353 = n781 ^ x37 ^ 1'b0 ;
  assign n3354 = n3353 ^ n2403 ^ n815 ;
  assign n3355 = n3352 & n3354 ;
  assign n3357 = n3356 ^ n3355 ^ 1'b0 ;
  assign n3358 = n1217 & n2906 ;
  assign n3359 = n3358 ^ n813 ^ 1'b0 ;
  assign n3360 = ~n937 & n2098 ;
  assign n3361 = n1164 | n3360 ;
  assign n3362 = n1495 | n1728 ;
  assign n3363 = ~n593 & n1901 ;
  assign n3364 = n601 & n3363 ;
  assign n3365 = n928 | n3364 ;
  assign n3366 = n563 & n3365 ;
  assign n3367 = n2292 ^ n2013 ^ n309 ;
  assign n3368 = n3367 ^ n2050 ^ 1'b0 ;
  assign n3369 = n498 & ~n2619 ;
  assign n3370 = n1701 | n3048 ;
  assign n3371 = n1505 | n1588 ;
  assign n3372 = n3371 ^ n563 ^ 1'b0 ;
  assign n3373 = n1304 | n1344 ;
  assign n3374 = n2936 & ~n3373 ;
  assign n3375 = n406 & ~n1331 ;
  assign n3376 = n3375 ^ n821 ^ 1'b0 ;
  assign n3377 = n556 & ~n2319 ;
  assign n3378 = n3377 ^ n2363 ^ 1'b0 ;
  assign n3379 = n1467 ^ n421 ^ 1'b0 ;
  assign n3380 = ~n1639 & n3379 ;
  assign n3381 = ( n875 & ~n2561 ) | ( n875 & n3380 ) | ( ~n2561 & n3380 ) ;
  assign n3382 = x98 | n167 ;
  assign n3383 = n3382 ^ n278 ^ 1'b0 ;
  assign n3385 = n2842 ^ n1691 ^ n978 ;
  assign n3384 = n1150 ^ n708 ^ 1'b0 ;
  assign n3386 = n3385 ^ n3384 ^ 1'b0 ;
  assign n3387 = ~n2697 & n3386 ;
  assign n3388 = ~n3383 & n3387 ;
  assign n3389 = n3027 ^ n1588 ^ 1'b0 ;
  assign n3390 = n159 | n1222 ;
  assign n3391 = ~n1056 & n3390 ;
  assign n3392 = n398 & n636 ;
  assign n3393 = n3392 ^ n324 ^ 1'b0 ;
  assign n3394 = n2652 ^ n143 ^ 1'b0 ;
  assign n3395 = n3393 & ~n3394 ;
  assign n3396 = ~n1787 & n2014 ;
  assign n3397 = n1143 & n3396 ;
  assign n3398 = ( x42 & n1853 ) | ( x42 & n3397 ) | ( n1853 & n3397 ) ;
  assign n3399 = n3398 ^ n2391 ^ 1'b0 ;
  assign n3400 = n2489 | n3399 ;
  assign n3401 = x21 & n3400 ;
  assign n3402 = n2742 ^ n1217 ^ 1'b0 ;
  assign n3406 = n2904 ^ n875 ^ 1'b0 ;
  assign n3407 = n1897 & n3406 ;
  assign n3408 = ~x79 & n3407 ;
  assign n3409 = x54 & ~n1065 ;
  assign n3410 = n3409 ^ n1186 ^ 1'b0 ;
  assign n3411 = n718 & n3410 ;
  assign n3412 = n3411 ^ n143 ^ 1'b0 ;
  assign n3413 = n3408 | n3412 ;
  assign n3403 = ( n293 & n297 ) | ( n293 & ~n620 ) | ( n297 & ~n620 ) ;
  assign n3404 = n3403 ^ x29 ^ 1'b0 ;
  assign n3405 = n3404 ^ n2704 ^ 1'b0 ;
  assign n3414 = n3413 ^ n3405 ^ 1'b0 ;
  assign n3415 = n1756 ^ n1271 ^ 1'b0 ;
  assign n3416 = n3415 ^ n475 ^ 1'b0 ;
  assign n3417 = n460 & ~n3416 ;
  assign n3418 = n2969 ^ n1455 ^ n258 ;
  assign n3419 = n3418 ^ n2644 ^ 1'b0 ;
  assign n3420 = n195 & ~n709 ;
  assign n3421 = x105 & n2477 ;
  assign n3422 = ~n3068 & n3421 ;
  assign n3423 = n935 | n939 ;
  assign n3424 = n1681 | n3423 ;
  assign n3425 = n1325 & ~n1485 ;
  assign n3426 = ~n1880 & n3425 ;
  assign n3427 = n560 & n2546 ;
  assign n3428 = n145 & n3427 ;
  assign n3429 = n3428 ^ n621 ^ 1'b0 ;
  assign n3430 = n373 & ~n1510 ;
  assign n3432 = n1340 ^ n920 ^ 1'b0 ;
  assign n3433 = n2414 & ~n3432 ;
  assign n3431 = n543 & n2901 ;
  assign n3434 = n3433 ^ n3431 ^ 1'b0 ;
  assign n3435 = n718 & ~n1840 ;
  assign n3436 = n2300 | n3435 ;
  assign n3437 = n3436 ^ n1491 ^ 1'b0 ;
  assign n3438 = x25 & n1398 ;
  assign n3439 = n175 & n3400 ;
  assign n3440 = n1891 ^ n305 ^ 1'b0 ;
  assign n3441 = n1560 | n3440 ;
  assign n3442 = n1406 & ~n2113 ;
  assign n3443 = n3441 | n3442 ;
  assign n3444 = n3443 ^ n2407 ^ 1'b0 ;
  assign n3445 = n523 | n1111 ;
  assign n3446 = n1330 & n3445 ;
  assign n3447 = ~n1765 & n3446 ;
  assign n3448 = n2331 & n3447 ;
  assign n3449 = n498 | n1264 ;
  assign n3450 = n1424 & ~n2531 ;
  assign n3451 = n1433 & n2847 ;
  assign n3452 = n1005 & n3451 ;
  assign n3453 = ( n489 & n2151 ) | ( n489 & n3452 ) | ( n2151 & n3452 ) ;
  assign n3454 = n2492 & ~n3418 ;
  assign n3455 = n3454 ^ n404 ^ 1'b0 ;
  assign n3456 = n1279 & ~n2462 ;
  assign n3457 = n3455 & ~n3456 ;
  assign n3458 = n3457 ^ n969 ^ 1'b0 ;
  assign n3459 = n362 & n541 ;
  assign n3460 = n1331 & n1457 ;
  assign n3461 = n3460 ^ n1562 ^ 1'b0 ;
  assign n3462 = n3461 ^ n1390 ^ 1'b0 ;
  assign n3463 = ~n3459 & n3462 ;
  assign n3464 = n1348 | n3426 ;
  assign n3465 = n3464 ^ n3119 ^ 1'b0 ;
  assign n3466 = n1993 & n2107 ;
  assign n3467 = n368 & n3466 ;
  assign n3468 = ~n203 & n3467 ;
  assign n3469 = n1782 ^ n1623 ^ 1'b0 ;
  assign n3470 = n210 & n296 ;
  assign n3471 = n1277 & n1687 ;
  assign n3472 = n3471 ^ n1627 ^ 1'b0 ;
  assign n3473 = ~n1250 & n3472 ;
  assign n3474 = ~n3470 & n3473 ;
  assign n3475 = x98 | n1485 ;
  assign n3476 = n3475 ^ n2188 ^ 1'b0 ;
  assign n3477 = n1084 & n1342 ;
  assign n3478 = ( n632 & ~n1748 ) | ( n632 & n2444 ) | ( ~n1748 & n2444 ) ;
  assign n3479 = n3478 ^ n2861 ^ 1'b0 ;
  assign n3480 = x61 & ~n2969 ;
  assign n3481 = n1083 & n3480 ;
  assign n3482 = n389 | n1581 ;
  assign n3483 = n3482 ^ n1089 ^ 1'b0 ;
  assign n3484 = ~n3481 & n3483 ;
  assign n3485 = n3484 ^ n3027 ^ 1'b0 ;
  assign n3486 = ( n1733 & n2378 ) | ( n1733 & ~n3369 ) | ( n2378 & ~n3369 ) ;
  assign n3487 = ( n640 & n1661 ) | ( n640 & n1956 ) | ( n1661 & n1956 ) ;
  assign n3488 = n2514 ^ n2059 ^ 1'b0 ;
  assign n3489 = n791 & ~n822 ;
  assign n3490 = n458 & ~n3489 ;
  assign n3491 = n3490 ^ n1785 ^ 1'b0 ;
  assign n3492 = n1317 & n2880 ;
  assign n3493 = n3401 & n3492 ;
  assign n3494 = n2575 ^ n824 ^ 1'b0 ;
  assign n3495 = n735 | n3422 ;
  assign n3496 = n3116 | n3447 ;
  assign n3497 = n3496 ^ n534 ^ 1'b0 ;
  assign n3498 = n679 & ~n1939 ;
  assign n3499 = n3498 ^ n2919 ^ 1'b0 ;
  assign n3500 = n1776 ^ n708 ^ 1'b0 ;
  assign n3501 = n1641 & ~n3500 ;
  assign n3502 = n643 ^ x67 ^ 1'b0 ;
  assign n3503 = n2673 ^ n2144 ^ n874 ;
  assign n3504 = n3503 ^ n1773 ^ n1184 ;
  assign n3505 = n200 ^ x102 ^ 1'b0 ;
  assign n3506 = n273 & n2746 ;
  assign n3507 = n182 & n3506 ;
  assign n3508 = n1947 ^ x83 ^ 1'b0 ;
  assign n3509 = n625 | n1617 ;
  assign n3510 = n278 & ~n3509 ;
  assign n3511 = ( n258 & ~n1237 ) | ( n258 & n2579 ) | ( ~n1237 & n2579 ) ;
  assign n3512 = n3510 | n3511 ;
  assign n3513 = n1819 ^ n1372 ^ 1'b0 ;
  assign n3514 = ~n3512 & n3513 ;
  assign n3515 = n3514 ^ n1939 ^ n217 ;
  assign n3516 = n2353 ^ n1914 ^ 1'b0 ;
  assign n3517 = n2497 | n3516 ;
  assign n3518 = ( n2281 & n3515 ) | ( n2281 & n3517 ) | ( n3515 & n3517 ) ;
  assign n3519 = ~n1128 & n2131 ;
  assign n3520 = ~n1009 & n3519 ;
  assign n3521 = n2359 | n3520 ;
  assign n3522 = n1511 & ~n2482 ;
  assign n3523 = ~n3521 & n3522 ;
  assign n3524 = n3523 ^ n762 ^ 1'b0 ;
  assign n3525 = ~n455 & n505 ;
  assign n3526 = n3524 & n3525 ;
  assign n3527 = n1878 ^ n150 ^ 1'b0 ;
  assign n3528 = n571 | n3527 ;
  assign n3529 = n3121 ^ n469 ^ 1'b0 ;
  assign n3530 = n580 & n2718 ;
  assign n3531 = n2328 ^ n430 ^ 1'b0 ;
  assign n3532 = n3531 ^ n811 ^ n797 ;
  assign n3533 = ( x123 & ~n1620 ) | ( x123 & n3035 ) | ( ~n1620 & n3035 ) ;
  assign n3534 = n2774 | n3533 ;
  assign n3535 = n3534 ^ n2792 ^ 1'b0 ;
  assign n3536 = n2288 & n3535 ;
  assign n3537 = n2512 | n3188 ;
  assign n3538 = n2207 ^ n255 ^ 1'b0 ;
  assign n3539 = x12 & n3538 ;
  assign n3540 = n2621 ^ n2397 ^ 1'b0 ;
  assign n3541 = n3233 ^ n1031 ^ 1'b0 ;
  assign n3542 = n1124 | n3541 ;
  assign n3543 = n753 ^ x92 ^ 1'b0 ;
  assign n3544 = n157 | n3473 ;
  assign n3545 = n1750 ^ n605 ^ 1'b0 ;
  assign n3546 = n3544 & n3545 ;
  assign n3547 = n1241 & n3540 ;
  assign n3548 = n3182 ^ n363 ^ 1'b0 ;
  assign n3550 = n1253 & ~n2160 ;
  assign n3549 = n949 & n1190 ;
  assign n3551 = n3550 ^ n3549 ^ 1'b0 ;
  assign n3554 = n1708 ^ n861 ^ 1'b0 ;
  assign n3555 = n1509 | n3554 ;
  assign n3556 = x69 | n3555 ;
  assign n3552 = n478 ^ n445 ^ 1'b0 ;
  assign n3553 = ~n1138 & n3552 ;
  assign n3557 = n3556 ^ n3553 ^ 1'b0 ;
  assign n3558 = n307 ^ n184 ^ 1'b0 ;
  assign n3559 = ( n709 & n1073 ) | ( n709 & n3558 ) | ( n1073 & n3558 ) ;
  assign n3560 = ( n145 & ~n344 ) | ( n145 & n1033 ) | ( ~n344 & n1033 ) ;
  assign n3561 = ~n2673 & n3560 ;
  assign n3562 = ~n875 & n1951 ;
  assign n3563 = n3562 ^ n1738 ^ 1'b0 ;
  assign n3564 = n2299 & ~n3563 ;
  assign n3565 = n2016 ^ n1641 ^ 1'b0 ;
  assign n3566 = n3565 ^ n3474 ^ 1'b0 ;
  assign n3567 = n985 & n3566 ;
  assign n3568 = n1309 ^ n982 ^ 1'b0 ;
  assign n3569 = n1266 & ~n3568 ;
  assign n3570 = n1972 ^ n389 ^ 1'b0 ;
  assign n3571 = n3570 ^ n414 ^ 1'b0 ;
  assign n3572 = ~n167 & n171 ;
  assign n3573 = x39 & n3572 ;
  assign n3574 = n143 & n1439 ;
  assign n3575 = n3574 ^ n611 ^ x25 ;
  assign n3576 = n3575 ^ n1452 ^ n589 ;
  assign n3577 = ( n587 & n2917 ) | ( n587 & ~n3576 ) | ( n2917 & ~n3576 ) ;
  assign n3578 = n481 | n1907 ;
  assign n3579 = n3578 ^ n842 ^ 1'b0 ;
  assign n3580 = n1074 & n3579 ;
  assign n3581 = n1120 & n1687 ;
  assign n3582 = n3581 ^ n476 ^ 1'b0 ;
  assign n3583 = n1510 & ~n3582 ;
  assign n3584 = x93 | n509 ;
  assign n3585 = n3584 ^ n1003 ^ 1'b0 ;
  assign n3586 = n143 & n3585 ;
  assign n3587 = n3586 ^ n2562 ^ 1'b0 ;
  assign n3588 = n3587 ^ n494 ^ 1'b0 ;
  assign n3589 = ~n499 & n3588 ;
  assign n3590 = ( n1191 & n1838 ) | ( n1191 & ~n2445 ) | ( n1838 & ~n2445 ) ;
  assign n3591 = x110 & ~n945 ;
  assign n3592 = ~n1209 & n3591 ;
  assign n3593 = n3592 ^ n679 ^ 1'b0 ;
  assign n3594 = n1674 & ~n3593 ;
  assign n3595 = ~n3590 & n3594 ;
  assign n3596 = n1898 & ~n2049 ;
  assign n3597 = n1085 | n3596 ;
  assign n3598 = n1313 & n3597 ;
  assign n3599 = ~n915 & n3598 ;
  assign n3600 = ~n283 & n1878 ;
  assign n3601 = ~n844 & n3600 ;
  assign n3602 = n1245 & ~n2392 ;
  assign n3604 = n421 ^ x26 ^ 1'b0 ;
  assign n3603 = n2605 ^ n2287 ^ n1044 ;
  assign n3605 = n3604 ^ n3603 ^ 1'b0 ;
  assign n3606 = n1863 & ~n3130 ;
  assign n3607 = n2466 ^ n1787 ^ 1'b0 ;
  assign n3608 = n3606 & n3607 ;
  assign n3609 = n1831 ^ n1054 ^ 1'b0 ;
  assign n3610 = n249 & n3609 ;
  assign n3611 = n3610 ^ n3147 ^ 1'b0 ;
  assign n3612 = n1509 ^ n959 ^ 1'b0 ;
  assign n3613 = n832 & n3612 ;
  assign n3614 = n3613 ^ n288 ^ 1'b0 ;
  assign n3615 = n305 & n3614 ;
  assign n3616 = n440 & ~n498 ;
  assign n3617 = n719 ^ x107 ^ 1'b0 ;
  assign n3618 = n3616 & n3617 ;
  assign n3619 = ~n1283 & n3618 ;
  assign n3620 = ~n3153 & n3619 ;
  assign n3621 = ~n875 & n953 ;
  assign n3622 = n3621 ^ n327 ^ 1'b0 ;
  assign n3623 = n3622 ^ n431 ^ 1'b0 ;
  assign n3624 = ~n1987 & n3087 ;
  assign n3625 = n3623 & n3624 ;
  assign n3626 = n2373 & ~n3625 ;
  assign n3628 = n1680 ^ n1601 ^ 1'b0 ;
  assign n3629 = ~n275 & n3628 ;
  assign n3630 = n3629 ^ n567 ^ 1'b0 ;
  assign n3627 = n1531 | n2497 ;
  assign n3631 = n3630 ^ n3627 ^ 1'b0 ;
  assign n3632 = n1120 ^ n435 ^ 1'b0 ;
  assign n3633 = n3632 ^ n2366 ^ n277 ;
  assign n3634 = n3631 & ~n3633 ;
  assign n3635 = ~n3626 & n3634 ;
  assign n3636 = n213 | n1382 ;
  assign n3637 = n1691 ^ n622 ^ 1'b0 ;
  assign n3638 = n3636 & ~n3637 ;
  assign n3639 = ~n645 & n3638 ;
  assign n3640 = n1311 ^ n1149 ^ 1'b0 ;
  assign n3641 = n3306 & ~n3640 ;
  assign n3642 = n276 | n3641 ;
  assign n3643 = n2471 ^ n1037 ^ 1'b0 ;
  assign n3644 = n1251 & ~n3643 ;
  assign n3645 = ~n625 & n2659 ;
  assign n3646 = ~n407 & n3645 ;
  assign n3647 = n442 | n3584 ;
  assign n3648 = ( n540 & n1553 ) | ( n540 & n3647 ) | ( n1553 & n3647 ) ;
  assign n3649 = ~n1380 & n2321 ;
  assign n3655 = ~n653 & n1661 ;
  assign n3656 = x33 & ~n3655 ;
  assign n3657 = n3009 & n3656 ;
  assign n3650 = x97 & ~n2831 ;
  assign n3651 = n1476 & n3650 ;
  assign n3652 = n225 & ~n3651 ;
  assign n3653 = n3652 ^ n2167 ^ 1'b0 ;
  assign n3654 = n2662 | n3653 ;
  assign n3658 = n3657 ^ n3654 ^ 1'b0 ;
  assign n3659 = ~n3649 & n3658 ;
  assign n3660 = n1766 | n2221 ;
  assign n3661 = n129 & n817 ;
  assign n3662 = n3661 ^ n1083 ^ 1'b0 ;
  assign n3663 = n3662 ^ n1003 ^ 1'b0 ;
  assign n3664 = ~n3660 & n3663 ;
  assign n3665 = n246 & n2170 ;
  assign n3666 = n468 ^ n368 ^ 1'b0 ;
  assign n3667 = n1555 & ~n3666 ;
  assign n3668 = n708 & n3667 ;
  assign n3669 = n3668 ^ n1888 ^ n1509 ;
  assign n3670 = n3665 & ~n3669 ;
  assign n3671 = n3670 ^ n3570 ^ 1'b0 ;
  assign n3672 = n1398 ^ x99 ^ 1'b0 ;
  assign n3673 = n1484 | n3672 ;
  assign n3674 = n2005 & n3140 ;
  assign n3675 = n3674 ^ n3584 ^ n754 ;
  assign n3676 = n3675 ^ n789 ^ 1'b0 ;
  assign n3677 = ~x6 & n1537 ;
  assign n3678 = x64 & ~n3626 ;
  assign n3679 = n3378 ^ n1115 ^ 1'b0 ;
  assign n3680 = n1597 & n3679 ;
  assign n3681 = n2659 ^ n1687 ^ n1254 ;
  assign n3683 = n831 ^ n303 ^ 1'b0 ;
  assign n3684 = n3683 ^ n334 ^ 1'b0 ;
  assign n3685 = n2207 & n3684 ;
  assign n3682 = ( n256 & ~n808 ) | ( n256 & n1120 ) | ( ~n808 & n1120 ) ;
  assign n3686 = n3685 ^ n3682 ^ 1'b0 ;
  assign n3687 = n288 & ~n3686 ;
  assign n3688 = n675 & n3687 ;
  assign n3689 = ~n3681 & n3688 ;
  assign n3690 = ( n3442 & n3680 ) | ( n3442 & ~n3689 ) | ( n3680 & ~n3689 ) ;
  assign n3691 = n1529 & n2028 ;
  assign n3692 = n595 | n3691 ;
  assign n3693 = x88 | n3692 ;
  assign n3694 = n2022 ^ n1779 ^ 1'b0 ;
  assign n3695 = ~n1219 & n3511 ;
  assign n3696 = n3695 ^ n3373 ^ 1'b0 ;
  assign n3697 = ~n548 & n3696 ;
  assign n3698 = n1458 ^ n853 ^ 1'b0 ;
  assign n3699 = n816 | n3237 ;
  assign n3700 = n3698 | n3699 ;
  assign n3701 = n1654 & n2880 ;
  assign n3702 = n3435 ^ n2425 ^ 1'b0 ;
  assign n3703 = n1746 ^ n494 ^ 1'b0 ;
  assign n3704 = n1774 & n3703 ;
  assign n3705 = n1351 & n3704 ;
  assign n3706 = n3705 ^ n1649 ^ 1'b0 ;
  assign n3707 = n2280 & n3706 ;
  assign n3708 = n1296 & n3707 ;
  assign n3709 = ~n3259 & n3708 ;
  assign n3710 = ~x75 & n3709 ;
  assign n3711 = n3710 ^ n2865 ^ 1'b0 ;
  assign n3712 = ~n3302 & n3711 ;
  assign n3713 = n3712 ^ n1026 ^ 1'b0 ;
  assign n3717 = n1691 ^ n1569 ^ 1'b0 ;
  assign n3718 = n2892 & n3717 ;
  assign n3719 = ~n2589 & n3718 ;
  assign n3716 = n2497 ^ n1322 ^ 1'b0 ;
  assign n3714 = n2153 & ~n3616 ;
  assign n3715 = n3714 ^ n1728 ^ 1'b0 ;
  assign n3720 = n3719 ^ n3716 ^ n3715 ;
  assign n3721 = n2410 ^ n1691 ^ n425 ;
  assign n3722 = n2090 ^ n513 ^ 1'b0 ;
  assign n3723 = ~n1491 & n3722 ;
  assign n3724 = ~n3721 & n3723 ;
  assign n3725 = n788 & n2091 ;
  assign n3726 = n3725 ^ n1186 ^ 1'b0 ;
  assign n3727 = x4 & ~n2670 ;
  assign n3728 = ~n355 & n2605 ;
  assign n3729 = n3728 ^ n699 ^ 1'b0 ;
  assign n3730 = n1568 & n3729 ;
  assign n3731 = n735 & n1805 ;
  assign n3732 = n2945 | n3731 ;
  assign n3733 = n3730 | n3732 ;
  assign n3734 = n2743 & n3733 ;
  assign n3735 = ( ~n177 & n277 ) | ( ~n177 & n2321 ) | ( n277 & n2321 ) ;
  assign n3736 = n577 | n3735 ;
  assign n3737 = ~n505 & n3269 ;
  assign n3738 = n767 ^ x90 ^ 1'b0 ;
  assign n3739 = n1308 & n1343 ;
  assign n3740 = ~n3738 & n3739 ;
  assign n3741 = n2183 & ~n3740 ;
  assign n3743 = n1853 ^ n1113 ^ 1'b0 ;
  assign n3744 = ~n1585 & n3743 ;
  assign n3742 = ~n835 & n1331 ;
  assign n3745 = n3744 ^ n3742 ^ 1'b0 ;
  assign n3746 = ( n1401 & n2796 ) | ( n1401 & n3745 ) | ( n2796 & n3745 ) ;
  assign n3751 = n1202 ^ n866 ^ 1'b0 ;
  assign n3748 = ( ~x46 & n220 ) | ( ~x46 & n2992 ) | ( n220 & n2992 ) ;
  assign n3749 = ~n1103 & n3748 ;
  assign n3747 = ~n1190 & n1507 ;
  assign n3750 = n3749 ^ n3747 ^ 1'b0 ;
  assign n3752 = n3751 ^ n3750 ^ n180 ;
  assign n3753 = ( n255 & ~n553 ) | ( n255 & n1093 ) | ( ~n553 & n1093 ) ;
  assign n3756 = ~n386 & n435 ;
  assign n3757 = n992 & n3756 ;
  assign n3754 = n915 ^ n865 ^ 1'b0 ;
  assign n3755 = n294 & n3754 ;
  assign n3758 = n3757 ^ n3755 ^ 1'b0 ;
  assign n3759 = n1510 & n3758 ;
  assign n3760 = ~n3753 & n3759 ;
  assign n3761 = ~n540 & n1948 ;
  assign n3762 = n3140 ^ n517 ^ 1'b0 ;
  assign n3763 = n799 & n2168 ;
  assign n3764 = n3763 ^ n2829 ^ 1'b0 ;
  assign n3765 = n2484 & ~n3764 ;
  assign n3766 = n931 & n3765 ;
  assign n3767 = n1814 ^ n180 ^ 1'b0 ;
  assign n3768 = n3045 | n3767 ;
  assign n3769 = n3768 ^ n2010 ^ 1'b0 ;
  assign n3770 = n2824 & n3769 ;
  assign n3771 = n1182 & n1277 ;
  assign n3772 = ~x102 & n3771 ;
  assign n3773 = n2165 | n3772 ;
  assign n3774 = n3773 ^ n1956 ^ 1'b0 ;
  assign n3775 = ~n425 & n3774 ;
  assign n3776 = ~n323 & n1188 ;
  assign n3777 = n1071 & n3698 ;
  assign n3778 = n2198 & n3777 ;
  assign n3779 = n1137 & ~n3778 ;
  assign n3780 = n3779 ^ n1510 ^ 1'b0 ;
  assign n3781 = n2726 ^ n732 ^ 1'b0 ;
  assign n3783 = x33 & n1244 ;
  assign n3784 = n3783 ^ n1092 ^ 1'b0 ;
  assign n3782 = n479 & ~n1550 ;
  assign n3785 = n3784 ^ n3782 ^ 1'b0 ;
  assign n3786 = ~x72 & n3785 ;
  assign n3787 = n1432 ^ n934 ^ 1'b0 ;
  assign n3788 = x48 & n3787 ;
  assign n3789 = n3709 ^ n986 ^ 1'b0 ;
  assign n3790 = n2905 ^ n1631 ^ 1'b0 ;
  assign n3793 = n257 ^ x61 ^ 1'b0 ;
  assign n3794 = n2211 ^ n801 ^ 1'b0 ;
  assign n3795 = n3793 & ~n3794 ;
  assign n3796 = n529 | n1231 ;
  assign n3797 = n3796 ^ n1221 ^ 1'b0 ;
  assign n3798 = n3795 | n3797 ;
  assign n3791 = n2955 ^ n1204 ^ 1'b0 ;
  assign n3792 = ~n1811 & n3791 ;
  assign n3799 = n3798 ^ n3792 ^ 1'b0 ;
  assign n3800 = n2340 ^ x48 ^ 1'b0 ;
  assign n3801 = ( x109 & n3535 ) | ( x109 & n3800 ) | ( n3535 & n3800 ) ;
  assign n3802 = n1235 ^ n627 ^ 1'b0 ;
  assign n3803 = n3801 & ~n3802 ;
  assign n3804 = n3803 ^ n2113 ^ 1'b0 ;
  assign n3805 = n1635 ^ x65 ^ 1'b0 ;
  assign n3806 = n642 & n3805 ;
  assign n3807 = n2647 | n2819 ;
  assign n3808 = n3806 | n3807 ;
  assign n3809 = n2529 & ~n3808 ;
  assign n3810 = n1956 & n2026 ;
  assign n3811 = ~n2957 & n3810 ;
  assign n3812 = n679 ^ x75 ^ 1'b0 ;
  assign n3813 = n481 | n3812 ;
  assign n3814 = n3813 ^ n2856 ^ 1'b0 ;
  assign n3815 = n3814 ^ n2172 ^ 1'b0 ;
  assign n3816 = n1753 ^ x50 ^ 1'b0 ;
  assign n3817 = n3816 ^ n3389 ^ 1'b0 ;
  assign n3818 = n3815 & n3817 ;
  assign n3819 = n1266 ^ n423 ^ 1'b0 ;
  assign n3820 = n1440 | n3819 ;
  assign n3821 = n2701 | n3097 ;
  assign n3822 = n3821 ^ n669 ^ 1'b0 ;
  assign n3823 = ( n959 & n3820 ) | ( n959 & n3822 ) | ( n3820 & n3822 ) ;
  assign n3824 = n1691 ^ n762 ^ 1'b0 ;
  assign n3825 = n904 & n3824 ;
  assign n3828 = ~n681 & n960 ;
  assign n3826 = n791 & ~n994 ;
  assign n3827 = n881 & n3826 ;
  assign n3829 = n3828 ^ n3827 ^ 1'b0 ;
  assign n3830 = n384 & ~n3829 ;
  assign n3831 = x42 & n3830 ;
  assign n3832 = n3831 ^ n1981 ^ 1'b0 ;
  assign n3833 = n179 | n3832 ;
  assign n3834 = n3833 ^ n3225 ^ 1'b0 ;
  assign n3835 = n1656 ^ n359 ^ 1'b0 ;
  assign n3836 = n2389 | n3835 ;
  assign n3837 = n1880 | n3836 ;
  assign n3840 = n784 & n959 ;
  assign n3841 = ~n387 & n1471 ;
  assign n3842 = n1182 | n3841 ;
  assign n3843 = ~n1138 & n2949 ;
  assign n3844 = n3842 & n3843 ;
  assign n3845 = n1666 ^ n664 ^ 1'b0 ;
  assign n3846 = n3113 | n3845 ;
  assign n3847 = n3846 ^ n1174 ^ 1'b0 ;
  assign n3848 = n3641 | n3847 ;
  assign n3849 = n2252 ^ n218 ^ 1'b0 ;
  assign n3850 = ~n3848 & n3849 ;
  assign n3851 = n3850 ^ n2637 ^ 1'b0 ;
  assign n3852 = n3844 | n3851 ;
  assign n3853 = n3840 & ~n3852 ;
  assign n3838 = ~n1913 & n2679 ;
  assign n3839 = n3838 ^ n1448 ^ 1'b0 ;
  assign n3854 = n3853 ^ n3839 ^ 1'b0 ;
  assign n3855 = ~x6 & n768 ;
  assign n3856 = ( ~n471 & n2317 ) | ( ~n471 & n3855 ) | ( n2317 & n3855 ) ;
  assign n3857 = n3856 ^ n987 ^ 1'b0 ;
  assign n3858 = n2670 ^ n1223 ^ 1'b0 ;
  assign n3859 = n3858 ^ n3278 ^ n2890 ;
  assign n3860 = n3145 ^ n651 ^ n147 ;
  assign n3861 = ~n1406 & n2417 ;
  assign n3862 = n3861 ^ n1899 ^ 1'b0 ;
  assign n3863 = x50 & ~n3862 ;
  assign n3864 = n3860 & n3863 ;
  assign n3865 = n2819 & n3864 ;
  assign n3866 = n2471 ^ n1840 ^ 1'b0 ;
  assign n3867 = ~n2710 & n3866 ;
  assign n3868 = n3867 ^ n2844 ^ 1'b0 ;
  assign n3869 = n1130 | n3146 ;
  assign n3870 = n3868 & ~n3869 ;
  assign n3871 = n1026 & n1442 ;
  assign n3872 = n3871 ^ n634 ^ 1'b0 ;
  assign n3873 = n3872 ^ n2587 ^ 1'b0 ;
  assign n3874 = n2490 & ~n3121 ;
  assign n3875 = x59 & n3874 ;
  assign n3876 = ~n1708 & n3875 ;
  assign n3877 = ~n1086 & n3876 ;
  assign n3878 = n1572 & ~n2281 ;
  assign n3879 = ~n2131 & n3878 ;
  assign n3880 = n152 & ~n1485 ;
  assign n3881 = n368 | n1385 ;
  assign n3884 = n632 ^ n472 ^ 1'b0 ;
  assign n3885 = ( n200 & ~n814 ) | ( n200 & n3884 ) | ( ~n814 & n3884 ) ;
  assign n3886 = n1565 ^ n1509 ^ 1'b0 ;
  assign n3887 = n3885 | n3886 ;
  assign n3882 = n1250 ^ n832 ^ 1'b0 ;
  assign n3883 = ~n1053 & n3882 ;
  assign n3888 = n3887 ^ n3883 ^ 1'b0 ;
  assign n3889 = n3881 & n3888 ;
  assign n3890 = ~n2501 & n3889 ;
  assign n3891 = n1943 | n3757 ;
  assign n3892 = n3592 & ~n3891 ;
  assign n3893 = n1241 ^ n243 ^ 1'b0 ;
  assign n3894 = n1606 & ~n3893 ;
  assign n3895 = n3894 ^ n1450 ^ n852 ;
  assign n3896 = ~n517 & n3895 ;
  assign n3897 = n2278 ^ n2116 ^ 1'b0 ;
  assign n3898 = ~n3896 & n3897 ;
  assign n3899 = ( n358 & n446 ) | ( n358 & ~n3898 ) | ( n446 & ~n3898 ) ;
  assign n3900 = n3892 | n3899 ;
  assign n3901 = n3890 & ~n3900 ;
  assign n3902 = n1651 ^ n1094 ^ 1'b0 ;
  assign n3903 = n1488 | n3902 ;
  assign n3904 = n1405 & n1476 ;
  assign n3905 = n3904 ^ n2278 ^ 1'b0 ;
  assign n3906 = n2436 & n3905 ;
  assign n3907 = n3903 & n3906 ;
  assign n3908 = n3907 ^ n468 ^ n190 ;
  assign n3909 = n406 & n585 ;
  assign n3910 = ~n3308 & n3909 ;
  assign n3911 = n2561 & n3596 ;
  assign n3912 = n3910 & n3911 ;
  assign n3920 = n194 & n2417 ;
  assign n3918 = n448 | n852 ;
  assign n3919 = n1308 & ~n3918 ;
  assign n3921 = n3920 ^ n3919 ^ 1'b0 ;
  assign n3913 = n2315 | n3622 ;
  assign n3914 = n1035 & ~n3913 ;
  assign n3915 = n2626 & ~n3914 ;
  assign n3916 = n2305 & n3915 ;
  assign n3917 = n1015 | n3916 ;
  assign n3922 = n3921 ^ n3917 ^ 1'b0 ;
  assign n3923 = n995 | n1657 ;
  assign n3924 = x20 | n3923 ;
  assign n3925 = n3924 ^ n3698 ^ 1'b0 ;
  assign n3926 = n709 | n1089 ;
  assign n3927 = n3926 ^ n1971 ^ 1'b0 ;
  assign n3928 = n288 & ~n2192 ;
  assign n3929 = n1095 ^ n133 ^ 1'b0 ;
  assign n3930 = ~n3928 & n3929 ;
  assign n3931 = n3603 ^ n290 ^ 1'b0 ;
  assign n3932 = n3576 ^ n1135 ^ 1'b0 ;
  assign n3933 = n674 & ~n3932 ;
  assign n3934 = ~n939 & n2927 ;
  assign n3935 = n3934 ^ n3056 ^ 1'b0 ;
  assign n3936 = n2170 | n3288 ;
  assign n3937 = n3257 ^ n2489 ^ 1'b0 ;
  assign n3938 = ~n1579 & n3625 ;
  assign n3939 = n3776 & ~n3938 ;
  assign n3940 = n3939 ^ n1688 ^ 1'b0 ;
  assign n3941 = n587 | n2878 ;
  assign n3942 = n3941 ^ x112 ^ 1'b0 ;
  assign n3943 = ~n2976 & n3942 ;
  assign n3944 = ~n194 & n1570 ;
  assign n3945 = n324 & n1081 ;
  assign n3946 = n3202 ^ n1385 ^ 1'b0 ;
  assign n3947 = n3159 & ~n3946 ;
  assign n3948 = n1231 ^ n456 ^ n147 ;
  assign n3949 = n1198 & n3948 ;
  assign n3950 = n2001 ^ n1121 ^ n874 ;
  assign n3951 = n2399 ^ n377 ^ 1'b0 ;
  assign n3956 = n1425 ^ n438 ^ 1'b0 ;
  assign n3957 = ( n200 & n1747 ) | ( n200 & ~n3956 ) | ( n1747 & ~n3956 ) ;
  assign n3952 = ~n730 & n2483 ;
  assign n3953 = n3952 ^ n1861 ^ 1'b0 ;
  assign n3954 = n478 | n3953 ;
  assign n3955 = n2822 | n3954 ;
  assign n3958 = n3957 ^ n3955 ^ n1517 ;
  assign n3960 = x72 & n1279 ;
  assign n3959 = x93 & ~n2728 ;
  assign n3961 = n3960 ^ n3959 ^ 1'b0 ;
  assign n3962 = ~n866 & n2715 ;
  assign n3963 = n1890 & ~n3463 ;
  assign n3964 = ~n3780 & n3963 ;
  assign n3965 = ( x122 & n565 ) | ( x122 & ~n954 ) | ( n565 & ~n954 ) ;
  assign n3966 = n2235 & n3965 ;
  assign n3967 = n868 | n2172 ;
  assign n3968 = x66 | n3967 ;
  assign n3969 = n3968 ^ n3606 ^ 1'b0 ;
  assign n3970 = ~n389 & n3969 ;
  assign n3971 = n2626 ^ n1794 ^ 1'b0 ;
  assign n3972 = n1308 & ~n3971 ;
  assign n3973 = n541 | n3972 ;
  assign n3974 = n3973 ^ n3483 ^ 1'b0 ;
  assign n3975 = ~n904 & n1746 ;
  assign n3976 = n446 & n1150 ;
  assign n3977 = n2715 ^ n407 ^ 1'b0 ;
  assign n3978 = n3976 & n3977 ;
  assign n3979 = n2022 & ~n3978 ;
  assign n3980 = n3245 & n3979 ;
  assign n3981 = n3980 ^ n3049 ^ 1'b0 ;
  assign n3982 = n913 | n1444 ;
  assign n3983 = ~n1832 & n3982 ;
  assign n3984 = ~n3738 & n3983 ;
  assign n3985 = n3984 ^ n2489 ^ 1'b0 ;
  assign n3986 = n419 | n3985 ;
  assign n3987 = n3986 ^ n1567 ^ 1'b0 ;
  assign n3991 = n620 & ~n1890 ;
  assign n3988 = n710 ^ n438 ^ 1'b0 ;
  assign n3989 = n2489 & n3988 ;
  assign n3990 = ~n1570 & n3989 ;
  assign n3992 = n3991 ^ n3990 ^ 1'b0 ;
  assign n3993 = n2218 & ~n3786 ;
  assign n3994 = n430 & ~n3962 ;
  assign n3995 = ~n3895 & n3994 ;
  assign n3996 = n3925 ^ n2066 ^ 1'b0 ;
  assign n3997 = n2137 & n3996 ;
  assign n3998 = n1336 ^ n575 ^ 1'b0 ;
  assign n3999 = n3998 ^ n1850 ^ 1'b0 ;
  assign n4000 = n3999 ^ n2510 ^ 1'b0 ;
  assign n4001 = n4000 ^ n2985 ^ n1502 ;
  assign n4002 = n4001 ^ n1363 ^ 1'b0 ;
  assign n4006 = n1209 ^ n468 ^ 1'b0 ;
  assign n4005 = ~n324 & n2083 ;
  assign n4004 = n3999 ^ n1992 ^ 1'b0 ;
  assign n4007 = n4006 ^ n4005 ^ n4004 ;
  assign n4003 = n1634 | n3813 ;
  assign n4008 = n4007 ^ n4003 ^ 1'b0 ;
  assign n4009 = n1136 & ~n4008 ;
  assign n4010 = n2806 ^ n204 ^ 1'b0 ;
  assign n4011 = ~n297 & n430 ;
  assign n4012 = n1433 ^ n871 ^ 1'b0 ;
  assign n4013 = n4011 | n4012 ;
  assign n4014 = n506 ^ n368 ^ 1'b0 ;
  assign n4015 = n442 & ~n4014 ;
  assign n4017 = n791 & ~n3056 ;
  assign n4018 = n4017 ^ n3147 ^ 1'b0 ;
  assign n4016 = n138 & n1357 ;
  assign n4019 = n4018 ^ n4016 ^ 1'b0 ;
  assign n4020 = n2201 ^ n2074 ^ 1'b0 ;
  assign n4021 = n741 & n1281 ;
  assign n4022 = n4021 ^ n2948 ^ n600 ;
  assign n4023 = n2639 | n4022 ;
  assign n4024 = n4023 ^ n2038 ^ 1'b0 ;
  assign n4025 = ~n215 & n1198 ;
  assign n4026 = n620 & ~n1620 ;
  assign n4027 = n4026 ^ n1701 ^ 1'b0 ;
  assign n4028 = ( n1933 & n4025 ) | ( n1933 & n4027 ) | ( n4025 & n4027 ) ;
  assign n4029 = ( n319 & ~n1377 ) | ( n319 & n1426 ) | ( ~n1377 & n1426 ) ;
  assign n4030 = n4029 ^ n2095 ^ x10 ;
  assign n4031 = n462 | n1300 ;
  assign n4032 = n4031 ^ n3289 ^ 1'b0 ;
  assign n4033 = ~n202 & n4032 ;
  assign n4034 = n373 | n586 ;
  assign n4035 = n866 | n4034 ;
  assign n4036 = ( n180 & ~n3048 ) | ( n180 & n4035 ) | ( ~n3048 & n4035 ) ;
  assign n4037 = n671 & ~n2441 ;
  assign n4038 = x24 | n4037 ;
  assign n4039 = n4036 | n4038 ;
  assign n4040 = n4039 ^ n1515 ^ 1'b0 ;
  assign n4041 = n4033 & ~n4040 ;
  assign n4046 = n2597 & ~n3885 ;
  assign n4047 = n279 & n4046 ;
  assign n4048 = n1661 & n4047 ;
  assign n4042 = x121 & n569 ;
  assign n4043 = ~x6 & n4042 ;
  assign n4044 = n4043 ^ n1576 ^ 1'b0 ;
  assign n4045 = n632 | n4044 ;
  assign n4049 = n4048 ^ n4045 ^ 1'b0 ;
  assign n4050 = n4041 & n4049 ;
  assign n4051 = n3651 ^ n1761 ^ 1'b0 ;
  assign n4052 = n2827 ^ n1476 ^ 1'b0 ;
  assign n4053 = n1077 ^ n774 ^ 1'b0 ;
  assign n4054 = n4053 ^ n3884 ^ 1'b0 ;
  assign n4055 = n3233 | n4054 ;
  assign n4056 = n1319 | n4055 ;
  assign n4057 = n4056 ^ n3021 ^ 1'b0 ;
  assign n4058 = n275 & ~n4057 ;
  assign n4059 = ~n878 & n3830 ;
  assign n4060 = n4059 ^ n531 ^ 1'b0 ;
  assign n4061 = ~n3921 & n4060 ;
  assign n4062 = n3529 ^ n1901 ^ 1'b0 ;
  assign n4063 = n134 & n4062 ;
  assign n4064 = ( x47 & n1254 ) | ( x47 & n4063 ) | ( n1254 & n4063 ) ;
  assign n4065 = n618 ^ x21 ^ 1'b0 ;
  assign n4066 = ( n157 & n882 ) | ( n157 & n943 ) | ( n882 & n943 ) ;
  assign n4067 = n2611 | n4066 ;
  assign n4068 = n4067 ^ x16 ^ 1'b0 ;
  assign n4069 = n4065 & ~n4068 ;
  assign n4070 = n759 & n2390 ;
  assign n4071 = n928 | n2373 ;
  assign n4072 = n2499 ^ n918 ^ 1'b0 ;
  assign n4073 = n4071 | n4072 ;
  assign n4074 = n458 & ~n513 ;
  assign n4075 = n4074 ^ n781 ^ 1'b0 ;
  assign n4076 = ( n852 & ~n1367 ) | ( n852 & n3217 ) | ( ~n1367 & n3217 ) ;
  assign n4077 = n4075 & n4076 ;
  assign n4080 = n3411 ^ n1765 ^ 1'b0 ;
  assign n4081 = n1797 | n4080 ;
  assign n4079 = x61 & ~n2108 ;
  assign n4082 = n4081 ^ n4079 ^ 1'b0 ;
  assign n4078 = ~n2508 & n2543 ;
  assign n4083 = n4082 ^ n4078 ^ 1'b0 ;
  assign n4086 = x70 & ~n926 ;
  assign n4087 = n3413 & n4086 ;
  assign n4088 = n4087 ^ n1012 ^ 1'b0 ;
  assign n4084 = n3145 ^ n379 ^ 1'b0 ;
  assign n4085 = n4084 ^ n1750 ^ 1'b0 ;
  assign n4089 = n4088 ^ n4085 ^ 1'b0 ;
  assign n4090 = ~n1470 & n1745 ;
  assign n4091 = ( n2647 & n2702 ) | ( n2647 & ~n2813 ) | ( n2702 & ~n2813 ) ;
  assign n4092 = n2464 ^ n2261 ^ 1'b0 ;
  assign n4093 = ~n737 & n4092 ;
  assign n4094 = x6 & ~n771 ;
  assign n4098 = x5 & ~n1040 ;
  assign n4095 = ~n319 & n3463 ;
  assign n4096 = n4095 ^ n3055 ^ 1'b0 ;
  assign n4097 = n3741 | n4096 ;
  assign n4099 = n4098 ^ n4097 ^ 1'b0 ;
  assign n4100 = n569 & ~n690 ;
  assign n4101 = n4100 ^ n3874 ^ 1'b0 ;
  assign n4102 = n1337 ^ n1254 ^ n256 ;
  assign n4103 = x100 & ~n1176 ;
  assign n4104 = n4103 ^ n1105 ^ 1'b0 ;
  assign n4105 = ~n1742 & n4104 ;
  assign n4106 = n3237 ^ n2085 ^ n315 ;
  assign n4107 = n3182 & ~n4106 ;
  assign n4108 = n267 & n3179 ;
  assign n4109 = ~n3898 & n4108 ;
  assign n4111 = n763 & n882 ;
  assign n4110 = n2484 & n3210 ;
  assign n4112 = n4111 ^ n4110 ^ 1'b0 ;
  assign n4113 = ~n615 & n2226 ;
  assign n4114 = n4113 ^ n3240 ^ 1'b0 ;
  assign n4115 = n166 | n4114 ;
  assign n4116 = ( n1953 & n3637 ) | ( n1953 & ~n4115 ) | ( n3637 & ~n4115 ) ;
  assign n4117 = n4112 & ~n4116 ;
  assign n4118 = n4087 ^ n3111 ^ 1'b0 ;
  assign n4119 = n4118 ^ n3786 ^ 1'b0 ;
  assign n4120 = ( n210 & n2866 ) | ( n210 & ~n3839 ) | ( n2866 & ~n3839 ) ;
  assign n4121 = n2659 ^ n1812 ^ 1'b0 ;
  assign n4122 = n849 | n1019 ;
  assign n4123 = n4037 ^ n588 ^ 1'b0 ;
  assign n4124 = n4122 | n4123 ;
  assign n4125 = x52 | n4124 ;
  assign n4126 = n869 ^ n575 ^ 1'b0 ;
  assign n4127 = ~n890 & n4126 ;
  assign n4128 = n1015 & n4127 ;
  assign n4129 = n3848 | n3885 ;
  assign n4130 = n4128 & ~n4129 ;
  assign n4131 = n519 & ~n4130 ;
  assign n4132 = n4131 ^ n2013 ^ 1'b0 ;
  assign n4133 = n4125 & n4132 ;
  assign n4134 = n4121 & n4133 ;
  assign n4135 = n1534 | n2823 ;
  assign n4136 = n3011 ^ n860 ^ 1'b0 ;
  assign n4137 = n4136 ^ n623 ^ 1'b0 ;
  assign n4138 = ~n468 & n2014 ;
  assign n4139 = n4138 ^ n446 ^ 1'b0 ;
  assign n4140 = n1698 & n4139 ;
  assign n4141 = n4140 ^ n3554 ^ 1'b0 ;
  assign n4142 = x64 & ~n1361 ;
  assign n4143 = ( n359 & n586 ) | ( n359 & ~n1134 ) | ( n586 & ~n1134 ) ;
  assign n4144 = n2656 ^ n2156 ^ 1'b0 ;
  assign n4145 = n4143 & n4144 ;
  assign n4146 = n4145 ^ n1722 ^ 1'b0 ;
  assign n4147 = n4142 | n4146 ;
  assign n4148 = n4147 ^ n3448 ^ n648 ;
  assign n4149 = n1788 & ~n4148 ;
  assign n4150 = n1535 | n3844 ;
  assign n4151 = n622 & n3561 ;
  assign n4152 = n3735 ^ n2692 ^ 1'b0 ;
  assign n4153 = ( n175 & n2525 ) | ( n175 & n4152 ) | ( n2525 & n4152 ) ;
  assign n4154 = n4153 ^ n613 ^ 1'b0 ;
  assign n4155 = x40 & ~n4154 ;
  assign n4156 = x23 | n3314 ;
  assign n4157 = n867 & n2419 ;
  assign n4158 = n1083 | n1876 ;
  assign n4159 = n4158 ^ n1935 ^ 1'b0 ;
  assign n4160 = n4159 ^ n305 ^ 1'b0 ;
  assign n4161 = ~n2396 & n4160 ;
  assign n4165 = x89 & n2545 ;
  assign n4166 = n633 & n4165 ;
  assign n4164 = ( ~n777 & n1469 ) | ( ~n777 & n1801 ) | ( n1469 & n1801 ) ;
  assign n4167 = n4166 ^ n4164 ^ 1'b0 ;
  assign n4168 = ( n560 & n1925 ) | ( n560 & n4167 ) | ( n1925 & n4167 ) ;
  assign n4162 = n3709 ^ n816 ^ n801 ;
  assign n4163 = ~n1017 & n4162 ;
  assign n4169 = n4168 ^ n4163 ^ 1'b0 ;
  assign n4170 = n1836 ^ n217 ^ 1'b0 ;
  assign n4171 = ~n1862 & n4170 ;
  assign n4172 = n3675 | n4006 ;
  assign n4173 = n4171 & n4172 ;
  assign n4174 = n4173 ^ n1497 ^ 1'b0 ;
  assign n4175 = n476 ^ n435 ^ 1'b0 ;
  assign n4176 = ( n1396 & n2491 ) | ( n1396 & ~n4175 ) | ( n2491 & ~n4175 ) ;
  assign n4177 = n4176 ^ n2869 ^ 1'b0 ;
  assign n4182 = n2991 ^ x123 ^ 1'b0 ;
  assign n4178 = n1311 & n2001 ;
  assign n4179 = ~n679 & n4178 ;
  assign n4180 = n1576 & ~n4179 ;
  assign n4181 = ~n2831 & n4180 ;
  assign n4183 = n4182 ^ n4181 ^ 1'b0 ;
  assign n4184 = ~n847 & n2170 ;
  assign n4185 = n336 & ~n1701 ;
  assign n4186 = ~n2176 & n4185 ;
  assign n4187 = n3706 & ~n4186 ;
  assign n4188 = n1337 ^ n330 ^ 1'b0 ;
  assign n4189 = x72 & ~n4188 ;
  assign n4190 = ( ~n571 & n673 ) | ( ~n571 & n4189 ) | ( n673 & n4189 ) ;
  assign n4191 = n3704 & n4190 ;
  assign n4192 = n3095 | n4089 ;
  assign n4193 = ( n728 & ~n1100 ) | ( n728 & n1448 ) | ( ~n1100 & n1448 ) ;
  assign n4194 = n3233 & ~n4193 ;
  assign n4195 = n2913 ^ n699 ^ 1'b0 ;
  assign n4196 = n2913 & ~n3138 ;
  assign n4197 = n4196 ^ x57 ^ 1'b0 ;
  assign n4198 = n732 | n2619 ;
  assign n4199 = n645 | n4198 ;
  assign n4200 = n3716 ^ n2479 ^ 1'b0 ;
  assign n4201 = n414 | n466 ;
  assign n4202 = n2776 & ~n2863 ;
  assign n4203 = n4202 ^ n3241 ^ 1'b0 ;
  assign n4204 = n983 | n4203 ;
  assign n4205 = n3741 ^ n2250 ^ 1'b0 ;
  assign n4206 = n3136 & ~n3336 ;
  assign n4207 = ~n3715 & n4206 ;
  assign n4208 = n3615 | n4007 ;
  assign n4209 = n884 & n1600 ;
  assign n4210 = n4209 ^ n732 ^ 1'b0 ;
  assign n4211 = n359 & n4210 ;
  assign n4212 = ~n672 & n4211 ;
  assign n4213 = n2740 & n4212 ;
  assign n4214 = n1937 & ~n2204 ;
  assign n4215 = n4214 ^ n2998 ^ 1'b0 ;
  assign n4216 = ( n1046 & n2839 ) | ( n1046 & n3828 ) | ( n2839 & n3828 ) ;
  assign n4217 = n4216 ^ n4159 ^ 1'b0 ;
  assign n4218 = n3240 & n4217 ;
  assign n4219 = n4215 & n4218 ;
  assign n4220 = n4213 | n4219 ;
  assign n4221 = n805 & ~n4220 ;
  assign n4222 = ~n3346 & n3953 ;
  assign n4223 = n706 | n2718 ;
  assign n4224 = n4223 ^ n815 ^ 1'b0 ;
  assign n4225 = n2021 & ~n4224 ;
  assign n4226 = ~n2426 & n3920 ;
  assign n4227 = n3233 & n4226 ;
  assign n4228 = ( n163 & n1333 ) | ( n163 & n1392 ) | ( n1333 & n1392 ) ;
  assign n4229 = n3006 ^ n3001 ^ 1'b0 ;
  assign n4230 = n4228 & n4229 ;
  assign n4231 = n1465 | n2054 ;
  assign n4232 = n4231 ^ n925 ^ 1'b0 ;
  assign n4233 = n2070 | n4232 ;
  assign n4234 = x86 & ~n3572 ;
  assign n4235 = n4234 ^ n2932 ^ 1'b0 ;
  assign n4236 = n468 & n3830 ;
  assign n4237 = n641 | n4236 ;
  assign n4238 = n1488 ^ n767 ^ 1'b0 ;
  assign n4239 = n4238 ^ n389 ^ 1'b0 ;
  assign n4240 = n4237 & n4239 ;
  assign n4241 = n3896 ^ n784 ^ 1'b0 ;
  assign n4242 = n3414 & ~n4241 ;
  assign n4243 = ( n1979 & n2551 ) | ( n1979 & n3237 ) | ( n2551 & n3237 ) ;
  assign n4244 = n420 & n3850 ;
  assign n4245 = x105 & ~n1005 ;
  assign n4246 = n4245 ^ x52 ^ 1'b0 ;
  assign n4247 = n4246 ^ n195 ^ 1'b0 ;
  assign n4248 = x103 & n1432 ;
  assign n4249 = n4248 ^ n3613 ^ 1'b0 ;
  assign n4250 = n2859 & ~n4249 ;
  assign n4251 = ~n220 & n4250 ;
  assign n4252 = n1553 | n3785 ;
  assign n4253 = n3792 & ~n4252 ;
  assign n4254 = n3687 ^ n820 ^ 1'b0 ;
  assign n4255 = n1439 & ~n4254 ;
  assign n4256 = n166 | n3973 ;
  assign n4257 = n4256 ^ n445 ^ 1'b0 ;
  assign n4258 = n900 & n4257 ;
  assign n4259 = n4258 ^ n738 ^ 1'b0 ;
  assign n4260 = n756 & n3546 ;
  assign n4261 = ( n3283 & n3937 ) | ( n3283 & ~n4139 ) | ( n3937 & ~n4139 ) ;
  assign n4262 = x34 | n745 ;
  assign n4263 = ~n3898 & n4262 ;
  assign n4264 = n1331 & ~n3869 ;
  assign n4265 = n1003 & ~n4264 ;
  assign n4266 = n1681 & ~n1853 ;
  assign n4267 = n562 & n884 ;
  assign n4268 = n1199 & n4267 ;
  assign n4269 = ( ~x64 & n213 ) | ( ~x64 & n1092 ) | ( n213 & n1092 ) ;
  assign n4270 = ~n152 & n4269 ;
  assign n4271 = ~n753 & n4270 ;
  assign n4272 = n539 | n2564 ;
  assign n4273 = n1266 & ~n4272 ;
  assign n4274 = n4122 | n4273 ;
  assign n4275 = n2626 | n4274 ;
  assign n4276 = ~n4271 & n4275 ;
  assign n4277 = n4276 ^ n2171 ^ 1'b0 ;
  assign n4278 = n281 | n4277 ;
  assign n4279 = n732 & ~n4278 ;
  assign n4280 = n1103 & ~n4279 ;
  assign n4281 = n1147 & n1680 ;
  assign n4282 = n238 | n3580 ;
  assign n4283 = n4281 & ~n4282 ;
  assign n4284 = n1567 & ~n2201 ;
  assign n4285 = ~n437 & n4284 ;
  assign n4286 = n1279 | n4285 ;
  assign n4287 = n231 & ~n4286 ;
  assign n4289 = ~n861 & n1526 ;
  assign n4288 = n2583 & ~n3006 ;
  assign n4290 = n4289 ^ n4288 ^ 1'b0 ;
  assign n4291 = n4290 ^ n2259 ^ 1'b0 ;
  assign n4292 = n166 | n4291 ;
  assign n4293 = n616 & ~n3631 ;
  assign n4294 = n597 & ~n3820 ;
  assign n4295 = ~x55 & n4294 ;
  assign n4296 = n2189 ^ n829 ^ 1'b0 ;
  assign n4297 = n3209 ^ n1154 ^ 1'b0 ;
  assign n4298 = n530 & n808 ;
  assign n4299 = ~n3998 & n4298 ;
  assign n4300 = ~x47 & n838 ;
  assign n4301 = n2401 ^ n1728 ^ n1199 ;
  assign n4302 = ( n1487 & n4216 ) | ( n1487 & ~n4301 ) | ( n4216 & ~n4301 ) ;
  assign n4303 = ~n1386 & n2567 ;
  assign n4304 = n213 & n2855 ;
  assign n4305 = n809 ^ n292 ^ 1'b0 ;
  assign n4306 = n4305 ^ n718 ^ 1'b0 ;
  assign n4307 = ~n1247 & n4306 ;
  assign n4308 = n4307 ^ n1615 ^ 1'b0 ;
  assign n4309 = n3166 ^ n2140 ^ 1'b0 ;
  assign n4310 = ~n3890 & n4309 ;
  assign n4311 = n1021 & ~n3918 ;
  assign n4312 = ~n4263 & n4311 ;
  assign n4313 = n2647 & n4312 ;
  assign n4314 = n2675 ^ n1353 ^ 1'b0 ;
  assign n4315 = ( n188 & n556 ) | ( n188 & ~n1109 ) | ( n556 & ~n1109 ) ;
  assign n4316 = n4315 ^ n1821 ^ 1'b0 ;
  assign n4317 = x31 & ~n1982 ;
  assign n4318 = n4316 & n4317 ;
  assign n4319 = n678 & ~n1097 ;
  assign n4320 = n4319 ^ n217 ^ 1'b0 ;
  assign n4321 = n1331 ^ n1295 ^ 1'b0 ;
  assign n4322 = n989 & ~n4321 ;
  assign n4323 = ~n2562 & n4322 ;
  assign n4324 = n455 | n4323 ;
  assign n4325 = ( ~n2474 & n3784 ) | ( ~n2474 & n4324 ) | ( n3784 & n4324 ) ;
  assign n4326 = n632 & ~n4150 ;
  assign n4327 = n4326 ^ n368 ^ 1'b0 ;
  assign n4328 = x103 & ~n3965 ;
  assign n4329 = n4328 ^ n1654 ^ 1'b0 ;
  assign n4330 = ( n506 & n3539 ) | ( n506 & n4329 ) | ( n3539 & n4329 ) ;
  assign n4331 = n3945 ^ n1152 ^ 1'b0 ;
  assign n4332 = n479 & n4106 ;
  assign n4333 = n4332 ^ n4205 ^ 1'b0 ;
  assign n4334 = n1692 | n2951 ;
  assign n4336 = n1865 ^ n1276 ^ 1'b0 ;
  assign n4335 = n1913 | n2828 ;
  assign n4337 = n4336 ^ n4335 ^ n3276 ;
  assign n4338 = n2853 & n3547 ;
  assign n4339 = n297 & ~n876 ;
  assign n4340 = n4339 ^ n1192 ^ 1'b0 ;
  assign n4341 = n4340 ^ n556 ^ 1'b0 ;
  assign n4342 = ~n657 & n4341 ;
  assign n4343 = n496 ^ x79 ^ 1'b0 ;
  assign n4344 = ~n299 & n4343 ;
  assign n4345 = ( n3162 & n4342 ) | ( n3162 & ~n4344 ) | ( n4342 & ~n4344 ) ;
  assign n4346 = n2095 ^ n2048 ^ 1'b0 ;
  assign n4347 = n3883 & ~n4346 ;
  assign n4348 = n1999 & n4347 ;
  assign n4352 = n2931 & n3400 ;
  assign n4349 = x111 & n1457 ;
  assign n4350 = n1761 & n4349 ;
  assign n4351 = n4350 ^ n1720 ^ n1562 ;
  assign n4353 = n4352 ^ n4351 ^ 1'b0 ;
  assign n4354 = ( ~x6 & n3419 ) | ( ~x6 & n3973 ) | ( n3419 & n3973 ) ;
  assign n4355 = n3257 ^ n384 ^ 1'b0 ;
  assign n4356 = x56 & n1033 ;
  assign n4357 = ~x16 & n4356 ;
  assign n4358 = n4357 ^ n1830 ^ 1'b0 ;
  assign n4359 = ~n1913 & n4358 ;
  assign n4360 = n4359 ^ n1370 ^ 1'b0 ;
  assign n4361 = n2412 ^ n1902 ^ 1'b0 ;
  assign n4362 = ~n682 & n4361 ;
  assign n4363 = n809 & n1188 ;
  assign n4364 = n4363 ^ n732 ^ 1'b0 ;
  assign n4365 = n2484 & ~n4364 ;
  assign n4366 = n3846 ^ n1162 ^ 1'b0 ;
  assign n4367 = ~n1631 & n1801 ;
  assign n4368 = n1895 & n4367 ;
  assign n4369 = n2618 & n4368 ;
  assign n4370 = n2370 & ~n3998 ;
  assign n4371 = n3062 | n4370 ;
  assign n4372 = n174 | n4371 ;
  assign n4373 = n4048 & ~n4372 ;
  assign n4374 = n4373 ^ n1526 ^ 1'b0 ;
  assign n4375 = ~n180 & n4374 ;
  assign n4376 = n250 | n299 ;
  assign n4377 = n4376 ^ x24 ^ 1'b0 ;
  assign n4378 = n675 & n4377 ;
  assign n4379 = n4378 ^ n2712 ^ 1'b0 ;
  assign n4380 = n2490 ^ n1641 ^ 1'b0 ;
  assign n4381 = n4380 ^ n2262 ^ 1'b0 ;
  assign n4382 = ( n3659 & ~n4379 ) | ( n3659 & n4381 ) | ( ~n4379 & n4381 ) ;
  assign n4383 = n1008 | n3239 ;
  assign n4384 = n4383 ^ n560 ^ 1'b0 ;
  assign n4385 = n4384 ^ n1788 ^ 1'b0 ;
  assign n4386 = n1529 & n4385 ;
  assign n4387 = ( n1910 & n3784 ) | ( n1910 & n4386 ) | ( n3784 & n4386 ) ;
  assign n4388 = n803 & ~n1747 ;
  assign n4389 = ~x35 & n232 ;
  assign n4390 = n4389 ^ n3294 ^ 1'b0 ;
  assign n4391 = n1086 | n4390 ;
  assign n4392 = n3938 ^ n2634 ^ 1'b0 ;
  assign n4393 = ~n1134 & n4392 ;
  assign n4394 = n1338 | n4314 ;
  assign n4395 = n287 & n640 ;
  assign n4396 = ~n721 & n4395 ;
  assign n4397 = x101 & n2913 ;
  assign n4398 = n1661 & n4397 ;
  assign n4399 = n4398 ^ n481 ^ 1'b0 ;
  assign n4400 = ~n755 & n4399 ;
  assign n4401 = ~n680 & n3246 ;
  assign n4402 = ~n4400 & n4401 ;
  assign n4403 = ( n835 & n2605 ) | ( n835 & ~n3582 ) | ( n2605 & ~n3582 ) ;
  assign n4404 = n4045 ^ n656 ^ 1'b0 ;
  assign n4405 = ~n4403 & n4404 ;
  assign n4406 = n2647 ^ n1556 ^ 1'b0 ;
  assign n4407 = n4405 & n4406 ;
  assign n4408 = n3554 ^ n1679 ^ 1'b0 ;
  assign n4409 = n4408 ^ n3571 ^ n708 ;
  assign n4410 = n2463 ^ n1028 ^ 1'b0 ;
  assign n4411 = n4159 | n4410 ;
  assign n4412 = n4411 ^ n3106 ^ 1'b0 ;
  assign n4413 = x5 & n1097 ;
  assign n4414 = n2250 & n4413 ;
  assign n4415 = n1136 & n4414 ;
  assign n4416 = n1124 & n2182 ;
  assign n4417 = n2896 & ~n4416 ;
  assign n4418 = n4417 ^ n1759 ^ 1'b0 ;
  assign n4419 = ( ~n1202 & n1867 ) | ( ~n1202 & n2442 ) | ( n1867 & n2442 ) ;
  assign n4420 = n4419 ^ n1993 ^ 1'b0 ;
  assign n4421 = n4420 ^ n2261 ^ 1'b0 ;
  assign n4422 = n4418 & n4421 ;
  assign n4423 = n1053 | n4422 ;
  assign n4424 = x14 & ~n4423 ;
  assign n4425 = n559 & n3733 ;
  assign n4426 = n4425 ^ n1174 ^ 1'b0 ;
  assign n4427 = n4426 ^ n1005 ^ 1'b0 ;
  assign n4428 = n2378 ^ n2130 ^ 1'b0 ;
  assign n4429 = n141 & ~n3304 ;
  assign n4430 = n900 | n4037 ;
  assign n4431 = n4430 ^ n2845 ^ 1'b0 ;
  assign n4432 = n4429 & n4431 ;
  assign n4433 = ~n3239 & n4432 ;
  assign n4434 = n4433 ^ n808 ^ 1'b0 ;
  assign n4435 = n277 & ~n2028 ;
  assign n4436 = n4435 ^ n487 ^ 1'b0 ;
  assign n4437 = ~n3364 & n3904 ;
  assign n4438 = n2146 | n4437 ;
  assign n4439 = n1656 ^ n1095 ^ 1'b0 ;
  assign n4440 = n1170 & ~n4439 ;
  assign n4441 = n4440 ^ n1631 ^ 1'b0 ;
  assign n4442 = n1304 | n3940 ;
  assign n4443 = n3240 | n4442 ;
  assign n4444 = n2270 & ~n3952 ;
  assign n4445 = n1488 & n4444 ;
  assign n4446 = n2049 ^ n786 ^ 1'b0 ;
  assign n4447 = n1189 & ~n4446 ;
  assign n4448 = n1527 & n4447 ;
  assign n4449 = n4448 ^ n1889 ^ n1369 ;
  assign n4450 = ~n2158 & n4449 ;
  assign n4451 = ( n1465 & ~n2656 ) | ( n1465 & n4450 ) | ( ~n2656 & n4450 ) ;
  assign n4452 = ~n1467 & n4215 ;
  assign n4453 = n2151 & n3583 ;
  assign n4454 = n3662 & n4453 ;
  assign n4455 = n1189 & n2963 ;
  assign n4456 = n4455 ^ n1390 ^ 1'b0 ;
  assign n4457 = n3046 ^ n1429 ^ 1'b0 ;
  assign n4458 = n459 & ~n4457 ;
  assign n4459 = x80 | n1759 ;
  assign n4460 = n1578 ^ n874 ^ 1'b0 ;
  assign n4461 = ~n1502 & n4460 ;
  assign n4462 = n2286 & n4461 ;
  assign n4463 = n4462 ^ n517 ^ 1'b0 ;
  assign n4464 = n4463 ^ n2396 ^ 1'b0 ;
  assign n4465 = n3113 | n4464 ;
  assign n4466 = n3304 ^ n680 ^ 1'b0 ;
  assign n4467 = ~n480 & n4466 ;
  assign n4468 = n2527 ^ n2484 ^ n1651 ;
  assign n4469 = n4468 ^ n1945 ^ 1'b0 ;
  assign n4470 = n4467 & ~n4469 ;
  assign n4471 = ~n278 & n2272 ;
  assign n4472 = n855 ^ n493 ^ 1'b0 ;
  assign n4473 = ~n1574 & n1748 ;
  assign n4474 = n4473 ^ n3198 ^ 1'b0 ;
  assign n4475 = n1120 & n4452 ;
  assign n4476 = n4475 ^ n1700 ^ 1'b0 ;
  assign n4477 = n175 | n3657 ;
  assign n4478 = n2098 ^ n222 ^ 1'b0 ;
  assign n4479 = n1743 & n3982 ;
  assign n4480 = ~n3982 & n4479 ;
  assign n4481 = n884 & n1627 ;
  assign n4482 = n1229 ^ n530 ^ 1'b0 ;
  assign n4483 = ~n1301 & n4482 ;
  assign n4484 = n4483 ^ n505 ^ 1'b0 ;
  assign n4485 = n1096 & ~n4484 ;
  assign n4486 = n2593 & n4485 ;
  assign n4487 = x54 & n642 ;
  assign n4488 = n4487 ^ n827 ^ 1'b0 ;
  assign n4489 = n2148 | n3868 ;
  assign n4490 = n4489 ^ n3099 ^ 1'b0 ;
  assign n4491 = n4488 | n4490 ;
  assign n4492 = n391 & n3514 ;
  assign n4493 = ~n1052 & n4492 ;
  assign n4496 = n541 & ~n1534 ;
  assign n4494 = n2537 ^ n498 ^ 1'b0 ;
  assign n4495 = n1600 & n4494 ;
  assign n4497 = n4496 ^ n4495 ^ 1'b0 ;
  assign n4498 = n3987 | n4497 ;
  assign n4501 = n1575 & n1754 ;
  assign n4502 = ~n1572 & n4501 ;
  assign n4500 = ~n1208 & n2221 ;
  assign n4503 = n4502 ^ n4500 ^ 1'b0 ;
  assign n4504 = ~n3601 & n4503 ;
  assign n4505 = n4504 ^ n2866 ^ 1'b0 ;
  assign n4506 = n815 ^ n276 ^ 1'b0 ;
  assign n4507 = n817 | n4506 ;
  assign n4508 = n4505 & n4507 ;
  assign n4509 = n4508 ^ n1697 ^ 1'b0 ;
  assign n4499 = n2270 & ~n2884 ;
  assign n4510 = n4509 ^ n4499 ^ 1'b0 ;
  assign n4511 = n1540 & ~n3033 ;
  assign n4512 = n487 | n3719 ;
  assign n4520 = ( n1711 & n2281 ) | ( n1711 & n2660 ) | ( n2281 & n2660 ) ;
  assign n4513 = n475 & ~n2782 ;
  assign n4514 = n4513 ^ n1776 ^ 1'b0 ;
  assign n4515 = n4126 & n4514 ;
  assign n4516 = n4515 ^ n421 ^ 1'b0 ;
  assign n4517 = ( ~n943 & n1772 ) | ( ~n943 & n3855 ) | ( n1772 & n3855 ) ;
  assign n4518 = n4516 & n4517 ;
  assign n4519 = ~n3709 & n4518 ;
  assign n4521 = n4520 ^ n4519 ^ 1'b0 ;
  assign n4522 = x34 & ~n3019 ;
  assign n4523 = n167 | n4522 ;
  assign n4524 = ~x59 & n2597 ;
  assign n4525 = n3701 & ~n4524 ;
  assign n4526 = n4525 ^ n362 ^ 1'b0 ;
  assign n4527 = n2900 ^ n2074 ^ 1'b0 ;
  assign n4528 = n678 ^ x8 ^ 1'b0 ;
  assign n4529 = n3321 ^ n1824 ^ 1'b0 ;
  assign n4530 = ~n4528 & n4529 ;
  assign n4531 = ( ~n876 & n1420 ) | ( ~n876 & n4530 ) | ( n1420 & n4530 ) ;
  assign n4532 = n2567 | n4531 ;
  assign n4533 = n4527 | n4532 ;
  assign n4534 = n675 | n4533 ;
  assign n4535 = n803 | n4043 ;
  assign n4536 = n4416 & ~n4535 ;
  assign n4537 = n3159 & ~n4536 ;
  assign n4538 = n841 & n4537 ;
  assign n4539 = n3744 & ~n4538 ;
  assign n4540 = ~n3982 & n4539 ;
  assign n4541 = n667 | n2991 ;
  assign n4542 = n496 | n3100 ;
  assign n4543 = n471 & n2091 ;
  assign n4544 = x72 & ~n1327 ;
  assign n4545 = ~n1623 & n4544 ;
  assign n4546 = n2674 & n4423 ;
  assign n4547 = n4545 & n4546 ;
  assign n4548 = n4351 ^ n3068 ^ 1'b0 ;
  assign n4549 = ~n2281 & n2580 ;
  assign n4550 = n2028 | n2224 ;
  assign n4551 = n836 & ~n4550 ;
  assign n4552 = ~n1390 & n1575 ;
  assign n4553 = n4551 & n4552 ;
  assign n4554 = n281 | n4553 ;
  assign n4555 = n978 & ~n1053 ;
  assign n4556 = n4555 ^ n3082 ^ n157 ;
  assign n4557 = ~n1831 & n4556 ;
  assign n4558 = n4557 ^ n1761 ^ 1'b0 ;
  assign n4559 = x4 & ~n2206 ;
  assign n4560 = n4559 ^ n397 ^ 1'b0 ;
  assign n4561 = x23 & ~n4560 ;
  assign n4562 = ( n4405 & n4558 ) | ( n4405 & n4561 ) | ( n4558 & n4561 ) ;
  assign n4566 = n2240 & ~n3840 ;
  assign n4563 = x24 & n792 ;
  assign n4564 = n4563 ^ n531 ^ 1'b0 ;
  assign n4565 = ~n1592 & n4564 ;
  assign n4567 = n4566 ^ n4565 ^ 1'b0 ;
  assign n4568 = n4567 ^ n1377 ^ n762 ;
  assign n4569 = n2949 ^ n2699 ^ 1'b0 ;
  assign n4570 = n1045 ^ x13 ^ 1'b0 ;
  assign n4571 = n1470 & n4570 ;
  assign n4572 = n1871 & ~n4571 ;
  assign n4573 = n1044 ^ n620 ^ 1'b0 ;
  assign n4574 = n4025 & ~n4573 ;
  assign n4575 = n4574 ^ n3839 ^ n188 ;
  assign n4576 = ~n1037 & n4575 ;
  assign n4577 = n2896 ^ n511 ^ 1'b0 ;
  assign n4578 = ~n4224 & n4577 ;
  assign n4579 = n1100 ^ n774 ^ 1'b0 ;
  assign n4580 = n4579 ^ n2751 ^ 1'b0 ;
  assign n4581 = n3445 & n4580 ;
  assign n4582 = n1066 & ~n1268 ;
  assign n4583 = n4582 ^ n725 ^ 1'b0 ;
  assign n4584 = n2031 ^ n588 ^ 1'b0 ;
  assign n4585 = n4583 | n4584 ;
  assign n4586 = ~n152 & n2442 ;
  assign n4587 = n2561 ^ n754 ^ 1'b0 ;
  assign n4588 = n4586 | n4587 ;
  assign n4589 = n1527 ^ n1192 ^ n719 ;
  assign n4590 = n947 ^ n382 ^ 1'b0 ;
  assign n4591 = n4590 ^ n3131 ^ 1'b0 ;
  assign n4592 = n3041 | n4591 ;
  assign n4593 = ~n4589 & n4592 ;
  assign n4597 = n601 & ~n2426 ;
  assign n4594 = x69 & ~n1884 ;
  assign n4595 = n4594 ^ x95 ^ 1'b0 ;
  assign n4596 = n4595 ^ x69 ^ x29 ;
  assign n4598 = n4597 ^ n4596 ^ 1'b0 ;
  assign n4599 = n205 & ~n2293 ;
  assign n4600 = n4599 ^ n4420 ^ 1'b0 ;
  assign n4601 = n1755 ^ n604 ^ 1'b0 ;
  assign n4602 = n4600 | n4601 ;
  assign n4603 = n2987 ^ n569 ^ 1'b0 ;
  assign n4604 = n3295 ^ n517 ^ 1'b0 ;
  assign n4605 = n4604 ^ n3872 ^ n276 ;
  assign n4606 = ~n391 & n2165 ;
  assign n4607 = n4477 ^ n1027 ^ 1'b0 ;
  assign n4608 = n4606 | n4607 ;
  assign n4609 = n143 | n1670 ;
  assign n4610 = ~n4354 & n4609 ;
  assign n4611 = n2886 ^ n2683 ^ 1'b0 ;
  assign n4612 = n4611 ^ n2647 ^ 1'b0 ;
  assign n4613 = n2486 ^ n2324 ^ 1'b0 ;
  assign n4614 = n2452 & n3637 ;
  assign n4615 = n808 & ~n4614 ;
  assign n4616 = n4615 ^ n1351 ^ 1'b0 ;
  assign n4617 = n239 & n2659 ;
  assign n4618 = n3295 & n4617 ;
  assign n4619 = n1491 & ~n4126 ;
  assign n4620 = n2419 | n4619 ;
  assign n4621 = n4620 ^ n660 ^ 1'b0 ;
  assign n4622 = n3048 ^ n2203 ^ n988 ;
  assign n4623 = n3546 & ~n4622 ;
  assign n4624 = n2758 | n4623 ;
  assign n4625 = n861 | n1202 ;
  assign n4626 = n4625 ^ n192 ^ 1'b0 ;
  assign n4627 = n143 & n4626 ;
  assign n4628 = n2240 & n4627 ;
  assign n4629 = n2287 ^ n930 ^ 1'b0 ;
  assign n4630 = ~n2456 & n4629 ;
  assign n4631 = n4628 | n4630 ;
  assign n4632 = n2953 ^ n225 ^ 1'b0 ;
  assign n4633 = x22 | n2824 ;
  assign n4634 = n1697 & n4633 ;
  assign n4635 = n4632 & n4634 ;
  assign n4636 = n479 | n1383 ;
  assign n4637 = ~n3114 & n4155 ;
  assign n4638 = n4636 & n4637 ;
  assign n4639 = ( n442 & ~n630 ) | ( n442 & n1077 ) | ( ~n630 & n1077 ) ;
  assign n4640 = n4279 | n4639 ;
  assign n4641 = n3678 ^ n1753 ^ 1'b0 ;
  assign n4642 = n814 & ~n1592 ;
  assign n4643 = ~n511 & n4642 ;
  assign n4644 = n4643 ^ x44 ^ 1'b0 ;
  assign n4645 = n4644 ^ n1973 ^ 1'b0 ;
  assign n4646 = n2515 & ~n4645 ;
  assign n4647 = n4641 & n4646 ;
  assign n4648 = n845 | n1410 ;
  assign n4649 = n530 & n4519 ;
  assign n4650 = n575 & n741 ;
  assign n4651 = n2560 ^ n2127 ^ 1'b0 ;
  assign n4652 = ~n3842 & n4651 ;
  assign n4653 = n2759 ^ n1616 ^ 1'b0 ;
  assign n4654 = n4073 | n4653 ;
  assign n4655 = n4652 | n4654 ;
  assign n4657 = n756 & ~n4595 ;
  assign n4658 = n4657 ^ n1904 ^ n469 ;
  assign n4659 = n1609 & n4658 ;
  assign n4660 = n3521 & ~n4659 ;
  assign n4661 = n4660 ^ n2566 ^ 1'b0 ;
  assign n4656 = n1147 & ~n4213 ;
  assign n4662 = n4661 ^ n4656 ^ 1'b0 ;
  assign n4663 = ~n1089 & n4662 ;
  assign n4664 = ~n3975 & n4663 ;
  assign n4665 = n3706 ^ n277 ^ 1'b0 ;
  assign n4666 = n1179 ^ n801 ^ 1'b0 ;
  assign n4667 = n1222 & ~n2656 ;
  assign n4668 = n4667 ^ n2131 ^ 1'b0 ;
  assign n4669 = n4418 & n4668 ;
  assign n4670 = n1566 | n2109 ;
  assign n4671 = n710 & ~n4670 ;
  assign n4672 = n1351 & n1858 ;
  assign n4673 = ~n1643 & n4672 ;
  assign n4674 = n585 & ~n4673 ;
  assign n4675 = n4671 & n4674 ;
  assign n4676 = n1411 ^ n404 ^ 1'b0 ;
  assign n4677 = n1266 ^ n865 ^ 1'b0 ;
  assign n4678 = ~n1201 & n4677 ;
  assign n4679 = x17 & n3179 ;
  assign n4680 = n973 | n1258 ;
  assign n4681 = n4680 ^ n531 ^ 1'b0 ;
  assign n4682 = ~n4679 & n4681 ;
  assign n4683 = n4678 & n4682 ;
  assign n4684 = n4281 & ~n4683 ;
  assign n4685 = n890 | n1714 ;
  assign n4686 = n4684 | n4685 ;
  assign n4687 = n1410 | n3869 ;
  assign n4688 = n4687 ^ n2312 ^ 1'b0 ;
  assign n4689 = n4688 ^ n266 ^ 1'b0 ;
  assign n4690 = ~n3120 & n4689 ;
  assign n4691 = n3590 ^ n2187 ^ 1'b0 ;
  assign n4692 = ~n2066 & n4691 ;
  assign n4693 = n4692 ^ n1191 ^ 1'b0 ;
  assign n4694 = n1642 | n4235 ;
  assign n4695 = n4255 ^ n1926 ^ 1'b0 ;
  assign n4696 = n1217 & ~n4695 ;
  assign n4697 = n983 & n4370 ;
  assign n4698 = ~n159 & n2608 ;
  assign n4700 = n2115 ^ n2011 ^ n642 ;
  assign n4701 = n294 & ~n4700 ;
  assign n4699 = n3716 & ~n4426 ;
  assign n4702 = n4701 ^ n4699 ^ 1'b0 ;
  assign n4703 = ( n143 & n417 ) | ( n143 & n3616 ) | ( n417 & n3616 ) ;
  assign n4704 = ~n863 & n4703 ;
  assign n4705 = ~n1361 & n4704 ;
  assign n4706 = n3461 | n4705 ;
  assign n4707 = n4702 | n4706 ;
  assign n4708 = n292 & n2254 ;
  assign n4709 = ~n1705 & n2793 ;
  assign n4710 = ~n1962 & n4709 ;
  assign n4711 = n4481 ^ n937 ^ 1'b0 ;
  assign n4712 = n4710 | n4711 ;
  assign n4713 = ~n2026 & n2373 ;
  assign n4714 = n4713 ^ n571 ^ 1'b0 ;
  assign n4715 = n1256 & n2568 ;
  assign n4716 = n4715 ^ n461 ^ 1'b0 ;
  assign n4717 = n3159 ^ n327 ^ 1'b0 ;
  assign n4718 = n4717 ^ n2031 ^ 1'b0 ;
  assign n4719 = n2026 | n4718 ;
  assign n4723 = n3128 & ~n4053 ;
  assign n4722 = n795 | n1853 ;
  assign n4720 = n1634 | n1750 ;
  assign n4721 = n4720 ^ n901 ^ 1'b0 ;
  assign n4724 = n4723 ^ n4722 ^ n4721 ;
  assign n4725 = n2543 & ~n2559 ;
  assign n4726 = n1661 & n4725 ;
  assign n4727 = n1828 ^ x75 ^ 1'b0 ;
  assign n4728 = n4727 ^ n256 ^ 1'b0 ;
  assign n4729 = n4726 & n4728 ;
  assign n4730 = ( n1840 & n1878 ) | ( n1840 & ~n1972 ) | ( n1878 & ~n1972 ) ;
  assign n4731 = n1433 ^ n1412 ^ 1'b0 ;
  assign n4733 = ( ~x74 & n2132 ) | ( ~x74 & n4727 ) | ( n2132 & n4727 ) ;
  assign n4732 = n496 & ~n2569 ;
  assign n4734 = n4733 ^ n4732 ^ 1'b0 ;
  assign n4737 = n587 & ~n2319 ;
  assign n4738 = n1761 & ~n4737 ;
  assign n4735 = n2492 & n2639 ;
  assign n4736 = ~n331 & n4735 ;
  assign n4739 = n4738 ^ n4736 ^ 1'b0 ;
  assign n4740 = n530 & n1479 ;
  assign n4742 = n3097 ^ x62 ^ 1'b0 ;
  assign n4741 = n358 | n398 ;
  assign n4743 = n4742 ^ n4741 ^ 1'b0 ;
  assign n4744 = ~n1761 & n2952 ;
  assign n4745 = n4744 ^ n3114 ^ 1'b0 ;
  assign n4746 = ~n4743 & n4745 ;
  assign n4747 = n4746 ^ n3908 ^ 1'b0 ;
  assign n4748 = n303 | n1174 ;
  assign n4749 = n2135 | n3953 ;
  assign n4750 = n2776 | n4749 ;
  assign n4751 = n762 & ~n3706 ;
  assign n4752 = ~n2266 & n4751 ;
  assign n4753 = n4752 ^ n575 ^ 1'b0 ;
  assign n4754 = n2412 ^ n1217 ^ 1'b0 ;
  assign n4755 = n2328 | n4754 ;
  assign n4756 = n4755 ^ n1722 ^ 1'b0 ;
  assign n4757 = ~n1454 & n4756 ;
  assign n4758 = n4528 ^ n1124 ^ 1'b0 ;
  assign n4759 = n296 | n4758 ;
  assign n4760 = n4759 ^ n4166 ^ 1'b0 ;
  assign n4761 = n4757 & n4760 ;
  assign n4762 = ~n1865 & n3993 ;
  assign n4763 = n4762 ^ n1412 ^ 1'b0 ;
  assign n4764 = n749 ^ n676 ^ 1'b0 ;
  assign n4765 = n3066 & ~n4764 ;
  assign n4766 = n2257 | n4765 ;
  assign n4767 = ~n1746 & n4766 ;
  assign n4770 = ~n1281 & n1623 ;
  assign n4771 = n2293 & n4770 ;
  assign n4768 = n1033 ^ n959 ^ 1'b0 ;
  assign n4769 = n3470 & n4768 ;
  assign n4772 = n4771 ^ n4769 ^ 1'b0 ;
  assign n4773 = ~n2349 & n4772 ;
  assign n4774 = n741 ^ n571 ^ 1'b0 ;
  assign n4775 = x9 & ~n308 ;
  assign n4776 = n4775 ^ n3869 ^ n1394 ;
  assign n4777 = n4398 & n4776 ;
  assign n4778 = n3547 ^ n530 ^ 1'b0 ;
  assign n4779 = n3998 ^ n3283 ^ 1'b0 ;
  assign n4780 = n4779 ^ n3424 ^ 1'b0 ;
  assign n4781 = n4004 & ~n4780 ;
  assign n4782 = n3916 & n4781 ;
  assign n4783 = x54 & ~n612 ;
  assign n4784 = n927 & n1228 ;
  assign n4785 = n1703 ^ n723 ^ 1'b0 ;
  assign n4786 = n4785 ^ n1725 ^ 1'b0 ;
  assign n4787 = n1067 ^ n942 ^ 1'b0 ;
  assign n4788 = n1390 | n4787 ;
  assign n4789 = n349 & ~n1882 ;
  assign n4790 = n890 & n4789 ;
  assign n4791 = n1413 ^ n369 ^ 1'b0 ;
  assign n4792 = n3772 ^ n829 ^ n814 ;
  assign n4793 = n1219 | n1476 ;
  assign n4795 = n1401 | n4579 ;
  assign n4796 = n4795 ^ n3577 ^ 1'b0 ;
  assign n4794 = n3982 ^ x116 ^ 1'b0 ;
  assign n4797 = n4796 ^ n4794 ^ 1'b0 ;
  assign n4798 = n1538 ^ n1198 ^ 1'b0 ;
  assign n4799 = n4798 ^ n569 ^ 1'b0 ;
  assign n4800 = n559 & n4799 ;
  assign n4801 = n4800 ^ n3279 ^ 1'b0 ;
  assign n4802 = n679 & n4801 ;
  assign n4803 = n150 | n1348 ;
  assign n4804 = x46 | n4803 ;
  assign n4805 = n1369 ^ n1325 ^ 1'b0 ;
  assign n4806 = ~n150 & n4805 ;
  assign n4807 = ~n1023 & n4806 ;
  assign n4808 = ~n4804 & n4807 ;
  assign n4809 = n3527 ^ n2993 ^ n662 ;
  assign n4810 = n4381 & ~n4488 ;
  assign n4811 = n3444 | n4810 ;
  assign n4812 = n662 | n1295 ;
  assign n4813 = n4812 ^ n1679 ^ 1'b0 ;
  assign n4814 = n3550 & ~n4813 ;
  assign n4815 = n4814 ^ n763 ^ 1'b0 ;
  assign n4816 = ~n1327 & n2214 ;
  assign n4817 = n4816 ^ n3575 ^ 1'b0 ;
  assign n4818 = x35 & ~n2153 ;
  assign n4819 = ~n4817 & n4818 ;
  assign n4820 = ~n137 & n4819 ;
  assign n4821 = n1925 ^ n1056 ^ 1'b0 ;
  assign n4822 = n2162 | n3635 ;
  assign n4823 = ~n2353 & n2865 ;
  assign n4824 = n1713 | n3289 ;
  assign n4825 = n2830 & n4824 ;
  assign n4826 = n4825 ^ n3227 ^ 1'b0 ;
  assign n4827 = n2839 ^ n1382 ^ 1'b0 ;
  assign n4828 = n4827 ^ n3200 ^ 1'b0 ;
  assign n4829 = ( x94 & n542 ) | ( x94 & ~n4828 ) | ( n542 & ~n4828 ) ;
  assign n4830 = n2648 ^ n2322 ^ 1'b0 ;
  assign n4831 = ~n357 & n4830 ;
  assign n4832 = n4831 ^ n4216 ^ n3006 ;
  assign n4833 = n1245 ^ x21 ^ 1'b0 ;
  assign n4834 = n4833 ^ n3532 ^ 1'b0 ;
  assign n4835 = n224 | n4139 ;
  assign n4836 = n4835 ^ n3346 ^ 1'b0 ;
  assign n4837 = ~n166 & n4836 ;
  assign n4838 = ~n488 & n1152 ;
  assign n4839 = n2235 ^ n420 ^ 1'b0 ;
  assign n4840 = ~n4838 & n4839 ;
  assign n4841 = ( ~n791 & n1922 ) | ( ~n791 & n4191 ) | ( n1922 & n4191 ) ;
  assign n4842 = n4841 ^ n3339 ^ 1'b0 ;
  assign n4843 = ~n2632 & n4842 ;
  assign n4847 = n2445 & n4652 ;
  assign n4848 = n4847 ^ n3921 ^ 1'b0 ;
  assign n4844 = n2807 ^ n423 ^ 1'b0 ;
  assign n4845 = n4632 ^ n722 ^ 1'b0 ;
  assign n4846 = n4844 & ~n4845 ;
  assign n4849 = n4848 ^ n4846 ^ 1'b0 ;
  assign n4850 = n953 ^ n620 ^ 1'b0 ;
  assign n4851 = ~n2559 & n4850 ;
  assign n4852 = ~n143 & n4851 ;
  assign n4853 = n2593 & n4852 ;
  assign n4854 = n3631 ^ n2718 ^ 1'b0 ;
  assign n4855 = ~n194 & n778 ;
  assign n4856 = n4855 ^ n455 ^ 1'b0 ;
  assign n4857 = ( ~n838 & n4854 ) | ( ~n838 & n4856 ) | ( n4854 & n4856 ) ;
  assign n4858 = n4824 ^ n2991 ^ 1'b0 ;
  assign n4859 = n4857 & ~n4858 ;
  assign n4860 = ( n2892 & ~n3297 ) | ( n2892 & n3978 ) | ( ~n3297 & n3978 ) ;
  assign n4861 = n4860 ^ n826 ^ 1'b0 ;
  assign n4862 = n2423 & ~n4370 ;
  assign n4863 = n4862 ^ n1978 ^ 1'b0 ;
  assign n4864 = n878 & n4863 ;
  assign n4865 = n971 & n4864 ;
  assign n4866 = n4865 ^ x21 ^ 1'b0 ;
  assign n4867 = n4866 ^ n1276 ^ 1'b0 ;
  assign n4868 = n2388 ^ n1740 ^ 1'b0 ;
  assign n4869 = n4868 ^ n1879 ^ 1'b0 ;
  assign n4870 = n4867 | n4869 ;
  assign n4871 = n4870 ^ n597 ^ 1'b0 ;
  assign n4872 = n3784 | n4871 ;
  assign n4873 = x98 | n391 ;
  assign n4874 = n4873 ^ n1661 ^ 1'b0 ;
  assign n4875 = n909 & ~n1799 ;
  assign n4876 = n2771 | n4875 ;
  assign n4877 = ( n208 & ~n4874 ) | ( n208 & n4876 ) | ( ~n4874 & n4876 ) ;
  assign n4878 = n2829 & ~n4877 ;
  assign n4879 = n4878 ^ n1192 ^ 1'b0 ;
  assign n4880 = n791 | n4540 ;
  assign n4881 = ( n1385 & n2458 ) | ( n1385 & n3007 ) | ( n2458 & n3007 ) ;
  assign n4882 = ~n1925 & n4881 ;
  assign n4883 = ~n2418 & n4882 ;
  assign n4884 = n1045 | n2967 ;
  assign n4885 = n2275 ^ n1437 ^ 1'b0 ;
  assign n4886 = n969 & ~n4885 ;
  assign n4887 = n4522 ^ n4521 ^ n2084 ;
  assign n4888 = n2829 ^ n2714 ^ 1'b0 ;
  assign n4889 = n1396 & n4888 ;
  assign n4890 = n2172 & n4889 ;
  assign n4891 = n2340 & ~n4890 ;
  assign n4892 = n4891 ^ n1560 ^ 1'b0 ;
  assign n4893 = n2794 ^ n2564 ^ 1'b0 ;
  assign n4894 = x98 ^ x90 ^ 1'b0 ;
  assign n4895 = n376 & n4894 ;
  assign n4896 = n3785 & n4895 ;
  assign n4897 = ~n1869 & n4896 ;
  assign n4898 = x79 & ~n4897 ;
  assign n4899 = n3414 ^ n2619 ^ 1'b0 ;
  assign n4900 = ~n2285 & n4453 ;
  assign n4901 = n4899 & n4900 ;
  assign n4902 = n1776 & n3385 ;
  assign n4903 = n344 | n1575 ;
  assign n4904 = x84 & ~n4903 ;
  assign n4905 = n4904 ^ n261 ^ 1'b0 ;
  assign n4906 = n3730 ^ n3219 ^ 1'b0 ;
  assign n4908 = n1111 | n1386 ;
  assign n4907 = n1346 | n2575 ;
  assign n4909 = n4908 ^ n4907 ^ 1'b0 ;
  assign n4910 = n4909 ^ n2373 ^ 1'b0 ;
  assign n4911 = n4496 ^ n999 ^ 1'b0 ;
  assign n4912 = n4578 & n4911 ;
  assign n4913 = n3955 ^ n1332 ^ 1'b0 ;
  assign n4914 = n1572 | n1804 ;
  assign n4915 = n2328 & ~n4914 ;
  assign n4916 = n260 | n4915 ;
  assign n4917 = n4913 | n4916 ;
  assign n4918 = x62 & ~n4355 ;
  assign n4920 = n4025 ^ n1983 ^ 1'b0 ;
  assign n4921 = n620 & n4920 ;
  assign n4922 = n1685 | n4921 ;
  assign n4923 = ~n875 & n4922 ;
  assign n4919 = n3879 ^ n2490 ^ n1794 ;
  assign n4924 = n4923 ^ n4919 ^ 1'b0 ;
  assign n4925 = n904 | n3378 ;
  assign n4926 = n1711 ^ n829 ^ 1'b0 ;
  assign n4927 = ~n307 & n4926 ;
  assign n4928 = n4025 ^ n3021 ^ 1'b0 ;
  assign n4929 = n4927 & n4928 ;
  assign n4930 = n3517 ^ n3445 ^ n493 ;
  assign n4931 = n1329 | n4930 ;
  assign n4932 = n4355 & ~n4931 ;
  assign n4933 = ~x59 & n4932 ;
  assign n4934 = n1164 | n1257 ;
  assign n4935 = n175 & n4934 ;
  assign n4936 = n775 ^ n613 ^ 1'b0 ;
  assign n4937 = n1919 & n4936 ;
  assign n4938 = n2193 & n4937 ;
  assign n4939 = n4371 ^ n374 ^ 1'b0 ;
  assign n4940 = n3486 & ~n4939 ;
  assign n4941 = n4736 ^ n3571 ^ 1'b0 ;
  assign n4942 = n2876 & n4517 ;
  assign n4943 = ~n1081 & n2261 ;
  assign n4944 = n4943 ^ n2890 ^ 1'b0 ;
  assign n4945 = ( ~n2362 & n2529 ) | ( ~n2362 & n2718 ) | ( n2529 & n2718 ) ;
  assign n4946 = n3087 ^ n1027 ^ 1'b0 ;
  assign n4947 = n1118 & ~n4946 ;
  assign n4948 = n527 & n648 ;
  assign n4949 = ~n4947 & n4948 ;
  assign n4950 = ~x27 & n876 ;
  assign n4951 = n4950 ^ n1902 ^ n317 ;
  assign n4952 = n4951 ^ n3890 ^ 1'b0 ;
  assign n4953 = x77 & ~n4952 ;
  assign n4954 = n4953 ^ n4168 ^ 1'b0 ;
  assign n4955 = n4949 | n4954 ;
  assign n4956 = n4151 & ~n4779 ;
  assign n4959 = n225 & ~n831 ;
  assign n4960 = n2458 & n4959 ;
  assign n4961 = n2652 ^ n2303 ^ 1'b0 ;
  assign n4962 = n3072 & ~n4961 ;
  assign n4963 = n4960 & n4962 ;
  assign n4957 = ( n744 & n802 ) | ( n744 & ~n1121 ) | ( n802 & ~n1121 ) ;
  assign n4958 = n4957 ^ n3940 ^ 1'b0 ;
  assign n4964 = n4963 ^ n4958 ^ 1'b0 ;
  assign n4965 = n4956 & n4964 ;
  assign n4966 = n709 & ~n878 ;
  assign n4967 = ~n1405 & n1844 ;
  assign n4968 = ~n1380 & n2906 ;
  assign n4969 = n4967 & n4968 ;
  assign n4970 = n2870 | n4041 ;
  assign n4971 = n144 & n392 ;
  assign n4972 = n477 & n4971 ;
  assign n4973 = n4972 ^ n3738 ^ 1'b0 ;
  assign n4974 = ~n1229 & n1242 ;
  assign n4975 = n4974 ^ x46 ^ 1'b0 ;
  assign n4976 = n419 & n1344 ;
  assign n4977 = n4976 ^ n208 ^ 1'b0 ;
  assign n4978 = n4975 | n4977 ;
  assign n4979 = x57 & n4266 ;
  assign n4980 = n3601 ^ n775 ^ 1'b0 ;
  assign n4981 = ~n1941 & n4980 ;
  assign n4982 = n4981 ^ n575 ^ 1'b0 ;
  assign n4983 = n2261 & n4982 ;
  assign n4984 = n1761 ^ n1334 ^ 1'b0 ;
  assign n4985 = n4983 & ~n4984 ;
  assign n4986 = n3665 & n4738 ;
  assign n4987 = n3166 & n4986 ;
  assign n4988 = n4657 | n4987 ;
  assign n4989 = n4988 ^ n574 ^ 1'b0 ;
  assign n4990 = n1793 & ~n4071 ;
  assign n4991 = n4897 ^ n225 ^ 1'b0 ;
  assign n4992 = n1878 & ~n4991 ;
  assign n4993 = ~x38 & n1831 ;
  assign n4994 = n4993 ^ n3087 ^ 1'b0 ;
  assign n4995 = ~n618 & n4994 ;
  assign n4996 = n4601 ^ n4069 ^ 1'b0 ;
  assign n4997 = ~n2993 & n4996 ;
  assign n4998 = n2364 ^ n326 ^ 1'b0 ;
  assign n4999 = n4998 ^ n4647 ^ n637 ;
  assign n5000 = n986 ^ n744 ^ n285 ;
  assign n5001 = n3087 & n5000 ;
  assign n5002 = ~n2535 & n5001 ;
  assign n5003 = n2662 | n4123 ;
  assign n5004 = n5003 ^ n3988 ^ 1'b0 ;
  assign n5005 = ( n821 & ~n1969 ) | ( n821 & n2172 ) | ( ~n1969 & n2172 ) ;
  assign n5006 = n3608 ^ n1698 ^ 1'b0 ;
  assign n5007 = x17 & n5006 ;
  assign n5008 = n2003 & n2127 ;
  assign n5009 = ~n2020 & n5008 ;
  assign n5010 = n3951 ^ n3251 ^ 1'b0 ;
  assign n5011 = n3884 | n5010 ;
  assign n5012 = n2378 & n4764 ;
  assign n5013 = n766 ^ n484 ^ 1'b0 ;
  assign n5014 = n1078 & n5013 ;
  assign n5015 = n5014 ^ n1067 ^ n430 ;
  assign n5016 = ( x14 & ~n4219 ) | ( x14 & n5015 ) | ( ~n4219 & n5015 ) ;
  assign n5017 = ( ~x77 & n1134 ) | ( ~x77 & n1429 ) | ( n1134 & n1429 ) ;
  assign n5018 = n702 ^ x121 ^ x97 ;
  assign n5019 = n4357 | n5018 ;
  assign n5020 = n5017 & ~n5019 ;
  assign n5021 = n3171 ^ n3089 ^ 1'b0 ;
  assign n5022 = n371 | n5021 ;
  assign n5023 = n5022 ^ n1863 ^ 1'b0 ;
  assign n5025 = n154 | n811 ;
  assign n5026 = x38 | n5025 ;
  assign n5027 = n2287 & ~n2756 ;
  assign n5028 = ~n5026 & n5027 ;
  assign n5024 = n2658 & ~n3107 ;
  assign n5029 = n5028 ^ n5024 ^ 1'b0 ;
  assign n5030 = n5029 ^ n4778 ^ 1'b0 ;
  assign n5031 = ~n4314 & n5030 ;
  assign n5032 = n2558 | n3855 ;
  assign n5033 = n5032 ^ n2405 ^ 1'b0 ;
  assign n5034 = n951 & ~n2123 ;
  assign n5035 = ~n5033 & n5034 ;
  assign n5036 = n3107 ^ n2026 ^ 1'b0 ;
  assign n5037 = n4207 & n5036 ;
  assign n5038 = n5035 & ~n5037 ;
  assign n5039 = n4132 ^ n3676 ^ 1'b0 ;
  assign n5040 = ~n2333 & n5039 ;
  assign n5043 = n190 | n283 ;
  assign n5044 = n5043 ^ n3323 ^ n2456 ;
  assign n5041 = n695 & n3539 ;
  assign n5042 = n5041 ^ n1750 ^ 1'b0 ;
  assign n5045 = n5044 ^ n5042 ^ 1'b0 ;
  assign n5046 = ~n1143 & n5045 ;
  assign n5047 = ~n377 & n515 ;
  assign n5048 = ~n4957 & n5047 ;
  assign n5049 = ( n487 & ~n3479 ) | ( n487 & n5048 ) | ( ~n3479 & n5048 ) ;
  assign n5050 = x110 & ~n4769 ;
  assign n5051 = ~n4867 & n5050 ;
  assign n5052 = n5051 ^ n1943 ^ 1'b0 ;
  assign n5053 = ~n999 & n1936 ;
  assign n5054 = n1190 ^ n487 ^ 1'b0 ;
  assign n5055 = x29 & n3892 ;
  assign n5056 = n1457 & ~n2073 ;
  assign n5057 = n5056 ^ n539 ^ 1'b0 ;
  assign n5058 = n4082 & n5057 ;
  assign n5059 = ~n5055 & n5058 ;
  assign n5060 = n1977 ^ n1545 ^ 1'b0 ;
  assign n5061 = n460 & ~n5060 ;
  assign n5062 = n3762 | n5061 ;
  assign n5063 = n4400 ^ n2943 ^ 1'b0 ;
  assign n5064 = n1981 | n3065 ;
  assign n5065 = n897 ^ n484 ^ 1'b0 ;
  assign n5066 = n2125 & n5065 ;
  assign n5067 = ~n5064 & n5066 ;
  assign n5068 = n701 ^ n699 ^ 1'b0 ;
  assign n5069 = ~n3411 & n5068 ;
  assign n5070 = n5069 ^ n1957 ^ 1'b0 ;
  assign n5071 = ~n1662 & n5070 ;
  assign n5072 = n1562 & n2449 ;
  assign n5073 = ~n3062 & n5072 ;
  assign n5074 = n5073 ^ n4287 ^ 1'b0 ;
  assign n5075 = n556 & ~n826 ;
  assign n5076 = n277 & ~n361 ;
  assign n5077 = ~n2674 & n5076 ;
  assign n5078 = n5077 ^ n358 ^ 1'b0 ;
  assign n5079 = n5075 & n5078 ;
  assign n5080 = ~n3234 & n3856 ;
  assign n5081 = x20 & ~n4957 ;
  assign n5082 = n5081 ^ n4224 ^ 1'b0 ;
  assign n5083 = n3295 & ~n3510 ;
  assign n5084 = n4409 ^ n560 ^ 1'b0 ;
  assign n5085 = n3212 ^ n1394 ^ 1'b0 ;
  assign n5086 = n2261 & ~n2612 ;
  assign n5087 = n2270 & n3246 ;
  assign n5088 = ~x126 & n5087 ;
  assign n5089 = n445 & ~n5088 ;
  assign n5090 = ~n5086 & n5089 ;
  assign n5091 = n5085 & ~n5090 ;
  assign n5092 = ~n989 & n1847 ;
  assign n5093 = n741 & n3644 ;
  assign n5094 = n2497 & ~n2779 ;
  assign n5095 = ~n1201 & n1735 ;
  assign n5096 = n509 & n5095 ;
  assign n5097 = n5094 | n5096 ;
  assign n5098 = n5093 | n5097 ;
  assign n5099 = ~n147 & n241 ;
  assign n5100 = n5099 ^ n1819 ^ 1'b0 ;
  assign n5101 = ~n444 & n4004 ;
  assign n5102 = n5101 ^ n438 ^ 1'b0 ;
  assign n5103 = n657 | n992 ;
  assign n5104 = n1439 | n5103 ;
  assign n5105 = n1505 ^ n540 ^ 1'b0 ;
  assign n5106 = x52 & ~n5105 ;
  assign n5107 = ( n1575 & ~n5104 ) | ( n1575 & n5106 ) | ( ~n5104 & n5106 ) ;
  assign n5108 = n355 ^ n302 ^ 1'b0 ;
  assign n5109 = ( n2774 & ~n3030 ) | ( n2774 & n5108 ) | ( ~n3030 & n5108 ) ;
  assign n5110 = n1167 & ~n5109 ;
  assign n5111 = ~n1062 & n5110 ;
  assign n5113 = n3041 | n3473 ;
  assign n5114 = n3473 & ~n5113 ;
  assign n5112 = n407 ^ n210 ^ 1'b0 ;
  assign n5115 = n5114 ^ n5112 ^ 1'b0 ;
  assign n5116 = n808 & ~n4095 ;
  assign n5117 = ~n2233 & n5116 ;
  assign n5119 = n657 & n3685 ;
  assign n5118 = n755 | n3502 ;
  assign n5120 = n5119 ^ n5118 ^ 1'b0 ;
  assign n5121 = ~n886 & n5120 ;
  assign n5122 = n5121 ^ n692 ^ 1'b0 ;
  assign n5126 = ~n960 & n1567 ;
  assign n5127 = n5126 ^ n1614 ^ 1'b0 ;
  assign n5128 = n2530 & ~n5127 ;
  assign n5129 = n5128 ^ n2720 ^ 1'b0 ;
  assign n5130 = n2014 | n5129 ;
  assign n5131 = n5130 ^ n395 ^ 1'b0 ;
  assign n5123 = n469 & n708 ;
  assign n5124 = ~n1147 & n5123 ;
  assign n5125 = n4138 & n5124 ;
  assign n5132 = n5131 ^ n5125 ^ 1'b0 ;
  assign n5133 = n4122 ^ n847 ^ 1'b0 ;
  assign n5134 = n2376 | n2486 ;
  assign n5135 = ( n2673 & ~n4145 ) | ( n2673 & n4318 ) | ( ~n4145 & n4318 ) ;
  assign n5136 = n642 | n765 ;
  assign n5137 = ( n1792 & n2949 ) | ( n1792 & ~n5136 ) | ( n2949 & ~n5136 ) ;
  assign n5138 = n1890 & n3499 ;
  assign n5139 = ~n3357 & n3696 ;
  assign n5140 = ~n3696 & n5139 ;
  assign n5141 = n2933 & ~n4893 ;
  assign n5142 = ~n1867 & n5141 ;
  assign n5143 = n4299 ^ n208 ^ 1'b0 ;
  assign n5144 = x24 & ~n1152 ;
  assign n5145 = n2140 & ~n5144 ;
  assign n5146 = n4189 ^ n1348 ^ 1'b0 ;
  assign n5147 = n821 ^ x79 ^ 1'b0 ;
  assign n5148 = n2012 | n5147 ;
  assign n5151 = n4148 ^ n673 ^ 1'b0 ;
  assign n5149 = ~n165 & n3577 ;
  assign n5150 = n5149 ^ n1853 ^ 1'b0 ;
  assign n5152 = n5151 ^ n5150 ^ n1060 ;
  assign n5153 = n993 & n2363 ;
  assign n5154 = n5153 ^ n3610 ^ 1'b0 ;
  assign n5155 = n2746 & ~n5154 ;
  assign n5156 = n5155 ^ n1512 ^ 1'b0 ;
  assign n5158 = ~n813 & n4981 ;
  assign n5159 = n5158 ^ n2903 ^ 1'b0 ;
  assign n5157 = n4628 ^ n4560 ^ 1'b0 ;
  assign n5160 = n5159 ^ n5157 ^ 1'b0 ;
  assign n5161 = ~n916 & n5160 ;
  assign n5162 = n2603 & n5161 ;
  assign n5163 = n5162 ^ n208 ^ 1'b0 ;
  assign n5164 = n1201 ^ n241 ^ 1'b0 ;
  assign n5165 = n5164 ^ n1446 ^ 1'b0 ;
  assign n5166 = n2224 ^ n1517 ^ 1'b0 ;
  assign n5167 = n2315 | n3757 ;
  assign n5168 = n3298 ^ n1819 ^ 1'b0 ;
  assign n5169 = n3013 ^ n195 ^ 1'b0 ;
  assign n5170 = ~n5168 & n5169 ;
  assign n5171 = n2878 & ~n3846 ;
  assign n5172 = n2778 & n4201 ;
  assign n5173 = x113 & ~n1134 ;
  assign n5174 = n5173 ^ n3704 ^ 1'b0 ;
  assign n5175 = ~n1398 & n5144 ;
  assign n5176 = n3139 & n5175 ;
  assign n5177 = n5174 & ~n5176 ;
  assign n5178 = n2987 ^ n1608 ^ 1'b0 ;
  assign n5179 = n5178 ^ n1068 ^ 1'b0 ;
  assign n5180 = x58 & n2444 ;
  assign n5181 = n5180 ^ n3064 ^ 1'b0 ;
  assign n5182 = n1882 | n4007 ;
  assign n5183 = n5182 ^ n615 ^ 1'b0 ;
  assign n5184 = n3162 | n5183 ;
  assign n5185 = n5181 | n5184 ;
  assign n5186 = ~n2450 & n4364 ;
  assign n5187 = ~n5185 & n5186 ;
  assign n5188 = n3327 | n3346 ;
  assign n5199 = ~n417 & n3433 ;
  assign n5200 = n5199 ^ n1625 ^ 1'b0 ;
  assign n5189 = n737 ^ x111 ^ 1'b0 ;
  assign n5190 = n1095 & n5189 ;
  assign n5191 = n5190 ^ n2215 ^ 1'b0 ;
  assign n5192 = ~n855 & n1175 ;
  assign n5193 = n5192 ^ n1693 ^ 1'b0 ;
  assign n5194 = n1031 & n5193 ;
  assign n5195 = n5194 ^ n2039 ^ 1'b0 ;
  assign n5196 = n5195 ^ n888 ^ 1'b0 ;
  assign n5197 = n5191 & n5196 ;
  assign n5198 = n2955 & n5197 ;
  assign n5201 = n5200 ^ n5198 ^ 1'b0 ;
  assign n5202 = n5188 & ~n5201 ;
  assign n5203 = n2938 ^ n1999 ^ 1'b0 ;
  assign n5204 = n224 | n2300 ;
  assign n5205 = n1337 | n5204 ;
  assign n5206 = n5205 ^ n1334 ^ n730 ;
  assign n5207 = n5206 ^ n2402 ^ 1'b0 ;
  assign n5213 = ~n1455 & n4149 ;
  assign n5214 = n5213 ^ n1899 ^ 1'b0 ;
  assign n5208 = n685 | n3828 ;
  assign n5209 = n1972 & ~n2581 ;
  assign n5210 = n3872 | n5209 ;
  assign n5211 = n5210 ^ x69 ^ 1'b0 ;
  assign n5212 = ~n5208 & n5211 ;
  assign n5215 = n5214 ^ n5212 ^ 1'b0 ;
  assign n5217 = x46 & ~n1386 ;
  assign n5218 = ~n3491 & n5217 ;
  assign n5216 = ~n1079 & n2466 ;
  assign n5219 = n5218 ^ n5216 ^ 1'b0 ;
  assign n5220 = ( ~x24 & n2421 ) | ( ~x24 & n2585 ) | ( n2421 & n2585 ) ;
  assign n5221 = n3179 & n5220 ;
  assign n5222 = ~n4461 & n5221 ;
  assign n5223 = n496 & ~n4166 ;
  assign n5224 = n5223 ^ n630 ^ 1'b0 ;
  assign n5225 = n249 & ~n1083 ;
  assign n5226 = ~x103 & n5225 ;
  assign n5227 = n3567 & n5226 ;
  assign n5228 = n1567 | n5227 ;
  assign n5229 = n1716 & ~n4876 ;
  assign n5230 = n5228 & n5229 ;
  assign n5231 = n3561 & n5144 ;
  assign n5232 = n4661 ^ n3699 ^ 1'b0 ;
  assign n5233 = n5048 ^ n3376 ^ 1'b0 ;
  assign n5234 = n2214 & n5233 ;
  assign n5235 = ( n2268 & ~n2861 ) | ( n2268 & n5234 ) | ( ~n2861 & n5234 ) ;
  assign n5237 = n737 | n4903 ;
  assign n5238 = n876 | n5237 ;
  assign n5239 = ~n355 & n5238 ;
  assign n5240 = n5239 ^ x44 ^ 1'b0 ;
  assign n5236 = n3577 ^ n1588 ^ 1'b0 ;
  assign n5241 = n5240 ^ n5236 ^ 1'b0 ;
  assign n5242 = n1243 ^ n388 ^ 1'b0 ;
  assign n5244 = n808 & ~n1664 ;
  assign n5243 = ~n867 & n2034 ;
  assign n5245 = n5244 ^ n5243 ^ 1'b0 ;
  assign n5246 = n468 | n5245 ;
  assign n5258 = n1947 ^ n412 ^ 1'b0 ;
  assign n5259 = n3631 ^ n1828 ^ 1'b0 ;
  assign n5260 = n5258 | n5259 ;
  assign n5247 = ~n2972 & n4718 ;
  assign n5248 = n5247 ^ n5093 ^ n1623 ;
  assign n5249 = n4389 ^ n2882 ^ 1'b0 ;
  assign n5250 = n5249 ^ n2882 ^ n1229 ;
  assign n5251 = ~n2374 & n5250 ;
  assign n5252 = n824 & n2473 ;
  assign n5253 = n5252 ^ n1107 ^ 1'b0 ;
  assign n5254 = n2543 & ~n5253 ;
  assign n5255 = n5251 & ~n5254 ;
  assign n5256 = n5255 ^ n3278 ^ 1'b0 ;
  assign n5257 = ~n5248 & n5256 ;
  assign n5261 = n5260 ^ n5257 ^ 1'b0 ;
  assign n5262 = n156 & ~n1505 ;
  assign n5265 = n1221 ^ n960 ^ 1'b0 ;
  assign n5263 = ~n1083 & n1167 ;
  assign n5264 = n5263 ^ n1026 ^ 1'b0 ;
  assign n5266 = n5265 ^ n5264 ^ 1'b0 ;
  assign n5267 = n5262 | n5266 ;
  assign n5268 = ( ~n351 & n863 ) | ( ~n351 & n866 ) | ( n863 & n866 ) ;
  assign n5269 = n5268 ^ n2070 ^ 1'b0 ;
  assign n5270 = n1473 & ~n5269 ;
  assign n5271 = n4671 & n5270 ;
  assign n5272 = n4203 | n5271 ;
  assign n5273 = n5267 & ~n5272 ;
  assign n5274 = ~n3413 & n3696 ;
  assign n5275 = x114 & n1325 ;
  assign n5276 = n5275 ^ n4868 ^ 1'b0 ;
  assign n5277 = n3343 ^ x39 ^ 1'b0 ;
  assign n5278 = n853 & n4766 ;
  assign n5279 = n5278 ^ x55 ^ 1'b0 ;
  assign n5280 = n241 & n2948 ;
  assign n5281 = n5280 ^ n1679 ^ 1'b0 ;
  assign n5282 = n3186 ^ n1943 ^ 1'b0 ;
  assign n5283 = n5281 & n5282 ;
  assign n5284 = n1300 ^ n904 ^ n475 ;
  assign n5285 = n849 | n1300 ;
  assign n5286 = n5285 ^ n892 ^ 1'b0 ;
  assign n5287 = n1404 & n5286 ;
  assign n5288 = n5267 | n5287 ;
  assign n5289 = n1629 | n5288 ;
  assign n5290 = x53 & ~n540 ;
  assign n5291 = n1945 | n5290 ;
  assign n5292 = n2016 ^ n1507 ^ 1'b0 ;
  assign n5293 = n5291 & ~n5292 ;
  assign n5294 = ~n3118 & n5293 ;
  assign n5297 = n1899 ^ x34 ^ 1'b0 ;
  assign n5295 = n3071 ^ n1975 ^ 1'b0 ;
  assign n5296 = n3474 & ~n5295 ;
  assign n5298 = n5297 ^ n5296 ^ n2448 ;
  assign n5299 = x114 & ~n1390 ;
  assign n5300 = n5299 ^ n3233 ^ 1'b0 ;
  assign n5301 = n5300 ^ n4299 ^ n198 ;
  assign n5302 = n5301 ^ n3662 ^ 1'b0 ;
  assign n5303 = n1801 & ~n4281 ;
  assign n5304 = n5303 ^ x29 ^ 1'b0 ;
  assign n5305 = n5119 ^ n2055 ^ 1'b0 ;
  assign n5306 = n3229 ^ n1015 ^ 1'b0 ;
  assign n5307 = n5306 ^ n2675 ^ 1'b0 ;
  assign n5308 = ~n287 & n5307 ;
  assign n5309 = n5308 ^ n2851 ^ 1'b0 ;
  assign n5310 = n5309 ^ n1386 ^ 1'b0 ;
  assign n5311 = n4978 ^ n4705 ^ 1'b0 ;
  assign n5312 = n1324 & ~n3572 ;
  assign n5313 = n5312 ^ n4963 ^ 1'b0 ;
  assign n5314 = n4122 | n5313 ;
  assign n5315 = n1205 | n5314 ;
  assign n5316 = n229 ^ n225 ^ 1'b0 ;
  assign n5317 = ( ~n1204 & n3622 ) | ( ~n1204 & n5316 ) | ( n3622 & n5316 ) ;
  assign n5318 = ~n2726 & n5193 ;
  assign n5321 = n5086 ^ n3648 ^ 1'b0 ;
  assign n5319 = n755 & n3037 ;
  assign n5320 = ~n4849 & n5319 ;
  assign n5322 = n5321 ^ n5320 ^ 1'b0 ;
  assign n5323 = n2302 & n5322 ;
  assign n5324 = n4043 ^ n1827 ^ 1'b0 ;
  assign n5325 = n5324 ^ n2380 ^ 1'b0 ;
  assign n5326 = n4829 | n5325 ;
  assign n5327 = ~n2330 & n4348 ;
  assign n5328 = n4513 ^ n902 ^ 1'b0 ;
  assign n5329 = n533 & n5328 ;
  assign n5330 = n3404 | n5329 ;
  assign n5331 = ~n2014 & n5330 ;
  assign n5338 = n675 & n1716 ;
  assign n5339 = n1467 & n5338 ;
  assign n5332 = n4152 ^ n2554 ^ 1'b0 ;
  assign n5333 = n3515 & n5332 ;
  assign n5334 = n3872 & n5333 ;
  assign n5335 = ~n2187 & n4082 ;
  assign n5336 = ~n331 & n5335 ;
  assign n5337 = n5334 | n5336 ;
  assign n5340 = n5339 ^ n5337 ^ 1'b0 ;
  assign n5341 = n2656 ^ n1672 ^ 1'b0 ;
  assign n5342 = n1850 & n5341 ;
  assign n5343 = x69 & ~n351 ;
  assign n5344 = ~n5342 & n5343 ;
  assign n5345 = n2481 ^ n569 ^ 1'b0 ;
  assign n5346 = n1330 & n5345 ;
  assign n5347 = n5346 ^ n3099 ^ 1'b0 ;
  assign n5348 = n2658 & ~n5312 ;
  assign n5349 = n808 & ~n1723 ;
  assign n5350 = n2409 & ~n3376 ;
  assign n5351 = n5350 ^ n1868 ^ n874 ;
  assign n5352 = ( n379 & ~n2376 ) | ( n379 & n3170 ) | ( ~n2376 & n3170 ) ;
  assign n5353 = n5108 ^ n1790 ^ 1'b0 ;
  assign n5354 = n5352 & ~n5353 ;
  assign n5355 = n1755 & ~n4022 ;
  assign n5356 = ( n915 & n2245 ) | ( n915 & n2853 ) | ( n2245 & n2853 ) ;
  assign n5357 = n5356 ^ n3017 ^ 1'b0 ;
  assign n5358 = n1077 ^ n357 ^ 1'b0 ;
  assign n5359 = n5358 ^ n2835 ^ 1'b0 ;
  assign n5360 = ~n5357 & n5359 ;
  assign n5361 = n3030 ^ n1363 ^ 1'b0 ;
  assign n5362 = x89 & ~n5361 ;
  assign n5363 = n1319 & ~n5362 ;
  assign n5364 = n3850 & n5363 ;
  assign n5365 = n1448 | n2187 ;
  assign n5366 = n5365 ^ n884 ^ 1'b0 ;
  assign n5367 = n3006 & ~n5366 ;
  assign n5368 = ( n745 & n4506 ) | ( n745 & n5367 ) | ( n4506 & n5367 ) ;
  assign n5369 = n2531 ^ n1623 ^ 1'b0 ;
  assign n5370 = n934 & n5369 ;
  assign n5371 = n3582 & ~n4055 ;
  assign n5372 = x69 & ~n2685 ;
  assign n5373 = n5372 ^ n2340 ^ 1'b0 ;
  assign n5374 = n5371 | n5373 ;
  assign n5375 = ( n3290 & n4820 ) | ( n3290 & n5374 ) | ( n4820 & n5374 ) ;
  assign n5376 = n1856 | n4183 ;
  assign n5377 = n595 ^ x78 ^ 1'b0 ;
  assign n5378 = n2948 | n5377 ;
  assign n5379 = n391 & n5378 ;
  assign n5380 = n1757 ^ n215 ^ 1'b0 ;
  assign n5381 = n5379 | n5380 ;
  assign n5382 = n2951 ^ n1526 ^ 1'b0 ;
  assign n5383 = ~n2792 & n5382 ;
  assign n5384 = n2504 ^ n709 ^ 1'b0 ;
  assign n5385 = n2969 & ~n5384 ;
  assign n5386 = n5385 ^ n2361 ^ 1'b0 ;
  assign n5387 = n5383 & n5386 ;
  assign n5388 = n1821 & ~n5231 ;
  assign n5389 = ~n1394 & n5388 ;
  assign n5390 = n1057 | n3955 ;
  assign n5391 = n5390 ^ n801 ^ 1'b0 ;
  assign n5392 = n1787 ^ n1639 ^ 1'b0 ;
  assign n5393 = n5392 ^ n861 ^ 1'b0 ;
  assign n5394 = ~n5391 & n5393 ;
  assign n5396 = ~n453 & n1263 ;
  assign n5397 = n3655 & n5396 ;
  assign n5398 = n1212 & ~n5397 ;
  assign n5395 = n501 & n1209 ;
  assign n5399 = n5398 ^ n5395 ^ 1'b0 ;
  assign n5400 = n4585 & ~n5399 ;
  assign n5401 = n3037 ^ n1552 ^ 1'b0 ;
  assign n5402 = n427 & n5401 ;
  assign n5403 = n2809 & ~n3814 ;
  assign n5404 = ~n1735 & n5403 ;
  assign n5405 = n1354 & n2287 ;
  assign n5406 = n5405 ^ n2182 ^ 1'b0 ;
  assign n5407 = n2542 ^ n2066 ^ 1'b0 ;
  assign n5408 = ~n5406 & n5407 ;
  assign n5409 = n4784 ^ n4215 ^ 1'b0 ;
  assign n5410 = n3979 & ~n5409 ;
  assign n5411 = x32 & ~n3284 ;
  assign n5412 = n5411 ^ n1412 ^ 1'b0 ;
  assign n5413 = n2615 | n5412 ;
  assign n5414 = n3565 ^ n1270 ^ n759 ;
  assign n5415 = n1281 ^ n172 ^ 1'b0 ;
  assign n5416 = n5415 ^ n3373 ^ n340 ;
  assign n5417 = n5416 ^ n1136 ^ 1'b0 ;
  assign n5418 = n4661 | n5417 ;
  assign n5419 = n5414 | n5418 ;
  assign n5420 = n518 & ~n1097 ;
  assign n5421 = n2947 ^ n874 ^ 1'b0 ;
  assign n5422 = n5420 & n5421 ;
  assign n5423 = n5422 ^ n4556 ^ 1'b0 ;
  assign n5425 = n3295 ^ n1953 ^ 1'b0 ;
  assign n5426 = x95 & n5425 ;
  assign n5424 = n4723 ^ n3925 ^ 1'b0 ;
  assign n5427 = n5426 ^ n5424 ^ 1'b0 ;
  assign n5428 = n740 & n2776 ;
  assign n5429 = ~x103 & n5428 ;
  assign n5430 = ~n5108 & n5429 ;
  assign n5431 = ( n481 & n1421 ) | ( n481 & n3975 ) | ( n1421 & n3975 ) ;
  assign n5432 = n1089 ^ x104 ^ 1'b0 ;
  assign n5433 = x86 & n3687 ;
  assign n5434 = ~n2127 & n5433 ;
  assign n5435 = n5434 ^ n2859 ^ n2014 ;
  assign n5436 = n2823 & n3792 ;
  assign n5437 = n2054 & n5436 ;
  assign n5438 = x34 & ~n851 ;
  assign n5439 = n5438 ^ x23 ^ 1'b0 ;
  assign n5440 = n448 | n5439 ;
  assign n5441 = n5440 ^ n4794 ^ 1'b0 ;
  assign n5442 = n5441 ^ n4745 ^ 1'b0 ;
  assign n5443 = n231 | n1662 ;
  assign n5444 = n3601 | n4043 ;
  assign n5445 = n5444 ^ n1773 ^ 1'b0 ;
  assign n5446 = n5443 | n5445 ;
  assign n5447 = ( n2319 & ~n2497 ) | ( n2319 & n3744 ) | ( ~n2497 & n3744 ) ;
  assign n5448 = ~n1444 & n5447 ;
  assign n5449 = n4303 | n5448 ;
  assign n5450 = n5449 ^ n2652 ^ 1'b0 ;
  assign n5451 = x43 & n4566 ;
  assign n5452 = n3808 & ~n4293 ;
  assign n5453 = n5452 ^ n857 ^ 1'b0 ;
  assign n5454 = n1509 | n2564 ;
  assign n5455 = n5454 ^ n2014 ^ 1'b0 ;
  assign n5458 = n1306 ^ x61 ^ 1'b0 ;
  assign n5456 = n3460 ^ n2946 ^ 1'b0 ;
  assign n5457 = n3590 | n5456 ;
  assign n5459 = n5458 ^ n5457 ^ 1'b0 ;
  assign n5460 = ~n5455 & n5459 ;
  assign n5461 = n5460 ^ n1209 ^ 1'b0 ;
  assign n5462 = n5029 & ~n5441 ;
  assign n5463 = n3286 | n3727 ;
  assign n5464 = n4350 ^ n157 ^ 1'b0 ;
  assign n5465 = n5463 | n5464 ;
  assign n5466 = n2591 & ~n5465 ;
  assign n5467 = n3997 ^ n2419 ^ 1'b0 ;
  assign n5468 = n3037 & n3772 ;
  assign n5469 = n4151 ^ x24 ^ 1'b0 ;
  assign n5470 = n1898 & ~n5469 ;
  assign n5471 = n2989 & ~n5470 ;
  assign n5472 = n493 & n1804 ;
  assign n5473 = n1432 & ~n5472 ;
  assign n5474 = n1138 | n2213 ;
  assign n5475 = n5474 ^ n5086 ^ 1'b0 ;
  assign n5476 = n2892 ^ n2462 ^ 1'b0 ;
  assign n5477 = n374 & n5476 ;
  assign n5478 = n5477 ^ n986 ^ 1'b0 ;
  assign n5479 = n5475 & n5478 ;
  assign n5480 = n2559 | n4753 ;
  assign n5481 = n1651 & ~n5480 ;
  assign n5482 = n1350 & n2170 ;
  assign n5483 = ~x79 & n5482 ;
  assign n5484 = n1392 & n5483 ;
  assign n5485 = ~n5136 & n5482 ;
  assign n5486 = n2289 & ~n4281 ;
  assign n5487 = ( n1077 & n1835 ) | ( n1077 & n5486 ) | ( n1835 & n5486 ) ;
  assign n5492 = n754 | n1450 ;
  assign n5493 = n4118 | n5492 ;
  assign n5489 = n1865 | n4007 ;
  assign n5490 = n5489 ^ n4827 ^ 1'b0 ;
  assign n5491 = n4344 & ~n5490 ;
  assign n5494 = n5493 ^ n5491 ^ 1'b0 ;
  assign n5488 = n1121 | n1652 ;
  assign n5495 = n5494 ^ n5488 ^ 1'b0 ;
  assign n5496 = ~n869 & n5312 ;
  assign n5497 = ~x84 & n5496 ;
  assign n5498 = ~n2328 & n2414 ;
  assign n5499 = n5498 ^ n3417 ^ 1'b0 ;
  assign n5500 = n3698 ^ n1289 ^ n446 ;
  assign n5501 = n238 & ~n3561 ;
  assign n5502 = n5501 ^ n2174 ^ 1'b0 ;
  assign n5503 = n5500 | n5502 ;
  assign n5504 = n2452 | n4793 ;
  assign n5505 = n3579 ^ n1758 ^ 1'b0 ;
  assign n5506 = n5505 ^ n1603 ^ 1'b0 ;
  assign n5507 = n3986 ^ n1675 ^ n1329 ;
  assign n5508 = n3400 ^ n747 ^ 1'b0 ;
  assign n5509 = n273 & n556 ;
  assign n5510 = n5509 ^ n4340 ^ 1'b0 ;
  assign n5511 = x13 & x95 ;
  assign n5512 = ~n1929 & n5511 ;
  assign n5513 = n916 & n5512 ;
  assign n5514 = n4155 ^ n475 ^ 1'b0 ;
  assign n5515 = n5513 | n5514 ;
  assign n5516 = n5515 ^ n4892 ^ 1'b0 ;
  assign n5517 = n5092 ^ n386 ^ 1'b0 ;
  assign n5518 = n2206 | n5517 ;
  assign n5519 = n5518 ^ n1895 ^ 1'b0 ;
  assign n5520 = x124 & ~n682 ;
  assign n5521 = ~n1177 & n5520 ;
  assign n5522 = n861 & ~n5521 ;
  assign n5523 = n1617 & ~n5522 ;
  assign n5524 = x85 & n2033 ;
  assign n5525 = x6 & ~n1842 ;
  assign n5526 = n5525 ^ n1754 ^ 1'b0 ;
  assign n5527 = n2427 | n5526 ;
  assign n5528 = n5527 ^ n2108 ^ 1'b0 ;
  assign n5529 = n3188 & ~n5528 ;
  assign n5530 = n5189 ^ n3527 ^ 1'b0 ;
  assign n5531 = ~n2412 & n5530 ;
  assign n5532 = n4567 ^ n913 ^ 1'b0 ;
  assign n5533 = n5531 & ~n5532 ;
  assign n5534 = ~n4973 & n5533 ;
  assign n5535 = n2697 & n5534 ;
  assign n5536 = n1233 & ~n3180 ;
  assign n5537 = n5536 ^ n4840 ^ n1803 ;
  assign n5538 = ~n3210 & n4007 ;
  assign n5539 = n2910 ^ n2816 ^ 1'b0 ;
  assign n5540 = n5539 ^ n293 ^ 1'b0 ;
  assign n5541 = n3653 ^ n147 ^ 1'b0 ;
  assign n5542 = n5540 & n5541 ;
  assign n5543 = n1176 ^ n632 ^ 1'b0 ;
  assign n5544 = n904 & ~n5543 ;
  assign n5545 = n472 | n869 ;
  assign n5546 = n195 | n5545 ;
  assign n5547 = n5546 ^ n2132 ^ 1'b0 ;
  assign n5548 = ~n2809 & n5547 ;
  assign n5549 = ( n1566 & n1973 ) | ( n1566 & ~n2536 ) | ( n1973 & ~n2536 ) ;
  assign n5550 = n640 & n5549 ;
  assign n5551 = n2159 & ~n5550 ;
  assign n5552 = n5551 ^ n3573 ^ 1'b0 ;
  assign n5553 = n5548 | n5552 ;
  assign n5554 = n2710 & ~n5553 ;
  assign n5555 = n384 & ~n1021 ;
  assign n5556 = ~x53 & n5555 ;
  assign n5557 = n5556 ^ n4413 ^ 1'b0 ;
  assign n5558 = n1052 & n5557 ;
  assign n5559 = n5558 ^ n2135 ^ 1'b0 ;
  assign n5560 = ~n5244 & n5559 ;
  assign n5561 = ~n1361 & n5560 ;
  assign n5562 = n2268 & ~n3404 ;
  assign n5563 = n2774 ^ n993 ^ 1'b0 ;
  assign n5564 = n1985 & n5563 ;
  assign n5565 = n986 & n5564 ;
  assign n5566 = n5565 ^ n2787 ^ 1'b0 ;
  assign n5567 = n5566 ^ n2925 ^ 1'b0 ;
  assign n5568 = ~n5562 & n5567 ;
  assign n5569 = n860 & n3949 ;
  assign n5571 = x18 & ~x54 ;
  assign n5570 = ~n1395 & n4440 ;
  assign n5572 = n5571 ^ n5570 ^ 1'b0 ;
  assign n5573 = n5572 ^ n3533 ^ 1'b0 ;
  assign n5574 = x101 | n1270 ;
  assign n5575 = n147 & n1271 ;
  assign n5576 = n3442 ^ n2910 ^ 1'b0 ;
  assign n5577 = n5576 ^ n941 ^ n351 ;
  assign n5578 = n3982 ^ x122 ^ 1'b0 ;
  assign n5579 = ~n1779 & n1838 ;
  assign n5580 = n4055 & n5579 ;
  assign n5581 = ~n506 & n4295 ;
  assign n5582 = n5580 & n5581 ;
  assign n5583 = x100 | n4560 ;
  assign n5584 = n5583 ^ x110 ^ 1'b0 ;
  assign n5585 = n767 & n954 ;
  assign n5586 = n5585 ^ n1581 ^ 1'b0 ;
  assign n5587 = n5586 ^ n1113 ^ 1'b0 ;
  assign n5588 = n5584 & ~n5587 ;
  assign n5589 = ~n732 & n1271 ;
  assign n5590 = n5589 ^ n538 ^ 1'b0 ;
  assign n5591 = n5590 ^ n4307 ^ 1'b0 ;
  assign n5592 = n1849 & ~n5591 ;
  assign n5593 = n769 | n1823 ;
  assign n5594 = ~n3498 & n5593 ;
  assign n5595 = n2450 & ~n5594 ;
  assign n5596 = n826 & ~n2274 ;
  assign n5597 = n4623 & n5596 ;
  assign n5598 = n2810 ^ x34 ^ 1'b0 ;
  assign n5599 = n4919 ^ n3986 ^ 1'b0 ;
  assign n5600 = n1240 & ~n5107 ;
  assign n5601 = ~n903 & n2735 ;
  assign n5602 = n5601 ^ n4142 ^ 1'b0 ;
  assign n5603 = n5602 ^ n2468 ^ 1'b0 ;
  assign n5604 = n697 & n1688 ;
  assign n5605 = ~n4335 & n5604 ;
  assign n5606 = ~n145 & n2712 ;
  assign n5607 = n2237 ^ n1523 ^ 1'b0 ;
  assign n5608 = n5223 & ~n5607 ;
  assign n5609 = n794 & n3972 ;
  assign n5610 = n2866 & n5609 ;
  assign n5611 = n5610 ^ n3397 ^ 1'b0 ;
  assign n5617 = n273 & n3476 ;
  assign n5618 = n5617 ^ n3965 ^ 1'b0 ;
  assign n5612 = n1983 ^ n538 ^ 1'b0 ;
  assign n5613 = x90 & n5612 ;
  assign n5614 = n5613 ^ n3685 ^ n3236 ;
  assign n5615 = n5614 ^ n3497 ^ n1380 ;
  assign n5616 = n5615 ^ n3135 ^ 1'b0 ;
  assign n5619 = n5618 ^ n5616 ^ 1'b0 ;
  assign n5620 = ~n3165 & n5619 ;
  assign n5621 = n1574 | n3921 ;
  assign n5622 = n3561 & ~n5621 ;
  assign n5623 = n3362 ^ n695 ^ 1'b0 ;
  assign n5624 = n632 ^ n466 ^ 1'b0 ;
  assign n5625 = n5624 ^ n205 ^ 1'b0 ;
  assign n5626 = ~n1686 & n5625 ;
  assign n5627 = n3165 & n5626 ;
  assign n5628 = n2938 & ~n5627 ;
  assign n5629 = n5628 ^ n2642 ^ 1'b0 ;
  assign n5630 = n4994 | n5629 ;
  assign n5631 = x69 | n754 ;
  assign n5632 = ~n517 & n1336 ;
  assign n5633 = n1538 | n3948 ;
  assign n5634 = n5633 ^ n4545 ^ 1'b0 ;
  assign n5635 = n2748 | n2909 ;
  assign n5636 = n2983 ^ n1750 ^ 1'b0 ;
  assign n5637 = n5635 & ~n5636 ;
  assign n5638 = n5637 ^ n643 ^ 1'b0 ;
  assign n5639 = n5634 | n5638 ;
  assign n5640 = n5639 ^ n1847 ^ 1'b0 ;
  assign n5641 = ~n5632 & n5640 ;
  assign n5642 = ~n5631 & n5641 ;
  assign n5643 = n4319 ^ n1237 ^ 1'b0 ;
  assign n5644 = n660 & ~n2987 ;
  assign n5645 = ~n215 & n2405 ;
  assign n5646 = ~n2821 & n5645 ;
  assign n5647 = n2020 ^ n1413 ^ 1'b0 ;
  assign n5648 = n5245 ^ n3632 ^ 1'b0 ;
  assign n5650 = n4112 ^ n1343 ^ n1192 ;
  assign n5649 = n1572 ^ n1040 ^ 1'b0 ;
  assign n5651 = n5650 ^ n5649 ^ 1'b0 ;
  assign n5652 = n2537 | n2648 ;
  assign n5653 = n2762 & n5652 ;
  assign n5654 = ~n1003 & n2270 ;
  assign n5655 = n5654 ^ n5033 ^ 1'b0 ;
  assign n5656 = n5655 ^ n2078 ^ 1'b0 ;
  assign n5657 = n5653 & n5656 ;
  assign n5658 = ~n950 & n1350 ;
  assign n5659 = ~n1350 & n5658 ;
  assign n5660 = n918 | n5659 ;
  assign n5661 = x66 | n5660 ;
  assign n5662 = ( n1070 & n1404 ) | ( n1070 & n3392 ) | ( n1404 & n3392 ) ;
  assign n5663 = n2067 ^ n1005 ^ 1'b0 ;
  assign n5664 = n5662 | n5663 ;
  assign n5665 = ( n362 & n411 ) | ( n362 & n5664 ) | ( n411 & n5664 ) ;
  assign n5666 = n5665 ^ x41 ^ 1'b0 ;
  assign n5667 = n4020 ^ n2645 ^ n896 ;
  assign n5668 = n5340 ^ n2685 ^ 1'b0 ;
  assign n5669 = ~n5667 & n5668 ;
  assign n5670 = n1252 & n5554 ;
  assign n5671 = n5473 ^ n1198 ^ 1'b0 ;
  assign n5672 = n2497 | n4432 ;
  assign n5673 = n3331 & n5672 ;
  assign n5674 = ~n2658 & n5673 ;
  assign n5675 = ~n2635 & n5470 ;
  assign n5676 = n5675 ^ n5290 ^ 1'b0 ;
  assign n5677 = n2455 | n5676 ;
  assign n5678 = n2516 ^ x75 ^ 1'b0 ;
  assign n5679 = n1722 | n5678 ;
  assign n5680 = n5679 ^ x105 ^ 1'b0 ;
  assign n5681 = n791 & n3118 ;
  assign n5682 = n3049 & n5681 ;
  assign n5683 = n4648 & n5682 ;
  assign n5684 = n1510 | n1861 ;
  assign n5685 = ( n1996 & n5026 ) | ( n1996 & n5684 ) | ( n5026 & n5684 ) ;
  assign n5686 = ~x103 & n5685 ;
  assign n5687 = n2937 & n5686 ;
  assign n5690 = x15 & ~n5018 ;
  assign n5691 = n345 & n5690 ;
  assign n5688 = n4992 ^ n1342 ^ 1'b0 ;
  assign n5689 = n2140 & n5688 ;
  assign n5692 = n5691 ^ n5689 ^ 1'b0 ;
  assign n5693 = ( x23 & ~n317 ) | ( x23 & n1804 ) | ( ~n317 & n1804 ) ;
  assign n5694 = ~n4786 & n5693 ;
  assign n5695 = ~n2840 & n2946 ;
  assign n5696 = n4292 & n5695 ;
  assign n5697 = n2717 & ~n5654 ;
  assign n5698 = n5697 ^ n318 ^ 1'b0 ;
  assign n5699 = n1325 | n2758 ;
  assign n5700 = ~n3186 & n3806 ;
  assign n5701 = n5700 ^ n5161 ^ 1'b0 ;
  assign n5702 = n1830 ^ n888 ^ x119 ;
  assign n5703 = n1053 | n1128 ;
  assign n5704 = n1012 & ~n5703 ;
  assign n5705 = ~n5702 & n5704 ;
  assign n5706 = n5151 | n5705 ;
  assign n5707 = n5701 & ~n5706 ;
  assign n5708 = n2561 & n5644 ;
  assign n5709 = n5708 ^ n759 ^ 1'b0 ;
  assign n5711 = n669 | n2434 ;
  assign n5712 = n505 & ~n3990 ;
  assign n5713 = ~n5711 & n5712 ;
  assign n5714 = n5713 ^ n2054 ^ 1'b0 ;
  assign n5715 = n822 & n5714 ;
  assign n5710 = n3717 ^ n900 ^ 1'b0 ;
  assign n5716 = n5715 ^ n5710 ^ n559 ;
  assign n5717 = x24 & n604 ;
  assign n5718 = n1421 & n5717 ;
  assign n5719 = ~n551 & n5637 ;
  assign n5720 = n5429 & n5719 ;
  assign n5721 = n414 ^ x38 ^ 1'b0 ;
  assign n5722 = n5577 ^ n4066 ^ 1'b0 ;
  assign n5723 = n1120 & ~n3237 ;
  assign n5724 = n1024 ^ n794 ^ 1'b0 ;
  assign n5725 = n1728 & n5724 ;
  assign n5726 = ~n5723 & n5725 ;
  assign n5727 = n254 ^ x32 ^ 1'b0 ;
  assign n5728 = n5727 ^ n4578 ^ 1'b0 ;
  assign n5729 = n1743 & n3978 ;
  assign n5730 = ~n4161 & n5729 ;
  assign n5731 = n2992 & n3283 ;
  assign n5732 = n3896 ^ n1261 ^ n292 ;
  assign n5733 = n4061 ^ n2014 ^ 1'b0 ;
  assign n5734 = ~n5732 & n5733 ;
  assign n5735 = n5734 ^ n825 ^ 1'b0 ;
  assign n5737 = n5342 ^ n2324 ^ 1'b0 ;
  assign n5736 = ~n1190 & n3336 ;
  assign n5738 = n5737 ^ n5736 ^ 1'b0 ;
  assign n5739 = ~n1042 & n3543 ;
  assign n5740 = n1317 ^ n1058 ^ 1'b0 ;
  assign n5741 = n190 & n4128 ;
  assign n5742 = n4917 ^ n809 ^ 1'b0 ;
  assign n5743 = x115 & n1898 ;
  assign n5744 = n5743 ^ n3404 ^ 1'b0 ;
  assign n5745 = ~x100 & n5744 ;
  assign n5746 = n4901 ^ n2484 ^ 1'b0 ;
  assign n5747 = n4308 | n5746 ;
  assign n5749 = n890 | n5443 ;
  assign n5750 = n559 | n5749 ;
  assign n5751 = n5750 ^ n2452 ^ n824 ;
  assign n5748 = n4203 | n4650 ;
  assign n5752 = n5751 ^ n5748 ^ 1'b0 ;
  assign n5758 = ~n760 & n2709 ;
  assign n5753 = x20 & n273 ;
  assign n5754 = ~n2499 & n5753 ;
  assign n5755 = n5754 ^ n2333 ^ 1'b0 ;
  assign n5756 = n3890 & ~n5755 ;
  assign n5757 = n5179 & n5756 ;
  assign n5759 = n5758 ^ n5757 ^ 1'b0 ;
  assign n5760 = n2153 | n4318 ;
  assign n5761 = n1152 | n1469 ;
  assign n5762 = n3887 & ~n5761 ;
  assign n5763 = ~n2635 & n3606 ;
  assign n5765 = ~n1703 & n2742 ;
  assign n5766 = n1718 & n5765 ;
  assign n5764 = n3236 ^ x37 ^ 1'b0 ;
  assign n5767 = n5766 ^ n5764 ^ 1'b0 ;
  assign n5768 = n3171 & ~n5767 ;
  assign n5769 = n3816 ^ n849 ^ 1'b0 ;
  assign n5770 = n600 | n5769 ;
  assign n5771 = n5770 ^ n2028 ^ 1'b0 ;
  assign n5772 = ~n1874 & n5771 ;
  assign n5781 = n2340 & ~n2444 ;
  assign n5782 = n5781 ^ n1166 ^ 1'b0 ;
  assign n5783 = ~n1579 & n5782 ;
  assign n5774 = ( x6 & n496 ) | ( x6 & ~n1159 ) | ( n496 & ~n1159 ) ;
  assign n5775 = n5774 ^ n305 ^ 1'b0 ;
  assign n5773 = n5015 | n5758 ;
  assign n5776 = n5775 ^ n5773 ^ 1'b0 ;
  assign n5777 = n3455 ^ n1748 ^ 1'b0 ;
  assign n5778 = n5776 & n5777 ;
  assign n5779 = n387 & n5778 ;
  assign n5780 = n2483 & n5779 ;
  assign n5784 = n5783 ^ n5780 ^ 1'b0 ;
  assign n5786 = ~x101 & n3246 ;
  assign n5787 = n5786 ^ n2662 ^ 1'b0 ;
  assign n5788 = n1757 & n5787 ;
  assign n5789 = ~n632 & n5788 ;
  assign n5785 = n709 ^ x62 ^ 1'b0 ;
  assign n5790 = n5789 ^ n5785 ^ 1'b0 ;
  assign n5791 = ~x8 & n1411 ;
  assign n5792 = n5791 ^ n1835 ^ 1'b0 ;
  assign n5793 = n1767 | n5651 ;
  assign n5794 = n1479 & ~n5793 ;
  assign n5795 = n1810 | n5208 ;
  assign n5796 = n486 | n5795 ;
  assign n5797 = n5563 & n5796 ;
  assign n5798 = ~n1790 & n5797 ;
  assign n5799 = n2658 ^ n2125 ^ x58 ;
  assign n5800 = n3017 | n5799 ;
  assign n5801 = n5800 ^ n1256 ^ 1'b0 ;
  assign n5802 = n2925 | n5801 ;
  assign n5803 = n3219 ^ n620 ^ n276 ;
  assign n5804 = n5803 ^ n749 ^ 1'b0 ;
  assign n5805 = n5804 ^ n2720 ^ 1'b0 ;
  assign n5806 = ~n499 & n4626 ;
  assign n5807 = n1794 | n2107 ;
  assign n5808 = n2949 & ~n5807 ;
  assign n5809 = n5806 & n5808 ;
  assign n5810 = ~n971 & n2078 ;
  assign n5811 = n540 & ~n5810 ;
  assign n5812 = n1285 & n5811 ;
  assign n5813 = ( n2313 & ~n2910 ) | ( n2313 & n3795 ) | ( ~n2910 & n3795 ) ;
  assign n5814 = ( x47 & ~n5812 ) | ( x47 & n5813 ) | ( ~n5812 & n5813 ) ;
  assign n5815 = n745 & n4694 ;
  assign n5816 = n4032 & n5815 ;
  assign n5817 = n2220 ^ x11 ^ 1'b0 ;
  assign n5818 = ~n3056 & n5817 ;
  assign n5819 = n5818 ^ n1107 ^ 1'b0 ;
  assign n5820 = n3059 & ~n5240 ;
  assign n5821 = n456 | n542 ;
  assign n5822 = n152 & ~n5821 ;
  assign n5823 = ~n1568 & n3395 ;
  assign n5824 = n5823 ^ n4628 ^ 1'b0 ;
  assign n5825 = n5822 | n5824 ;
  assign n5826 = ~n925 & n1917 ;
  assign n5827 = n5826 ^ n5739 ^ n3884 ;
  assign n5828 = ~n4653 & n4820 ;
  assign n5829 = n3824 ^ n2492 ^ n1115 ;
  assign n5830 = ( n157 & ~n4420 ) | ( n157 & n5829 ) | ( ~n4420 & n5829 ) ;
  assign n5831 = n888 & ~n3167 ;
  assign n5832 = n5831 ^ n2515 ^ 1'b0 ;
  assign n5833 = n5832 ^ n4768 ^ 1'b0 ;
  assign n5834 = n5830 & ~n5833 ;
  assign n5835 = n4210 ^ n3142 ^ 1'b0 ;
  assign n5836 = n1212 & ~n5835 ;
  assign n5837 = ~n239 & n2529 ;
  assign n5839 = n5092 ^ n150 ^ 1'b0 ;
  assign n5838 = n2885 & n3717 ;
  assign n5840 = n5839 ^ n5838 ^ 1'b0 ;
  assign n5841 = n5837 | n5840 ;
  assign n5842 = n3575 ^ n415 ^ n256 ;
  assign n5844 = n1495 ^ n702 ^ 1'b0 ;
  assign n5843 = n2185 ^ n2087 ^ 1'b0 ;
  assign n5845 = n5844 ^ n5843 ^ 1'b0 ;
  assign n5846 = n138 & ~n1719 ;
  assign n5847 = n4990 ^ n4800 ^ 1'b0 ;
  assign n5848 = n5846 & ~n5847 ;
  assign n5849 = n876 & ~n2823 ;
  assign n5850 = n3790 ^ n3439 ^ 1'b0 ;
  assign n5851 = n3606 ^ n1612 ^ 1'b0 ;
  assign n5852 = n2010 | n5851 ;
  assign n5853 = ( ~n4867 & n5779 ) | ( ~n4867 & n5852 ) | ( n5779 & n5852 ) ;
  assign n5854 = n5853 ^ x97 ^ 1'b0 ;
  assign n5855 = ~n145 & n147 ;
  assign n5856 = n484 | n2068 ;
  assign n5857 = n5855 | n5856 ;
  assign n5858 = n5857 ^ n175 ^ 1'b0 ;
  assign n5859 = n2000 | n4708 ;
  assign n5860 = n1176 ^ n632 ^ n327 ;
  assign n5861 = n5315 ^ n4168 ^ 1'b0 ;
  assign n5862 = n5860 & n5861 ;
  assign n5863 = n2694 | n2989 ;
  assign n5864 = n5863 ^ n498 ^ 1'b0 ;
  assign n5865 = n2810 | n5864 ;
  assign n5866 = n2597 & n4742 ;
  assign n5867 = ~n2200 & n5866 ;
  assign n5868 = n3485 ^ n1545 ^ 1'b0 ;
  assign n5869 = n2518 & ~n5868 ;
  assign n5870 = n5869 ^ n323 ^ 1'b0 ;
  assign n5871 = n4279 ^ n2961 ^ n1719 ;
  assign n5872 = ( n1705 & n5365 ) | ( n1705 & n5871 ) | ( n5365 & n5871 ) ;
  assign n5873 = n933 & ~n1469 ;
  assign n5874 = n5873 ^ n813 ^ 1'b0 ;
  assign n5875 = n4230 & n5544 ;
  assign n5876 = ~n5874 & n5875 ;
  assign n5877 = x107 & n355 ;
  assign n5878 = n5877 ^ n5093 ^ 1'b0 ;
  assign n5879 = n406 & n5878 ;
  assign n5884 = n2361 & n3039 ;
  assign n5885 = n5884 ^ n587 ^ 1'b0 ;
  assign n5881 = n1737 & n1893 ;
  assign n5882 = n1867 & n5881 ;
  assign n5880 = n1046 | n3999 ;
  assign n5883 = n5882 ^ n5880 ^ 1'b0 ;
  assign n5886 = n5885 ^ n5883 ^ 1'b0 ;
  assign n5887 = n1931 ^ n202 ^ 1'b0 ;
  assign n5888 = n5887 ^ n1372 ^ 1'b0 ;
  assign n5889 = n3136 | n5888 ;
  assign n5890 = n1865 & ~n5889 ;
  assign n5891 = n5890 ^ n2116 ^ 1'b0 ;
  assign n5892 = n882 & ~n2323 ;
  assign n5893 = n3408 & n5892 ;
  assign n5894 = n5863 ^ n642 ^ n161 ;
  assign n5895 = n5894 ^ n5613 ^ 1'b0 ;
  assign n5896 = n349 & ~n5895 ;
  assign n5897 = n5893 | n5896 ;
  assign n5898 = n2246 | n5897 ;
  assign n5899 = n5898 ^ n4901 ^ 1'b0 ;
  assign n5900 = n238 ^ x59 ^ 1'b0 ;
  assign n5901 = n3698 & ~n5900 ;
  assign n5902 = n931 | n5901 ;
  assign n5903 = ~n3601 & n5902 ;
  assign n5904 = n4448 & n5903 ;
  assign n5905 = n2499 | n2946 ;
  assign n5906 = n1758 | n5011 ;
  assign n5907 = n1842 ^ n417 ^ 1'b0 ;
  assign n5908 = n740 & n5907 ;
  assign n5909 = n5908 ^ n2777 ^ 1'b0 ;
  assign n5910 = ~n1133 & n2724 ;
  assign n5911 = n5910 ^ n3456 ^ 1'b0 ;
  assign n5913 = n4236 ^ n1642 ^ 1'b0 ;
  assign n5914 = n3350 & n5913 ;
  assign n5912 = n2378 & ~n4357 ;
  assign n5915 = n5914 ^ n5912 ^ 1'b0 ;
  assign n5918 = ~n1953 & n5260 ;
  assign n5916 = n172 & ~n3503 ;
  assign n5917 = n5916 ^ n4251 ^ n3279 ;
  assign n5919 = n5918 ^ n5917 ^ 1'b0 ;
  assign n5920 = n5915 | n5919 ;
  assign n5921 = n5351 & n5536 ;
  assign n5922 = n3948 ^ n196 ^ 1'b0 ;
  assign n5923 = n3587 & ~n5922 ;
  assign n5924 = n3839 & n5923 ;
  assign n5925 = ~n4927 & n5924 ;
  assign n5926 = ~n3533 & n3795 ;
  assign n5927 = ~n1433 & n5926 ;
  assign n5928 = n387 & ~n5927 ;
  assign n5929 = n973 ^ x31 ^ 1'b0 ;
  assign n5930 = ~n1880 & n5929 ;
  assign n5931 = n4134 ^ n2869 ^ n1481 ;
  assign n5932 = ~n2455 & n2527 ;
  assign n5933 = ~n675 & n5932 ;
  assign n5934 = ~n147 & n4697 ;
  assign n5935 = n4960 & n5191 ;
  assign n5936 = n5569 ^ n923 ^ 1'b0 ;
  assign n5937 = n5935 & ~n5936 ;
  assign n5938 = ~n2167 & n3991 ;
  assign n5939 = n5938 ^ n3858 ^ 1'b0 ;
  assign n5940 = n5939 ^ n2523 ^ 1'b0 ;
  assign n5941 = n533 | n5940 ;
  assign n5942 = ( n882 & ~n2172 ) | ( n882 & n5277 ) | ( ~n2172 & n5277 ) ;
  assign n5943 = n886 | n5566 ;
  assign n5944 = n5943 ^ n2154 ^ 1'b0 ;
  assign n5945 = n1132 & ~n5944 ;
  assign n5946 = n2961 ^ n174 ^ 1'b0 ;
  assign n5947 = n4359 ^ n845 ^ 1'b0 ;
  assign n5948 = n796 | n5947 ;
  assign n5949 = n5948 ^ n2339 ^ 1'b0 ;
  assign n5950 = ( n1662 & n5946 ) | ( n1662 & ~n5949 ) | ( n5946 & ~n5949 ) ;
  assign n5951 = n138 | n3017 ;
  assign n5952 = ~n256 & n1192 ;
  assign n5953 = n5684 ^ n3112 ^ 1'b0 ;
  assign n5954 = ~n725 & n5953 ;
  assign n5957 = ~n2419 & n4171 ;
  assign n5955 = n642 & ~n2075 ;
  assign n5956 = ~n1527 & n5955 ;
  assign n5958 = n5957 ^ n5956 ^ 1'b0 ;
  assign n5959 = n1103 | n5958 ;
  assign n5960 = ~n667 & n1497 ;
  assign n5961 = n5960 ^ n1391 ^ 1'b0 ;
  assign n5962 = n2551 ^ n2003 ^ n1767 ;
  assign n5963 = n5962 ^ n976 ^ 1'b0 ;
  assign n5964 = n540 & n3431 ;
  assign n5965 = n5964 ^ n4076 ^ 1'b0 ;
  assign n5966 = n1956 & ~n5965 ;
  assign n5967 = ~n506 & n1469 ;
  assign n5968 = n3998 & n4661 ;
  assign n5969 = n2324 & ~n5968 ;
  assign n5970 = n1647 & ~n3415 ;
  assign n5971 = ~n3809 & n5970 ;
  assign n5972 = n1111 & n5971 ;
  assign n5973 = ( n997 & n1167 ) | ( n997 & ~n5193 ) | ( n1167 & ~n5193 ) ;
  assign n5974 = n347 | n5973 ;
  assign n5975 = n1743 ^ n1726 ^ 1'b0 ;
  assign n5976 = ~n2782 & n5975 ;
  assign n5977 = n5974 & ~n5976 ;
  assign n5980 = x39 | n1038 ;
  assign n5978 = n1412 | n5855 ;
  assign n5979 = n3933 & n5978 ;
  assign n5981 = n5980 ^ n5979 ^ 1'b0 ;
  assign n5982 = n459 & n5981 ;
  assign n5983 = n364 & n5982 ;
  assign n5984 = n5274 ^ n1046 ^ 1'b0 ;
  assign n5985 = n2883 & n5984 ;
  assign n5986 = ( n915 & n1270 ) | ( n915 & n1809 ) | ( n1270 & n1809 ) ;
  assign n5987 = n4542 & n4953 ;
  assign n5988 = n5987 ^ n3287 ^ 1'b0 ;
  assign n5989 = n5986 | n5988 ;
  assign n5990 = ~n400 & n3616 ;
  assign n5991 = n5990 ^ n2274 ^ 1'b0 ;
  assign n5992 = n2513 & ~n5991 ;
  assign n5993 = n1396 & n4215 ;
  assign n5994 = n319 & n4364 ;
  assign n5995 = n5994 ^ n4408 ^ 1'b0 ;
  assign n5996 = n1912 & ~n5995 ;
  assign n5997 = ( ~n409 & n5207 ) | ( ~n409 & n5996 ) | ( n5207 & n5996 ) ;
  assign n5998 = n5703 ^ n355 ^ 1'b0 ;
  assign n5999 = ~n1390 & n5998 ;
  assign n6000 = n642 & n939 ;
  assign n6001 = n5908 & ~n6000 ;
  assign n6002 = ~n5999 & n6001 ;
  assign n6003 = n1620 ^ n509 ^ 1'b0 ;
  assign n6004 = n660 & ~n4833 ;
  assign n6005 = ( x52 & n2575 ) | ( x52 & ~n6004 ) | ( n2575 & ~n6004 ) ;
  assign n6006 = n6005 ^ n4175 ^ 1'b0 ;
  assign n6007 = n559 ^ x6 ^ 1'b0 ;
  assign n6008 = ~n2293 & n2617 ;
  assign n6009 = n6008 ^ n3982 ^ 1'b0 ;
  assign n6013 = n1575 ^ n256 ^ 1'b0 ;
  assign n6010 = x113 & n139 ;
  assign n6011 = ~n1745 & n6010 ;
  assign n6012 = n388 & ~n6011 ;
  assign n6014 = n6013 ^ n6012 ^ 1'b0 ;
  assign n6015 = n6009 | n6014 ;
  assign n6016 = n6007 & ~n6015 ;
  assign n6017 = n6016 ^ n5040 ^ 1'b0 ;
  assign n6018 = ( n2768 & ~n2846 ) | ( n2768 & n3310 ) | ( ~n2846 & n3310 ) ;
  assign n6019 = n3025 & n6018 ;
  assign n6020 = n3372 & n3687 ;
  assign n6022 = n1291 & ~n3249 ;
  assign n6021 = n838 ^ x98 ^ 1'b0 ;
  assign n6023 = n6022 ^ n6021 ^ n4238 ;
  assign n6024 = ~n1024 & n4963 ;
  assign n6025 = ~n4389 & n6024 ;
  assign n6026 = n440 | n2652 ;
  assign n6027 = n6026 ^ n4311 ^ 1'b0 ;
  assign n6028 = n2759 ^ n2324 ^ 1'b0 ;
  assign n6029 = n6027 & n6028 ;
  assign n6030 = n1134 ^ n400 ^ n362 ;
  assign n6031 = n548 ^ x110 ^ 1'b0 ;
  assign n6032 = n2091 & ~n6031 ;
  assign n6033 = n6032 ^ n1953 ^ 1'b0 ;
  assign n6034 = n6030 | n6033 ;
  assign n6035 = n3138 ^ n425 ^ 1'b0 ;
  assign n6036 = n6035 ^ n2084 ^ 1'b0 ;
  assign n6037 = n3226 ^ n2233 ^ n1279 ;
  assign n6038 = n3048 & n6037 ;
  assign n6039 = n3806 & n5226 ;
  assign n6040 = n634 & ~n2193 ;
  assign n6041 = n6040 ^ n425 ^ 1'b0 ;
  assign n6042 = n6039 & n6041 ;
  assign n6043 = ~n4702 & n6042 ;
  assign n6044 = n892 | n2832 ;
  assign n6045 = n529 | n4171 ;
  assign n6046 = n4541 ^ n1432 ^ 1'b0 ;
  assign n6047 = n3339 & n6046 ;
  assign n6051 = n351 | n3165 ;
  assign n6048 = n5877 ^ n4890 ^ n3956 ;
  assign n6049 = n5539 ^ n2694 ^ 1'b0 ;
  assign n6050 = n6048 & n6049 ;
  assign n6052 = n6051 ^ n6050 ^ 1'b0 ;
  assign n6053 = n4583 ^ n3539 ^ 1'b0 ;
  assign n6054 = n2886 ^ n254 ^ 1'b0 ;
  assign n6055 = n4792 & n6054 ;
  assign n6056 = n1680 ^ n973 ^ 1'b0 ;
  assign n6057 = n649 & n1835 ;
  assign n6058 = ~n4824 & n6057 ;
  assign n6059 = n3606 & n6058 ;
  assign n6060 = n1733 & ~n1929 ;
  assign n6061 = n2060 | n3590 ;
  assign n6062 = n1623 & n6061 ;
  assign n6063 = x13 & ~n3010 ;
  assign n6064 = n6063 ^ n4053 ^ 1'b0 ;
  assign n6065 = n1189 & ~n6064 ;
  assign n6066 = ~n2499 & n6065 ;
  assign n6067 = n4430 ^ n2124 ^ x55 ;
  assign n6068 = n5883 | n6067 ;
  assign n6069 = n6068 ^ n3672 ^ 1'b0 ;
  assign n6070 = n4340 & n6069 ;
  assign n6071 = ~n471 & n6070 ;
  assign n6072 = n6071 ^ n2210 ^ n175 ;
  assign n6073 = n2948 ^ n2150 ^ 1'b0 ;
  assign n6074 = n589 | n2754 ;
  assign n6075 = ( n1594 & n3410 ) | ( n1594 & ~n6074 ) | ( n3410 & ~n6074 ) ;
  assign n6076 = n6075 ^ n3104 ^ 1'b0 ;
  assign n6077 = n6073 & ~n6076 ;
  assign n6078 = n6077 ^ n1057 ^ 1'b0 ;
  assign n6079 = n456 | n2276 ;
  assign n6080 = ~n2655 & n5550 ;
  assign n6081 = n1988 & n2806 ;
  assign n6082 = n6081 ^ n4678 ^ 1'b0 ;
  assign n6083 = n3518 | n6082 ;
  assign n6084 = n6083 ^ n971 ^ 1'b0 ;
  assign n6085 = n6080 & ~n6084 ;
  assign n6086 = n6079 & n6085 ;
  assign n6087 = ( ~n455 & n959 ) | ( ~n455 & n1758 ) | ( n959 & n1758 ) ;
  assign n6088 = n6087 ^ n4265 ^ 1'b0 ;
  assign n6089 = n1461 ^ n708 ^ 1'b0 ;
  assign n6090 = ~n1510 & n6089 ;
  assign n6091 = n6090 ^ n5511 ^ n1776 ;
  assign n6092 = n194 | n6091 ;
  assign n6093 = n3704 ^ n2144 ^ n1198 ;
  assign n6094 = n4088 & ~n6093 ;
  assign n6095 = n988 & n2213 ;
  assign n6096 = n6095 ^ x17 ^ 1'b0 ;
  assign n6097 = n1232 & n6096 ;
  assign n6098 = n4266 ^ n260 ^ 1'b0 ;
  assign n6099 = n3940 | n6098 ;
  assign n6100 = ~n851 & n2892 ;
  assign n6101 = n2917 & n6100 ;
  assign n6102 = n5855 ^ n808 ^ 1'b0 ;
  assign n6103 = ~n6101 & n6102 ;
  assign n6104 = ~n487 & n6103 ;
  assign n6105 = n4180 ^ n2070 ^ 1'b0 ;
  assign n6106 = n1386 | n6105 ;
  assign n6107 = n6106 ^ n4751 ^ 1'b0 ;
  assign n6108 = n1319 ^ n327 ^ 1'b0 ;
  assign n6109 = n6108 ^ n5549 ^ n3180 ;
  assign n6110 = n6109 ^ n2537 ^ 1'b0 ;
  assign n6111 = n3476 | n4329 ;
  assign n6114 = n1467 | n4319 ;
  assign n6112 = n5238 ^ n3140 ^ 1'b0 ;
  assign n6113 = n2715 & ~n6112 ;
  assign n6115 = n6114 ^ n6113 ^ 1'b0 ;
  assign n6116 = n2417 ^ n1920 ^ 1'b0 ;
  assign n6117 = ~n3226 & n6116 ;
  assign n6118 = n6117 ^ n3289 ^ 1'b0 ;
  assign n6119 = n2812 | n2886 ;
  assign n6120 = n1862 & ~n6119 ;
  assign n6121 = n775 | n6120 ;
  assign n6122 = ( n633 & ~n1046 ) | ( n633 & n6121 ) | ( ~n1046 & n6121 ) ;
  assign n6124 = n1541 | n2931 ;
  assign n6123 = ~n639 & n5879 ;
  assign n6125 = n6124 ^ n6123 ^ 1'b0 ;
  assign n6126 = n3921 | n6125 ;
  assign n6127 = n3171 ^ n892 ^ 1'b0 ;
  assign n6128 = ~n820 & n2330 ;
  assign n6129 = ~n6127 & n6128 ;
  assign n6130 = n4800 ^ x36 ^ 1'b0 ;
  assign n6131 = ~n1079 & n6130 ;
  assign n6132 = ~n637 & n2635 ;
  assign n6133 = ~n1672 & n6132 ;
  assign n6134 = ~n609 & n4352 ;
  assign n6135 = ~n6133 & n6134 ;
  assign n6136 = n6131 | n6135 ;
  assign n6137 = n4703 ^ n3674 ^ n1359 ;
  assign n6138 = n6137 ^ x31 ^ 1'b0 ;
  assign n6139 = n2905 ^ n977 ^ 1'b0 ;
  assign n6140 = ( n1405 & n2697 ) | ( n1405 & ~n6139 ) | ( n2697 & ~n6139 ) ;
  assign n6141 = n2556 ^ n675 ^ 1'b0 ;
  assign n6142 = n1225 | n6141 ;
  assign n6143 = n6142 ^ x62 ^ 1'b0 ;
  assign n6144 = n442 & ~n6143 ;
  assign n6151 = n5775 ^ n1520 ^ 1'b0 ;
  assign n6150 = n915 & n6139 ;
  assign n6152 = n6151 ^ n6150 ^ 1'b0 ;
  assign n6147 = n3174 ^ n2531 ^ 1'b0 ;
  assign n6145 = n198 & ~n2153 ;
  assign n6146 = ~n609 & n6145 ;
  assign n6148 = n6147 ^ n6146 ^ 1'b0 ;
  assign n6149 = n1026 & ~n6148 ;
  assign n6153 = n6152 ^ n6149 ^ 1'b0 ;
  assign n6154 = n6144 & ~n6153 ;
  assign n6155 = n6154 ^ n5191 ^ 1'b0 ;
  assign n6156 = n6155 ^ n1635 ^ 1'b0 ;
  assign n6157 = n1895 & n2158 ;
  assign n6158 = n3001 & ~n6087 ;
  assign n6159 = n1015 & n1623 ;
  assign n6160 = n6158 | n6159 ;
  assign n6161 = n6157 | n6160 ;
  assign n6164 = n311 & ~n4448 ;
  assign n6165 = ~n1524 & n6164 ;
  assign n6162 = n1140 & ~n2568 ;
  assign n6163 = n6162 ^ n2318 ^ 1'b0 ;
  assign n6166 = n6165 ^ n6163 ^ 1'b0 ;
  assign n6167 = n1601 & n3262 ;
  assign n6168 = ( ~n2319 & n2558 ) | ( ~n2319 & n6167 ) | ( n2558 & n6167 ) ;
  assign n6169 = n605 & n1426 ;
  assign n6170 = n4519 | n6169 ;
  assign n6171 = n6168 | n6170 ;
  assign n6172 = n299 & n1786 ;
  assign n6173 = n671 & n1067 ;
  assign n6174 = ~n6172 & n6173 ;
  assign n6175 = n4382 & n6163 ;
  assign n6176 = n6175 ^ n1128 ^ 1'b0 ;
  assign n6177 = n6174 | n6176 ;
  assign n6178 = n1969 & n2302 ;
  assign n6179 = n6178 ^ n6080 ^ 1'b0 ;
  assign n6180 = n5962 ^ n5549 ^ 1'b0 ;
  assign n6181 = ~n1190 & n6180 ;
  assign n6182 = n6032 | n6181 ;
  assign n6183 = n3719 ^ n1662 ^ 1'b0 ;
  assign n6184 = ~n414 & n6183 ;
  assign n6185 = n391 & n6184 ;
  assign n6186 = n3241 & n3749 ;
  assign n6187 = ~n2447 & n6186 ;
  assign n6188 = n945 & n5901 ;
  assign n6189 = ( n5857 & n6187 ) | ( n5857 & ~n6188 ) | ( n6187 & ~n6188 ) ;
  assign n6190 = x58 & ~n6189 ;
  assign n6191 = n2387 | n3402 ;
  assign n6192 = n427 & n857 ;
  assign n6193 = ~n6191 & n6192 ;
  assign n6194 = n2908 ^ n1219 ^ 1'b0 ;
  assign n6195 = n2772 | n6194 ;
  assign n6196 = n6195 ^ n3856 ^ 1'b0 ;
  assign n6197 = n332 & n6196 ;
  assign n6198 = n1761 | n1941 ;
  assign n6199 = n930 | n6198 ;
  assign n6200 = ~n5260 & n6199 ;
  assign n6201 = ~n6197 & n6200 ;
  assign n6202 = ( n1481 & n1791 ) | ( n1481 & ~n2146 ) | ( n1791 & ~n2146 ) ;
  assign n6203 = ~n2788 & n3816 ;
  assign n6204 = n6203 ^ n2188 ^ 1'b0 ;
  assign n6205 = n4833 ^ n664 ^ 1'b0 ;
  assign n6206 = n4330 ^ n3628 ^ 1'b0 ;
  assign n6208 = ( ~x123 & n883 ) | ( ~x123 & n2014 ) | ( n883 & n2014 ) ;
  assign n6209 = n1935 | n6075 ;
  assign n6210 = n6208 & ~n6209 ;
  assign n6207 = ( ~n589 & n926 ) | ( ~n589 & n933 ) | ( n926 & n933 ) ;
  assign n6211 = n6210 ^ n6207 ^ n2031 ;
  assign n6212 = ~n3361 & n6211 ;
  assign n6213 = n1711 | n6212 ;
  assign n6214 = n716 ^ n565 ^ 1'b0 ;
  assign n6215 = ~n2006 & n6214 ;
  assign n6216 = ~n6109 & n6215 ;
  assign n6217 = n1147 & n3055 ;
  assign n6218 = n6217 ^ n210 ^ 1'b0 ;
  assign n6219 = n1957 | n6218 ;
  assign n6220 = n6216 & ~n6219 ;
  assign n6221 = n1909 | n3000 ;
  assign n6222 = n3850 | n6221 ;
  assign n6223 = n6222 ^ n4519 ^ 1'b0 ;
  assign n6224 = x62 & ~n6223 ;
  assign n6225 = x90 ^ x42 ^ 1'b0 ;
  assign n6226 = n139 & n6225 ;
  assign n6227 = n2198 | n3101 ;
  assign n6228 = ~n4788 & n6227 ;
  assign n6229 = ~n6226 & n6228 ;
  assign n6230 = n5316 ^ n2295 ^ n1169 ;
  assign n6231 = n6147 ^ n2460 ^ 1'b0 ;
  assign n6232 = ~n3925 & n6231 ;
  assign n6233 = ( n5595 & ~n6230 ) | ( n5595 & n6232 ) | ( ~n6230 & n6232 ) ;
  assign n6234 = n1785 ^ n1552 ^ 1'b0 ;
  assign n6235 = ~n3675 & n6234 ;
  assign n6236 = n884 & n6235 ;
  assign n6237 = x13 | n3253 ;
  assign n6238 = n5054 & n6237 ;
  assign n6239 = n4007 | n4083 ;
  assign n6240 = n6239 ^ x124 ^ 1'b0 ;
  assign n6241 = ~n313 & n5774 ;
  assign n6242 = ~n6240 & n6241 ;
  assign n6243 = n6242 ^ n257 ^ 1'b0 ;
  assign n6244 = ~n2285 & n6243 ;
  assign n6245 = ~n6082 & n6244 ;
  assign n6246 = n3615 ^ n3339 ^ 1'b0 ;
  assign n6247 = n6246 ^ n6041 ^ n2353 ;
  assign n6248 = n3062 | n3762 ;
  assign n6249 = n3413 & n6248 ;
  assign n6250 = x85 & n3140 ;
  assign n6251 = ~n2854 & n6250 ;
  assign n6252 = n1414 ^ n945 ^ 1'b0 ;
  assign n6253 = n5234 & n6252 ;
  assign n6254 = n6253 ^ n735 ^ 1'b0 ;
  assign n6256 = n3873 ^ n1402 ^ 1'b0 ;
  assign n6255 = ( ~n1353 & n3214 ) | ( ~n1353 & n4513 ) | ( n3214 & n4513 ) ;
  assign n6257 = n6256 ^ n6255 ^ n4753 ;
  assign n6258 = n6257 ^ n2869 ^ 1'b0 ;
  assign n6259 = n1099 | n1794 ;
  assign n6260 = n676 & ~n6259 ;
  assign n6261 = ~n3672 & n6260 ;
  assign n6262 = n4616 | n6261 ;
  assign n6263 = n1728 | n6262 ;
  assign n6266 = n1710 ^ n1074 ^ 1'b0 ;
  assign n6267 = n6266 ^ n4448 ^ 1'b0 ;
  assign n6268 = ~n3000 & n6267 ;
  assign n6264 = ~n1769 & n3030 ;
  assign n6265 = n2717 & ~n6264 ;
  assign n6269 = n6268 ^ n6265 ^ 1'b0 ;
  assign n6273 = n1435 ^ n950 ^ 1'b0 ;
  assign n6270 = ~n2636 & n3483 ;
  assign n6271 = x19 & n6270 ;
  assign n6272 = n5586 & n6271 ;
  assign n6274 = n6273 ^ n6272 ^ 1'b0 ;
  assign n6275 = n6274 ^ n5797 ^ 1'b0 ;
  assign n6276 = n5193 & n5637 ;
  assign n6277 = n6276 ^ n2931 ^ 1'b0 ;
  assign n6278 = n488 & n4644 ;
  assign n6279 = ( n5275 & n6013 ) | ( n5275 & ~n6278 ) | ( n6013 & ~n6278 ) ;
  assign n6280 = n1510 & ~n2427 ;
  assign n6281 = n6279 & n6280 ;
  assign n6282 = n460 ^ n319 ^ 1'b0 ;
  assign n6283 = ~n6281 & n6282 ;
  assign n6284 = n1369 & ~n6283 ;
  assign n6285 = n1849 & ~n6284 ;
  assign n6286 = ~n6073 & n6285 ;
  assign n6287 = n2601 ^ n1183 ^ 1'b0 ;
  assign n6288 = ~n2006 & n6287 ;
  assign n6289 = n5859 ^ n335 ^ 1'b0 ;
  assign n6291 = n2013 ^ n147 ^ 1'b0 ;
  assign n6290 = n2504 ^ n1568 ^ 1'b0 ;
  assign n6292 = n6291 ^ n6290 ^ 1'b0 ;
  assign n6293 = n6292 ^ n2728 ^ n1150 ;
  assign n6294 = ~n1296 & n2937 ;
  assign n6295 = n2844 | n6294 ;
  assign n6296 = n4895 & n6295 ;
  assign n6297 = ~n2949 & n6296 ;
  assign n6298 = n6297 ^ n5973 ^ 1'b0 ;
  assign n6299 = n5344 | n6298 ;
  assign n6300 = ( ~n1211 & n2274 ) | ( ~n1211 & n3945 ) | ( n2274 & n3945 ) ;
  assign n6301 = n2312 & ~n6300 ;
  assign n6302 = n157 & ~n2151 ;
  assign n6303 = n6302 ^ n5477 ^ 1'b0 ;
  assign n6304 = n6303 ^ n2869 ^ 1'b0 ;
  assign n6305 = n6301 | n6304 ;
  assign n6306 = n3957 ^ n803 ^ 1'b0 ;
  assign n6307 = n1755 & ~n6306 ;
  assign n6308 = n4065 ^ n1446 ^ 1'b0 ;
  assign n6309 = n3494 | n6308 ;
  assign n6310 = ( n2917 & n3685 ) | ( n2917 & n4989 ) | ( n3685 & n4989 ) ;
  assign n6311 = n2278 & n6310 ;
  assign n6313 = n1827 ^ n371 ^ 1'b0 ;
  assign n6314 = n1485 | n6313 ;
  assign n6312 = ~n723 & n1738 ;
  assign n6315 = n6314 ^ n6312 ^ 1'b0 ;
  assign n6316 = n6315 ^ n3072 ^ 1'b0 ;
  assign n6317 = n3200 | n6316 ;
  assign n6318 = ~n3234 & n5033 ;
  assign n6319 = n6318 ^ n6112 ^ n922 ;
  assign n6320 = n1261 ^ x0 ^ 1'b0 ;
  assign n6321 = n1560 | n6320 ;
  assign n6322 = n6321 ^ n2115 ^ n1981 ;
  assign n6323 = ~n1483 & n6322 ;
  assign n6324 = n2494 & n3124 ;
  assign n6325 = n4727 ^ n3855 ^ 1'b0 ;
  assign n6326 = n1068 & n6325 ;
  assign n6329 = n1084 & ~n2604 ;
  assign n6330 = n6329 ^ n290 ^ 1'b0 ;
  assign n6327 = n2192 ^ n871 ^ 1'b0 ;
  assign n6328 = n5138 & ~n6327 ;
  assign n6331 = n6330 ^ n6328 ^ 1'b0 ;
  assign n6332 = n3806 & n5385 ;
  assign n6333 = n6332 ^ n3140 ^ 1'b0 ;
  assign n6334 = n3142 ^ n2476 ^ x11 ;
  assign n6335 = n874 & n6137 ;
  assign n6336 = ~n6334 & n6335 ;
  assign n6337 = n5638 ^ n4717 ^ 1'b0 ;
  assign n6338 = ~n2144 & n3019 ;
  assign n6339 = ~n277 & n6338 ;
  assign n6340 = n6337 | n6339 ;
  assign n6341 = n1661 | n5983 ;
  assign n6342 = n3625 & ~n6341 ;
  assign n6343 = n616 ^ x114 ^ 1'b0 ;
  assign n6344 = n5649 ^ n2647 ^ 1'b0 ;
  assign n6345 = ~n1581 & n6344 ;
  assign n6346 = n5857 & n6345 ;
  assign n6347 = n6346 ^ n5665 ^ 1'b0 ;
  assign n6348 = n3554 ^ x54 ^ 1'b0 ;
  assign n6349 = x17 & n2847 ;
  assign n6350 = n6349 ^ n174 ^ 1'b0 ;
  assign n6356 = n3914 ^ n930 ^ 1'b0 ;
  assign n6351 = n2684 & n2851 ;
  assign n6352 = ~n902 & n6351 ;
  assign n6353 = x35 & n575 ;
  assign n6354 = n6353 ^ n1642 ^ 1'b0 ;
  assign n6355 = n6352 & ~n6354 ;
  assign n6357 = n6356 ^ n6355 ^ 1'b0 ;
  assign n6358 = n4657 | n6357 ;
  assign n6359 = n6358 ^ n2991 ^ 1'b0 ;
  assign n6360 = n364 | n2183 ;
  assign n6361 = x98 & ~n6360 ;
  assign n6362 = n2419 | n2829 ;
  assign n6363 = n6362 ^ n4143 ^ 1'b0 ;
  assign n6364 = n2615 | n6363 ;
  assign n6365 = n6361 | n6364 ;
  assign n6366 = n3314 & ~n6365 ;
  assign n6367 = n444 | n3811 ;
  assign n6368 = ( ~n147 & n690 ) | ( ~n147 & n2137 ) | ( n690 & n2137 ) ;
  assign n6369 = n224 & ~n6368 ;
  assign n6370 = n6369 ^ n5579 ^ n1811 ;
  assign n6371 = n6370 ^ n2409 ^ n1880 ;
  assign n6372 = n6371 ^ n4019 ^ 1'b0 ;
  assign n6373 = n179 & n2165 ;
  assign n6374 = n6373 ^ n3795 ^ 1'b0 ;
  assign n6375 = n6374 ^ n4844 ^ 1'b0 ;
  assign n6376 = n3334 & ~n6375 ;
  assign n6377 = n2028 ^ n536 ^ 1'b0 ;
  assign n6378 = n989 & n6377 ;
  assign n6382 = n1609 ^ n1089 ^ n959 ;
  assign n6380 = ~n928 & n2174 ;
  assign n6381 = ~n1720 & n6380 ;
  assign n6383 = n6382 ^ n6381 ^ 1'b0 ;
  assign n6384 = n1303 & n6383 ;
  assign n6379 = n725 & n844 ;
  assign n6385 = n6384 ^ n6379 ^ 1'b0 ;
  assign n6386 = n6385 ^ n442 ^ 1'b0 ;
  assign n6387 = n4454 & ~n6386 ;
  assign n6388 = ~n6378 & n6387 ;
  assign n6389 = n2376 & n6388 ;
  assign n6390 = ~n1306 & n2985 ;
  assign n6391 = n1933 & n6390 ;
  assign n6392 = n6391 ^ n438 ^ 1'b0 ;
  assign n6393 = n1211 & ~n4128 ;
  assign n6394 = ~n1865 & n6393 ;
  assign n6395 = n4961 ^ n3411 ^ 1'b0 ;
  assign n6396 = ~n6394 & n6395 ;
  assign n6397 = ~n4125 & n5350 ;
  assign n6401 = n400 | n733 ;
  assign n6398 = n2338 & ~n5014 ;
  assign n6399 = n2951 | n6398 ;
  assign n6400 = n6399 ^ n6348 ^ n4299 ;
  assign n6402 = n6401 ^ n6400 ^ 1'b0 ;
  assign n6403 = n5120 & n6402 ;
  assign n6407 = n1250 & ~n6214 ;
  assign n6406 = n2771 & ~n2832 ;
  assign n6408 = n6407 ^ n6406 ^ 1'b0 ;
  assign n6404 = n3868 ^ n3062 ^ 1'b0 ;
  assign n6405 = n1353 | n6404 ;
  assign n6409 = n6408 ^ n6405 ^ 1'b0 ;
  assign n6410 = n1201 ^ n652 ^ 1'b0 ;
  assign n6411 = ( n1898 & n4936 ) | ( n1898 & ~n6410 ) | ( n4936 & ~n6410 ) ;
  assign n6412 = n2299 ^ n1155 ^ 1'b0 ;
  assign n6413 = ~n2556 & n6412 ;
  assign n6414 = n2819 & n6413 ;
  assign n6415 = n6411 | n6414 ;
  assign n6416 = n907 & ~n1028 ;
  assign n6417 = n2792 | n4344 ;
  assign n6418 = n6416 & ~n6417 ;
  assign n6419 = n2178 & ~n6418 ;
  assign n6420 = n4095 ^ n2697 ^ 1'b0 ;
  assign n6421 = n985 & ~n6420 ;
  assign n6422 = n1089 | n1113 ;
  assign n6423 = n2235 | n6422 ;
  assign n6424 = n6423 ^ n2159 ^ 1'b0 ;
  assign n6425 = n1537 & n5813 ;
  assign n6426 = n6425 ^ n530 ^ 1'b0 ;
  assign n6427 = n6426 ^ n5159 ^ n4798 ;
  assign n6428 = n6427 ^ n692 ^ 1'b0 ;
  assign n6429 = n1332 | n5129 ;
  assign n6430 = n3067 & ~n6429 ;
  assign n6431 = n4901 | n6430 ;
  assign n6432 = n6431 ^ n4451 ^ 1'b0 ;
  assign n6433 = ~n577 & n6432 ;
  assign n6434 = n2556 & n6433 ;
  assign n6435 = n6434 ^ n821 ^ 1'b0 ;
  assign n6436 = n6062 & ~n6435 ;
  assign n6437 = n2833 & ~n4972 ;
  assign n6438 = n574 & ~n6437 ;
  assign n6440 = n620 & n3764 ;
  assign n6439 = n1392 | n4024 ;
  assign n6441 = n6440 ^ n6439 ^ 1'b0 ;
  assign n6442 = n695 ^ n292 ^ 1'b0 ;
  assign n6443 = n6442 ^ n675 ^ 1'b0 ;
  assign n6444 = ~n6441 & n6443 ;
  assign n6445 = n2434 ^ n395 ^ n326 ;
  assign n6446 = n539 | n1766 ;
  assign n6447 = ~n2759 & n6446 ;
  assign n6448 = ~n1223 & n6447 ;
  assign n6449 = n6448 ^ n5674 ^ 1'b0 ;
  assign n6450 = n1645 & n1889 ;
  assign n6451 = n1021 | n2556 ;
  assign n6452 = n6451 ^ n4902 ^ 1'b0 ;
  assign n6453 = n6151 ^ n2264 ^ 1'b0 ;
  assign n6454 = n2299 & n6453 ;
  assign n6455 = ( n299 & n6440 ) | ( n299 & n6454 ) | ( n6440 & n6454 ) ;
  assign n6456 = n4705 | n6455 ;
  assign n6457 = n6456 ^ n556 ^ 1'b0 ;
  assign n6458 = n6457 ^ n2826 ^ 1'b0 ;
  assign n6459 = n4213 | n6458 ;
  assign n6460 = n3615 ^ n3476 ^ 1'b0 ;
  assign n6461 = ( n1079 & n1429 ) | ( n1079 & n5655 ) | ( n1429 & n5655 ) ;
  assign n6462 = n6460 | n6461 ;
  assign n6463 = n6462 ^ n1787 ^ 1'b0 ;
  assign n6464 = n4863 ^ n161 ^ 1'b0 ;
  assign n6467 = n3957 ^ n2455 ^ n710 ;
  assign n6465 = n959 | n1847 ;
  assign n6466 = ~n1620 & n6465 ;
  assign n6468 = n6467 ^ n6466 ^ 1'b0 ;
  assign n6469 = n2823 ^ n1691 ^ 1'b0 ;
  assign n6470 = n5840 & n6469 ;
  assign n6471 = n315 & n3895 ;
  assign n6472 = ~n559 & n6471 ;
  assign n6473 = n6472 ^ n2546 ^ n1500 ;
  assign n6477 = ~n656 & n2067 ;
  assign n6474 = n1512 | n2951 ;
  assign n6475 = n6137 & ~n6187 ;
  assign n6476 = n6474 & n6475 ;
  assign n6478 = n6477 ^ n6476 ^ n1217 ;
  assign n6479 = ( n1380 & ~n3204 ) | ( n1380 & n4125 ) | ( ~n3204 & n4125 ) ;
  assign n6480 = x20 & n1642 ;
  assign n6481 = ~n6479 & n6480 ;
  assign n6482 = n1350 & n4100 ;
  assign n6483 = n6482 ^ n152 ^ 1'b0 ;
  assign n6484 = n5324 | n6483 ;
  assign n6485 = n1457 & ~n2486 ;
  assign n6486 = n6485 ^ n3508 ^ 1'b0 ;
  assign n6487 = ~n1955 & n3287 ;
  assign n6488 = n6039 ^ n2504 ^ 1'b0 ;
  assign n6489 = n3278 | n6000 ;
  assign n6490 = n6489 ^ n5953 ^ 1'b0 ;
  assign n6491 = ( n2714 & n6488 ) | ( n2714 & n6490 ) | ( n6488 & n6490 ) ;
  assign n6492 = n3165 | n4008 ;
  assign n6493 = n6492 ^ n1972 ^ 1'b0 ;
  assign n6494 = n6493 ^ n2754 ^ 1'b0 ;
  assign n6495 = n6224 ^ n5364 ^ 1'b0 ;
  assign n6496 = n2382 & n4289 ;
  assign n6497 = ~n5684 & n6496 ;
  assign n6498 = n6497 ^ n5770 ^ 1'b0 ;
  assign n6499 = n6498 ^ n2076 ^ 1'b0 ;
  assign n6500 = n6348 & n6499 ;
  assign n6501 = ~n1838 & n3147 ;
  assign n6502 = ~n1929 & n6501 ;
  assign n6503 = n913 & n6502 ;
  assign n6504 = n6503 ^ n2248 ^ 1'b0 ;
  assign n6505 = n2307 & ~n3238 ;
  assign n6506 = ~n3636 & n6505 ;
  assign n6507 = n6506 ^ n4806 ^ 1'b0 ;
  assign n6508 = n3859 | n6507 ;
  assign n6509 = ~n5365 & n6508 ;
  assign n6510 = ~n770 & n1970 ;
  assign n6511 = n6510 ^ n677 ^ 1'b0 ;
  assign n6512 = n4950 ^ n1250 ^ x21 ;
  assign n6513 = n4662 ^ n4215 ^ n265 ;
  assign n6514 = n6512 & ~n6513 ;
  assign n6515 = n6511 & n6514 ;
  assign n6516 = ~n2327 & n5511 ;
  assign n6517 = n3438 ^ n1687 ^ 1'b0 ;
  assign n6518 = ~n6516 & n6517 ;
  assign n6519 = n311 & ~n3140 ;
  assign n6520 = n6387 & n6519 ;
  assign n6521 = ~x6 & n5813 ;
  assign n6522 = n6521 ^ n5188 ^ 1'b0 ;
  assign n6523 = ~n1293 & n1761 ;
  assign n6524 = n6523 ^ n3300 ^ 1'b0 ;
  assign n6525 = n6522 | n6524 ;
  assign n6526 = ~n2516 & n4906 ;
  assign n6527 = n5044 ^ n1329 ^ 1'b0 ;
  assign n6528 = n814 & n3629 ;
  assign n6529 = n6528 ^ n3813 ^ 1'b0 ;
  assign n6530 = n6529 ^ n4279 ^ 1'b0 ;
  assign n6531 = n5106 & ~n6530 ;
  assign n6532 = x1 & n6531 ;
  assign n6533 = n4243 ^ n1334 ^ 1'b0 ;
  assign n6534 = n6532 | n6533 ;
  assign n6535 = n3348 & ~n6534 ;
  assign n6537 = n1038 | n2619 ;
  assign n6538 = n6537 ^ n4868 ^ 1'b0 ;
  assign n6539 = n6538 ^ n3986 ^ 1'b0 ;
  assign n6536 = n2599 | n4815 ;
  assign n6540 = n6539 ^ n6536 ^ 1'b0 ;
  assign n6541 = ~n1634 & n3608 ;
  assign n6542 = ~n143 & n6541 ;
  assign n6543 = n5057 & ~n6542 ;
  assign n6544 = n6543 ^ x43 ^ 1'b0 ;
  assign n6545 = n784 & n3856 ;
  assign n6546 = n4693 ^ n2346 ^ 1'b0 ;
  assign n6547 = ~n6545 & n6546 ;
  assign n6548 = n143 & n1850 ;
  assign n6549 = n6548 ^ n1569 ^ 1'b0 ;
  assign n6550 = n294 & n2228 ;
  assign n6551 = n2924 & ~n3903 ;
  assign n6552 = n3298 | n6551 ;
  assign n6553 = n4107 | n6552 ;
  assign n6554 = n2720 & n3822 ;
  assign n6555 = ~n2533 & n6554 ;
  assign n6556 = ~n387 & n3237 ;
  assign n6557 = ~n2949 & n6556 ;
  assign n6558 = ( n4488 & ~n6555 ) | ( n4488 & n6557 ) | ( ~n6555 & n6557 ) ;
  assign n6559 = ( ~n1079 & n3883 ) | ( ~n1079 & n6558 ) | ( n3883 & n6558 ) ;
  assign n6560 = n6559 ^ n3727 ^ 1'b0 ;
  assign n6561 = n6553 & n6560 ;
  assign n6562 = n3098 & n6561 ;
  assign n6563 = n6562 ^ n4616 ^ 1'b0 ;
  assign n6564 = n4053 & ~n6474 ;
  assign n6565 = n6564 ^ n515 ^ 1'b0 ;
  assign n6566 = n5064 | n6565 ;
  assign n6576 = n1892 ^ n1805 ^ 1'b0 ;
  assign n6577 = n3314 | n6576 ;
  assign n6578 = n6109 ^ n1629 ^ 1'b0 ;
  assign n6579 = ~n6577 & n6578 ;
  assign n6572 = n1256 & ~n1281 ;
  assign n6573 = n775 & n6572 ;
  assign n6567 = x126 & n2696 ;
  assign n6568 = n5978 & n6567 ;
  assign n6569 = n1425 & n1792 ;
  assign n6570 = n6569 ^ n1353 ^ 1'b0 ;
  assign n6571 = ~n6568 & n6570 ;
  assign n6574 = n6573 ^ n6571 ^ n5499 ;
  assign n6575 = ( n983 & ~n1926 ) | ( n983 & n6574 ) | ( ~n1926 & n6574 ) ;
  assign n6580 = n6579 ^ n6575 ^ n2366 ;
  assign n6581 = n2153 & ~n3925 ;
  assign n6582 = n2914 & n6581 ;
  assign n6583 = n1801 & n2794 ;
  assign n6584 = ~n2461 & n6583 ;
  assign n6585 = n6584 ^ n1133 ^ 1'b0 ;
  assign n6586 = n983 & ~n5354 ;
  assign n6587 = n775 & ~n1469 ;
  assign n6588 = n6587 ^ n3799 ^ 1'b0 ;
  assign n6589 = ~n218 & n5198 ;
  assign n6590 = n2312 & n6589 ;
  assign n6591 = n6040 ^ n709 ^ 1'b0 ;
  assign n6592 = n1882 & n6591 ;
  assign n6593 = ~n531 & n883 ;
  assign n6594 = n6593 ^ n386 ^ 1'b0 ;
  assign n6595 = ( n2102 & n3113 ) | ( n2102 & ~n6594 ) | ( n3113 & ~n6594 ) ;
  assign n6596 = ~n2068 & n4671 ;
  assign n6597 = n6595 & ~n6596 ;
  assign n6598 = n3558 ^ n3391 ^ 1'b0 ;
  assign n6599 = n1359 & n6598 ;
  assign n6600 = ~n1021 & n4380 ;
  assign n6601 = ~n1062 & n6600 ;
  assign n6602 = n1797 | n6601 ;
  assign n6603 = n6599 & ~n6602 ;
  assign n6604 = n709 & ~n5176 ;
  assign n6605 = ~n716 & n4149 ;
  assign n6606 = ~n1851 & n4292 ;
  assign n6607 = n4618 & n5178 ;
  assign n6608 = ~n2381 & n6607 ;
  assign n6609 = n5829 ^ n4796 ^ 1'b0 ;
  assign n6610 = ~n179 & n366 ;
  assign n6611 = n6610 ^ n3021 ^ 1'b0 ;
  assign n6612 = n2066 & n2235 ;
  assign n6613 = n673 ^ n421 ^ 1'b0 ;
  assign n6614 = n2931 | n6613 ;
  assign n6615 = n3150 ^ n382 ^ 1'b0 ;
  assign n6616 = ~n1708 & n2218 ;
  assign n6617 = ( ~n468 & n2397 ) | ( ~n468 & n2733 ) | ( n2397 & n2733 ) ;
  assign n6618 = n4765 | n6617 ;
  assign n6619 = x82 | n4715 ;
  assign n6620 = x103 & n6619 ;
  assign n6621 = n2618 & ~n3107 ;
  assign n6622 = n1473 ^ n150 ^ 1'b0 ;
  assign n6623 = x108 & ~n6622 ;
  assign n6624 = n6623 ^ n3009 ^ 1'b0 ;
  assign n6625 = n5645 & ~n6624 ;
  assign n6626 = ( n826 & n1854 ) | ( n826 & n3424 ) | ( n1854 & n3424 ) ;
  assign n6628 = ~n709 & n1017 ;
  assign n6627 = n3696 & n3792 ;
  assign n6629 = n6628 ^ n6627 ^ 1'b0 ;
  assign n6630 = n6629 ^ n6237 ^ n710 ;
  assign n6631 = n2497 ^ n803 ^ 1'b0 ;
  assign n6632 = ~n657 & n6631 ;
  assign n6633 = n6632 ^ n2940 ^ 1'b0 ;
  assign n6634 = n1270 & ~n6633 ;
  assign n6637 = n208 & n3210 ;
  assign n6638 = n2978 & n6637 ;
  assign n6636 = n815 & n2821 ;
  assign n6639 = n6638 ^ n6636 ^ 1'b0 ;
  assign n6640 = n3579 ^ n1647 ^ 1'b0 ;
  assign n6641 = ( n1553 & n5330 ) | ( n1553 & ~n6640 ) | ( n5330 & ~n6640 ) ;
  assign n6642 = n6639 & ~n6641 ;
  assign n6643 = n6642 ^ x94 ^ 1'b0 ;
  assign n6635 = n1390 | n3162 ;
  assign n6644 = n6643 ^ n6635 ^ 1'b0 ;
  assign n6645 = n4233 | n6644 ;
  assign n6646 = n6645 ^ n5054 ^ 1'b0 ;
  assign n6647 = n2772 ^ n241 ^ 1'b0 ;
  assign n6648 = n3022 & n6647 ;
  assign n6649 = n1790 & ~n3279 ;
  assign n6650 = n2621 & ~n6649 ;
  assign n6651 = n1079 | n3533 ;
  assign n6652 = n3677 | n6651 ;
  assign n6653 = n6652 ^ n1973 ^ 1'b0 ;
  assign n6654 = n1084 & ~n3761 ;
  assign n6655 = ~n6653 & n6654 ;
  assign n6656 = n842 ^ n745 ^ 1'b0 ;
  assign n6657 = n208 | n6656 ;
  assign n6658 = n6612 & ~n6657 ;
  assign n6659 = n4273 ^ n947 ^ 1'b0 ;
  assign n6661 = n3955 ^ n2454 ^ 1'b0 ;
  assign n6660 = ~n2458 & n5390 ;
  assign n6662 = n6661 ^ n6660 ^ 1'b0 ;
  assign n6663 = n6662 ^ n6484 ^ 1'b0 ;
  assign n6664 = n530 & ~n615 ;
  assign n6665 = n6664 ^ n925 ^ 1'b0 ;
  assign n6666 = n6064 ^ n254 ^ 1'b0 ;
  assign n6667 = ~n6665 & n6666 ;
  assign n6668 = n622 ^ n406 ^ 1'b0 ;
  assign n6669 = n1862 & n6668 ;
  assign n6670 = n6669 ^ n2905 ^ 1'b0 ;
  assign n6671 = n2010 | n6670 ;
  assign n6672 = ~n177 & n2608 ;
  assign n6673 = n1965 & n2746 ;
  assign n6674 = n3410 & n6673 ;
  assign n6675 = n6291 ^ n2405 ^ 1'b0 ;
  assign n6676 = ~n569 & n6675 ;
  assign n6677 = ~n4398 & n6410 ;
  assign n6678 = ~n813 & n2070 ;
  assign n6679 = n2333 ^ n154 ^ 1'b0 ;
  assign n6680 = ~n490 & n6679 ;
  assign n6681 = ( n1219 & ~n6678 ) | ( n1219 & n6680 ) | ( ~n6678 & n6680 ) ;
  assign n6682 = x9 & n2180 ;
  assign n6683 = n6681 & n6682 ;
  assign n6684 = n2751 | n6683 ;
  assign n6685 = n2899 & ~n3495 ;
  assign n6686 = n6685 ^ n1722 ^ 1'b0 ;
  assign n6687 = ~n1324 & n6686 ;
  assign n6688 = n6687 ^ n680 ^ 1'b0 ;
  assign n6689 = n898 ^ n560 ^ 1'b0 ;
  assign n6690 = n3641 ^ n2034 ^ n1853 ;
  assign n6691 = ~n215 & n1987 ;
  assign n6692 = n6169 | n6691 ;
  assign n6693 = n3535 & ~n6692 ;
  assign n6694 = n3482 ^ n501 ^ 1'b0 ;
  assign n6695 = n4667 & ~n6694 ;
  assign n6696 = n133 | n215 ;
  assign n6697 = ( n988 & n1711 ) | ( n988 & ~n6696 ) | ( n1711 & ~n6696 ) ;
  assign n6698 = n6697 ^ n4488 ^ 1'b0 ;
  assign n6699 = ~n1008 & n1726 ;
  assign n6700 = ~n753 & n6699 ;
  assign n6701 = n6700 ^ n1244 ^ 1'b0 ;
  assign n6702 = n2228 & ~n6701 ;
  assign n6711 = n3748 ^ n1463 ^ 1'b0 ;
  assign n6712 = n2520 | n6711 ;
  assign n6710 = n3266 | n6691 ;
  assign n6713 = n6712 ^ n6710 ^ 1'b0 ;
  assign n6706 = n1785 | n2105 ;
  assign n6707 = n6270 | n6706 ;
  assign n6703 = n1145 & n2014 ;
  assign n6704 = n6703 ^ n519 ^ 1'b0 ;
  assign n6705 = n3504 | n6704 ;
  assign n6708 = n6707 ^ n6705 ^ 1'b0 ;
  assign n6709 = n3193 & n6708 ;
  assign n6714 = n6713 ^ n6709 ^ 1'b0 ;
  assign n6715 = n1823 & ~n3840 ;
  assign n6716 = n296 & ~n6715 ;
  assign n6717 = n6716 ^ n4451 ^ 1'b0 ;
  assign n6718 = n6040 | n6717 ;
  assign n6719 = n6718 ^ n3945 ^ 1'b0 ;
  assign n6720 = n2998 ^ n992 ^ 1'b0 ;
  assign n6721 = n6720 ^ n2378 ^ 1'b0 ;
  assign n6722 = n2188 | n3091 ;
  assign n6723 = ~n1898 & n6722 ;
  assign n6724 = ~n1788 & n6723 ;
  assign n6725 = n6724 ^ n5043 ^ 1'b0 ;
  assign n6726 = n1365 & n6157 ;
  assign n6727 = n643 & n6726 ;
  assign n6728 = n4784 ^ n437 ^ 1'b0 ;
  assign n6729 = n5693 ^ n794 ^ 1'b0 ;
  assign n6733 = n272 | n2361 ;
  assign n6730 = n1300 ^ n507 ^ 1'b0 ;
  assign n6731 = n3153 & n6730 ;
  assign n6732 = n884 & n6731 ;
  assign n6734 = n6733 ^ n6732 ^ 1'b0 ;
  assign n6735 = ~x81 & n6734 ;
  assign n6736 = n6252 ^ n3616 ^ 1'b0 ;
  assign n6737 = x47 & n6736 ;
  assign n6738 = x10 & n6608 ;
  assign n6739 = n4316 & n6738 ;
  assign n6742 = n1483 ^ n876 ^ 1'b0 ;
  assign n6740 = n403 & ~n1367 ;
  assign n6741 = ~n2921 & n6740 ;
  assign n6743 = n6742 ^ n6741 ^ 1'b0 ;
  assign n6744 = n3814 | n6743 ;
  assign n6745 = ~n1199 & n1836 ;
  assign n6746 = ~n1624 & n6745 ;
  assign n6747 = n4648 ^ n3861 ^ 1'b0 ;
  assign n6748 = n4147 ^ n709 ^ 1'b0 ;
  assign n6749 = n5860 ^ n2724 ^ 1'b0 ;
  assign n6750 = n3373 & ~n5754 ;
  assign n6751 = ~x29 & n2433 ;
  assign n6752 = ~n4233 & n6751 ;
  assign n6753 = n6752 ^ n855 ^ 1'b0 ;
  assign n6754 = n3241 & n6753 ;
  assign n6755 = ( ~n6749 & n6750 ) | ( ~n6749 & n6754 ) | ( n6750 & n6754 ) ;
  assign n6756 = x0 & n1592 ;
  assign n6757 = n6756 ^ n5728 ^ n959 ;
  assign n6758 = n1201 & ~n4671 ;
  assign n6759 = n3975 ^ n330 ^ 1'b0 ;
  assign n6760 = ( n1334 & n2639 ) | ( n1334 & ~n6759 ) | ( n2639 & ~n6759 ) ;
  assign n6764 = n3601 & ~n4560 ;
  assign n6765 = n338 | n6764 ;
  assign n6766 = n5962 & ~n6765 ;
  assign n6767 = n1955 | n3858 ;
  assign n6768 = n6766 & ~n6767 ;
  assign n6769 = n6768 ^ n977 ^ 1'b0 ;
  assign n6770 = n5356 & n6769 ;
  assign n6761 = n1683 & ~n1770 ;
  assign n6762 = n6761 ^ n903 ^ 1'b0 ;
  assign n6763 = n6762 ^ n559 ^ 1'b0 ;
  assign n6771 = n6770 ^ n6763 ^ 1'b0 ;
  assign n6773 = ~n326 & n517 ;
  assign n6774 = n3574 & ~n6773 ;
  assign n6775 = n1479 & n6774 ;
  assign n6772 = n2644 | n6372 ;
  assign n6776 = n6775 ^ n6772 ^ 1'b0 ;
  assign n6779 = ~n489 & n791 ;
  assign n6780 = n6779 ^ n1426 ^ 1'b0 ;
  assign n6781 = n4190 | n6780 ;
  assign n6782 = n6781 ^ n374 ^ 1'b0 ;
  assign n6783 = n2312 | n6782 ;
  assign n6777 = n3404 ^ n2882 ^ 1'b0 ;
  assign n6778 = n489 & ~n6777 ;
  assign n6784 = n6783 ^ n6778 ^ n3834 ;
  assign n6785 = n742 | n2424 ;
  assign n6786 = n2874 & n5676 ;
  assign n6787 = ~n6785 & n6786 ;
  assign n6788 = ~n1484 & n4069 ;
  assign n6789 = ~n3098 & n6788 ;
  assign n6790 = n2221 ^ n266 ^ 1'b0 ;
  assign n6791 = n6254 | n6790 ;
  assign n6792 = n4408 ^ x49 ^ 1'b0 ;
  assign n6793 = n6792 ^ n3076 ^ 1'b0 ;
  assign n6794 = n3724 | n5209 ;
  assign n6795 = n999 | n1562 ;
  assign n6796 = n6795 ^ n5791 ^ 1'b0 ;
  assign n6797 = n6757 ^ n3150 ^ 1'b0 ;
  assign n6799 = n1162 ^ n317 ^ 1'b0 ;
  assign n6798 = n949 & n3683 ;
  assign n6800 = n6799 ^ n6798 ^ 1'b0 ;
  assign n6801 = ~n2010 & n6629 ;
  assign n6802 = n5138 & n6043 ;
  assign n6803 = n601 | n852 ;
  assign n6804 = n3482 & ~n6803 ;
  assign n6805 = ( n1624 & ~n2834 ) | ( n1624 & n3215 ) | ( ~n2834 & n3215 ) ;
  assign n6806 = ~n593 & n3249 ;
  assign n6807 = ~n1308 & n6806 ;
  assign n6808 = n1142 & ~n6807 ;
  assign n6809 = n344 & n6808 ;
  assign n6810 = ~n4408 & n4597 ;
  assign n6811 = ~n301 & n6810 ;
  assign n6812 = n5508 | n6811 ;
  assign n6813 = n6812 ^ n628 ^ 1'b0 ;
  assign n6814 = ( n1847 & n4875 ) | ( n1847 & ~n6610 ) | ( n4875 & ~n6610 ) ;
  assign n6815 = n6814 ^ n1250 ^ 1'b0 ;
  assign n6816 = ~n1410 & n5064 ;
  assign n6817 = ~n4575 & n6816 ;
  assign n6818 = n3717 | n6817 ;
  assign n6819 = n5550 ^ n5429 ^ 1'b0 ;
  assign n6820 = n1109 | n6819 ;
  assign n6821 = n2605 & ~n6820 ;
  assign n6822 = n1761 | n6470 ;
  assign n6823 = n6821 & ~n6822 ;
  assign n6824 = n722 & n1558 ;
  assign n6825 = ~x123 & n6824 ;
  assign n6826 = n6825 ^ n3226 ^ 1'b0 ;
  assign n6827 = ~n3601 & n6826 ;
  assign n6828 = n3302 | n5479 ;
  assign n6831 = n4098 & n5625 ;
  assign n6832 = n6831 ^ n1600 ^ 1'b0 ;
  assign n6829 = n1467 | n4001 ;
  assign n6830 = n3758 & n6829 ;
  assign n6833 = n6832 ^ n6830 ^ 1'b0 ;
  assign n6834 = n3738 ^ n3064 ^ 1'b0 ;
  assign n6835 = ~n1588 & n5022 ;
  assign n6836 = ( ~n978 & n3587 ) | ( ~n978 & n3682 ) | ( n3587 & n3682 ) ;
  assign n6837 = n1581 ^ n369 ^ 1'b0 ;
  assign n6838 = n2874 & n6837 ;
  assign n6839 = n6612 & n6838 ;
  assign n6840 = n2421 | n3772 ;
  assign n6841 = n3369 & ~n5652 ;
  assign n6842 = n1325 & n6841 ;
  assign n6843 = n3411 & n6842 ;
  assign n6844 = n3393 | n6843 ;
  assign n6845 = ~n3234 & n6844 ;
  assign n6846 = n6845 ^ n138 ^ 1'b0 ;
  assign n6847 = n2075 | n6846 ;
  assign n6848 = n6847 ^ n557 ^ 1'b0 ;
  assign n6849 = n1327 ^ n851 ^ 1'b0 ;
  assign n6850 = n3629 & n6849 ;
  assign n6851 = n6850 ^ n3230 ^ 1'b0 ;
  assign n6852 = n1720 & ~n6851 ;
  assign n6853 = n4143 & n4315 ;
  assign n6854 = ~n6852 & n6853 ;
  assign n6855 = n5973 ^ n188 ^ 1'b0 ;
  assign n6856 = ~n6086 & n6855 ;
  assign n6857 = n3637 & n6856 ;
  assign n6858 = n3603 ^ n2214 ^ n1095 ;
  assign n6859 = n1438 | n5804 ;
  assign n6860 = n6858 & ~n6859 ;
  assign n6861 = ( n480 & n559 ) | ( n480 & n5298 ) | ( n559 & n5298 ) ;
  assign n6862 = n1939 & n2551 ;
  assign n6863 = n4145 & n6862 ;
  assign n6864 = ~n459 & n2490 ;
  assign n6865 = n6864 ^ n1424 ^ 1'b0 ;
  assign n6866 = n6865 ^ n2014 ^ 1'b0 ;
  assign n6867 = n6863 & ~n6866 ;
  assign n6868 = n4436 ^ n2976 ^ 1'b0 ;
  assign n6869 = ~n4087 & n6868 ;
  assign n6870 = ~n1933 & n5981 ;
  assign n6871 = n6870 ^ n813 ^ 1'b0 ;
  assign n6872 = n1281 | n6432 ;
  assign n6873 = n3533 ^ n1672 ^ 1'b0 ;
  assign n6874 = ~n1545 & n5431 ;
  assign n6875 = n6874 ^ n4809 ^ 1'b0 ;
  assign n6876 = n6875 ^ n3982 ^ 1'b0 ;
  assign n6881 = n971 | n3691 ;
  assign n6882 = n5281 | n6881 ;
  assign n6877 = n1737 ^ n1250 ^ n256 ;
  assign n6878 = n6877 ^ n2394 ^ 1'b0 ;
  assign n6879 = n2399 | n6878 ;
  assign n6880 = n3236 | n6879 ;
  assign n6883 = n6882 ^ n6880 ^ 1'b0 ;
  assign n6885 = n5908 ^ n2290 ^ 1'b0 ;
  assign n6884 = ~n3512 & n4172 ;
  assign n6886 = n6885 ^ n6884 ^ 1'b0 ;
  assign n6887 = x113 & ~n754 ;
  assign n6888 = n6887 ^ x24 ^ 1'b0 ;
  assign n6889 = ~n943 & n2389 ;
  assign n6890 = n4355 ^ n1217 ^ 1'b0 ;
  assign n6891 = ~n4606 & n6890 ;
  assign n6892 = n6891 ^ n538 ^ 1'b0 ;
  assign n6893 = n4981 & n6892 ;
  assign n6894 = n4827 & n6893 ;
  assign n6895 = ~n3699 & n6894 ;
  assign n6896 = ~n6889 & n6895 ;
  assign n6897 = n5167 ^ n3083 ^ 1'b0 ;
  assign n6898 = n2298 & ~n6897 ;
  assign n6899 = n6166 ^ n1932 ^ n595 ;
  assign n6900 = n6676 ^ n3146 ^ 1'b0 ;
  assign n6904 = n1221 & n4186 ;
  assign n6901 = ~n1374 & n1672 ;
  assign n6902 = ~n1396 & n4215 ;
  assign n6903 = ~n6901 & n6902 ;
  assign n6905 = n6904 ^ n6903 ^ 1'b0 ;
  assign n6906 = n3257 | n6368 ;
  assign n6907 = n1487 | n6906 ;
  assign n6908 = n6907 ^ n2319 ^ 1'b0 ;
  assign n6909 = n4724 | n6908 ;
  assign n6910 = n215 & n321 ;
  assign n6911 = n1124 & n5092 ;
  assign n6912 = n6910 | n6911 ;
  assign n6913 = n4380 | n6912 ;
  assign n6914 = n533 & ~n6392 ;
  assign n6915 = n208 & n1354 ;
  assign n6916 = n6915 ^ n1223 ^ 1'b0 ;
  assign n6917 = n4530 & ~n5285 ;
  assign n6918 = ~n3119 & n6821 ;
  assign n6919 = n6918 ^ n832 ^ 1'b0 ;
  assign n6920 = n6917 & ~n6919 ;
  assign n6921 = n6920 ^ n4405 ^ 1'b0 ;
  assign n6922 = n4125 & ~n5672 ;
  assign n6923 = n2798 | n4614 ;
  assign n6924 = n1150 | n2724 ;
  assign n6925 = n1895 | n2878 ;
  assign n6926 = n6925 ^ n4551 ^ 1'b0 ;
  assign n6927 = n261 & ~n4950 ;
  assign n6928 = n6927 ^ n4564 ^ 1'b0 ;
  assign n6929 = n810 ^ x5 ^ 1'b0 ;
  assign n6930 = n2802 & n4575 ;
  assign n6931 = n6929 & n6930 ;
  assign n6932 = n6931 ^ n3365 ^ 1'b0 ;
  assign n6933 = n6932 ^ n6550 ^ 1'b0 ;
  assign n6934 = n784 & ~n5513 ;
  assign n6935 = n2919 ^ n1011 ^ 1'b0 ;
  assign n6936 = n1232 & ~n6935 ;
  assign n6937 = n1888 & n6384 ;
  assign n6938 = ~n5093 & n6937 ;
  assign n6939 = n1143 & n1211 ;
  assign n6940 = ~x103 & n6939 ;
  assign n6941 = n915 & ~n929 ;
  assign n6942 = n5373 ^ n4091 ^ 1'b0 ;
  assign n6943 = ~n2426 & n6942 ;
  assign n6944 = n4605 & ~n6943 ;
  assign n6948 = n2915 & ~n5571 ;
  assign n6945 = n1136 ^ x107 ^ 1'b0 ;
  assign n6946 = n3998 & ~n6945 ;
  assign n6947 = ~n1668 & n6946 ;
  assign n6949 = n6948 ^ n6947 ^ 1'b0 ;
  assign n6950 = n2365 & n3004 ;
  assign n6951 = n3574 & n6950 ;
  assign n6952 = n2050 ^ n760 ^ 1'b0 ;
  assign n6953 = n583 & n6952 ;
  assign n6954 = ( n1867 & ~n6029 ) | ( n1867 & n6953 ) | ( ~n6029 & n6953 ) ;
  assign n6955 = n3982 ^ n3533 ^ 1'b0 ;
  assign n6956 = n2384 & ~n6955 ;
  assign n6957 = ( ~n3310 & n3706 ) | ( ~n3310 & n4104 ) | ( n3706 & n4104 ) ;
  assign n6958 = n6957 ^ n1217 ^ 1'b0 ;
  assign n6959 = n3153 & n6958 ;
  assign n6960 = n3825 & n6959 ;
  assign n6961 = n3844 & n6960 ;
  assign n6962 = n2336 | n4547 ;
  assign n6963 = n283 & ~n6962 ;
  assign n6964 = x56 & ~n4046 ;
  assign n6965 = n4912 & n6212 ;
  assign n6966 = n5976 ^ n2949 ^ 1'b0 ;
  assign n6967 = n2286 ^ n1967 ^ 1'b0 ;
  assign n6968 = n4729 | n6967 ;
  assign n6969 = n3249 | n6968 ;
  assign n6970 = n3542 ^ n1147 ^ 1'b0 ;
  assign n6971 = n2458 ^ n344 ^ 1'b0 ;
  assign n6972 = n4411 ^ n1578 ^ 1'b0 ;
  assign n6973 = n1912 ^ n827 ^ 1'b0 ;
  assign n6974 = n5345 ^ n971 ^ n559 ;
  assign n6975 = n2450 | n5593 ;
  assign n6976 = n1277 & ~n2024 ;
  assign n6977 = n6976 ^ n3537 ^ 1'b0 ;
  assign n6978 = n1102 ^ x122 ^ 1'b0 ;
  assign n6979 = ~n1247 & n6978 ;
  assign n6980 = n1695 | n1708 ;
  assign n6981 = n6980 ^ n321 ^ 1'b0 ;
  assign n6982 = n6981 ^ n433 ^ 1'b0 ;
  assign n6983 = n6982 ^ n5618 ^ 1'b0 ;
  assign n6984 = n6861 & n6983 ;
  assign n6985 = n5616 ^ n3139 ^ 1'b0 ;
  assign n6986 = ~n2308 & n6531 ;
  assign n6987 = n6986 ^ n3083 ^ 1'b0 ;
  assign n6988 = ~n4187 & n6987 ;
  assign n6989 = n5004 ^ n2835 ^ 1'b0 ;
  assign n6990 = n437 & n1681 ;
  assign n6991 = ( ~n225 & n533 ) | ( ~n225 & n6990 ) | ( n533 & n6990 ) ;
  assign n6992 = n3884 | n3949 ;
  assign n6993 = n6991 & n6992 ;
  assign n6994 = n6993 ^ n2689 ^ 1'b0 ;
  assign n6995 = n3441 | n4305 ;
  assign n6996 = x110 & n3269 ;
  assign n6997 = n533 & ~n2126 ;
  assign n6998 = n901 & ~n4638 ;
  assign n6999 = ( n609 & n1586 ) | ( n609 & ~n4413 ) | ( n1586 & ~n4413 ) ;
  assign n7000 = n6999 ^ n6628 ^ 1'b0 ;
  assign n7001 = n2402 & n5948 ;
  assign n7002 = n4899 ^ n1433 ^ 1'b0 ;
  assign n7003 = n949 & n3546 ;
  assign n7004 = n2310 & n7003 ;
  assign n7005 = n3266 ^ n2468 ^ 1'b0 ;
  assign n7006 = n7004 | n7005 ;
  assign n7007 = ( ~n1672 & n4960 ) | ( ~n1672 & n6080 ) | ( n4960 & n6080 ) ;
  assign n7008 = x49 & ~x67 ;
  assign n7009 = n651 | n6259 ;
  assign n7010 = n2435 | n7009 ;
  assign n7011 = n5422 ^ n2435 ^ 1'b0 ;
  assign n7012 = n3272 ^ n2013 ^ n1491 ;
  assign n7013 = n5371 & ~n7012 ;
  assign n7014 = n7013 ^ n6259 ^ 1'b0 ;
  assign n7015 = n934 & n7014 ;
  assign n7016 = ~n4391 & n7015 ;
  assign n7020 = n708 & ~n3846 ;
  assign n7021 = n7020 ^ n4084 ^ 1'b0 ;
  assign n7017 = n1217 ^ n884 ^ 1'b0 ;
  assign n7018 = ~n357 & n7017 ;
  assign n7019 = n726 | n7018 ;
  assign n7022 = n7021 ^ n7019 ^ n4753 ;
  assign n7023 = n1804 & ~n7022 ;
  assign n7024 = n2780 & n7023 ;
  assign n7025 = n3334 & n6733 ;
  assign n7026 = n7025 ^ n2494 ^ n613 ;
  assign n7027 = n1437 ^ n611 ^ 1'b0 ;
  assign n7028 = ~n7026 & n7027 ;
  assign n7029 = n4212 ^ n885 ^ 1'b0 ;
  assign n7030 = n1899 & n7029 ;
  assign n7031 = ~n541 & n3076 ;
  assign n7032 = n6862 & n6929 ;
  assign n7033 = n4597 & n7032 ;
  assign n7034 = n3899 ^ n1311 ^ 1'b0 ;
  assign n7035 = n3316 & ~n7034 ;
  assign n7036 = n7033 & n7035 ;
  assign n7037 = n3704 & n7036 ;
  assign n7038 = ( n157 & ~n3404 ) | ( n157 & n3757 ) | ( ~n3404 & n3757 ) ;
  assign n7039 = ~n3681 & n6742 ;
  assign n7040 = n935 & ~n4832 ;
  assign n7041 = n6004 ^ n4304 ^ 1'b0 ;
  assign n7042 = n1038 & ~n1056 ;
  assign n7043 = n7042 ^ n2953 ^ 1'b0 ;
  assign n7044 = n6055 ^ n2395 ^ 1'b0 ;
  assign n7045 = ~n5701 & n7044 ;
  assign n7046 = ~n3460 & n7045 ;
  assign n7047 = ~n7043 & n7046 ;
  assign n7048 = n2733 & ~n5726 ;
  assign n7049 = n1649 & n5631 ;
  assign n7050 = n7049 ^ n1616 ^ 1'b0 ;
  assign n7051 = n3488 ^ n299 ^ 1'b0 ;
  assign n7052 = n355 & ~n695 ;
  assign n7053 = n2561 & n7052 ;
  assign n7054 = n7053 ^ n2886 ^ 1'b0 ;
  assign n7055 = ( n1250 & n1549 ) | ( n1250 & ~n1732 ) | ( n1549 & ~n1732 ) ;
  assign n7056 = n3908 ^ n1836 ^ 1'b0 ;
  assign n7057 = n7055 & n7056 ;
  assign n7058 = ~n3846 & n3998 ;
  assign n7059 = n3846 & n7058 ;
  assign n7060 = n7059 ^ n3056 ^ 1'b0 ;
  assign n7061 = n427 & n763 ;
  assign n7062 = ~n763 & n7061 ;
  assign n7063 = n438 & n2983 ;
  assign n7064 = n7062 & n7063 ;
  assign n7065 = n7064 ^ n4472 ^ 1'b0 ;
  assign n7066 = n7060 | n7065 ;
  assign n7067 = n1166 | n4549 ;
  assign n7068 = n7067 ^ n3910 ^ 1'b0 ;
  assign n7069 = n1805 | n3248 ;
  assign n7070 = n4467 | n7069 ;
  assign n7071 = n7070 ^ n718 ^ n157 ;
  assign n7079 = n1723 | n3365 ;
  assign n7072 = n1479 | n2877 ;
  assign n7073 = n1044 & n1758 ;
  assign n7074 = n7072 & n7073 ;
  assign n7075 = n7074 ^ n5052 ^ 1'b0 ;
  assign n7076 = ~n928 & n7075 ;
  assign n7077 = n2150 & n4112 ;
  assign n7078 = n7076 & ~n7077 ;
  assign n7080 = n7079 ^ n7078 ^ 1'b0 ;
  assign n7082 = n444 | n1581 ;
  assign n7083 = n7082 ^ n1229 ^ 1'b0 ;
  assign n7084 = n7083 ^ n1253 ^ 1'b0 ;
  assign n7085 = x23 & ~n7084 ;
  assign n7081 = n1705 | n5804 ;
  assign n7086 = n7085 ^ n7081 ^ 1'b0 ;
  assign n7089 = n412 & n3386 ;
  assign n7090 = n7089 ^ n4250 ^ 1'b0 ;
  assign n7091 = n1285 | n7090 ;
  assign n7087 = n4359 ^ n1990 ^ 1'b0 ;
  assign n7088 = ~n2315 & n7087 ;
  assign n7092 = n7091 ^ n7088 ^ 1'b0 ;
  assign n7093 = ~n4616 & n7092 ;
  assign n7094 = n2010 | n3062 ;
  assign n7095 = n7094 ^ n556 ^ 1'b0 ;
  assign n7096 = n6871 & n7095 ;
  assign n7097 = n6680 ^ n1346 ^ 1'b0 ;
  assign n7098 = n7097 ^ n234 ^ 1'b0 ;
  assign n7099 = n6771 & n7098 ;
  assign n7100 = ( ~n278 & n897 ) | ( ~n278 & n6366 ) | ( n897 & n6366 ) ;
  assign n7101 = n920 & ~n2318 ;
  assign n7102 = n2128 ^ x75 ^ 1'b0 ;
  assign n7103 = n5332 ^ n3391 ^ 1'b0 ;
  assign n7104 = n7103 ^ n3486 ^ 1'b0 ;
  assign n7105 = x20 & n7104 ;
  assign n7106 = ( x20 & n1413 ) | ( x20 & ~n1847 ) | ( n1413 & ~n1847 ) ;
  assign n7107 = n1563 & n7106 ;
  assign n7108 = n7107 ^ n1228 ^ 1'b0 ;
  assign n7109 = n2543 ^ n920 ^ 1'b0 ;
  assign n7110 = ~n1019 & n7109 ;
  assign n7111 = n7110 ^ n5826 ^ n3982 ;
  assign n7112 = n7111 ^ n4702 ^ n2837 ;
  assign n7113 = n2172 ^ n258 ^ 1'b0 ;
  assign n7114 = n2694 | n7113 ;
  assign n7115 = n545 | n6599 ;
  assign n7116 = n2946 | n7115 ;
  assign n7117 = n3041 ^ n1270 ^ 1'b0 ;
  assign n7118 = n551 | n7117 ;
  assign n7119 = n1867 ^ x49 ^ 1'b0 ;
  assign n7120 = n5131 ^ n2760 ^ 1'b0 ;
  assign n7121 = n6062 ^ n3515 ^ 1'b0 ;
  assign n7122 = x57 & n3856 ;
  assign n7123 = n3328 | n7122 ;
  assign n7124 = n1612 | n7123 ;
  assign n7125 = n2021 ^ n1385 ^ 1'b0 ;
  assign n7126 = n3156 & ~n7125 ;
  assign n7127 = n227 & ~n7126 ;
  assign n7128 = ~n2629 & n7127 ;
  assign n7129 = n883 & ~n7128 ;
  assign n7130 = n7124 & n7129 ;
  assign n7131 = n5713 & ~n7130 ;
  assign n7132 = n832 & ~n1611 ;
  assign n7133 = n2268 & n7132 ;
  assign n7134 = ( n411 & n6308 ) | ( n411 & ~n7133 ) | ( n6308 & ~n7133 ) ;
  assign n7135 = n2915 ^ n344 ^ 1'b0 ;
  assign n7136 = n3131 & ~n7135 ;
  assign n7137 = ~n6211 & n7136 ;
  assign n7140 = n771 & n901 ;
  assign n7141 = n861 & n7140 ;
  assign n7138 = n3238 ^ n759 ^ 1'b0 ;
  assign n7139 = n7138 ^ n1890 ^ 1'b0 ;
  assign n7142 = n7141 ^ n7139 ^ 1'b0 ;
  assign n7143 = n7137 & n7142 ;
  assign n7144 = n4420 ^ x67 ^ 1'b0 ;
  assign n7145 = n1285 & n7144 ;
  assign n7146 = n7145 ^ n1877 ^ 1'b0 ;
  assign n7147 = n2564 ^ n1596 ^ 1'b0 ;
  assign n7148 = n7146 | n7147 ;
  assign n7149 = n1703 ^ n241 ^ 1'b0 ;
  assign n7150 = n627 & ~n7149 ;
  assign n7153 = n3481 ^ n674 ^ 1'b0 ;
  assign n7154 = n1871 & n7153 ;
  assign n7152 = n1357 & ~n2010 ;
  assign n7155 = n7154 ^ n7152 ^ 1'b0 ;
  assign n7151 = ~n745 & n1939 ;
  assign n7156 = n7155 ^ n7151 ^ 1'b0 ;
  assign n7157 = ( n1596 & n1819 ) | ( n1596 & ~n4528 ) | ( n1819 & ~n4528 ) ;
  assign n7158 = n5415 | n7157 ;
  assign n7159 = n3514 ^ n2865 ^ 1'b0 ;
  assign n7160 = n1714 | n7159 ;
  assign n7161 = n4527 & ~n7160 ;
  assign n7162 = n3717 & n3974 ;
  assign n7163 = n7162 ^ n5593 ^ 1'b0 ;
  assign n7164 = ~n861 & n3606 ;
  assign n7165 = n7164 ^ n1849 ^ 1'b0 ;
  assign n7166 = n7163 | n7165 ;
  assign n7167 = n2021 & ~n7166 ;
  assign n7169 = n3368 & ~n4905 ;
  assign n7170 = n7169 ^ n4589 ^ 1'b0 ;
  assign n7168 = n931 | n4022 ;
  assign n7171 = n7170 ^ n7168 ^ 1'b0 ;
  assign n7172 = x26 & n900 ;
  assign n7173 = ~n144 & n7172 ;
  assign n7174 = n7173 ^ n6515 ^ 1'b0 ;
  assign n7175 = n6542 | n7174 ;
  assign n7176 = n6634 & ~n7175 ;
  assign n7177 = n7176 ^ x24 ^ 1'b0 ;
  assign n7178 = ( n1008 & n2322 ) | ( n1008 & ~n2821 ) | ( n2322 & ~n2821 ) ;
  assign n7180 = n2286 & ~n3641 ;
  assign n7181 = ~n1529 & n7180 ;
  assign n7182 = n5352 & n7181 ;
  assign n7179 = ~n728 & n5953 ;
  assign n7183 = n7182 ^ n7179 ^ 1'b0 ;
  assign n7184 = n5092 ^ n2790 ^ 1'b0 ;
  assign n7185 = n7183 & ~n7184 ;
  assign n7187 = ~n549 & n675 ;
  assign n7188 = n3590 & ~n7187 ;
  assign n7186 = n2107 & n5302 ;
  assign n7189 = n7188 ^ n7186 ^ 1'b0 ;
  assign n7190 = ( ~n1759 & n5911 ) | ( ~n1759 & n6019 ) | ( n5911 & n6019 ) ;
  assign n7191 = n5801 ^ n1484 ^ 1'b0 ;
  assign n7192 = n2513 & ~n2583 ;
  assign n7193 = n1487 & ~n3527 ;
  assign n7194 = n7193 ^ n5315 ^ 1'b0 ;
  assign n7195 = n3960 & n7165 ;
  assign n7196 = n182 & n3465 ;
  assign n7197 = ~n5336 & n5394 ;
  assign n7198 = n7197 ^ n4875 ^ 1'b0 ;
  assign n7203 = n324 & ~n1077 ;
  assign n7199 = n2103 & n3806 ;
  assign n7200 = n949 & n1878 ;
  assign n7201 = n7200 ^ n3217 ^ 1'b0 ;
  assign n7202 = ~n7199 & n7201 ;
  assign n7204 = n7203 ^ n7202 ^ 1'b0 ;
  assign n7205 = n2496 & n5461 ;
  assign n7206 = ~n2131 & n4531 ;
  assign n7207 = n252 | n3988 ;
  assign n7208 = n3575 ^ n1811 ^ 1'b0 ;
  assign n7210 = n1911 & n2474 ;
  assign n7211 = n3308 & ~n6879 ;
  assign n7212 = ~n874 & n7211 ;
  assign n7213 = ~n7210 & n7212 ;
  assign n7209 = n4527 ^ n2553 ^ n2454 ;
  assign n7214 = n7213 ^ n7209 ^ 1'b0 ;
  assign n7215 = ~n7208 & n7214 ;
  assign n7216 = ~n3615 & n7215 ;
  assign n7217 = ( n400 & n1831 ) | ( n400 & n5375 ) | ( n1831 & n5375 ) ;
  assign n7218 = ( n4755 & n4784 ) | ( n4755 & n7217 ) | ( n4784 & n7217 ) ;
  assign n7219 = n3198 ^ n2293 ^ n1263 ;
  assign n7220 = n4682 & ~n7219 ;
  assign n7224 = ~n1235 & n2613 ;
  assign n7225 = n7224 ^ n2508 ^ 1'b0 ;
  assign n7221 = ~n645 & n1369 ;
  assign n7222 = n2611 | n7221 ;
  assign n7223 = ~n1079 & n7222 ;
  assign n7226 = n7225 ^ n7223 ^ 1'b0 ;
  assign n7227 = x6 | n587 ;
  assign n7228 = n7227 ^ n1978 ^ 1'b0 ;
  assign n7229 = n7228 ^ n1419 ^ 1'b0 ;
  assign n7230 = n3154 ^ n1252 ^ 1'b0 ;
  assign n7231 = n445 ^ n224 ^ 1'b0 ;
  assign n7232 = n7231 ^ n152 ^ 1'b0 ;
  assign n7233 = n4814 & n7232 ;
  assign n7234 = n4039 ^ n3827 ^ 1'b0 ;
  assign n7235 = n7234 ^ n6002 ^ 1'b0 ;
  assign n7236 = n556 & n2055 ;
  assign n7237 = n580 & n3136 ;
  assign n7238 = n4471 & n7237 ;
  assign n7239 = ( ~n3816 & n4467 ) | ( ~n3816 & n7238 ) | ( n4467 & n7238 ) ;
  assign n7240 = n1348 | n3903 ;
  assign n7241 = n6159 & ~n7240 ;
  assign n7242 = n5533 & n7241 ;
  assign n7243 = ~n1469 & n2853 ;
  assign n7244 = n625 & n2660 ;
  assign n7245 = n4755 | n6634 ;
  assign n7246 = n2091 & ~n4204 ;
  assign n7247 = ~n5052 & n7246 ;
  assign n7248 = n6529 ^ n3469 ^ 1'b0 ;
  assign n7249 = n229 & ~n2414 ;
  assign n7250 = n542 & n2585 ;
  assign n7251 = n279 & n7250 ;
  assign n7252 = ~n954 & n7251 ;
  assign n7253 = n7249 & ~n7252 ;
  assign n7254 = ~n656 & n3924 ;
  assign n7255 = n7254 ^ n5074 ^ 1'b0 ;
  assign n7256 = n1723 ^ n1615 ^ 1'b0 ;
  assign n7257 = n1898 & n7256 ;
  assign n7258 = n7257 ^ n4269 ^ 1'b0 ;
  assign n7259 = n628 ^ x65 ^ 1'b0 ;
  assign n7260 = ( n1231 & n7258 ) | ( n1231 & n7259 ) | ( n7258 & n7259 ) ;
  assign n7261 = n2111 | n5264 ;
  assign n7262 = n1123 | n7261 ;
  assign n7263 = n7262 ^ n2380 ^ 1'b0 ;
  assign n7266 = ~n679 & n6467 ;
  assign n7267 = n7266 ^ n1890 ^ 1'b0 ;
  assign n7264 = ~n2220 & n3308 ;
  assign n7265 = ~n3542 & n7264 ;
  assign n7268 = n7267 ^ n7265 ^ 1'b0 ;
  assign n7269 = ~n1540 & n1625 ;
  assign n7270 = ~n2222 & n7269 ;
  assign n7271 = n2967 ^ n204 ^ 1'b0 ;
  assign n7272 = n7270 | n7271 ;
  assign n7273 = ( ~n5308 & n7268 ) | ( ~n5308 & n7272 ) | ( n7268 & n7272 ) ;
  assign n7274 = n3179 & n6653 ;
  assign n7275 = n7274 ^ n1880 ^ 1'b0 ;
  assign n7276 = n1635 ^ n1211 ^ 1'b0 ;
  assign n7277 = n1182 & n7276 ;
  assign n7278 = x107 & ~n1933 ;
  assign n7279 = n7278 ^ n1747 ^ 1'b0 ;
  assign n7280 = ~n7277 & n7279 ;
  assign n7281 = ~n3419 & n7280 ;
  assign n7282 = n7281 ^ n4112 ^ 1'b0 ;
  assign n7283 = x36 & ~n260 ;
  assign n7284 = n7283 ^ n7137 ^ 1'b0 ;
  assign n7285 = ( ~n4065 & n5178 ) | ( ~n4065 & n5517 ) | ( n5178 & n5517 ) ;
  assign n7286 = n5783 ^ n2095 ^ 1'b0 ;
  assign n7287 = ~n3214 & n7286 ;
  assign n7288 = n3335 & n7287 ;
  assign n7289 = n6720 ^ n3543 ^ x27 ;
  assign n7290 = ~n5551 & n7289 ;
  assign n7291 = n7288 & n7290 ;
  assign n7292 = n7291 ^ n1408 ^ 1'b0 ;
  assign n7293 = ~n2804 & n7292 ;
  assign n7294 = n4359 ^ n601 ^ 1'b0 ;
  assign n7295 = n7293 & ~n7294 ;
  assign n7296 = ~n1973 & n4171 ;
  assign n7297 = n7296 ^ n4737 ^ 1'b0 ;
  assign n7298 = n5321 & ~n5870 ;
  assign n7299 = n5826 ^ n4064 ^ n417 ;
  assign n7303 = n3669 ^ n1562 ^ 1'b0 ;
  assign n7304 = n5776 & ~n7303 ;
  assign n7305 = n7304 ^ x31 ^ 1'b0 ;
  assign n7300 = x69 & ~n1507 ;
  assign n7301 = n7300 ^ n636 ^ 1'b0 ;
  assign n7302 = n2504 & n7301 ;
  assign n7306 = n7305 ^ n7302 ^ 1'b0 ;
  assign n7307 = n7306 ^ n1925 ^ 1'b0 ;
  assign n7308 = n565 & n708 ;
  assign n7309 = n7308 ^ n2164 ^ 1'b0 ;
  assign n7310 = n993 & n7309 ;
  assign n7311 = ( n1296 & n3073 ) | ( n1296 & ~n7310 ) | ( n3073 & ~n7310 ) ;
  assign n7312 = n7311 ^ n2587 ^ 1'b0 ;
  assign n7313 = n4766 & n7312 ;
  assign n7314 = n6147 ^ n4182 ^ 1'b0 ;
  assign n7315 = ~n2814 & n7314 ;
  assign n7316 = x47 & n4809 ;
  assign n7317 = ~n1932 & n3603 ;
  assign n7318 = n646 & n7317 ;
  assign n7319 = ~n531 & n7318 ;
  assign n7320 = n7319 ^ n5850 ^ 1'b0 ;
  assign n7321 = x47 | n4793 ;
  assign n7322 = ~n5618 & n7321 ;
  assign n7323 = ~n1116 & n6667 ;
  assign n7324 = n7323 ^ n5887 ^ 1'b0 ;
  assign n7325 = n5026 & n7324 ;
  assign n7326 = n1853 & ~n6519 ;
  assign n7327 = n983 ^ n175 ^ 1'b0 ;
  assign n7328 = n4979 & ~n7327 ;
  assign n7329 = ~n2357 & n6000 ;
  assign n7330 = ( n5539 & ~n6763 ) | ( n5539 & n7329 ) | ( ~n6763 & n7329 ) ;
  assign n7331 = n6557 ^ n3327 ^ 1'b0 ;
  assign n7332 = n296 & ~n1097 ;
  assign n7333 = n1398 | n7332 ;
  assign n7336 = n480 | n1250 ;
  assign n7335 = n1813 & n5836 ;
  assign n7337 = n7336 ^ n7335 ^ 1'b0 ;
  assign n7334 = n1264 & ~n5978 ;
  assign n7338 = n7337 ^ n7334 ^ 1'b0 ;
  assign n7339 = n3511 ^ n983 ^ 1'b0 ;
  assign n7340 = n2504 ^ n1420 ^ 1'b0 ;
  assign n7341 = n1844 & ~n7340 ;
  assign n7342 = n4068 & ~n6135 ;
  assign n7343 = n7342 ^ n3677 ^ 1'b0 ;
  assign n7344 = n7343 ^ n4354 ^ 1'b0 ;
  assign n7345 = n5962 ^ n3289 ^ 1'b0 ;
  assign n7346 = n7345 ^ n5650 ^ 1'b0 ;
  assign n7347 = n956 ^ n838 ^ 1'b0 ;
  assign n7348 = ~x83 & n7347 ;
  assign n7349 = n2957 ^ n293 ^ 1'b0 ;
  assign n7350 = n7348 | n7349 ;
  assign n7351 = n1572 & n7350 ;
  assign n7353 = n767 & n2085 ;
  assign n7352 = n327 & ~n2192 ;
  assign n7354 = n7353 ^ n7352 ^ 1'b0 ;
  assign n7355 = n2248 & ~n2993 ;
  assign n7356 = n3426 ^ n2323 ^ 1'b0 ;
  assign n7357 = ~n1329 & n7356 ;
  assign n7358 = ~n7355 & n7357 ;
  assign n7359 = ~n6136 & n7358 ;
  assign n7360 = n5262 & ~n7160 ;
  assign n7361 = n7360 ^ n2861 ^ 1'b0 ;
  assign n7362 = n7361 ^ n6848 ^ n3041 ;
  assign n7363 = n2993 | n3580 ;
  assign n7364 = n7363 ^ n6649 ^ 1'b0 ;
  assign n7365 = ~n250 & n6929 ;
  assign n7366 = n7365 ^ n1842 ^ 1'b0 ;
  assign n7367 = n5371 ^ n1582 ^ 1'b0 ;
  assign n7368 = ~n681 & n4273 ;
  assign n7369 = n530 ^ n180 ^ 1'b0 ;
  assign n7370 = n1578 & n7369 ;
  assign n7371 = n3709 & n7370 ;
  assign n7372 = n6877 & n7371 ;
  assign n7373 = n7372 ^ n6988 ^ 1'b0 ;
  assign n7375 = n496 & n2295 ;
  assign n7374 = n2953 & n3744 ;
  assign n7376 = n7375 ^ n7374 ^ 1'b0 ;
  assign n7377 = n260 & n4409 ;
  assign n7378 = n7377 ^ n3237 ^ n368 ;
  assign n7380 = n765 & n7029 ;
  assign n7379 = n3965 | n4883 ;
  assign n7381 = n7380 ^ n7379 ^ 1'b0 ;
  assign n7382 = n2628 ^ n511 ^ 1'b0 ;
  assign n7384 = ~n559 & n1529 ;
  assign n7385 = n7384 ^ n2427 ^ n166 ;
  assign n7386 = n7385 ^ n2463 ^ 1'b0 ;
  assign n7391 = ( n1537 & n2021 ) | ( n1537 & n3641 ) | ( n2021 & n3641 ) ;
  assign n7388 = ~n882 & n5209 ;
  assign n7387 = n2057 & n4050 ;
  assign n7389 = n7388 ^ n7387 ^ 1'b0 ;
  assign n7390 = n5830 & n7389 ;
  assign n7392 = n7391 ^ n7390 ^ 1'b0 ;
  assign n7393 = n7386 & n7392 ;
  assign n7383 = n3269 ^ n1689 ^ n481 ;
  assign n7394 = n7393 ^ n7383 ^ 1'b0 ;
  assign n7395 = n386 | n1037 ;
  assign n7396 = n7395 ^ n2596 ^ 1'b0 ;
  assign n7399 = n2461 ^ n1608 ^ 1'b0 ;
  assign n7398 = n4506 | n5152 ;
  assign n7400 = n7399 ^ n7398 ^ 1'b0 ;
  assign n7397 = n3009 | n4909 ;
  assign n7401 = n7400 ^ n7397 ^ 1'b0 ;
  assign n7402 = ~n3135 & n3685 ;
  assign n7403 = n7402 ^ n2520 ^ 1'b0 ;
  assign n7404 = ~n3070 & n3615 ;
  assign n7405 = n5075 & n7404 ;
  assign n7406 = ~n1331 & n7405 ;
  assign n7407 = x50 & n4840 ;
  assign n7408 = ~n628 & n7407 ;
  assign n7409 = n4863 ^ n975 ^ 1'b0 ;
  assign n7410 = ~n7408 & n7409 ;
  assign n7411 = x34 & ~n1761 ;
  assign n7412 = n7411 ^ n4503 ^ 1'b0 ;
  assign n7413 = n1997 ^ n1774 ^ 1'b0 ;
  assign n7414 = n6446 ^ n1089 ^ 1'b0 ;
  assign n7415 = n7413 | n7414 ;
  assign n7422 = x90 | n468 ;
  assign n7416 = n1992 ^ n1842 ^ 1'b0 ;
  assign n7417 = n1311 ^ n605 ^ 1'b0 ;
  assign n7418 = n1005 | n7417 ;
  assign n7419 = n7418 ^ n681 ^ 1'b0 ;
  assign n7420 = ~n3264 & n7419 ;
  assign n7421 = ( n1154 & ~n7416 ) | ( n1154 & n7420 ) | ( ~n7416 & n7420 ) ;
  assign n7423 = n7422 ^ n7421 ^ 1'b0 ;
  assign n7424 = n4190 & ~n6728 ;
  assign n7425 = n2591 ^ n975 ^ 1'b0 ;
  assign n7426 = ( ~n613 & n1233 ) | ( ~n613 & n3338 ) | ( n1233 & n3338 ) ;
  assign n7427 = n806 | n4736 ;
  assign n7428 = n7427 ^ n6837 ^ 1'b0 ;
  assign n7429 = n4345 & n7428 ;
  assign n7430 = ( n7425 & n7426 ) | ( n7425 & ~n7429 ) | ( n7426 & ~n7429 ) ;
  assign n7431 = n2321 ^ n967 ^ 1'b0 ;
  assign n7432 = ( n1166 & n2471 ) | ( n1166 & n5978 ) | ( n2471 & n5978 ) ;
  assign n7433 = ~n2120 & n7432 ;
  assign n7434 = n7036 | n7433 ;
  assign n7437 = n2438 | n2905 ;
  assign n7435 = n511 & ~n2865 ;
  assign n7436 = n3745 & n7435 ;
  assign n7438 = n7437 ^ n7436 ^ n340 ;
  assign n7439 = ( n2013 & n5131 ) | ( n2013 & n7438 ) | ( n5131 & n7438 ) ;
  assign n7440 = n5554 ^ n2107 ^ 1'b0 ;
  assign n7441 = ~n5002 & n7440 ;
  assign n7442 = x88 & n2778 ;
  assign n7443 = n7029 & n7442 ;
  assign n7444 = n7443 ^ n2261 ^ 1'b0 ;
  assign n7445 = n673 | n6190 ;
  assign n7446 = n7445 ^ n4205 ^ 1'b0 ;
  assign n7447 = n407 & n7394 ;
  assign n7448 = n4564 ^ n2730 ^ 1'b0 ;
  assign n7449 = n210 & n7448 ;
  assign n7450 = n5805 & n7449 ;
  assign n7451 = n3410 ^ n1817 ^ n313 ;
  assign n7452 = n369 | n1612 ;
  assign n7453 = n885 | n7452 ;
  assign n7454 = n7453 ^ n2470 ^ 1'b0 ;
  assign n7455 = n4373 | n7454 ;
  assign n7456 = ( n1845 & ~n2630 ) | ( n1845 & n4125 ) | ( ~n2630 & n4125 ) ;
  assign n7457 = n297 & n1816 ;
  assign n7458 = n7457 ^ n1433 ^ 1'b0 ;
  assign n7459 = ~n7456 & n7458 ;
  assign n7460 = n4551 ^ n464 ^ 1'b0 ;
  assign n7461 = n4759 | n7460 ;
  assign n7462 = x112 & ~n3620 ;
  assign n7463 = n7462 ^ n1097 ^ 1'b0 ;
  assign n7464 = ( n618 & ~n5632 ) | ( n618 & n6167 ) | ( ~n5632 & n6167 ) ;
  assign n7465 = ( n4541 & n7463 ) | ( n4541 & n7464 ) | ( n7463 & n7464 ) ;
  assign n7466 = n2892 ^ n2382 ^ x5 ;
  assign n7467 = n7466 ^ n1325 ^ 1'b0 ;
  assign n7468 = n7465 & n7467 ;
  assign n7469 = n5152 & ~n7160 ;
  assign n7470 = ~n2754 & n5521 ;
  assign n7471 = n2685 ^ n1338 ^ 1'b0 ;
  assign n7472 = n7470 & ~n7471 ;
  assign n7473 = n7472 ^ n4686 ^ 1'b0 ;
  assign n7474 = n2619 ^ n1230 ^ 1'b0 ;
  assign n7475 = ~n258 & n5840 ;
  assign n7476 = n7474 | n7475 ;
  assign n7477 = n4899 | n6818 ;
  assign n7478 = n7477 ^ n6376 ^ 1'b0 ;
  assign n7479 = n3353 | n5868 ;
  assign n7480 = n308 & n402 ;
  assign n7481 = n1761 & n7480 ;
  assign n7482 = n1740 | n7481 ;
  assign n7483 = n5453 & ~n7482 ;
  assign n7484 = n5801 ^ n5640 ^ 1'b0 ;
  assign n7485 = ( n5109 & n7483 ) | ( n5109 & ~n7484 ) | ( n7483 & ~n7484 ) ;
  assign n7486 = ~n662 & n4221 ;
  assign n7487 = n1507 & ~n2395 ;
  assign n7488 = ~n1325 & n7487 ;
  assign n7489 = n2945 | n7488 ;
  assign n7490 = n2051 | n7489 ;
  assign n7491 = n7490 ^ n521 ^ 1'b0 ;
  assign n7492 = n3579 & ~n7491 ;
  assign n7493 = n5018 ^ n1520 ^ 1'b0 ;
  assign n7494 = ( n2071 & ~n6000 ) | ( n2071 & n7493 ) | ( ~n6000 & n7493 ) ;
  assign n7495 = ~n2899 & n7494 ;
  assign n7496 = n4893 ^ n2450 ^ 1'b0 ;
  assign n7497 = n3001 ^ n163 ^ 1'b0 ;
  assign n7498 = n2055 & n7497 ;
  assign n7499 = n5015 ^ n419 ^ 1'b0 ;
  assign n7500 = n6990 & n7499 ;
  assign n7501 = n5038 ^ n2382 ^ n683 ;
  assign n7503 = n3848 | n5374 ;
  assign n7504 = n7503 ^ n4325 ^ 1'b0 ;
  assign n7502 = n941 | n6401 ;
  assign n7505 = n7504 ^ n7502 ^ 1'b0 ;
  assign n7506 = n1812 ^ n1193 ^ 1'b0 ;
  assign n7507 = ~n2428 & n6636 ;
  assign n7508 = n7506 & n7507 ;
  assign n7509 = n7508 ^ n5420 ^ 1'b0 ;
  assign n7510 = n6189 | n7509 ;
  assign n7511 = n7510 ^ n3067 ^ 1'b0 ;
  assign n7512 = n1908 ^ n636 ^ 1'b0 ;
  assign n7513 = ~n3485 & n7512 ;
  assign n7514 = n2740 | n2760 ;
  assign n7515 = n7514 ^ n2812 ^ 1'b0 ;
  assign n7516 = n3348 | n7515 ;
  assign n7517 = n2561 & ~n2647 ;
  assign n7518 = ~n2286 & n7517 ;
  assign n7519 = n2529 & n4315 ;
  assign n7520 = ~n4808 & n7519 ;
  assign n7521 = n7518 & n7520 ;
  assign n7523 = n192 & n1121 ;
  assign n7524 = n7523 ^ n2710 ^ 1'b0 ;
  assign n7522 = n1351 & ~n3295 ;
  assign n7525 = n7524 ^ n7522 ^ 1'b0 ;
  assign n7526 = n7521 & ~n7525 ;
  assign n7527 = ~n2324 & n2433 ;
  assign n7528 = n7527 ^ n2733 ^ 1'b0 ;
  assign n7529 = n468 & n1343 ;
  assign n7531 = n4857 ^ n1142 ^ 1'b0 ;
  assign n7530 = n1493 & n2034 ;
  assign n7532 = n7531 ^ n7530 ^ 1'b0 ;
  assign n7533 = n2142 & ~n7532 ;
  assign n7534 = n2506 & n7533 ;
  assign n7535 = ~n4606 & n7534 ;
  assign n7536 = n5390 ^ n4331 ^ 1'b0 ;
  assign n7537 = n1988 & n4912 ;
  assign n7538 = n7537 ^ n4613 ^ 1'b0 ;
  assign n7539 = ( ~n4953 & n7536 ) | ( ~n4953 & n7538 ) | ( n7536 & n7538 ) ;
  assign n7540 = n7539 ^ n147 ^ 1'b0 ;
  assign n7541 = n6454 ^ n488 ^ 1'b0 ;
  assign n7542 = n3721 & ~n7541 ;
  assign n7543 = n1213 & n7542 ;
  assign n7544 = n1169 & ~n3623 ;
  assign n7545 = n7544 ^ n5189 ^ 1'b0 ;
  assign n7546 = ~n5503 & n7545 ;
  assign n7547 = n4090 ^ n1193 ^ 1'b0 ;
  assign n7548 = n2373 & n7547 ;
  assign n7549 = n5722 ^ n1659 ^ 1'b0 ;
  assign n7551 = n3731 ^ n2792 ^ 1'b0 ;
  assign n7552 = n3773 & ~n4219 ;
  assign n7553 = ~n7551 & n7552 ;
  assign n7550 = n577 | n3470 ;
  assign n7554 = n7553 ^ n7550 ^ 1'b0 ;
  assign n7555 = n2425 & ~n3121 ;
  assign n7556 = n2206 & n7555 ;
  assign n7557 = n7556 ^ n5371 ^ 1'b0 ;
  assign n7558 = n4152 & ~n6377 ;
  assign n7559 = n7558 ^ n5586 ^ 1'b0 ;
  assign n7560 = x120 & n134 ;
  assign n7561 = ~x120 & n7560 ;
  assign n7562 = n213 & n1154 ;
  assign n7563 = n7561 & n7562 ;
  assign n7564 = n5055 & ~n7563 ;
  assign n7565 = n7564 ^ n637 ^ 1'b0 ;
  assign n7566 = ~n1105 & n7565 ;
  assign n7567 = n1270 | n2823 ;
  assign n7568 = n1661 & ~n7567 ;
  assign n7569 = n7568 ^ n6264 ^ 1'b0 ;
  assign n7570 = n5571 ^ n4781 ^ 1'b0 ;
  assign n7571 = n942 ^ n756 ^ 1'b0 ;
  assign n7572 = n7022 ^ n1116 ^ 1'b0 ;
  assign n7573 = n7571 & ~n7572 ;
  assign n7574 = ~n3881 & n7573 ;
  assign n7580 = n4408 ^ n2278 ^ 1'b0 ;
  assign n7581 = ~n2349 & n7580 ;
  assign n7575 = n1365 ^ n1176 ^ n922 ;
  assign n7576 = n7575 ^ n3982 ^ 1'b0 ;
  assign n7577 = x97 & ~n7576 ;
  assign n7578 = ( n4944 & ~n6059 ) | ( n4944 & n7577 ) | ( ~n6059 & n7577 ) ;
  assign n7579 = n1537 & ~n7578 ;
  assign n7582 = n7581 ^ n7579 ^ 1'b0 ;
  assign n7583 = ~n1383 & n6675 ;
  assign n7584 = n7583 ^ n6863 ^ 1'b0 ;
  assign n7585 = ( n4690 & ~n6132 ) | ( n4690 & n7584 ) | ( ~n6132 & n7584 ) ;
  assign n7586 = n808 & ~n7029 ;
  assign n7587 = n3193 & ~n5014 ;
  assign n7588 = ~n2794 & n3140 ;
  assign n7589 = n2267 | n2380 ;
  assign n7590 = n1941 & n7589 ;
  assign n7591 = n7590 ^ n7245 ^ 1'b0 ;
  assign n7592 = n7588 & n7591 ;
  assign n7593 = n309 | n3009 ;
  assign n7594 = n7593 ^ n2476 ^ 1'b0 ;
  assign n7599 = n5806 ^ n808 ^ 1'b0 ;
  assign n7600 = n2699 & n7599 ;
  assign n7601 = n3430 ^ n1149 ^ 1'b0 ;
  assign n7602 = n7600 & n7601 ;
  assign n7595 = ~n874 & n3824 ;
  assign n7596 = n5063 & n7595 ;
  assign n7597 = n5368 & n7596 ;
  assign n7598 = n710 | n7597 ;
  assign n7603 = n7602 ^ n7598 ^ 1'b0 ;
  assign n7604 = n4966 ^ n2148 ^ 1'b0 ;
  assign n7605 = n4115 ^ n2270 ^ 1'b0 ;
  assign n7606 = n2438 & ~n7605 ;
  assign n7607 = n2829 ^ n2765 ^ 1'b0 ;
  assign n7608 = n7607 ^ n4777 ^ 1'b0 ;
  assign n7609 = n7606 & ~n7608 ;
  assign n7610 = n3092 & ~n7609 ;
  assign n7611 = n879 & n5352 ;
  assign n7612 = n7611 ^ n2829 ^ 1'b0 ;
  assign n7613 = n1224 | n2763 ;
  assign n7614 = n5816 & ~n7613 ;
  assign n7615 = n7527 ^ n6932 ^ n5038 ;
  assign n7616 = x110 | n1616 ;
  assign n7617 = n1331 & ~n7616 ;
  assign n7618 = n4152 ^ n384 ^ 1'b0 ;
  assign n7619 = ~n1526 & n7618 ;
  assign n7620 = n2810 | n6004 ;
  assign n7621 = n7620 ^ n5293 ^ 1'b0 ;
  assign n7622 = ( n351 & n7619 ) | ( n351 & ~n7621 ) | ( n7619 & ~n7621 ) ;
  assign n7623 = n5950 ^ x47 ^ 1'b0 ;
  assign n7624 = n2499 ^ n1281 ^ n521 ;
  assign n7625 = n3109 & n7099 ;
  assign n7626 = ~n3768 & n6191 ;
  assign n7627 = n7626 ^ n4661 ^ 1'b0 ;
  assign n7628 = n4094 ^ n677 ^ 1'b0 ;
  assign n7629 = ~n5168 & n7628 ;
  assign n7630 = n4055 ^ n2300 ^ 1'b0 ;
  assign n7631 = n7457 & n7630 ;
  assign n7632 = n3940 ^ n2635 ^ 1'b0 ;
  assign n7633 = n7631 & n7632 ;
  assign n7634 = n2026 & n2949 ;
  assign n7635 = n7634 ^ n861 ^ 1'b0 ;
  assign n7636 = x78 & n7635 ;
  assign n7637 = n7636 ^ n5852 ^ 1'b0 ;
  assign n7638 = n7633 & ~n7637 ;
  assign n7639 = ~n7629 & n7638 ;
  assign n7640 = n7524 ^ n5157 ^ 1'b0 ;
  assign n7641 = n4268 | n7640 ;
  assign n7642 = ~n1767 & n5931 ;
  assign n7643 = n7642 ^ n6366 ^ 1'b0 ;
  assign n7644 = n5889 ^ x51 ^ 1'b0 ;
  assign n7645 = n7644 ^ n3234 ^ 1'b0 ;
  assign n7646 = ~n2577 & n2751 ;
  assign n7647 = n1725 ^ x97 ^ 1'b0 ;
  assign n7648 = n7646 & ~n7647 ;
  assign n7649 = n5364 | n7648 ;
  assign n7650 = n4290 ^ n1617 ^ 1'b0 ;
  assign n7651 = n1015 | n4755 ;
  assign n7652 = n732 | n7651 ;
  assign n7653 = n7652 ^ n6879 ^ 1'b0 ;
  assign n7654 = n949 ^ n533 ^ n336 ;
  assign n7655 = n5764 & n7654 ;
  assign n7656 = ~n1191 & n1790 ;
  assign n7657 = n3272 & ~n4128 ;
  assign n7658 = x52 | n7657 ;
  assign n7659 = n2323 | n2659 ;
  assign n7660 = x48 & n6235 ;
  assign n7661 = n7659 & n7660 ;
  assign n7662 = n477 & ~n2113 ;
  assign n7663 = n5466 | n7662 ;
  assign n7664 = n7663 ^ n3733 ^ 1'b0 ;
  assign n7665 = n7501 ^ n7175 ^ 1'b0 ;
  assign n7667 = ~n2240 & n2705 ;
  assign n7668 = n2240 & n7667 ;
  assign n7669 = n4352 & ~n7668 ;
  assign n7670 = ~n4352 & n7669 ;
  assign n7666 = n377 | n588 ;
  assign n7671 = n7670 ^ n7666 ^ n1581 ;
  assign n7672 = n5062 & ~n5526 ;
  assign n7673 = n7672 ^ n809 ^ 1'b0 ;
  assign n7674 = ( n1718 & n2676 ) | ( n1718 & ~n5775 ) | ( n2676 & ~n5775 ) ;
  assign n7675 = n4935 & ~n7674 ;
  assign n7676 = n7675 ^ n815 ^ 1'b0 ;
  assign n7677 = n7673 | n7676 ;
  assign n7678 = n1698 & ~n5195 ;
  assign n7679 = x81 & n7678 ;
  assign n7680 = n849 & n7679 ;
  assign n7681 = n2306 ^ n1419 ^ 1'b0 ;
  assign n7682 = n1914 & n7681 ;
  assign n7683 = ~n796 & n3386 ;
  assign n7684 = n5109 & n7683 ;
  assign n7685 = ~n3968 & n5435 ;
  assign n7690 = n2207 & ~n6112 ;
  assign n7686 = n2928 ^ n377 ^ 1'b0 ;
  assign n7687 = n664 & n7686 ;
  assign n7688 = n7687 ^ n2573 ^ 1'b0 ;
  assign n7689 = n645 & n7688 ;
  assign n7691 = n7690 ^ n7689 ^ 1'b0 ;
  assign n7692 = n2221 & ~n7691 ;
  assign n7693 = n7692 ^ n1009 ^ 1'b0 ;
  assign n7694 = n1145 ^ n867 ^ 1'b0 ;
  assign n7695 = n3806 & n7694 ;
  assign n7696 = ~n556 & n7695 ;
  assign n7697 = n7696 ^ n1495 ^ 1'b0 ;
  assign n7698 = n6629 | n7697 ;
  assign n7699 = n3004 & n6055 ;
  assign n7701 = n1028 | n1064 ;
  assign n7702 = n7701 ^ n5244 ^ 1'b0 ;
  assign n7700 = x10 & n7548 ;
  assign n7703 = n7702 ^ n7700 ^ 1'b0 ;
  assign n7704 = ~x2 & n2265 ;
  assign n7705 = n7704 ^ n5768 ^ 1'b0 ;
  assign n7706 = n2409 & n3511 ;
  assign n7707 = n3359 ^ n3162 ^ n1115 ;
  assign n7708 = n2953 ^ n1338 ^ 1'b0 ;
  assign n7709 = ( n1686 & ~n2760 ) | ( n1686 & n3910 ) | ( ~n2760 & n3910 ) ;
  assign n7710 = n1147 & ~n7301 ;
  assign n7711 = n7709 & ~n7710 ;
  assign n7712 = n7711 ^ n5728 ^ n179 ;
  assign n7713 = ~n852 & n4774 ;
  assign n7714 = n5014 & n7713 ;
  assign n7715 = ~x107 & n7714 ;
  assign n7716 = n6905 ^ n2389 ^ 1'b0 ;
  assign n7717 = n4433 ^ n1687 ^ 1'b0 ;
  assign n7718 = n361 | n7717 ;
  assign n7719 = n2261 & n2354 ;
  assign n7720 = ~n1066 & n3792 ;
  assign n7721 = n1225 | n5290 ;
  assign n7722 = n3158 & ~n7721 ;
  assign n7723 = n415 & n7722 ;
  assign n7725 = ~n3350 & n4490 ;
  assign n7726 = ~n5778 & n7725 ;
  assign n7724 = n3340 & n4453 ;
  assign n7727 = n7726 ^ n7724 ^ 1'b0 ;
  assign n7728 = n2355 ^ n852 ^ 1'b0 ;
  assign n7729 = n1457 & ~n7728 ;
  assign n7730 = ~n553 & n7729 ;
  assign n7731 = n2213 & n7730 ;
  assign n7732 = n3501 & ~n4978 ;
  assign n7733 = n4877 | n7674 ;
  assign n7734 = n7733 ^ n3879 ^ 1'b0 ;
  assign n7735 = n7734 ^ n6211 ^ n2959 ;
  assign n7736 = n4159 & ~n7735 ;
  assign n7737 = ( n3481 & n3540 ) | ( n3481 & ~n7736 ) | ( n3540 & ~n7736 ) ;
  assign n7738 = n4388 ^ n2961 ^ 1'b0 ;
  assign n7741 = n4717 ^ n446 ^ 1'b0 ;
  assign n7739 = n6112 ^ n3951 ^ 1'b0 ;
  assign n7740 = n688 & ~n7739 ;
  assign n7742 = n7741 ^ n7740 ^ 1'b0 ;
  assign n7743 = ~n5539 & n6307 ;
  assign n7745 = n138 & n1193 ;
  assign n7746 = n7745 ^ n466 ^ 1'b0 ;
  assign n7744 = n1747 & n3424 ;
  assign n7747 = n7746 ^ n7744 ^ n2520 ;
  assign n7748 = n7747 ^ n5566 ^ 1'b0 ;
  assign n7749 = n7743 & n7748 ;
  assign n7750 = n1695 | n6407 ;
  assign n7751 = n7750 ^ n545 ^ 1'b0 ;
  assign n7752 = n2243 ^ n468 ^ 1'b0 ;
  assign n7753 = n2632 & n7752 ;
  assign n7754 = n4734 ^ n478 ^ 1'b0 ;
  assign n7755 = n7753 & ~n7754 ;
  assign n7756 = n7755 ^ n2479 ^ 1'b0 ;
  assign n7757 = ( n3367 & n7751 ) | ( n3367 & n7756 ) | ( n7751 & n7756 ) ;
  assign n7758 = x21 & n2896 ;
  assign n7759 = n7758 ^ n551 ^ 1'b0 ;
  assign n7760 = ~n507 & n5944 ;
  assign n7761 = ( n1858 & ~n7759 ) | ( n1858 & n7760 ) | ( ~n7759 & n7760 ) ;
  assign n7762 = n7713 ^ n2673 ^ 1'b0 ;
  assign n7765 = n3531 ^ n538 ^ 1'b0 ;
  assign n7763 = n468 & n7241 ;
  assign n7764 = n7763 ^ n2210 ^ 1'b0 ;
  assign n7766 = n7765 ^ n7764 ^ 1'b0 ;
  assign n7770 = n3255 & n5907 ;
  assign n7771 = n7770 ^ n392 ^ 1'b0 ;
  assign n7772 = n7771 ^ n5152 ^ n1898 ;
  assign n7767 = n2872 & ~n3430 ;
  assign n7768 = n7767 ^ n1293 ^ 1'b0 ;
  assign n7769 = n4496 | n7768 ;
  assign n7773 = n7772 ^ n7769 ^ n6854 ;
  assign n7774 = n669 | n3411 ;
  assign n7775 = n2448 | n3512 ;
  assign n7776 = n7775 ^ n3620 ^ 1'b0 ;
  assign n7777 = n6982 & n7776 ;
  assign n7778 = ~n556 & n6561 ;
  assign n7779 = ~n2890 & n3410 ;
  assign n7780 = n5840 ^ n1939 ^ 1'b0 ;
  assign n7782 = ( n229 & ~n2906 ) | ( n229 & n4037 ) | ( ~n2906 & n4037 ) ;
  assign n7781 = n3550 ^ n2494 ^ 1'b0 ;
  assign n7783 = n7782 ^ n7781 ^ n4777 ;
  assign n7784 = ( ~n811 & n5991 ) | ( ~n811 & n6342 ) | ( n5991 & n6342 ) ;
  assign n7785 = n3389 & ~n7213 ;
  assign n7786 = n231 & n7785 ;
  assign n7787 = n7786 ^ n2116 ^ 1'b0 ;
  assign n7788 = ~n1483 & n4853 ;
  assign n7789 = n7788 ^ n4666 ^ 1'b0 ;
  assign n7790 = n3437 | n7789 ;
  assign n7791 = n679 & ~n7790 ;
  assign n7797 = ~n1361 & n1608 ;
  assign n7795 = n1420 | n2333 ;
  assign n7796 = n4520 & ~n7795 ;
  assign n7798 = n7797 ^ n7796 ^ n2948 ;
  assign n7792 = n464 & ~n894 ;
  assign n7793 = n7792 ^ n2652 ^ 1'b0 ;
  assign n7794 = n3914 & n7793 ;
  assign n7799 = n7798 ^ n7794 ^ 1'b0 ;
  assign n7800 = n5691 ^ n3308 ^ 1'b0 ;
  assign n7801 = n523 & ~n7800 ;
  assign n7802 = n2022 & ~n6273 ;
  assign n7803 = n7802 ^ n533 ^ 1'b0 ;
  assign n7804 = n369 | n7803 ;
  assign n7805 = n6477 ^ n1322 ^ 1'b0 ;
  assign n7806 = ~x7 & n7606 ;
  assign n7807 = ~n1510 & n3459 ;
  assign n7808 = n349 & ~n7807 ;
  assign n7809 = n7808 ^ n1919 ^ 1'b0 ;
  assign n7810 = n7806 & ~n7809 ;
  assign n7811 = n7805 & n7810 ;
  assign n7815 = ~n3320 & n6181 ;
  assign n7812 = n1432 ^ x32 ^ 1'b0 ;
  assign n7813 = ~n3298 & n7812 ;
  assign n7814 = ~n5490 & n7813 ;
  assign n7816 = n7815 ^ n7814 ^ 1'b0 ;
  assign n7817 = ~n5720 & n7816 ;
  assign n7818 = ~n3550 & n7817 ;
  assign n7819 = n6704 ^ x41 ^ 1'b0 ;
  assign n7820 = n2497 | n7819 ;
  assign n7821 = ~n490 & n7820 ;
  assign n7822 = ~n5649 & n7662 ;
  assign n7823 = n1903 ^ n876 ^ 1'b0 ;
  assign n7824 = n7822 & ~n7823 ;
  assign n7825 = n632 & ~n5220 ;
  assign n7826 = ~n2979 & n7825 ;
  assign n7827 = ~n1261 & n1757 ;
  assign n7828 = n7827 ^ n1847 ^ 1'b0 ;
  assign n7829 = ( n3150 & ~n7826 ) | ( n3150 & n7828 ) | ( ~n7826 & n7828 ) ;
  assign n7830 = ~n4319 & n7829 ;
  assign n7831 = n1658 & ~n7483 ;
  assign n7832 = n7274 ^ n5050 ^ 1'b0 ;
  assign n7833 = n779 | n7832 ;
  assign n7834 = n7615 & ~n7833 ;
  assign n7835 = ~n1497 & n3160 ;
  assign n7836 = n7835 ^ n319 ^ 1'b0 ;
  assign n7837 = n2464 & n7836 ;
  assign n7838 = n6809 & n7416 ;
  assign n7839 = n7052 ^ n1452 ^ 1'b0 ;
  assign n7840 = n7839 ^ n2470 ^ 1'b0 ;
  assign n7841 = n4463 & n7712 ;
  assign n7842 = n7841 ^ n2870 ^ 1'b0 ;
  assign n7844 = n2644 & ~n2809 ;
  assign n7845 = n3982 & n7844 ;
  assign n7846 = ~n4463 & n7845 ;
  assign n7843 = ~n5347 & n7391 ;
  assign n7847 = n7846 ^ n7843 ^ 1'b0 ;
  assign n7848 = n5974 ^ n1692 ^ 1'b0 ;
  assign n7849 = n171 & ~n7848 ;
  assign n7850 = n1537 & n6222 ;
  assign n7851 = n7850 ^ n1182 ^ 1'b0 ;
  assign n7852 = n1943 ^ n1498 ^ x23 ;
  assign n7853 = n3319 & ~n6036 ;
  assign n7854 = n7852 & n7853 ;
  assign n7855 = n4866 & n7767 ;
  assign n7856 = n2448 ^ n2324 ^ 1'b0 ;
  assign n7857 = n4621 | n7856 ;
  assign n7858 = n7362 ^ n1664 ^ 1'b0 ;
  assign n7859 = ~n1832 & n2979 ;
  assign n7860 = n7859 ^ n2527 ^ 1'b0 ;
  assign n7866 = n4009 & n5085 ;
  assign n7861 = n6879 ^ n3632 ^ n2639 ;
  assign n7862 = n6152 & ~n6362 ;
  assign n7863 = n7861 & n7862 ;
  assign n7864 = n7050 | n7863 ;
  assign n7865 = n5261 | n7864 ;
  assign n7867 = n7866 ^ n7865 ^ 1'b0 ;
  assign n7868 = n6675 ^ n801 ^ 1'b0 ;
  assign n7869 = ~n4671 & n7868 ;
  assign n7870 = ~n1574 & n4342 ;
  assign n7871 = ~n2750 & n7870 ;
  assign n7872 = n7270 | n7871 ;
  assign n7873 = n7872 ^ n1500 ^ 1'b0 ;
  assign n7874 = ~n6058 & n7873 ;
  assign n7875 = n3659 ^ n3346 ^ 1'b0 ;
  assign n7876 = n5550 & n7875 ;
  assign n7877 = n3154 ^ n2697 ^ 1'b0 ;
  assign n7878 = ~n327 & n7877 ;
  assign n7879 = n1446 | n7878 ;
  assign n7880 = n5355 ^ n4095 ^ 1'b0 ;
  assign n7881 = ( n1629 & ~n2022 ) | ( n1629 & n3424 ) | ( ~n2022 & n3424 ) ;
  assign n7882 = ( ~n1083 & n2237 ) | ( ~n1083 & n7881 ) | ( n2237 & n7881 ) ;
  assign n7883 = ~n7880 & n7882 ;
  assign n7884 = n7883 ^ n4139 ^ 1'b0 ;
  assign n7886 = x6 & ~n4832 ;
  assign n7887 = ~n679 & n7886 ;
  assign n7885 = n2451 & ~n5928 ;
  assign n7888 = n7887 ^ n7885 ^ 1'b0 ;
  assign n7889 = x58 & n1047 ;
  assign n7890 = n7889 ^ n5557 ^ 1'b0 ;
  assign n7891 = n6646 ^ n999 ^ 1'b0 ;
  assign n7892 = n1691 ^ n959 ^ 1'b0 ;
  assign n7893 = x62 & ~n7892 ;
  assign n7894 = n509 & n7893 ;
  assign n7895 = n754 | n3557 ;
  assign n7896 = n7895 ^ n2342 ^ 1'b0 ;
  assign n7897 = ( n900 & ~n5593 ) | ( n900 & n7896 ) | ( ~n5593 & n7896 ) ;
  assign n7898 = ~n2983 & n7897 ;
  assign n7899 = ~n577 & n6695 ;
  assign n7900 = n7899 ^ n3255 ^ 1'b0 ;
  assign n7901 = n2627 & ~n4736 ;
  assign n7902 = n2861 & n7901 ;
  assign n7903 = ( ~n1361 & n3395 ) | ( ~n1361 & n6652 ) | ( n3395 & n6652 ) ;
  assign n7904 = ~n5111 & n7903 ;
  assign n7905 = ~n738 & n7904 ;
  assign n7906 = n371 | n1079 ;
  assign n7907 = n1067 & n1399 ;
  assign n7908 = ~n1067 & n7907 ;
  assign n7909 = n1252 & ~n7908 ;
  assign n7910 = n7908 & n7909 ;
  assign n7911 = n3729 & ~n4554 ;
  assign n7912 = n7910 & n7911 ;
  assign n7913 = n5397 ^ n2012 ^ 1'b0 ;
  assign n7914 = n2196 & n7913 ;
  assign n7915 = n6145 & n7914 ;
  assign n7916 = n7915 ^ n373 ^ 1'b0 ;
  assign n7917 = n4965 & n7916 ;
  assign n7918 = n7912 & n7917 ;
  assign n7922 = n3936 ^ n177 ^ 1'b0 ;
  assign n7919 = n3209 ^ n2362 ^ 1'b0 ;
  assign n7920 = n2969 & ~n7919 ;
  assign n7921 = n2014 & n7920 ;
  assign n7923 = n7922 ^ n7921 ^ 1'b0 ;
  assign n7924 = n3916 | n6187 ;
  assign n7925 = n7924 ^ n4320 ^ 1'b0 ;
  assign n7926 = ~n1179 & n2302 ;
  assign n7927 = ~n3583 & n7926 ;
  assign n7928 = n7927 ^ n4612 ^ 1'b0 ;
  assign n7929 = ~n7925 & n7928 ;
  assign n7930 = n6087 ^ n1735 ^ 1'b0 ;
  assign n7931 = n7930 ^ n456 ^ 1'b0 ;
  assign n7932 = n1847 ^ n775 ^ 1'b0 ;
  assign n7933 = ~n358 & n7932 ;
  assign n7934 = n7933 ^ n3399 ^ 1'b0 ;
  assign n7935 = n2477 & n7934 ;
  assign n7936 = n7935 ^ n879 ^ 1'b0 ;
  assign n7937 = n3641 ^ n2869 ^ 1'b0 ;
  assign n7938 = n1222 & ~n7937 ;
  assign n7939 = n7938 ^ n6181 ^ 1'b0 ;
  assign n7940 = n5371 ^ n5033 ^ 1'b0 ;
  assign n7941 = x5 & ~n6448 ;
  assign n7945 = ~n2386 & n3968 ;
  assign n7946 = n1832 & n7945 ;
  assign n7942 = n5119 ^ n232 ^ 1'b0 ;
  assign n7943 = n4116 ^ n3696 ^ 1'b0 ;
  assign n7944 = n7942 | n7943 ;
  assign n7947 = n7946 ^ n7944 ^ 1'b0 ;
  assign n7948 = n7941 & n7947 ;
  assign n7949 = n5310 ^ n3603 ^ 1'b0 ;
  assign n7950 = n6013 & ~n7949 ;
  assign n7951 = n2542 & n7950 ;
  assign n7952 = ~n3724 & n4892 ;
  assign n7953 = ~n3383 & n7952 ;
  assign n7954 = n273 & ~n7953 ;
  assign n7955 = n2898 ^ n1138 ^ 1'b0 ;
  assign n7956 = n7955 ^ n6206 ^ n3853 ;
  assign n7957 = n129 & n3302 ;
  assign n7958 = n192 & n3262 ;
  assign n7959 = n613 & n2470 ;
  assign n7960 = n1121 ^ n613 ^ 1'b0 ;
  assign n7961 = n7960 ^ n7394 ^ n2976 ;
  assign n7962 = x115 & ~n1136 ;
  assign n7963 = n858 & n7962 ;
  assign n7964 = n4238 ^ n2064 ^ 1'b0 ;
  assign n7965 = n533 & ~n5655 ;
  assign n7966 = ~n725 & n7965 ;
  assign n7967 = n902 & n1439 ;
  assign n7968 = ~n2790 & n4004 ;
  assign n7969 = n7607 ^ n3536 ^ 1'b0 ;
  assign n7970 = ~n7968 & n7969 ;
  assign n7971 = n4727 ^ n3022 ^ 1'b0 ;
  assign n7972 = n1130 | n7971 ;
  assign n7973 = ~n163 & n2217 ;
  assign n7974 = n7973 ^ n3404 ^ 1'b0 ;
  assign n7980 = ( ~n1587 & n1978 ) | ( ~n1587 & n2986 ) | ( n1978 & n2986 ) ;
  assign n7981 = n7980 ^ n6639 ^ 1'b0 ;
  assign n7975 = n4222 & ~n7532 ;
  assign n7976 = n147 & n3237 ;
  assign n7977 = n7976 ^ n3266 ^ 1'b0 ;
  assign n7978 = n2610 & n7977 ;
  assign n7979 = ~n7975 & n7978 ;
  assign n7982 = n7981 ^ n7979 ^ 1'b0 ;
  assign n7987 = n929 | n1509 ;
  assign n7983 = n861 ^ n455 ^ 1'b0 ;
  assign n7984 = n1570 & n7983 ;
  assign n7985 = n7984 ^ n2813 ^ n994 ;
  assign n7986 = n7985 ^ n1398 ^ 1'b0 ;
  assign n7988 = n7987 ^ n7986 ^ 1'b0 ;
  assign n7991 = n1250 | n2341 ;
  assign n7992 = n7991 ^ n368 ^ 1'b0 ;
  assign n7989 = n455 | n7880 ;
  assign n7990 = n4806 | n7989 ;
  assign n7993 = n7992 ^ n7990 ^ 1'b0 ;
  assign n7994 = n5915 | n7493 ;
  assign n7995 = n7993 & ~n7994 ;
  assign n7996 = n759 & ~n7584 ;
  assign n7997 = ~n4295 & n7996 ;
  assign n8001 = n269 & ~n2967 ;
  assign n8002 = n504 & n8001 ;
  assign n7998 = n2883 | n3000 ;
  assign n7999 = ~n6766 & n7998 ;
  assign n8000 = n7999 ^ n4804 ^ 1'b0 ;
  assign n8003 = n8002 ^ n8000 ^ n7456 ;
  assign n8004 = ~n147 & n269 ;
  assign n8005 = n8004 ^ n6225 ^ 1'b0 ;
  assign n8006 = n8005 ^ n6995 ^ n843 ;
  assign n8007 = n960 & ~n3193 ;
  assign n8008 = n1832 & n7345 ;
  assign n8009 = n8008 ^ n5897 ^ 1'b0 ;
  assign n8010 = n3072 & ~n5507 ;
  assign n8011 = ~x93 & n8010 ;
  assign n8012 = n1599 & ~n8011 ;
  assign n8013 = n7249 & ~n7604 ;
  assign n8014 = n7818 ^ n947 ^ 1'b0 ;
  assign n8015 = n1578 & n8014 ;
  assign n8018 = n1235 ^ n338 ^ 1'b0 ;
  assign n8019 = n930 & ~n8018 ;
  assign n8016 = n384 & ~n729 ;
  assign n8017 = ~n5837 & n8016 ;
  assign n8020 = n8019 ^ n8017 ^ 1'b0 ;
  assign n8021 = n643 | n8020 ;
  assign n8022 = n6009 ^ n4352 ^ 1'b0 ;
  assign n8023 = n1955 | n8022 ;
  assign n8024 = n6477 & ~n8023 ;
  assign n8025 = n8024 ^ n1917 ^ 1'b0 ;
  assign n8026 = n2922 ^ x98 ^ 1'b0 ;
  assign n8027 = n7288 ^ n2337 ^ 1'b0 ;
  assign n8028 = n2151 & n7538 ;
  assign n8029 = n8027 & n8028 ;
  assign n8030 = n2806 & n6449 ;
  assign n8031 = ~n2510 & n2848 ;
  assign n8032 = ~n2364 & n5637 ;
  assign n8033 = n8032 ^ n2866 ^ 1'b0 ;
  assign n8034 = n8033 ^ n7920 ^ 1'b0 ;
  assign n8035 = n2371 | n8034 ;
  assign n8036 = n6210 ^ n3195 ^ 1'b0 ;
  assign n8037 = n8036 ^ n4463 ^ 1'b0 ;
  assign n8038 = n458 & ~n8037 ;
  assign n8039 = ~n1410 & n2673 ;
  assign n8040 = n8039 ^ n1225 ^ 1'b0 ;
  assign n8041 = n4927 ^ n1369 ^ 1'b0 ;
  assign n8050 = n751 | n1138 ;
  assign n8051 = n8050 ^ n6657 ^ n1205 ;
  assign n8052 = n8051 ^ n386 ^ 1'b0 ;
  assign n8042 = ~n4087 & n5253 ;
  assign n8043 = n1955 & n8042 ;
  assign n8044 = n1651 & n5860 ;
  assign n8045 = n8044 ^ n4350 ^ 1'b0 ;
  assign n8046 = ~n5595 & n8045 ;
  assign n8047 = n8043 & n8046 ;
  assign n8048 = n5610 | n6497 ;
  assign n8049 = n8047 | n8048 ;
  assign n8053 = n8052 ^ n8049 ^ 1'b0 ;
  assign n8054 = n5310 ^ n311 ^ 1'b0 ;
  assign n8055 = n4408 | n5443 ;
  assign n8056 = n8055 ^ n7089 ^ 1'b0 ;
  assign n8060 = n3354 & ~n6840 ;
  assign n8061 = n8060 ^ n3350 ^ 1'b0 ;
  assign n8062 = n3389 & ~n8061 ;
  assign n8059 = n1406 | n2022 ;
  assign n8057 = n2922 & ~n4597 ;
  assign n8058 = n8057 ^ x41 ^ 1'b0 ;
  assign n8063 = n8062 ^ n8059 ^ n8058 ;
  assign n8064 = n331 & ~n373 ;
  assign n8065 = n8064 ^ n2048 ^ 1'b0 ;
  assign n8066 = n2121 & ~n7203 ;
  assign n8067 = n4375 & n8066 ;
  assign n8068 = ~n2845 & n8067 ;
  assign n8069 = ~n5152 & n5808 ;
  assign n8070 = n8069 ^ n4767 ^ 1'b0 ;
  assign n8071 = n7695 & n8008 ;
  assign n8074 = n7425 ^ n3780 ^ 1'b0 ;
  assign n8072 = ~n452 & n1697 ;
  assign n8073 = ~n2020 & n8072 ;
  assign n8075 = n8074 ^ n8073 ^ 1'b0 ;
  assign n8076 = n4430 ^ n2986 ^ 1'b0 ;
  assign n8077 = ~n1383 & n8076 ;
  assign n8078 = n339 & ~n1093 ;
  assign n8079 = n3813 ^ x2 ^ 1'b0 ;
  assign n8080 = ~n3510 & n8079 ;
  assign n8081 = n4661 & n8080 ;
  assign n8082 = n685 & n1647 ;
  assign n8083 = n4857 & ~n8082 ;
  assign n8084 = n3159 ^ n1716 ^ 1'b0 ;
  assign n8085 = ~n2189 & n8084 ;
  assign n8086 = n5220 & ~n8085 ;
  assign n8087 = n8086 ^ n1988 ^ 1'b0 ;
  assign n8088 = n3529 & n6742 ;
  assign n8089 = n8087 & n8088 ;
  assign n8090 = n4530 ^ n816 ^ 1'b0 ;
  assign n8091 = n196 & n4997 ;
  assign n8092 = n8091 ^ n1394 ^ 1'b0 ;
  assign n8093 = n8092 ^ n6423 ^ 1'b0 ;
  assign n8094 = n5832 & ~n8093 ;
  assign n8096 = n5638 ^ n2712 ^ n459 ;
  assign n8095 = n1888 & n2731 ;
  assign n8097 = n8096 ^ n8095 ^ 1'b0 ;
  assign n8098 = n8097 ^ n4467 ^ 1'b0 ;
  assign n8099 = ( ~x96 & n1771 ) | ( ~x96 & n3006 ) | ( n1771 & n3006 ) ;
  assign n8100 = n8099 ^ n1076 ^ n324 ;
  assign n8101 = ( n1867 & ~n4327 ) | ( n1867 & n6532 ) | ( ~n4327 & n6532 ) ;
  assign n8102 = n3789 ^ n2414 ^ 1'b0 ;
  assign n8103 = n1988 & ~n8102 ;
  assign n8104 = ~x98 & n8103 ;
  assign n8105 = n1067 & n3391 ;
  assign n8106 = n1465 & n8105 ;
  assign n8107 = n8106 ^ n5228 ^ n2142 ;
  assign n8108 = ( n1211 & n2057 ) | ( n1211 & ~n5843 ) | ( n2057 & ~n5843 ) ;
  assign n8109 = n5050 & n8108 ;
  assign n8110 = n8109 ^ n5273 ^ n3559 ;
  assign n8111 = n8110 ^ n3048 ^ n2458 ;
  assign n8112 = n4556 ^ n143 ^ 1'b0 ;
  assign n8113 = n8112 ^ n4396 ^ 1'b0 ;
  assign n8114 = n4095 & ~n7182 ;
  assign n8115 = n947 ^ x49 ^ 1'b0 ;
  assign n8116 = n281 | n8115 ;
  assign n8117 = n4011 & ~n8116 ;
  assign n8118 = n8117 ^ n5423 ^ 1'b0 ;
  assign n8119 = n2502 & n6421 ;
  assign n8120 = n4113 ^ x39 ^ 1'b0 ;
  assign n8121 = n2106 | n8120 ;
  assign n8122 = n3986 & ~n8121 ;
  assign n8123 = n4048 & n6246 ;
  assign n8124 = n6423 ^ n762 ^ 1'b0 ;
  assign n8125 = n1489 & ~n8124 ;
  assign n8126 = n8125 ^ n1624 ^ 1'b0 ;
  assign n8127 = n8126 ^ n1687 ^ 1'b0 ;
  assign n8128 = n6802 | n7857 ;
  assign n8129 = n3390 & n8066 ;
  assign n8130 = ~n639 & n8129 ;
  assign n8131 = n8130 ^ n5797 ^ 1'b0 ;
  assign n8132 = n4325 ^ n551 ^ 1'b0 ;
  assign n8133 = n8132 ^ n3368 ^ 1'b0 ;
  assign n8134 = n401 | n8133 ;
  assign n8137 = n336 & n8019 ;
  assign n8138 = ~n1433 & n8137 ;
  assign n8135 = ~n2701 & n4774 ;
  assign n8136 = ~n1394 & n8135 ;
  assign n8139 = n8138 ^ n8136 ^ 1'b0 ;
  assign n8140 = n4998 | n6783 ;
  assign n8141 = n6418 ^ n2922 ^ 1'b0 ;
  assign n8142 = n1639 & ~n8141 ;
  assign n8143 = n3575 | n4120 ;
  assign n8144 = n867 | n8143 ;
  assign n8145 = ~n2106 & n8144 ;
  assign n8146 = ~n2416 & n8145 ;
  assign n8147 = ~n3110 & n8146 ;
  assign n8148 = n2628 ^ x6 ^ 1'b0 ;
  assign n8149 = n7086 ^ n5517 ^ n5079 ;
  assign n8150 = n2733 | n2838 ;
  assign n8151 = n8150 ^ n4455 ^ 1'b0 ;
  assign n8152 = n4456 & ~n8151 ;
  assign n8153 = n8152 ^ n741 ^ 1'b0 ;
  assign n8154 = n1803 & ~n4292 ;
  assign n8155 = ~n530 & n8154 ;
  assign n8156 = ~n3458 & n8155 ;
  assign n8160 = ~n3360 & n5084 ;
  assign n8161 = n8160 ^ n4150 ^ 1'b0 ;
  assign n8157 = ~n2865 & n2992 ;
  assign n8158 = ~x125 & n8157 ;
  assign n8159 = n5634 & ~n8158 ;
  assign n8162 = n8161 ^ n8159 ^ 1'b0 ;
  assign n8163 = n1334 & n4171 ;
  assign n8164 = n8163 ^ n309 ^ 1'b0 ;
  assign n8165 = ( x99 & ~n2176 ) | ( x99 & n8164 ) | ( ~n2176 & n8164 ) ;
  assign n8166 = n4717 & ~n8119 ;
  assign n8167 = ~n8165 & n8166 ;
  assign n8169 = n5416 ^ n2159 ^ 1'b0 ;
  assign n8170 = n2903 & n8169 ;
  assign n8168 = n6109 ^ n1402 ^ n1250 ;
  assign n8171 = n8170 ^ n8168 ^ n2235 ;
  assign n8172 = ( n1750 & n4182 ) | ( n1750 & ~n6636 ) | ( n4182 & ~n6636 ) ;
  assign n8173 = n7800 & ~n8172 ;
  assign n8174 = n8173 ^ n5970 ^ 1'b0 ;
  assign n8175 = ( n2084 & n3859 ) | ( n2084 & n5852 ) | ( n3859 & n5852 ) ;
  assign n8176 = ( n2638 & ~n6126 ) | ( n2638 & n8175 ) | ( ~n6126 & n8175 ) ;
  assign n8177 = n8176 ^ x68 ^ 1'b0 ;
  assign n8178 = ( n2076 & ~n2131 ) | ( n2076 & n2832 ) | ( ~n2131 & n2832 ) ;
  assign n8179 = n1635 | n6716 ;
  assign n8180 = n8179 ^ n3192 ^ 1'b0 ;
  assign n8181 = n8178 | n8180 ;
  assign n8182 = n708 & n4269 ;
  assign n8183 = n373 & n8182 ;
  assign n8184 = n8183 ^ n241 ^ 1'b0 ;
  assign n8185 = n1285 & n1396 ;
  assign n8186 = n2022 & ~n8185 ;
  assign n8187 = n8186 ^ n2470 ^ 1'b0 ;
  assign n8188 = n1084 & ~n5067 ;
  assign n8189 = n8188 ^ n6187 ^ 1'b0 ;
  assign n8190 = n7045 ^ n5277 ^ 1'b0 ;
  assign n8191 = n8189 & ~n8190 ;
  assign n8193 = n851 | n1574 ;
  assign n8194 = n8193 ^ n1756 ^ 1'b0 ;
  assign n8192 = n425 | n6846 ;
  assign n8195 = n8194 ^ n8192 ^ 1'b0 ;
  assign n8196 = n8191 & ~n8195 ;
  assign n8197 = n2206 & n8196 ;
  assign n8198 = n4436 | n4676 ;
  assign n8199 = n6511 ^ n2685 ^ 1'b0 ;
  assign n8200 = n876 & n2650 ;
  assign n8201 = ( x65 & ~n4199 ) | ( x65 & n8200 ) | ( ~n4199 & n8200 ) ;
  assign n8202 = n2413 & n4936 ;
  assign n8203 = n8202 ^ n3273 ^ 1'b0 ;
  assign n8204 = n1193 ^ n231 ^ 1'b0 ;
  assign n8205 = ( n725 & n1851 ) | ( n725 & ~n3795 ) | ( n1851 & ~n3795 ) ;
  assign n8206 = n8205 ^ n6038 ^ 1'b0 ;
  assign n8207 = n4018 & n6237 ;
  assign n8208 = n4811 & n8207 ;
  assign n8209 = n5908 | n6165 ;
  assign n8210 = n754 | n4590 ;
  assign n8211 = n4929 & n6315 ;
  assign n8212 = n8211 ^ n4412 ^ 1'b0 ;
  assign n8213 = n8210 & ~n8212 ;
  assign n8214 = n8213 ^ n5067 ^ 1'b0 ;
  assign n8215 = n3122 & n8214 ;
  assign n8216 = n4630 & n5980 ;
  assign n8217 = n7012 & n8216 ;
  assign n8218 = n2109 & n6116 ;
  assign n8219 = n7736 & n8218 ;
  assign n8220 = n6573 ^ n5163 ^ 1'b0 ;
  assign n8221 = ( n1094 & n3714 ) | ( n1094 & ~n5455 ) | ( n3714 & ~n5455 ) ;
  assign n8222 = n6998 ^ n888 ^ 1'b0 ;
  assign n8223 = n6858 | n8222 ;
  assign n8224 = n4542 & n5412 ;
  assign n8225 = n180 | n6416 ;
  assign n8226 = n8225 ^ n6667 ^ 1'b0 ;
  assign n8227 = n5440 & n8226 ;
  assign n8228 = ~n5889 & n8227 ;
  assign n8229 = ~n8224 & n8228 ;
  assign n8230 = n5813 & ~n7085 ;
  assign n8231 = ~n7202 & n8230 ;
  assign n8232 = ~n1079 & n4597 ;
  assign n8233 = ~n6932 & n8232 ;
  assign n8234 = x111 & ~n8233 ;
  assign n8235 = n8234 ^ n5206 ^ 1'b0 ;
  assign n8236 = n7688 ^ n5463 ^ n2392 ;
  assign n8237 = n3321 & n4897 ;
  assign n8238 = n8236 & n8237 ;
  assign n8239 = n8238 ^ n1470 ^ 1'b0 ;
  assign n8240 = ( n2441 & n2774 ) | ( n2441 & ~n7734 ) | ( n2774 & ~n7734 ) ;
  assign n8241 = n5352 ^ n3438 ^ 1'b0 ;
  assign n8242 = ~n6259 & n8241 ;
  assign n8243 = n1996 & n8242 ;
  assign n8244 = n5571 ^ n4219 ^ 1'b0 ;
  assign n8245 = n8244 ^ n5119 ^ n3037 ;
  assign n8246 = ( n1052 & n2886 ) | ( n1052 & ~n5530 ) | ( n2886 & ~n5530 ) ;
  assign n8248 = n1769 ^ n1464 ^ n303 ;
  assign n8247 = n1261 & n1599 ;
  assign n8249 = n8248 ^ n8247 ^ n609 ;
  assign n8250 = n7071 & n8249 ;
  assign n8251 = ~n4630 & n8250 ;
  assign n8252 = ~x6 & n6579 ;
  assign n8253 = x6 & n8252 ;
  assign n8254 = n332 & ~n8253 ;
  assign n8255 = n2066 & n8254 ;
  assign n8259 = n475 & n3270 ;
  assign n8260 = n382 & n8259 ;
  assign n8261 = n4368 | n8260 ;
  assign n8262 = n8261 ^ n1790 ^ 1'b0 ;
  assign n8263 = ~n2275 & n8262 ;
  assign n8264 = n8263 ^ n7540 ^ 1'b0 ;
  assign n8256 = x16 & n5538 ;
  assign n8257 = n8256 ^ n1229 ^ 1'b0 ;
  assign n8258 = n4403 | n8257 ;
  assign n8265 = n8264 ^ n8258 ^ 1'b0 ;
  assign n8266 = n3848 ^ n1279 ^ 1'b0 ;
  assign n8267 = n1878 & n8266 ;
  assign n8268 = ~n1340 & n8267 ;
  assign n8269 = n2297 | n8268 ;
  assign n8270 = n163 & n3221 ;
  assign n8271 = n8269 & n8270 ;
  assign n8272 = n6238 ^ n5836 ^ 1'b0 ;
  assign n8273 = n1625 & n8272 ;
  assign n8274 = n1553 ^ x126 ^ 1'b0 ;
  assign n8275 = x69 & n8274 ;
  assign n8276 = n8275 ^ n1344 ^ 1'b0 ;
  assign n8277 = n8276 ^ n6382 ^ 1'b0 ;
  assign n8278 = n4596 & n8277 ;
  assign n8279 = x44 & ~n789 ;
  assign n8280 = n8279 ^ n628 ^ 1'b0 ;
  assign n8281 = n7033 | n8280 ;
  assign n8282 = n1361 | n8281 ;
  assign n8283 = ~n701 & n8282 ;
  assign n8284 = n8283 ^ n2564 ^ 1'b0 ;
  assign n8285 = n8284 ^ x48 ^ 1'b0 ;
  assign n8286 = ~n172 & n4084 ;
  assign n8287 = n8286 ^ n3206 ^ 1'b0 ;
  assign n8288 = n5501 | n8249 ;
  assign n8289 = ~n726 & n7500 ;
  assign n8290 = ~n8288 & n8289 ;
  assign n8291 = x127 & n634 ;
  assign n8292 = n1064 & n8291 ;
  assign n8293 = n1881 | n8292 ;
  assign n8294 = ~n1271 & n3246 ;
  assign n8295 = ( n2046 & ~n2746 ) | ( n2046 & n3641 ) | ( ~n2746 & n3641 ) ;
  assign n8296 = n577 & n8295 ;
  assign n8297 = n8296 ^ n2645 ^ 1'b0 ;
  assign n8298 = n3701 ^ n2924 ^ 1'b0 ;
  assign n8299 = n6005 ^ n898 ^ 1'b0 ;
  assign n8300 = n2371 | n8299 ;
  assign n8301 = n8300 ^ n4661 ^ 1'b0 ;
  assign n8302 = n1903 & n2116 ;
  assign n8303 = n8302 ^ n4751 ^ n1092 ;
  assign n8305 = n1102 ^ n941 ^ 1'b0 ;
  assign n8306 = n3292 & ~n8305 ;
  assign n8307 = ~n1527 & n8306 ;
  assign n8308 = ~n2624 & n8307 ;
  assign n8304 = ~n1334 & n2730 ;
  assign n8309 = n8308 ^ n8304 ^ 1'b0 ;
  assign n8310 = n8309 ^ n421 ^ 1'b0 ;
  assign n8311 = n240 & n2583 ;
  assign n8312 = n8311 ^ n6165 ^ 1'b0 ;
  assign n8313 = n446 & ~n2670 ;
  assign n8314 = n8313 ^ n954 ^ 1'b0 ;
  assign n8315 = n519 & ~n1680 ;
  assign n8316 = n4206 & n8315 ;
  assign n8317 = n8314 & n8316 ;
  assign n8318 = n616 & ~n4507 ;
  assign n8319 = n8318 ^ n2176 ^ 1'b0 ;
  assign n8320 = n2445 & ~n2925 ;
  assign n8321 = n4872 & n8320 ;
  assign n8322 = ( ~n3224 & n3287 ) | ( ~n3224 & n5852 ) | ( n3287 & n5852 ) ;
  assign n8323 = n6662 | n8322 ;
  assign n8324 = ~n152 & n6493 ;
  assign n8325 = n2599 & n8324 ;
  assign n8326 = n7054 ^ n2234 ^ 1'b0 ;
  assign n8327 = n6479 & n8326 ;
  assign n8328 = n2985 ^ n2412 ^ n2009 ;
  assign n8329 = n425 | n3418 ;
  assign n8330 = n8329 ^ n4557 ^ 1'b0 ;
  assign n8331 = ( x75 & n6911 ) | ( x75 & ~n7245 ) | ( n6911 & ~n7245 ) ;
  assign n8332 = n3261 ^ n985 ^ 1'b0 ;
  assign n8333 = n784 & n8332 ;
  assign n8334 = x0 & n1174 ;
  assign n8335 = ~n163 & n8334 ;
  assign n8336 = n4841 & ~n5461 ;
  assign n8337 = n8335 & n8336 ;
  assign n8338 = ~n3470 & n6295 ;
  assign n8339 = ~n1790 & n8338 ;
  assign n8340 = n154 | n8339 ;
  assign n8341 = n395 & ~n8340 ;
  assign n8342 = n4419 ^ n2754 ^ 1'b0 ;
  assign n8343 = ( n866 & ~n3316 ) | ( n866 & n8342 ) | ( ~n3316 & n8342 ) ;
  assign n8344 = n8341 | n8343 ;
  assign n8345 = n4927 ^ n1793 ^ 1'b0 ;
  assign n8346 = ~n8344 & n8345 ;
  assign n8347 = n503 & ~n625 ;
  assign n8348 = n3460 & n8347 ;
  assign n8349 = n8348 ^ x3 ^ 1'b0 ;
  assign n8350 = n8349 ^ n3569 ^ 1'b0 ;
  assign n8351 = n7213 & n8350 ;
  assign n8352 = n2906 ^ n2053 ^ 1'b0 ;
  assign n8353 = n5231 ^ n1782 ^ 1'b0 ;
  assign n8354 = n3356 & ~n5958 ;
  assign n8355 = ~n7987 & n8354 ;
  assign n8356 = n4918 & ~n7085 ;
  assign n8357 = n8356 ^ n8074 ^ 1'b0 ;
  assign n8358 = ~n5807 & n7988 ;
  assign n8359 = x27 & ~n806 ;
  assign n8360 = n806 & n8359 ;
  assign n8361 = n5345 & ~n8360 ;
  assign n8362 = n2341 & n8361 ;
  assign n8363 = n1862 | n7238 ;
  assign n8364 = n8363 ^ n8317 ^ 1'b0 ;
  assign n8365 = n3746 | n8364 ;
  assign n8372 = n3039 ^ n2648 ^ 1'b0 ;
  assign n8373 = x11 & n8372 ;
  assign n8370 = n3385 ^ x69 ^ 1'b0 ;
  assign n8371 = n4370 | n8370 ;
  assign n8374 = n8373 ^ n8371 ^ 1'b0 ;
  assign n8375 = n456 | n8374 ;
  assign n8366 = n1134 & n4806 ;
  assign n8367 = n2086 & ~n3635 ;
  assign n8368 = n973 & n8367 ;
  assign n8369 = n8366 | n8368 ;
  assign n8376 = n8375 ^ n8369 ^ 1'b0 ;
  assign n8377 = n3894 & ~n6636 ;
  assign n8378 = n4155 ^ n3009 ^ 1'b0 ;
  assign n8379 = n3140 & ~n8378 ;
  assign n8380 = n8377 & n8379 ;
  assign n8381 = n8007 & n8380 ;
  assign n8383 = ~n1005 & n6214 ;
  assign n8382 = ~n2520 & n5958 ;
  assign n8384 = n8383 ^ n8382 ^ 1'b0 ;
  assign n8385 = n1579 & n1654 ;
  assign n8386 = n8385 ^ n894 ^ 1'b0 ;
  assign n8387 = n5836 ^ n290 ^ 1'b0 ;
  assign n8388 = n8386 | n8387 ;
  assign n8395 = ( n368 & ~n389 ) | ( n368 & n683 ) | ( ~n389 & n683 ) ;
  assign n8394 = ~n1077 & n1596 ;
  assign n8396 = n8395 ^ n8394 ^ n4071 ;
  assign n8389 = n1230 & n1576 ;
  assign n8390 = n6829 ^ n3147 ^ 1'b0 ;
  assign n8391 = ~n8389 & n8390 ;
  assign n8392 = ~x79 & n8391 ;
  assign n8393 = n6821 & n8392 ;
  assign n8397 = n8396 ^ n8393 ^ 1'b0 ;
  assign n8403 = x34 & n400 ;
  assign n8398 = n3963 & n7820 ;
  assign n8399 = n531 | n4190 ;
  assign n8400 = n8399 ^ n3306 ^ 1'b0 ;
  assign n8401 = n8398 | n8400 ;
  assign n8402 = n5928 | n8401 ;
  assign n8404 = n8403 ^ n8402 ^ 1'b0 ;
  assign n8405 = n3367 ^ n3126 ^ 1'b0 ;
  assign n8406 = ~n319 & n5516 ;
  assign n8407 = n8406 ^ n2702 ^ 1'b0 ;
  assign n8408 = n6148 ^ n3856 ^ 1'b0 ;
  assign n8409 = n2996 & ~n8408 ;
  assign n8410 = n8409 ^ n1268 ^ 1'b0 ;
  assign n8411 = n8410 ^ n8027 ^ 1'b0 ;
  assign n8412 = n6893 ^ n5787 ^ n699 ;
  assign n8413 = n894 ^ n751 ^ 1'b0 ;
  assign n8414 = n8413 ^ n4344 ^ 1'b0 ;
  assign n8415 = n1602 & ~n2300 ;
  assign n8416 = n2697 & n8415 ;
  assign n8417 = ~n472 & n6027 ;
  assign n8418 = n7763 & n8417 ;
  assign n8419 = n431 | n3278 ;
  assign n8420 = n8419 ^ n2561 ^ 1'b0 ;
  assign n8422 = ~n1602 & n2503 ;
  assign n8423 = n8422 ^ n4987 ^ n299 ;
  assign n8421 = n437 & ~n499 ;
  assign n8424 = n8423 ^ n8421 ^ 1'b0 ;
  assign n8425 = n423 & ~n2802 ;
  assign n8426 = n3179 ^ n3100 ^ 1'b0 ;
  assign n8427 = n4776 & ~n8426 ;
  assign n8428 = n3283 ^ x81 ^ 1'b0 ;
  assign n8429 = ~n1228 & n1856 ;
  assign n8430 = x47 & ~n8429 ;
  assign n8431 = n8430 ^ n825 ^ 1'b0 ;
  assign n8432 = ( ~n3861 & n8428 ) | ( ~n3861 & n8431 ) | ( n8428 & n8431 ) ;
  assign n8433 = n3574 ^ n359 ^ 1'b0 ;
  assign n8434 = ~n7187 & n8433 ;
  assign n8435 = n8434 ^ n4902 ^ 1'b0 ;
  assign n8436 = n4183 & n7281 ;
  assign n8437 = n3270 | n8436 ;
  assign n8438 = n6382 ^ n4018 ^ 1'b0 ;
  assign n8439 = n1186 & n3215 ;
  assign n8440 = ( ~n1233 & n4380 ) | ( ~n1233 & n8439 ) | ( n4380 & n8439 ) ;
  assign n8441 = n5549 | n8440 ;
  assign n8442 = n8438 & ~n8441 ;
  assign n8443 = n1496 ^ n1053 ^ n754 ;
  assign n8444 = ( n6827 & n7163 ) | ( n6827 & ~n8443 ) | ( n7163 & ~n8443 ) ;
  assign n8445 = n8444 ^ n2054 ^ 1'b0 ;
  assign n8446 = n1943 & n6207 ;
  assign n8447 = n6751 ^ n305 ^ 1'b0 ;
  assign n8448 = n6538 & ~n8447 ;
  assign n8449 = n3251 ^ n1500 ^ n209 ;
  assign n8450 = n7997 | n8449 ;
  assign n8451 = n7734 & ~n8450 ;
  assign n8452 = n6318 ^ n5547 ^ 1'b0 ;
  assign n8453 = n489 & n5033 ;
  assign n8454 = n8453 ^ n1150 ^ 1'b0 ;
  assign n8455 = n8452 & n8454 ;
  assign n8456 = n8455 ^ x23 ^ 1'b0 ;
  assign n8457 = ~n1741 & n3140 ;
  assign n8458 = n6292 & ~n8457 ;
  assign n8459 = ~n732 & n993 ;
  assign n8460 = n8459 ^ n2621 ^ 1'b0 ;
  assign n8461 = ~n6587 & n8460 ;
  assign n8462 = n4727 & n8461 ;
  assign n8463 = n5613 & ~n6261 ;
  assign n8464 = ~n8306 & n8463 ;
  assign n8465 = n6964 | n8464 ;
  assign n8466 = n8462 & ~n8465 ;
  assign n8467 = n7345 ^ n7221 ^ 1'b0 ;
  assign n8468 = ~n588 & n8467 ;
  assign n8469 = n3689 ^ n371 ^ 1'b0 ;
  assign n8470 = ~n5832 & n6159 ;
  assign n8471 = n8470 ^ n1241 ^ 1'b0 ;
  assign n8472 = n4325 & n5281 ;
  assign n8474 = n3655 ^ n1960 ^ 1'b0 ;
  assign n8475 = n4011 & ~n8474 ;
  assign n8473 = n1252 & n6538 ;
  assign n8476 = n8475 ^ n8473 ^ 1'b0 ;
  assign n8477 = n1713 | n8476 ;
  assign n8478 = n6233 ^ n3391 ^ 1'b0 ;
  assign n8479 = n1062 & n8478 ;
  assign n8480 = n8477 & n8479 ;
  assign n8481 = ~n1962 & n8480 ;
  assign n8482 = ( n3006 & n3458 ) | ( n3006 & ~n8045 ) | ( n3458 & ~n8045 ) ;
  assign n8483 = n4578 ^ n1556 ^ 1'b0 ;
  assign n8484 = n3389 | n6189 ;
  assign n8485 = n3188 & ~n8484 ;
  assign n8486 = ~n4800 & n8485 ;
  assign n8487 = n6080 ^ n2180 ^ 1'b0 ;
  assign n8488 = n1470 & n4859 ;
  assign n8489 = n8264 & n8488 ;
  assign n8490 = n1951 & n5571 ;
  assign n8491 = n3479 & n6734 ;
  assign n8492 = n3255 & n5207 ;
  assign n8493 = ~n2222 & n8492 ;
  assign n8494 = ~n3084 & n8493 ;
  assign n8495 = n1658 & n8494 ;
  assign n8496 = x102 & ~n2998 ;
  assign n8497 = n3797 | n8496 ;
  assign n8498 = n6027 | n8497 ;
  assign n8499 = n6490 ^ n3333 ^ 1'b0 ;
  assign n8500 = ~n2204 & n3729 ;
  assign n8501 = ( ~n493 & n4447 ) | ( ~n493 & n8500 ) | ( n4447 & n8500 ) ;
  assign n8502 = n1133 & n5974 ;
  assign n8503 = n8502 ^ n1204 ^ 1'b0 ;
  assign n8504 = n2861 & ~n3582 ;
  assign n8505 = n8295 & ~n8504 ;
  assign n8506 = n8505 ^ n3866 ^ 1'b0 ;
  assign n8509 = x6 & n1878 ;
  assign n8507 = n7597 ^ n4021 ^ 1'b0 ;
  assign n8508 = ~n2283 & n8507 ;
  assign n8510 = n8509 ^ n8508 ^ 1'b0 ;
  assign n8511 = n5792 ^ n5015 ^ 1'b0 ;
  assign n8512 = n7678 & n8511 ;
  assign n8513 = n4700 & n6030 ;
  assign n8514 = x24 & ~n1223 ;
  assign n8516 = n2673 ^ n1620 ^ 1'b0 ;
  assign n8517 = n3558 | n8516 ;
  assign n8515 = ~n1909 & n2854 ;
  assign n8518 = n8517 ^ n8515 ^ 1'b0 ;
  assign n8519 = n1112 & n3269 ;
  assign n8520 = n8519 ^ n1128 ^ 1'b0 ;
  assign n8521 = n7753 & n8520 ;
  assign n8522 = ( n330 & n1088 ) | ( n330 & n5834 ) | ( n1088 & n5834 ) ;
  assign n8523 = n2510 & ~n4910 ;
  assign n8524 = n8523 ^ n1658 ^ 1'b0 ;
  assign n8525 = n8469 ^ n3120 ^ 1'b0 ;
  assign n8526 = n5459 ^ n1051 ^ 1'b0 ;
  assign n8527 = n6334 | n8526 ;
  assign n8529 = n1024 & n2515 ;
  assign n8528 = n362 & n6118 ;
  assign n8530 = n8529 ^ n8528 ^ 1'b0 ;
  assign n8531 = ( n7118 & ~n8527 ) | ( n7118 & n8530 ) | ( ~n8527 & n8530 ) ;
  assign n8532 = n1920 ^ n1031 ^ 1'b0 ;
  assign n8533 = n5434 ^ n1792 ^ 1'b0 ;
  assign n8534 = n1674 & ~n8533 ;
  assign n8535 = ~n8532 & n8534 ;
  assign n8536 = n728 | n8535 ;
  assign n8537 = n8059 & ~n8536 ;
  assign n8538 = n3424 & n3806 ;
  assign n8539 = n8538 ^ n2302 ^ 1'b0 ;
  assign n8547 = n172 & n4025 ;
  assign n8540 = n5664 ^ n2839 ^ 1'b0 ;
  assign n8541 = x101 & n8540 ;
  assign n8542 = ~n3405 & n8541 ;
  assign n8543 = n8542 ^ n2515 ^ 1'b0 ;
  assign n8544 = n4423 & ~n8543 ;
  assign n8545 = ~n645 & n8544 ;
  assign n8546 = n2758 & ~n8545 ;
  assign n8548 = n8547 ^ n8546 ^ 1'b0 ;
  assign n8549 = ~n3868 & n6088 ;
  assign n8550 = n8549 ^ n2102 ^ 1'b0 ;
  assign n8551 = n3348 ^ n2935 ^ 1'b0 ;
  assign n8552 = n3978 & ~n8551 ;
  assign n8553 = n3460 ^ n2486 ^ 1'b0 ;
  assign n8554 = ( n2394 & n5487 ) | ( n2394 & ~n8553 ) | ( n5487 & ~n8553 ) ;
  assign n8555 = ~n3166 & n8443 ;
  assign n8556 = ( n2071 & n4182 ) | ( n2071 & n8555 ) | ( n4182 & n8555 ) ;
  assign n8557 = ~n2558 & n3574 ;
  assign n8558 = n5590 & n8557 ;
  assign n8559 = n6753 & ~n8558 ;
  assign n8560 = n3062 & n8559 ;
  assign n8561 = ~n1444 & n8560 ;
  assign n8562 = n1295 | n4908 ;
  assign n8563 = n1454 | n1649 ;
  assign n8564 = n1511 & ~n8563 ;
  assign n8565 = n8564 ^ n1588 ^ 1'b0 ;
  assign n8566 = n8565 ^ n7090 ^ n6547 ;
  assign n8567 = n1296 | n2433 ;
  assign n8568 = n4923 ^ n4876 ^ 1'b0 ;
  assign n8569 = x75 & n6044 ;
  assign n8570 = n7425 ^ x4 ^ 1'b0 ;
  assign n8571 = ~n8569 & n8570 ;
  assign n8580 = n2416 & ~n6720 ;
  assign n8572 = n3894 ^ x54 ^ 1'b0 ;
  assign n8573 = ~n1229 & n8572 ;
  assign n8574 = ~n640 & n8573 ;
  assign n8575 = ( ~n4733 & n5120 ) | ( ~n4733 & n8043 ) | ( n5120 & n8043 ) ;
  assign n8576 = n1134 ^ n1105 ^ 1'b0 ;
  assign n8577 = ~n6929 & n8576 ;
  assign n8578 = ( n287 & n8575 ) | ( n287 & ~n8577 ) | ( n8575 & ~n8577 ) ;
  assign n8579 = ~n8574 & n8578 ;
  assign n8581 = n8580 ^ n8579 ^ 1'b0 ;
  assign n8582 = n8171 ^ n708 ^ 1'b0 ;
  assign n8583 = n4416 ^ n311 ^ 1'b0 ;
  assign n8584 = n8583 ^ n6614 ^ 1'b0 ;
  assign n8585 = n186 | n2330 ;
  assign n8586 = n755 | n4616 ;
  assign n8587 = n8586 ^ n637 ^ 1'b0 ;
  assign n8588 = n5637 ^ n1769 ^ 1'b0 ;
  assign n8589 = n5647 & n5872 ;
  assign n8590 = n8588 & n8589 ;
  assign n8591 = ~n1469 & n7171 ;
  assign n8592 = n8590 & n8591 ;
  assign n8593 = n1510 ^ n539 ^ 1'b0 ;
  assign n8594 = n3326 & ~n5955 ;
  assign n8595 = x74 & ~n2521 ;
  assign n8596 = n1865 | n2978 ;
  assign n8597 = n8595 & ~n8596 ;
  assign n8598 = n5067 & ~n8597 ;
  assign n8599 = n4921 ^ n797 ^ 1'b0 ;
  assign n8600 = n8599 ^ n1973 ^ 1'b0 ;
  assign n8601 = n634 & n8600 ;
  assign n8602 = n4771 & n8601 ;
  assign n8603 = n3179 | n4398 ;
  assign n8604 = n8603 ^ n4176 ^ 1'b0 ;
  assign n8605 = n8604 ^ n5083 ^ n1816 ;
  assign n8608 = n789 | n2436 ;
  assign n8609 = n3288 & ~n8608 ;
  assign n8610 = n1491 & n8609 ;
  assign n8606 = n4195 ^ n468 ^ 1'b0 ;
  assign n8607 = ~n1215 & n8606 ;
  assign n8611 = n8610 ^ n8607 ^ n308 ;
  assign n8612 = ~n5294 & n5564 ;
  assign n8613 = n4747 & n8612 ;
  assign n8614 = n8062 & ~n8613 ;
  assign n8615 = ~n4843 & n8614 ;
  assign n8616 = n5551 ^ n5402 ^ 1'b0 ;
  assign n8617 = n3824 & ~n8616 ;
  assign n8618 = n4013 & ~n4779 ;
  assign n8619 = n8618 ^ n5860 ^ 1'b0 ;
  assign n8620 = n8619 ^ n1553 ^ 1'b0 ;
  assign n8621 = n8236 ^ n2010 ^ 1'b0 ;
  assign n8622 = n8620 & ~n8621 ;
  assign n8623 = n2130 | n8622 ;
  assign n8624 = n8623 ^ n8429 ^ 1'b0 ;
  assign n8625 = n8617 & n8624 ;
  assign n8626 = n2639 | n8231 ;
  assign n8627 = n8626 ^ n2433 ^ 1'b0 ;
  assign n8628 = n815 & ~n8466 ;
  assign n8629 = x69 & ~n6352 ;
  assign n8630 = ~n1271 & n8629 ;
  assign n8631 = n8630 ^ n5434 ^ 1'b0 ;
  assign n8632 = n4856 & n8631 ;
  assign n8633 = ~n1805 & n6323 ;
  assign n8634 = n6827 ^ n6434 ^ n3356 ;
  assign n8635 = n3597 ^ n3210 ^ 1'b0 ;
  assign n8636 = ~n695 & n8635 ;
  assign n8637 = n8634 & n8636 ;
  assign n8638 = n5523 ^ n5014 ^ 1'b0 ;
  assign n8639 = ~n977 & n4064 ;
  assign n8640 = n4073 & n5064 ;
  assign n8641 = n8640 ^ n1132 ^ 1'b0 ;
  assign n8642 = n6382 ^ x54 ^ 1'b0 ;
  assign n8643 = n1681 | n8642 ;
  assign n8644 = n8641 | n8643 ;
  assign n8645 = n2948 ^ x20 ^ 1'b0 ;
  assign n8646 = n8645 ^ n632 ^ 1'b0 ;
  assign n8647 = n2396 ^ n362 ^ 1'b0 ;
  assign n8648 = n166 | n8647 ;
  assign n8649 = n530 & n1399 ;
  assign n8650 = ~n234 & n8649 ;
  assign n8651 = n8650 ^ n5992 ^ 1'b0 ;
  assign n8655 = n2243 & n5530 ;
  assign n8656 = ~n733 & n8655 ;
  assign n8652 = n3700 ^ n1244 ^ 1'b0 ;
  assign n8653 = n7264 & n8652 ;
  assign n8654 = n8653 ^ n3393 ^ 1'b0 ;
  assign n8657 = n8656 ^ n8654 ^ n3903 ;
  assign n8658 = n3204 ^ n1927 ^ 1'b0 ;
  assign n8659 = n6448 & ~n8658 ;
  assign n8660 = n628 & ~n1643 ;
  assign n8661 = n8660 ^ n4973 ^ 1'b0 ;
  assign n8662 = n5701 | n8661 ;
  assign n8663 = n8662 ^ n855 ^ 1'b0 ;
  assign n8664 = ~n2138 & n8663 ;
  assign n8665 = n8377 ^ n4707 ^ 1'b0 ;
  assign n8666 = n2124 & n8665 ;
  assign n8667 = n3752 | n6613 ;
  assign n8668 = n2525 & ~n8667 ;
  assign n8669 = n607 | n1346 ;
  assign n8670 = ~n1129 & n1170 ;
  assign n8671 = ~n1710 & n8670 ;
  assign n8672 = n7237 ^ n5236 ^ 1'b0 ;
  assign n8673 = ~n852 & n8672 ;
  assign n8674 = ~n8671 & n8673 ;
  assign n8675 = n5988 & ~n8128 ;
  assign n8676 = n7861 & n8675 ;
  assign n8677 = n3524 | n6191 ;
  assign n8678 = n930 & n6411 ;
  assign n8679 = ~n8677 & n8678 ;
  assign n8680 = ( n1129 & n4678 ) | ( n1129 & n8679 ) | ( n4678 & n8679 ) ;
  assign n8681 = n4960 ^ n1987 ^ 1'b0 ;
  assign n8682 = n8377 & n8681 ;
  assign n8683 = n3400 & ~n5610 ;
  assign n8684 = ~n3068 & n8683 ;
  assign n8685 = n8684 ^ n2529 ^ 1'b0 ;
  assign n8686 = ~n4186 & n8685 ;
  assign n8687 = ~n699 & n1967 ;
  assign n8688 = n6700 | n8687 ;
  assign n8696 = n7114 ^ n4204 ^ 1'b0 ;
  assign n8689 = n469 & n1540 ;
  assign n8690 = ~n257 & n1891 ;
  assign n8691 = n8690 ^ n3138 ^ 1'b0 ;
  assign n8692 = ~n1830 & n8691 ;
  assign n8693 = ~n8689 & n8692 ;
  assign n8694 = n6242 | n8693 ;
  assign n8695 = n1546 & ~n8694 ;
  assign n8697 = n8696 ^ n8695 ^ n7811 ;
  assign n8699 = n2107 | n7483 ;
  assign n8698 = n4796 | n6759 ;
  assign n8700 = n8699 ^ n8698 ^ 1'b0 ;
  assign n8701 = n2421 ^ n2231 ^ 1'b0 ;
  assign n8702 = ~n4969 & n8701 ;
  assign n8703 = n1281 ^ n313 ^ 1'b0 ;
  assign n8704 = n4428 ^ n697 ^ 1'b0 ;
  assign n8705 = ( n5797 & ~n8703 ) | ( n5797 & n8704 ) | ( ~n8703 & n8704 ) ;
  assign n8706 = n3498 & n3910 ;
  assign n8707 = n1553 & n1945 ;
  assign n8708 = n8706 | n8707 ;
  assign n8709 = x4 & ~n8708 ;
  assign n8710 = n1770 ^ n1279 ^ 1'b0 ;
  assign n8711 = n542 & n8710 ;
  assign n8712 = ( ~n551 & n4231 ) | ( ~n551 & n7820 ) | ( n4231 & n7820 ) ;
  assign n8713 = ( ~n2187 & n6708 ) | ( ~n2187 & n8712 ) | ( n6708 & n8712 ) ;
  assign n8714 = x23 & n1687 ;
  assign n8715 = n8714 ^ n1697 ^ 1'b0 ;
  assign n8716 = n8713 & n8715 ;
  assign n8718 = ( n729 & n5486 ) | ( n729 & ~n5811 ) | ( n5486 & ~n5811 ) ;
  assign n8717 = n3472 & n4467 ;
  assign n8719 = n8718 ^ n8717 ^ 1'b0 ;
  assign n8720 = n3630 ^ n1337 ^ n905 ;
  assign n8721 = n557 & ~n8720 ;
  assign n8722 = n8721 ^ n1500 ^ 1'b0 ;
  assign n8723 = n313 | n8722 ;
  assign n8724 = n8723 ^ n6126 ^ 1'b0 ;
  assign n8725 = n8719 & n8724 ;
  assign n8726 = n4019 & n5403 ;
  assign n8727 = n6415 ^ n6082 ^ 1'b0 ;
  assign n8728 = n3953 | n8727 ;
  assign n8729 = ~n1518 & n6227 ;
  assign n8730 = n2912 & n8729 ;
  assign n8731 = n3982 & ~n8730 ;
  assign n8732 = n8731 ^ n4771 ^ 1'b0 ;
  assign n8733 = n2487 | n8732 ;
  assign n8734 = n3950 & ~n8733 ;
  assign n8735 = n8734 ^ n1496 ^ 1'b0 ;
  assign n8736 = n2013 ^ n290 ^ 1'b0 ;
  assign n8737 = x52 & n8736 ;
  assign n8738 = n4972 ^ n1605 ^ 1'b0 ;
  assign n8739 = n8738 ^ n6207 ^ 1'b0 ;
  assign n8740 = ( ~n1847 & n2053 ) | ( ~n1847 & n6438 ) | ( n2053 & n6438 ) ;
  assign n8741 = n8740 ^ n490 ^ 1'b0 ;
  assign n8742 = n2622 & ~n2800 ;
  assign n8743 = ~n2123 & n4678 ;
  assign n8744 = n2096 & n8743 ;
  assign n8745 = n8267 ^ n4938 ^ 1'b0 ;
  assign n8746 = n4244 & ~n8745 ;
  assign n8747 = ( n2483 & ~n3990 ) | ( n2483 & n8746 ) | ( ~n3990 & n8746 ) ;
  assign n8748 = ~n1467 & n2515 ;
  assign n8749 = n8748 ^ n3404 ^ 1'b0 ;
  assign n8750 = n8749 ^ n7143 ^ 1'b0 ;
  assign n8751 = n8385 ^ n5028 ^ 1'b0 ;
  assign n8752 = ~n243 & n8751 ;
  assign n8753 = n2288 & n8752 ;
  assign n8754 = n673 & n1313 ;
  assign n8755 = n8754 ^ n5245 ^ 1'b0 ;
  assign n8756 = n2451 & n8755 ;
  assign n8757 = n7028 ^ n217 ^ 1'b0 ;
  assign n8758 = n1003 | n8757 ;
  assign n8761 = n1620 | n4216 ;
  assign n8762 = n8761 ^ n687 ^ 1'b0 ;
  assign n8763 = n4389 ^ n4175 ^ 1'b0 ;
  assign n8764 = n8762 | n8763 ;
  assign n8759 = n6112 | n7504 ;
  assign n8760 = n3032 & ~n8759 ;
  assign n8765 = n8764 ^ n8760 ^ 1'b0 ;
  assign n8766 = ~n6901 & n8765 ;
  assign n8767 = n5111 | n7367 ;
  assign n8768 = n844 & ~n3415 ;
  assign n8769 = n1394 & n4490 ;
  assign n8770 = x1 & n8769 ;
  assign n8771 = n2153 | n8770 ;
  assign n8772 = n8768 | n8771 ;
  assign n8773 = n1047 & ~n8772 ;
  assign n8774 = x34 & n2413 ;
  assign n8775 = ~n3687 & n8774 ;
  assign n8776 = ~n7412 & n8775 ;
  assign n8778 = n4921 ^ n4738 ^ 1'b0 ;
  assign n8779 = ~n2723 & n8778 ;
  assign n8780 = n7012 | n8779 ;
  assign n8777 = n2466 & n8746 ;
  assign n8781 = n8780 ^ n8777 ^ 1'b0 ;
  assign n8782 = n1370 ^ x100 ^ 1'b0 ;
  assign n8783 = n1999 & n8782 ;
  assign n8784 = n8783 ^ n3039 ^ 1'b0 ;
  assign n8785 = n8784 ^ n741 ^ 1'b0 ;
  assign n8786 = ~n4688 & n8785 ;
  assign n8787 = ( ~n4477 & n6155 ) | ( ~n4477 & n8786 ) | ( n6155 & n8786 ) ;
  assign n8788 = n1469 & ~n6211 ;
  assign n8789 = ~n1621 & n7071 ;
  assign n8790 = n505 & ~n745 ;
  assign n8791 = n1169 & n8790 ;
  assign n8792 = n8791 ^ n2694 ^ 1'b0 ;
  assign n8793 = n3800 & n8792 ;
  assign n8794 = n8630 & n8793 ;
  assign n8795 = n1348 & ~n3495 ;
  assign n8796 = n8656 ^ n1247 ^ 1'b0 ;
  assign n8797 = ~n1587 & n8796 ;
  assign n8798 = x46 & ~n243 ;
  assign n8799 = ~n1259 & n8798 ;
  assign n8800 = n8799 ^ n3395 ^ n1225 ;
  assign n8801 = n8800 ^ n2191 ^ 1'b0 ;
  assign n8802 = ( n4723 & n8797 ) | ( n4723 & n8801 ) | ( n8797 & n8801 ) ;
  assign n8803 = ~n1176 & n1370 ;
  assign n8804 = n3119 ^ n411 ^ 1'b0 ;
  assign n8805 = n7666 | n8804 ;
  assign n8806 = ~n1261 & n7052 ;
  assign n8807 = ~n513 & n8806 ;
  assign n8808 = ( n5653 & n5732 ) | ( n5653 & n8195 ) | ( n5732 & n8195 ) ;
  assign n8809 = ~n1641 & n4802 ;
  assign n8810 = n4310 ^ n3272 ^ n2376 ;
  assign n8811 = n1776 & n8810 ;
  assign n8812 = n8811 ^ n5995 ^ 1'b0 ;
  assign n8813 = n2198 & ~n8643 ;
  assign n8814 = ( n2731 & n5236 ) | ( n2731 & n7371 ) | ( n5236 & n7371 ) ;
  assign n8815 = ~n3711 & n4452 ;
  assign n8816 = n484 & n1993 ;
  assign n8817 = n3625 ^ n1908 ^ x103 ;
  assign n8818 = n666 | n2687 ;
  assign n8819 = n8818 ^ n2656 ^ 1'b0 ;
  assign n8820 = ( n8816 & n8817 ) | ( n8816 & n8819 ) | ( n8817 & n8819 ) ;
  assign n8821 = n1342 ^ n719 ^ 1'b0 ;
  assign n8822 = n3968 & ~n4183 ;
  assign n8823 = n1008 & n8822 ;
  assign n8824 = n3848 | n8823 ;
  assign n8825 = n1594 ^ n992 ^ 1'b0 ;
  assign n8826 = ~n1479 & n8825 ;
  assign n8827 = ~n658 & n8826 ;
  assign n8828 = n8827 ^ n2772 ^ n799 ;
  assign n8829 = n3586 ^ n1761 ^ 1'b0 ;
  assign n8830 = n737 & ~n2448 ;
  assign n8831 = n8830 ^ n5345 ^ 1'b0 ;
  assign n8832 = n8829 & ~n8831 ;
  assign n8833 = n437 | n7241 ;
  assign n8834 = ~n5429 & n8833 ;
  assign n8835 = ~n5410 & n8834 ;
  assign n8836 = n8543 ^ n4605 ^ 1'b0 ;
  assign n8837 = n709 | n7483 ;
  assign n8838 = n1979 ^ n674 ^ 1'b0 ;
  assign n8839 = n2568 | n4484 ;
  assign n8840 = n8839 ^ n1217 ^ 1'b0 ;
  assign n8841 = n8838 & n8840 ;
  assign n8842 = n8841 ^ n2445 ^ 1'b0 ;
  assign n8843 = n8142 ^ n4793 ^ 1'b0 ;
  assign n8844 = n1750 & ~n3266 ;
  assign n8845 = n8844 ^ n2835 ^ 1'b0 ;
  assign n8846 = n8845 ^ n8066 ^ 1'b0 ;
  assign n8847 = n6555 ^ n4870 ^ 1'b0 ;
  assign n8848 = n8846 & n8847 ;
  assign n8849 = n2802 | n5326 ;
  assign n8850 = n2566 ^ n792 ^ 1'b0 ;
  assign n8851 = n4303 ^ n3818 ^ 1'b0 ;
  assign n8852 = n8850 | n8851 ;
  assign n8853 = n556 ^ n296 ^ 1'b0 ;
  assign n8854 = n559 & ~n8431 ;
  assign n8855 = ( ~n4105 & n6529 ) | ( ~n4105 & n8854 ) | ( n6529 & n8854 ) ;
  assign n8856 = n8853 | n8855 ;
  assign n8857 = n1049 & ~n1929 ;
  assign n8858 = n455 & n8857 ;
  assign n8859 = n4045 & n8858 ;
  assign n8860 = ~n2046 & n2889 ;
  assign n8862 = n3009 ^ n1123 ^ n741 ;
  assign n8863 = n8862 ^ n6680 ^ 1'b0 ;
  assign n8864 = n7955 & ~n8863 ;
  assign n8861 = n4315 & n8101 ;
  assign n8865 = n8864 ^ n8861 ^ 1'b0 ;
  assign n8866 = n266 | n6979 ;
  assign n8867 = ( n2131 & n3369 ) | ( n2131 & ~n8718 ) | ( n3369 & ~n8718 ) ;
  assign n8868 = ( n496 & n2788 ) | ( n496 & ~n2976 ) | ( n2788 & ~n2976 ) ;
  assign n8869 = n8868 ^ n4132 ^ n3532 ;
  assign n8870 = n2255 & n4662 ;
  assign n8871 = n8869 & n8870 ;
  assign n8872 = n2681 | n8871 ;
  assign n8873 = n7527 | n8872 ;
  assign n8874 = n8873 ^ n423 ^ 1'b0 ;
  assign n8875 = ~n3027 & n3492 ;
  assign n8876 = ~n5031 & n8875 ;
  assign n8877 = ~n2470 & n5997 ;
  assign n8878 = n435 & ~n754 ;
  assign n8879 = n8349 ^ n6242 ^ 1'b0 ;
  assign n8880 = n8878 & n8879 ;
  assign n8881 = ~n6597 & n8880 ;
  assign n8882 = ( n1129 & n3303 ) | ( n1129 & ~n3921 ) | ( n3303 & ~n3921 ) ;
  assign n8883 = n8881 & ~n8882 ;
  assign n8884 = n3334 & n6097 ;
  assign n8885 = n8884 ^ n2000 ^ 1'b0 ;
  assign n8886 = n3350 & ~n6950 ;
  assign n8887 = ~n2262 & n2720 ;
  assign n8888 = n7007 ^ n404 ^ 1'b0 ;
  assign n8889 = n2405 & n4336 ;
  assign n8890 = ~n1411 & n4237 ;
  assign n8891 = n1510 ^ n1117 ^ 1'b0 ;
  assign n8892 = n6669 ^ n5289 ^ 1'b0 ;
  assign n8893 = ~n8891 & n8892 ;
  assign n8894 = ~n2462 & n3918 ;
  assign n8895 = n3614 & n8894 ;
  assign n8896 = n7368 ^ n4024 ^ 1'b0 ;
  assign n8897 = ~n3376 & n8896 ;
  assign n8898 = ~n7375 & n8638 ;
  assign n8899 = n3229 ^ n1060 ^ n648 ;
  assign n8900 = n8899 ^ n5423 ^ 1'b0 ;
  assign n8901 = ~n7245 & n8900 ;
  assign n8902 = ~n6661 & n8901 ;
  assign n8903 = n4013 ^ n2006 ^ n1056 ;
  assign n8904 = n8903 ^ n692 ^ 1'b0 ;
  assign n8905 = n3623 & n6493 ;
  assign n8906 = ~n8904 & n8905 ;
  assign n8907 = n796 | n3204 ;
  assign n8908 = n8907 ^ n4141 ^ 1'b0 ;
  assign n8909 = n8908 ^ n8384 ^ 1'b0 ;
  assign n8910 = ( n391 & ~n545 ) | ( n391 & n2533 ) | ( ~n545 & n2533 ) ;
  assign n8911 = n172 & ~n458 ;
  assign n8912 = n8911 ^ n1128 ^ 1'b0 ;
  assign n8913 = n8910 & n8912 ;
  assign n8914 = n8913 ^ n8784 ^ n7408 ;
  assign n8915 = n8914 ^ n3709 ^ 1'b0 ;
  assign n8916 = n1758 ^ x19 ^ 1'b0 ;
  assign n8917 = n4738 & n5620 ;
  assign n8918 = ~n969 & n8917 ;
  assign n8919 = n7743 & ~n8918 ;
  assign n8921 = n4056 | n8002 ;
  assign n8922 = n8921 ^ n2687 ^ 1'b0 ;
  assign n8923 = n196 | n8922 ;
  assign n8920 = n3595 ^ n1257 ^ 1'b0 ;
  assign n8924 = n8923 ^ n8920 ^ 1'b0 ;
  assign n8925 = ~n3460 & n8924 ;
  assign n8926 = ~n7271 & n8925 ;
  assign n8927 = n1615 | n4255 ;
  assign n8928 = n8927 ^ n808 ^ 1'b0 ;
  assign n8929 = n860 & ~n8837 ;
  assign n8930 = n1359 & n4624 ;
  assign n8931 = ~n6907 & n8930 ;
  assign n8932 = n3565 & ~n6967 ;
  assign n8933 = ~n2412 & n6295 ;
  assign n8934 = ~n5390 & n8933 ;
  assign n8935 = n3278 ^ n1523 ^ 1'b0 ;
  assign n8936 = n2763 & n4448 ;
  assign n8937 = n1733 & n8936 ;
  assign n8938 = n8935 & n8937 ;
  assign n8939 = n3186 & n5953 ;
  assign n8940 = n1926 & n8939 ;
  assign n8941 = n1638 ^ n1285 ^ 1'b0 ;
  assign n8942 = ~n5556 & n8941 ;
  assign n8943 = n2668 & ~n8942 ;
  assign n8944 = n5863 & n8943 ;
  assign n8945 = n8944 ^ n519 ^ 1'b0 ;
  assign n8946 = x104 & ~n1033 ;
  assign n8947 = n2508 ^ n2098 ^ n1138 ;
  assign n8948 = ( n2759 & ~n4285 ) | ( n2759 & n4919 ) | ( ~n4285 & n4919 ) ;
  assign n8949 = n8947 | n8948 ;
  assign n8950 = n8946 & ~n8949 ;
  assign n8951 = n4377 & ~n4927 ;
  assign n8952 = ( ~n1132 & n5747 ) | ( ~n1132 & n7131 ) | ( n5747 & n7131 ) ;
  assign n8953 = ~n1064 & n2829 ;
  assign n8954 = ~n4578 & n8953 ;
  assign n8955 = n8872 & ~n8954 ;
  assign n8956 = n8955 ^ n6095 ^ 1'b0 ;
  assign n8957 = n3696 ^ n3222 ^ 1'b0 ;
  assign n8958 = n810 & n8957 ;
  assign n8959 = ~n1115 & n7646 ;
  assign n8960 = n1948 & ~n8959 ;
  assign n8961 = ~n138 & n1365 ;
  assign n8962 = n8961 ^ n560 ^ 1'b0 ;
  assign n8963 = n4927 & ~n8962 ;
  assign n8964 = ~n2150 & n8963 ;
  assign n8965 = n2088 & ~n7678 ;
  assign n8966 = n8965 ^ n2160 ^ 1'b0 ;
  assign n8967 = n8966 ^ n6532 ^ 1'b0 ;
  assign n8968 = n2445 & n8967 ;
  assign n8969 = n5305 ^ n3336 ^ 1'b0 ;
  assign n8970 = n6252 ^ n4355 ^ 1'b0 ;
  assign n8971 = ~n6323 & n6339 ;
  assign n8972 = n1719 ^ n1077 ^ 1'b0 ;
  assign n8973 = ~n3508 & n8972 ;
  assign n8974 = n8973 ^ n6634 ^ 1'b0 ;
  assign n8975 = n4423 ^ n3039 ^ 1'b0 ;
  assign n8976 = n1567 & n8975 ;
  assign n8977 = n5297 & n8976 ;
  assign n8978 = n8974 & n8977 ;
  assign n8979 = n6708 ^ n1120 ^ 1'b0 ;
  assign n8980 = n4516 ^ n2170 ^ 1'b0 ;
  assign n8981 = n8980 ^ n6188 ^ 1'b0 ;
  assign n8982 = n231 & ~n8981 ;
  assign n8983 = ~n4753 & n8982 ;
  assign n8984 = n8983 ^ n901 ^ 1'b0 ;
  assign n8985 = ( n3625 & n4729 ) | ( n3625 & ~n5978 ) | ( n4729 & ~n5978 ) ;
  assign n8987 = ~n2911 & n3592 ;
  assign n8986 = ~n2413 & n2886 ;
  assign n8988 = n8987 ^ n8986 ^ n7289 ;
  assign n8989 = n3067 ^ n459 ^ 1'b0 ;
  assign n8990 = n8989 ^ n6858 ^ 1'b0 ;
  assign n8991 = n8990 ^ n4139 ^ 1'b0 ;
  assign n8992 = ~n147 & n4576 ;
  assign n8993 = n6821 ^ n3408 ^ 1'b0 ;
  assign n8994 = n8993 ^ n7348 ^ 1'b0 ;
  assign n8995 = n7308 & ~n8994 ;
  assign n8996 = n4344 ^ x118 ^ 1'b0 ;
  assign n8997 = n3429 & n8996 ;
  assign n8998 = n8997 ^ n3540 ^ 1'b0 ;
  assign n8999 = n7420 | n8998 ;
  assign n9000 = n494 | n8999 ;
  assign n9001 = n9000 ^ n8413 ^ n6721 ;
  assign n9002 = ~n2170 & n2289 ;
  assign n9003 = ~n1189 & n9002 ;
  assign n9004 = n9003 ^ n8689 ^ n6423 ;
  assign n9005 = n8490 ^ n3714 ^ 1'b0 ;
  assign n9006 = n6127 ^ n1070 ^ 1'b0 ;
  assign n9010 = x35 & n838 ;
  assign n9011 = ~n3364 & n9010 ;
  assign n9008 = n147 ^ x6 ^ 1'b0 ;
  assign n9007 = n368 | n2777 ;
  assign n9009 = n9008 ^ n9007 ^ 1'b0 ;
  assign n9012 = n9011 ^ n9009 ^ n1603 ;
  assign n9013 = n4206 | n5997 ;
  assign n9014 = n9013 ^ n7956 ^ 1'b0 ;
  assign n9015 = n1444 & ~n9014 ;
  assign n9016 = n2412 & n9015 ;
  assign n9017 = n1799 & ~n3653 ;
  assign n9018 = n7764 ^ n7089 ^ 1'b0 ;
  assign n9019 = n3580 | n9018 ;
  assign n9020 = n7729 ^ n7346 ^ 1'b0 ;
  assign n9021 = n556 & ~n9020 ;
  assign n9022 = n5260 ^ n2087 ^ 1'b0 ;
  assign n9023 = n1206 & n9022 ;
  assign n9024 = n9023 ^ n3403 ^ 1'b0 ;
  assign n9025 = n5970 & n9024 ;
  assign n9026 = n9025 ^ n3342 ^ 1'b0 ;
  assign n9027 = n4136 ^ n1603 ^ 1'b0 ;
  assign n9028 = n9027 ^ n6084 ^ 1'b0 ;
  assign n9029 = ~n3904 & n9028 ;
  assign n9030 = n9029 ^ n1028 ^ 1'b0 ;
  assign n9031 = n6115 ^ n4316 ^ 1'b0 ;
  assign n9032 = n7838 & ~n9031 ;
  assign n9033 = n1421 & ~n4682 ;
  assign n9034 = ( ~x33 & n672 ) | ( ~x33 & n9033 ) | ( n672 & n9033 ) ;
  assign n9035 = x84 & ~n6506 ;
  assign n9036 = n9035 ^ n2903 ^ 1'b0 ;
  assign n9037 = n675 & ~n6634 ;
  assign n9038 = n6857 | n9037 ;
  assign n9039 = n9038 ^ n8935 ^ 1'b0 ;
  assign n9040 = n2424 & ~n5481 ;
  assign n9041 = n8796 ^ n3019 ^ n1046 ;
  assign n9042 = n6382 ^ n1832 ^ 1'b0 ;
  assign n9043 = ~n9041 & n9042 ;
  assign n9044 = n368 | n3441 ;
  assign n9045 = n5580 & ~n9044 ;
  assign n9046 = ~n7122 & n9045 ;
  assign n9047 = n5549 | n6519 ;
  assign n9048 = n4437 & ~n9047 ;
  assign n9049 = ( n3709 & n7532 ) | ( n3709 & n9048 ) | ( n7532 & n9048 ) ;
  assign n9050 = ( n468 & ~n1943 ) | ( n468 & n2481 ) | ( ~n1943 & n2481 ) ;
  assign n9051 = ( ~n6323 & n6511 ) | ( ~n6323 & n9050 ) | ( n6511 & n9050 ) ;
  assign n9052 = n3343 ^ n2745 ^ 1'b0 ;
  assign n9053 = n2502 | n9052 ;
  assign n9054 = n2235 & ~n9053 ;
  assign n9055 = ~n2261 & n9054 ;
  assign n9056 = n8738 | n9055 ;
  assign n9057 = n5220 & ~n9056 ;
  assign n9058 = n4834 & n7116 ;
  assign n9059 = n7734 ^ n7281 ^ n4465 ;
  assign n9060 = n769 | n9059 ;
  assign n9061 = n2621 & n3869 ;
  assign n9063 = n3274 & n5447 ;
  assign n9064 = n9063 ^ n2138 ^ 1'b0 ;
  assign n9062 = n4046 & ~n6418 ;
  assign n9065 = n9064 ^ n9062 ^ 1'b0 ;
  assign n9066 = x8 & ~n2921 ;
  assign n9067 = n9066 ^ n8159 ^ 1'b0 ;
  assign n9068 = n4012 ^ n1120 ^ 1'b0 ;
  assign n9069 = n2302 & n5970 ;
  assign n9070 = n9069 ^ n8903 ^ 1'b0 ;
  assign n9071 = n143 & n2168 ;
  assign n9072 = ~n2020 & n9071 ;
  assign n9073 = ( n3304 & ~n3530 ) | ( n3304 & n5000 ) | ( ~n3530 & n5000 ) ;
  assign n9074 = n3313 & n6205 ;
  assign n9075 = n2604 & n9074 ;
  assign n9076 = n2012 | n2656 ;
  assign n9077 = n9076 ^ n694 ^ 1'b0 ;
  assign n9078 = n1780 | n4737 ;
  assign n9079 = n7554 & ~n9078 ;
  assign n9080 = n8099 ^ n2078 ^ 1'b0 ;
  assign n9081 = n9080 ^ n6888 ^ 1'b0 ;
  assign n9082 = n313 | n9081 ;
  assign n9085 = n255 | n2525 ;
  assign n9083 = n5172 ^ n2463 ^ 1'b0 ;
  assign n9084 = n5308 & ~n9083 ;
  assign n9086 = n9085 ^ n9084 ^ 1'b0 ;
  assign n9087 = n4126 & ~n8514 ;
  assign n9088 = ~n1038 & n2462 ;
  assign n9089 = n9088 ^ n2619 ^ 1'b0 ;
  assign n9090 = n5583 ^ n3450 ^ 1'b0 ;
  assign n9091 = ~n9089 & n9090 ;
  assign n9092 = n7846 ^ n4765 ^ n2912 ;
  assign n9093 = ( n2671 & n2845 ) | ( n2671 & n2949 ) | ( n2845 & n2949 ) ;
  assign n9094 = n930 | n7481 ;
  assign n9095 = n9093 & n9094 ;
  assign n9096 = ~n8078 & n9095 ;
  assign n9097 = n4517 ^ n3916 ^ 1'b0 ;
  assign n9098 = ~n9096 & n9097 ;
  assign n9099 = n3975 ^ n2014 ^ 1'b0 ;
  assign n9100 = n7291 ^ n6963 ^ 1'b0 ;
  assign n9101 = n8947 ^ n208 ^ 1'b0 ;
  assign n9102 = n849 | n9101 ;
  assign n9103 = n6254 & ~n9102 ;
  assign n9104 = n5759 | n9103 ;
  assign n9105 = n4800 | n9104 ;
  assign n9106 = ( n1771 & ~n2336 ) | ( n1771 & n4357 ) | ( ~n2336 & n4357 ) ;
  assign n9107 = n1361 & ~n7901 ;
  assign n9108 = n5967 & n9107 ;
  assign n9109 = n4973 & n9108 ;
  assign n9110 = x94 & n574 ;
  assign n9111 = ~n184 & n9110 ;
  assign n9112 = n9111 ^ n676 ^ 1'b0 ;
  assign n9113 = x16 & ~n8442 ;
  assign n9114 = n3592 & n9113 ;
  assign n9115 = x10 | n7704 ;
  assign n9116 = n9115 ^ n2042 ^ x70 ;
  assign n9117 = ~n5077 & n8730 ;
  assign n9118 = n9117 ^ n6350 ^ 1'b0 ;
  assign n9119 = ~n2192 & n9118 ;
  assign n9120 = n2554 & ~n3651 ;
  assign n9121 = ~n3815 & n9120 ;
  assign n9122 = n9121 ^ n3279 ^ 1'b0 ;
  assign n9123 = n5730 | n9122 ;
  assign n9124 = n5557 ^ n2829 ^ n573 ;
  assign n9125 = n2183 & n8187 ;
  assign n9126 = n4797 ^ n4394 ^ 1'b0 ;
  assign n9127 = n2885 & n9126 ;
  assign n9128 = n3303 & n9127 ;
  assign n9129 = n2994 & ~n6013 ;
  assign n9130 = n7103 ^ n4113 ^ 1'b0 ;
  assign n9131 = n9130 ^ n5069 ^ 1'b0 ;
  assign n9132 = n3195 ^ x81 ^ 1'b0 ;
  assign n9133 = ~n358 & n9132 ;
  assign n9134 = n7570 & n9133 ;
  assign n9135 = n3855 | n6977 ;
  assign n9136 = n4303 & ~n9135 ;
  assign n9137 = n2357 ^ n1675 ^ 1'b0 ;
  assign n9138 = ~n4524 & n9137 ;
  assign n9139 = n4987 | n9138 ;
  assign n9140 = x89 & ~n4357 ;
  assign n9141 = n545 & n9140 ;
  assign n9142 = n9141 ^ n7666 ^ 1'b0 ;
  assign n9143 = n7170 & n9142 ;
  assign n9144 = n718 & ~n7417 ;
  assign n9145 = n2348 ^ n1824 ^ 1'b0 ;
  assign n9146 = n901 & n9145 ;
  assign n9147 = n9146 ^ n6127 ^ 1'b0 ;
  assign n9148 = ( n376 & n1526 ) | ( n376 & n2946 ) | ( n1526 & n2946 ) ;
  assign n9149 = n1862 & n2042 ;
  assign n9150 = n3542 & n9149 ;
  assign n9151 = n9150 ^ n8074 ^ 1'b0 ;
  assign n9153 = n3761 | n7261 ;
  assign n9152 = n5881 | n6407 ;
  assign n9154 = n9153 ^ n9152 ^ 1'b0 ;
  assign n9155 = n7303 | n9154 ;
  assign n9156 = n9155 ^ n5583 ^ 1'b0 ;
  assign n9157 = n7506 ^ n2483 ^ 1'b0 ;
  assign n9158 = n9156 & n9157 ;
  assign n9160 = n1550 & ~n8349 ;
  assign n9159 = n2235 | n7358 ;
  assign n9161 = n9160 ^ n9159 ^ 1'b0 ;
  assign n9162 = n5954 ^ n2232 ^ 1'b0 ;
  assign n9164 = n1073 & ~n1078 ;
  assign n9163 = n2624 & ~n6099 ;
  assign n9165 = n9164 ^ n9163 ^ n1329 ;
  assign n9169 = n3580 ^ n2596 ^ 1'b0 ;
  assign n9166 = n180 | n2146 ;
  assign n9167 = n3162 | n9166 ;
  assign n9168 = n4068 & n9167 ;
  assign n9170 = n9169 ^ n9168 ^ 1'b0 ;
  assign n9171 = n3405 & ~n7394 ;
  assign n9172 = n6120 ^ n4257 ^ n1073 ;
  assign n9173 = n5844 | n6558 ;
  assign n9174 = n9173 ^ n2012 ^ 1'b0 ;
  assign n9175 = n2589 & ~n9174 ;
  assign n9176 = n3458 & n9175 ;
  assign n9177 = n6172 ^ n1844 ^ n775 ;
  assign n9178 = ~n9176 & n9177 ;
  assign n9179 = n9178 ^ n6565 ^ 1'b0 ;
  assign n9180 = n9172 & ~n9179 ;
  assign n9181 = n4910 ^ n4884 ^ 1'b0 ;
  assign n9182 = n2832 | n9181 ;
  assign n9183 = n3824 ^ n928 ^ 1'b0 ;
  assign n9184 = n9182 & ~n9183 ;
  assign n9185 = n9184 ^ n6995 ^ 1'b0 ;
  assign n9186 = ~n1761 & n9185 ;
  assign n9187 = n1545 | n9186 ;
  assign n9188 = n641 ^ n209 ^ 1'b0 ;
  assign n9189 = n1565 & n9188 ;
  assign n9190 = n2893 & n7373 ;
  assign n9191 = n9189 & ~n9190 ;
  assign n9195 = n6934 ^ n3898 ^ 1'b0 ;
  assign n9192 = ~n643 & n3229 ;
  assign n9193 = n1308 | n1324 ;
  assign n9194 = ~n9192 & n9193 ;
  assign n9196 = n9195 ^ n9194 ^ 1'b0 ;
  assign n9197 = ( n4148 & n4502 ) | ( n4148 & n8810 ) | ( n4502 & n8810 ) ;
  assign n9198 = n661 & n3327 ;
  assign n9199 = n9198 ^ n203 ^ 1'b0 ;
  assign n9200 = x52 & n9199 ;
  assign n9201 = n4097 & ~n4611 ;
  assign n9202 = n3788 & n9201 ;
  assign n9203 = n7746 ^ n4997 ^ 1'b0 ;
  assign n9204 = n3544 & n3653 ;
  assign n9205 = n9204 ^ n1083 ^ 1'b0 ;
  assign n9206 = x94 & n9205 ;
  assign n9207 = ~n1200 & n9206 ;
  assign n9208 = n3528 & ~n9207 ;
  assign n9209 = n5492 & n9208 ;
  assign n9210 = ~x6 & n2823 ;
  assign n9211 = n9210 ^ n5207 ^ 1'b0 ;
  assign n9212 = n9211 ^ n838 ^ 1'b0 ;
  assign n9213 = n9212 ^ n8693 ^ 1'b0 ;
  assign n9214 = ( x30 & n2484 ) | ( x30 & n4032 ) | ( n2484 & n4032 ) ;
  assign n9215 = n9214 ^ n476 ^ n175 ;
  assign n9216 = n4548 & ~n7514 ;
  assign n9217 = n3558 | n9060 ;
  assign n9218 = n138 & n620 ;
  assign n9219 = ~n620 & n9218 ;
  assign n9220 = n861 | n9219 ;
  assign n9221 = n861 & ~n9220 ;
  assign n9222 = n9221 ^ n1353 ^ 1'b0 ;
  assign n9223 = n8958 & ~n9222 ;
  assign n9224 = n6759 ^ n3806 ^ 1'b0 ;
  assign n9225 = ~n8248 & n9224 ;
  assign n9226 = ~n3102 & n9225 ;
  assign n9227 = n9226 ^ x122 ^ 1'b0 ;
  assign n9228 = n1840 ^ n878 ^ 1'b0 ;
  assign n9229 = n9228 ^ n3884 ^ n556 ;
  assign n9230 = ~n958 & n1959 ;
  assign n9231 = n1861 & n9230 ;
  assign n9232 = n9231 ^ x117 ^ 1'b0 ;
  assign n9233 = n3887 | n9232 ;
  assign n9234 = n9233 ^ x120 ^ 1'b0 ;
  assign n9235 = n2699 & n2705 ;
  assign n9236 = n9235 ^ n8650 ^ 1'b0 ;
  assign n9237 = n9236 ^ n3690 ^ 1'b0 ;
  assign n9238 = ~n4788 & n9237 ;
  assign n9239 = n9238 ^ n6511 ^ 1'b0 ;
  assign n9240 = n9234 & n9239 ;
  assign n9245 = n1865 ^ x24 ^ 1'b0 ;
  assign n9244 = n3013 & ~n5535 ;
  assign n9246 = n9245 ^ n9244 ^ 1'b0 ;
  assign n9241 = n8144 ^ n6928 ^ 1'b0 ;
  assign n9242 = n3869 | n9241 ;
  assign n9243 = n9242 ^ n1908 ^ 1'b0 ;
  assign n9247 = n9246 ^ n9243 ^ 1'b0 ;
  assign n9248 = n7476 | n9247 ;
  assign n9249 = n4353 & n7646 ;
  assign n9250 = n3789 | n5127 ;
  assign n9251 = n6455 | n9250 ;
  assign n9252 = n4296 | n9251 ;
  assign n9253 = ~n1009 & n9252 ;
  assign n9254 = n902 & ~n4327 ;
  assign n9255 = n7617 & n9254 ;
  assign n9256 = n157 & ~n2334 ;
  assign n9257 = ~n1769 & n4352 ;
  assign n9258 = ~n9256 & n9257 ;
  assign n9259 = n9258 ^ n3744 ^ 1'b0 ;
  assign n9260 = n459 & n4076 ;
  assign n9261 = n9260 ^ n5776 ^ n5575 ;
  assign n9262 = n143 | n6481 ;
  assign n9263 = ( n611 & ~n1340 ) | ( n611 & n2655 ) | ( ~n1340 & n2655 ) ;
  assign n9264 = n6381 | n9263 ;
  assign n9265 = n9264 ^ n3897 ^ 1'b0 ;
  assign n9266 = n1473 & ~n5989 ;
  assign n9267 = n9265 & ~n9266 ;
  assign n9274 = n3294 & n3610 ;
  assign n9275 = ~n3673 & n9274 ;
  assign n9268 = n775 | n2370 ;
  assign n9269 = n344 & ~n9268 ;
  assign n9270 = ~n2563 & n9269 ;
  assign n9271 = n4547 | n5915 ;
  assign n9272 = n6137 | n9271 ;
  assign n9273 = n9270 & n9272 ;
  assign n9276 = n9275 ^ n9273 ^ 1'b0 ;
  assign n9277 = n614 ^ x44 ^ 1'b0 ;
  assign n9278 = n7399 ^ n5797 ^ 1'b0 ;
  assign n9279 = ~n2777 & n4989 ;
  assign n9280 = n4880 & n7753 ;
  assign n9281 = n6450 & n9280 ;
  assign n9282 = x3 & ~n9281 ;
  assign n9283 = ~n636 & n9282 ;
  assign n9284 = n2668 & n5415 ;
  assign n9285 = ~n3574 & n9284 ;
  assign n9286 = n9285 ^ n6355 ^ 1'b0 ;
  assign n9287 = n7284 ^ n458 ^ 1'b0 ;
  assign n9288 = n9262 ^ n3460 ^ n2608 ;
  assign n9289 = n1180 & ~n4498 ;
  assign n9290 = ~n1250 & n9289 ;
  assign n9291 = ~n3604 & n8772 ;
  assign n9292 = n8464 | n9291 ;
  assign n9293 = n4112 & ~n9292 ;
  assign n9294 = n593 | n2988 ;
  assign n9295 = n1615 & ~n9294 ;
  assign n9296 = n5365 | n9295 ;
  assign n9297 = n5138 | n9296 ;
  assign n9298 = n8226 ^ n6716 ^ 1'b0 ;
  assign n9299 = ~n2082 & n3795 ;
  assign n9301 = n4191 ^ n2687 ^ n2172 ;
  assign n9300 = ~n2448 & n3145 ;
  assign n9302 = n9301 ^ n9300 ^ 1'b0 ;
  assign n9303 = ~n1009 & n1200 ;
  assign n9304 = n9303 ^ n3066 ^ 1'b0 ;
  assign n9305 = n4257 ^ n3961 ^ 1'b0 ;
  assign n9306 = n3616 & n6108 ;
  assign n9307 = n1143 & ~n9306 ;
  assign n9311 = n4645 & n7588 ;
  assign n9308 = n6662 ^ n4650 ^ 1'b0 ;
  assign n9309 = n5107 & ~n9308 ;
  assign n9310 = ~n1390 & n9309 ;
  assign n9312 = n9311 ^ n9310 ^ 1'b0 ;
  assign n9313 = n2499 | n3517 ;
  assign n9314 = n2328 & n4831 ;
  assign n9315 = ( ~n571 & n3704 ) | ( ~n571 & n9314 ) | ( n3704 & n9314 ) ;
  assign n9316 = n2992 | n8260 ;
  assign n9317 = n1202 & ~n9316 ;
  assign n9318 = ~n2632 & n4667 ;
  assign n9319 = ~n3356 & n9318 ;
  assign n9320 = n9319 ^ n3226 ^ n1017 ;
  assign n9321 = ~n5146 & n9320 ;
  assign n9322 = ~n977 & n9321 ;
  assign n9323 = n838 & ~n5352 ;
  assign n9324 = n3304 & n9323 ;
  assign n9325 = n9324 ^ n6439 ^ 1'b0 ;
  assign n9327 = n131 | n778 ;
  assign n9328 = n9327 ^ n4063 ^ n3781 ;
  assign n9326 = n3565 & n4334 ;
  assign n9329 = n9328 ^ n9326 ^ 1'b0 ;
  assign n9330 = ( ~n5829 & n9319 ) | ( ~n5829 & n9329 ) | ( n9319 & n9329 ) ;
  assign n9331 = n1659 ^ n1606 ^ 1'b0 ;
  assign n9332 = ~n555 & n9331 ;
  assign n9333 = n163 & ~n9332 ;
  assign n9334 = ~n6410 & n9333 ;
  assign n9335 = n3102 | n9334 ;
  assign n9336 = n9335 ^ n3975 ^ 1'b0 ;
  assign n9337 = n6487 | n7332 ;
  assign n9338 = n9336 & n9337 ;
  assign n9339 = n3526 ^ n2502 ^ 1'b0 ;
  assign n9340 = n6591 & n9339 ;
  assign n9341 = n262 & n9340 ;
  assign n9342 = n9341 ^ n5392 ^ 1'b0 ;
  assign n9343 = ( ~n2265 & n4180 ) | ( ~n2265 & n9342 ) | ( n4180 & n9342 ) ;
  assign n9344 = n8716 & ~n9343 ;
  assign n9347 = n5102 | n6620 ;
  assign n9348 = n8960 & ~n9347 ;
  assign n9345 = n1790 & n2039 ;
  assign n9346 = n2708 | n9345 ;
  assign n9349 = n9348 ^ n9346 ^ 1'b0 ;
  assign n9350 = n3463 ^ n687 ^ 1'b0 ;
  assign n9351 = ( ~n4352 & n5170 ) | ( ~n4352 & n8026 ) | ( n5170 & n8026 ) ;
  assign n9352 = n9350 | n9351 ;
  assign n9353 = n9352 ^ n6609 ^ 1'b0 ;
  assign n9354 = n1243 ^ n148 ^ 1'b0 ;
  assign n9355 = n814 & n9354 ;
  assign n9356 = x123 & n9355 ;
  assign n9357 = n420 | n3135 ;
  assign n9358 = n9357 ^ n6457 ^ 1'b0 ;
  assign n9359 = n4693 & ~n8496 ;
  assign n9360 = ~n8617 & n9359 ;
  assign n9361 = n3164 & ~n5776 ;
  assign n9362 = ( n5500 & ~n8959 ) | ( n5500 & n9361 ) | ( ~n8959 & n9361 ) ;
  assign n9363 = n7453 ^ n722 ^ 1'b0 ;
  assign n9364 = n2234 & ~n9363 ;
  assign n9365 = n1089 & n9364 ;
  assign n9366 = ~n9080 & n9365 ;
  assign n9367 = n1169 & ~n3940 ;
  assign n9368 = ~n1701 & n9367 ;
  assign n9369 = n2024 & ~n3225 ;
  assign n9370 = n9369 ^ n3023 ^ 1'b0 ;
  assign n9371 = n4514 & n6133 ;
  assign n9372 = ~n198 & n9371 ;
  assign n9373 = x23 & ~n2438 ;
  assign n9374 = n5845 ^ n4002 ^ 1'b0 ;
  assign n9375 = n6827 & ~n9374 ;
  assign n9376 = n5934 ^ n4416 ^ 1'b0 ;
  assign n9377 = n2709 | n9376 ;
  assign n9378 = ~n2942 & n5901 ;
  assign n9379 = n6862 & n9378 ;
  assign n9380 = ( n1363 & ~n3331 ) | ( n1363 & n3529 ) | ( ~n3331 & n3529 ) ;
  assign n9381 = ( n3122 & ~n9234 ) | ( n3122 & n9380 ) | ( ~n9234 & n9380 ) ;
  assign n9387 = n1230 & n1442 ;
  assign n9388 = n9387 ^ n1102 ^ 1'b0 ;
  assign n9384 = n3270 & ~n4021 ;
  assign n9385 = ~x29 & n9384 ;
  assign n9386 = n7751 | n9385 ;
  assign n9389 = n9388 ^ n9386 ^ 1'b0 ;
  assign n9382 = n1681 ^ n614 ^ n417 ;
  assign n9383 = n4829 | n9382 ;
  assign n9390 = n9389 ^ n9383 ^ 1'b0 ;
  assign n9391 = n8819 ^ n8032 ^ 1'b0 ;
  assign n9392 = ~n3420 & n4997 ;
  assign n9393 = n3382 ^ n1344 ^ x116 ;
  assign n9394 = n3512 | n9393 ;
  assign n9395 = n5354 & ~n9394 ;
  assign n9396 = ~n9392 & n9395 ;
  assign n9397 = ~n5650 & n9396 ;
  assign n9398 = n4921 & n5394 ;
  assign n9399 = n9398 ^ n8496 ^ 1'b0 ;
  assign n9400 = n8489 ^ n1785 ^ 1'b0 ;
  assign n9401 = n3986 ^ n1009 ^ 1'b0 ;
  assign n9402 = n1334 & ~n9401 ;
  assign n9403 = n2119 & n9402 ;
  assign n9404 = ~n5711 & n9403 ;
  assign n9405 = n8194 | n9404 ;
  assign n9406 = n1060 | n9405 ;
  assign n9407 = n6207 & n9406 ;
  assign n9408 = n4320 | n9407 ;
  assign n9409 = ~n6268 & n9408 ;
  assign n9410 = ~n2996 & n5783 ;
  assign n9411 = ( n1901 & ~n6214 ) | ( n1901 & n9410 ) | ( ~n6214 & n9410 ) ;
  assign n9412 = n9411 ^ n5232 ^ 1'b0 ;
  assign n9413 = n2053 | n6067 ;
  assign n9414 = n9413 ^ x81 ^ 1'b0 ;
  assign n9415 = n6061 & n9414 ;
  assign n9416 = ~n7828 & n9415 ;
  assign n9417 = n2903 | n9416 ;
  assign n9418 = n4250 ^ n630 ^ 1'b0 ;
  assign n9419 = n6115 & ~n8282 ;
  assign n9420 = n2000 & ~n4491 ;
  assign n9421 = ~n2106 & n9420 ;
  assign n9422 = n8541 & n9421 ;
  assign n9423 = n9419 | n9422 ;
  assign n9424 = n8410 ^ n7737 ^ 1'b0 ;
  assign n9425 = ~n8393 & n9424 ;
  assign n9426 = n1223 & ~n1756 ;
  assign n9427 = n9426 ^ n5020 ^ 1'b0 ;
  assign n9428 = n563 ^ n540 ^ 1'b0 ;
  assign n9429 = n3594 ^ n428 ^ 1'b0 ;
  assign n9430 = n4972 ^ n397 ^ 1'b0 ;
  assign n9431 = n4832 | n9430 ;
  assign n9432 = n6858 | n9431 ;
  assign n9433 = n9432 ^ n7230 ^ 1'b0 ;
  assign n9434 = n4029 & ~n8920 ;
  assign n9435 = ~n9433 & n9434 ;
  assign n9436 = n9435 ^ n7400 ^ 1'b0 ;
  assign n9438 = n6649 ^ n3970 ^ 1'b0 ;
  assign n9437 = n1642 & ~n5419 ;
  assign n9439 = n9438 ^ n9437 ^ 1'b0 ;
  assign n9440 = ~n1874 & n4216 ;
  assign n9441 = n9440 ^ n5705 ^ 1'b0 ;
  assign n9442 = n1418 & n5871 ;
  assign n9443 = n3120 | n3222 ;
  assign n9444 = n7800 | n9443 ;
  assign n9445 = n5973 & ~n9444 ;
  assign n9446 = n5240 ^ n4905 ^ 1'b0 ;
  assign n9447 = n1240 ^ n747 ^ 1'b0 ;
  assign n9448 = ( n2718 & n6460 ) | ( n2718 & n9160 ) | ( n6460 & n9160 ) ;
  assign n9449 = x48 & ~n9448 ;
  assign n9450 = ~n9447 & n9449 ;
  assign n9451 = n6311 ^ n6059 ^ 1'b0 ;
  assign n9452 = n1163 & ~n4976 ;
  assign n9453 = ~n3789 & n9452 ;
  assign n9454 = n180 & n2834 ;
  assign n9455 = ~n4969 & n9454 ;
  assign n9456 = ~n6494 & n9143 ;
  assign n9457 = n2217 & n4936 ;
  assign n9458 = n9457 ^ n3011 ^ 1'b0 ;
  assign n9459 = n2340 & ~n4422 ;
  assign n9460 = n9459 ^ n679 ^ 1'b0 ;
  assign n9461 = n5134 | n5649 ;
  assign n9462 = n4684 | n9461 ;
  assign n9463 = n9462 ^ n8111 ^ n2151 ;
  assign n9464 = n7258 ^ n5505 ^ 1'b0 ;
  assign n9465 = ~n3116 & n9464 ;
  assign n9466 = ~n2474 & n4100 ;
  assign n9467 = ~x107 & n9466 ;
  assign n9468 = x13 & n2696 ;
  assign n9469 = n9467 & n9468 ;
  assign n9470 = n2807 & n4630 ;
  assign n9471 = n3681 & n9470 ;
  assign n9472 = n3314 ^ n1001 ^ 1'b0 ;
  assign n9473 = n4463 ^ n2608 ^ 1'b0 ;
  assign n9478 = ~n1691 & n6013 ;
  assign n9474 = n533 | n575 ;
  assign n9475 = n3327 & ~n9474 ;
  assign n9476 = ~n632 & n9475 ;
  assign n9477 = n6907 & ~n9476 ;
  assign n9479 = n9478 ^ n9477 ^ 1'b0 ;
  assign n9480 = n688 & n9350 ;
  assign n9481 = n6158 | n9480 ;
  assign n9482 = ~n3858 & n9481 ;
  assign n9483 = n6850 & ~n9482 ;
  assign n9484 = n9483 ^ n6024 ^ 1'b0 ;
  assign n9485 = n5398 ^ n5312 ^ n4761 ;
  assign n9486 = n1401 | n9485 ;
  assign n9487 = ~n1616 & n2361 ;
  assign n9488 = ~n827 & n4543 ;
  assign n9489 = n9487 & n9488 ;
  assign n9490 = n301 & n9489 ;
  assign n9494 = n2512 ^ n2305 ^ 1'b0 ;
  assign n9491 = n3948 ^ n1836 ^ 1'b0 ;
  assign n9492 = n272 | n9491 ;
  assign n9493 = n5036 & ~n9492 ;
  assign n9495 = n9494 ^ n9493 ^ 1'b0 ;
  assign n9496 = n4474 ^ n879 ^ 1'b0 ;
  assign n9497 = ~n5881 & n9496 ;
  assign n9498 = n8406 ^ n2229 ^ 1'b0 ;
  assign n9499 = n1124 & ~n4345 ;
  assign n9500 = n9499 ^ n811 ^ 1'b0 ;
  assign n9504 = n3011 ^ n2930 ^ n1507 ;
  assign n9501 = n1992 & n5860 ;
  assign n9502 = n890 & n9501 ;
  assign n9503 = n9502 ^ x110 ^ 1'b0 ;
  assign n9505 = n9504 ^ n9503 ^ n2648 ;
  assign n9506 = n5112 & n9505 ;
  assign n9507 = n1024 | n9506 ;
  assign n9508 = n9500 | n9507 ;
  assign n9509 = n5138 & n7988 ;
  assign n9510 = n5505 & n9509 ;
  assign n9511 = n2240 ^ n660 ^ 1'b0 ;
  assign n9512 = n630 | n9511 ;
  assign n9513 = n3082 & ~n3746 ;
  assign n9514 = n7203 ^ n879 ^ 1'b0 ;
  assign n9515 = n4798 & n9514 ;
  assign n9516 = n1377 & n2580 ;
  assign n9517 = n3869 & n9516 ;
  assign n9518 = n9517 ^ n3527 ^ 1'b0 ;
  assign n9519 = n3169 & n6678 ;
  assign n9520 = n1612 & n9519 ;
  assign n9521 = n2090 | n3210 ;
  assign n9522 = n8876 | n9521 ;
  assign n9523 = n8896 ^ n8080 ^ 1'b0 ;
  assign n9524 = n1529 ^ n766 ^ 1'b0 ;
  assign n9525 = n9524 ^ n1750 ^ 1'b0 ;
  assign n9526 = n7373 & ~n9525 ;
  assign n9527 = n9526 ^ n3931 ^ 1'b0 ;
  assign n9536 = n898 ^ x126 ^ 1'b0 ;
  assign n9537 = n971 | n9536 ;
  assign n9529 = ~n243 & n6321 ;
  assign n9530 = n4373 & ~n9529 ;
  assign n9531 = n4831 & n5332 ;
  assign n9532 = ~n4184 & n9531 ;
  assign n9533 = n9532 ^ n3450 ^ 1'b0 ;
  assign n9534 = n3051 | n9533 ;
  assign n9535 = n9530 | n9534 ;
  assign n9528 = n591 & n851 ;
  assign n9538 = n9537 ^ n9535 ^ n9528 ;
  assign n9539 = ~n2371 & n8878 ;
  assign n9540 = ~n3758 & n9539 ;
  assign n9541 = n7544 ^ n732 ^ 1'b0 ;
  assign n9542 = ( n5721 & n7270 ) | ( n5721 & ~n9541 ) | ( n7270 & ~n9541 ) ;
  assign n9543 = n2892 & n5557 ;
  assign n9544 = n950 & n9543 ;
  assign n9545 = n3390 & ~n9544 ;
  assign n9546 = n9545 ^ n1003 ^ 1'b0 ;
  assign n9548 = n601 | n2048 ;
  assign n9549 = n3030 & ~n9548 ;
  assign n9547 = ~n6055 & n8562 ;
  assign n9550 = n9549 ^ n9547 ^ 1'b0 ;
  assign n9551 = n7025 ^ n6992 ^ 1'b0 ;
  assign n9552 = n8784 & n8894 ;
  assign n9553 = ~n6066 & n6615 ;
  assign n9554 = n9553 ^ n5832 ^ 1'b0 ;
  assign n9555 = n7877 & ~n9554 ;
  assign n9556 = ~n7676 & n8781 ;
  assign n9557 = n562 & n2667 ;
  assign n9558 = n5556 ^ n3081 ^ 1'b0 ;
  assign n9559 = n2006 | n9558 ;
  assign n9560 = ~n5290 & n5652 ;
  assign n9561 = n9560 ^ n4216 ^ 1'b0 ;
  assign n9562 = n953 & n9561 ;
  assign n9563 = n8276 & n9562 ;
  assign n9564 = n9563 ^ n272 ^ 1'b0 ;
  assign n9565 = n9564 ^ n4516 ^ 1'b0 ;
  assign n9566 = n9139 & ~n9565 ;
  assign n9567 = n6237 | n8555 ;
  assign n9568 = n5592 & n9567 ;
  assign n9569 = n3430 | n4493 ;
  assign n9570 = n4261 & ~n9569 ;
  assign n9571 = n9570 ^ n2193 ^ 1'b0 ;
  assign n9572 = ~n8588 & n9571 ;
  assign n9573 = n9537 & n9572 ;
  assign n9576 = ~n851 & n7863 ;
  assign n9574 = n8349 ^ n8249 ^ n5253 ;
  assign n9575 = n166 & n9574 ;
  assign n9577 = n9576 ^ n9575 ^ 1'b0 ;
  assign n9578 = n9573 ^ n2412 ^ 1'b0 ;
  assign n9579 = n7181 ^ n5150 ^ 1'b0 ;
  assign n9580 = n1992 | n9579 ;
  assign n9581 = n7683 | n9580 ;
  assign n9583 = n3628 ^ n2087 ^ 1'b0 ;
  assign n9582 = ~n3602 & n5995 ;
  assign n9584 = n9583 ^ n9582 ^ 1'b0 ;
  assign n9585 = n1697 & n3376 ;
  assign n9586 = n5854 | n9585 ;
  assign n9589 = n1512 ^ n1179 ^ 1'b0 ;
  assign n9590 = n2088 | n9589 ;
  assign n9591 = ~n6712 & n9590 ;
  assign n9587 = n6785 ^ n5808 ^ 1'b0 ;
  assign n9588 = n1695 | n9587 ;
  assign n9592 = n9591 ^ n9588 ^ 1'b0 ;
  assign n9593 = ~n1560 & n9592 ;
  assign n9594 = n9586 & n9593 ;
  assign n9595 = n7038 ^ n5487 ^ 1'b0 ;
  assign n9596 = ~n5503 & n9595 ;
  assign n9597 = n2621 | n2896 ;
  assign n9598 = ~n7351 & n9597 ;
  assign n9600 = ~n1045 & n8509 ;
  assign n9599 = n675 & n4773 ;
  assign n9601 = n9600 ^ n9599 ^ 1'b0 ;
  assign n9602 = n5577 ^ n3906 ^ 1'b0 ;
  assign n9603 = n3221 & n9602 ;
  assign n9604 = n1891 & ~n9603 ;
  assign n9605 = n2204 & n2720 ;
  assign n9606 = n9605 ^ n7690 ^ 1'b0 ;
  assign n9607 = n4370 | n9606 ;
  assign n9608 = ( n858 & ~n3369 ) | ( n858 & n6246 ) | ( ~n3369 & n6246 ) ;
  assign n9609 = n1549 | n5235 ;
  assign n9610 = n9608 & ~n9609 ;
  assign n9611 = ( n4252 & n4859 ) | ( n4252 & ~n9610 ) | ( n4859 & ~n9610 ) ;
  assign n9612 = n7137 & n9611 ;
  assign n9613 = n4640 & n9612 ;
  assign n9614 = n6659 ^ n4453 ^ 1'b0 ;
  assign n9615 = n4342 & ~n9614 ;
  assign n9616 = n6636 ^ n4983 ^ 1'b0 ;
  assign n9617 = n8510 & ~n9616 ;
  assign n9618 = n9617 ^ n788 ^ 1'b0 ;
  assign n9619 = n458 & ~n4779 ;
  assign n9620 = n4021 & n9619 ;
  assign n9621 = n9620 ^ n2777 ^ 1'b0 ;
  assign n9623 = n3148 & ~n5443 ;
  assign n9624 = n9623 ^ n5248 ^ 1'b0 ;
  assign n9622 = ~n802 & n1578 ;
  assign n9625 = n9624 ^ n9622 ^ 1'b0 ;
  assign n9626 = n9621 | n9625 ;
  assign n9627 = n9626 ^ n2397 ^ 1'b0 ;
  assign n9629 = n1337 ^ n218 ^ 1'b0 ;
  assign n9630 = n2979 & ~n9629 ;
  assign n9628 = n7042 ^ n3049 ^ 1'b0 ;
  assign n9631 = n9630 ^ n9628 ^ 1'b0 ;
  assign n9632 = n2924 & ~n9631 ;
  assign n9633 = ~n243 & n9378 ;
  assign n9634 = n9633 ^ n6784 ^ 1'b0 ;
  assign n9635 = n7631 & n9634 ;
  assign n9636 = n7419 ^ n658 ^ 1'b0 ;
  assign n9637 = n3952 | n9636 ;
  assign n9638 = ~n257 & n7259 ;
  assign n9639 = n1917 & n5243 ;
  assign n9640 = n9639 ^ n3558 ^ 1'b0 ;
  assign n9641 = n3160 & ~n9640 ;
  assign n9642 = ~n9638 & n9641 ;
  assign n9643 = n1388 ^ n478 ^ 1'b0 ;
  assign n9644 = n9611 & n9643 ;
  assign n9645 = ( x92 & ~n277 ) | ( x92 & n1743 ) | ( ~n277 & n1743 ) ;
  assign n9646 = ~n6442 & n9645 ;
  assign n9647 = n8632 & n8952 ;
  assign n9648 = ~n1136 & n6369 ;
  assign n9649 = n4819 & n9648 ;
  assign n9650 = ( n3597 & n6760 ) | ( n3597 & n9649 ) | ( n6760 & n9649 ) ;
  assign n9651 = n2330 & n2742 ;
  assign n9652 = n9651 ^ n7822 ^ 1'b0 ;
  assign n9653 = n1177 | n8194 ;
  assign n9654 = n456 | n9653 ;
  assign n9655 = n5320 | n9654 ;
  assign n9656 = n9655 ^ x84 ^ 1'b0 ;
  assign n9657 = n4899 | n9656 ;
  assign n9658 = n3997 ^ n2142 ^ 1'b0 ;
  assign n9659 = ~n6599 & n9658 ;
  assign n9660 = ~n5931 & n9659 ;
  assign n9661 = n4357 | n9167 ;
  assign n9662 = n3214 & n4351 ;
  assign n9663 = n593 & n3521 ;
  assign n9664 = n674 & ~n9663 ;
  assign n9665 = n2787 & n3483 ;
  assign n9666 = n6559 ^ n1619 ^ n1065 ;
  assign n9667 = n5613 & ~n6331 ;
  assign n9668 = n9666 & n9667 ;
  assign n9669 = n5843 & ~n9668 ;
  assign n9670 = ~n2798 & n9669 ;
  assign n9671 = n4843 & ~n7849 ;
  assign n9672 = n6889 ^ n5578 ^ n3696 ;
  assign n9673 = n371 | n8247 ;
  assign n9674 = n894 | n6372 ;
  assign n9675 = n9673 & ~n9674 ;
  assign n9676 = n3259 ^ n3066 ^ n2948 ;
  assign n9677 = n723 & ~n9676 ;
  assign n9678 = n5038 & ~n5457 ;
  assign n9679 = n2168 & ~n8123 ;
  assign n9680 = ~n2973 & n9679 ;
  assign n9683 = n3614 & ~n5482 ;
  assign n9684 = n4217 & ~n9683 ;
  assign n9685 = ( n478 & n3866 ) | ( n478 & ~n9684 ) | ( n3866 & ~n9684 ) ;
  assign n9681 = n2745 ^ n1854 ^ 1'b0 ;
  assign n9682 = ~n220 & n9681 ;
  assign n9686 = n9685 ^ n9682 ^ 1'b0 ;
  assign n9688 = n4429 & n4562 ;
  assign n9687 = n2176 & n9151 ;
  assign n9689 = n9688 ^ n9687 ^ 1'b0 ;
  assign n9690 = n9328 ^ n7734 ^ n1030 ;
  assign n9691 = n2470 ^ n640 ^ 1'b0 ;
  assign n9692 = ( ~n4095 & n6361 ) | ( ~n4095 & n9691 ) | ( n6361 & n9691 ) ;
  assign n9693 = n9645 | n9692 ;
  assign n9694 = ~n2560 & n9693 ;
  assign n9695 = n559 ^ n404 ^ 1'b0 ;
  assign n9696 = n5473 ^ n3894 ^ 1'b0 ;
  assign n9697 = x21 & n1429 ;
  assign n9698 = n9697 ^ n4063 ^ 1'b0 ;
  assign n9699 = n1973 ^ n953 ^ n621 ;
  assign n9700 = n5909 & ~n9699 ;
  assign n9701 = ~n4557 & n9700 ;
  assign n9702 = n789 | n4813 ;
  assign n9703 = n2911 & ~n9702 ;
  assign n9704 = n1343 & n6271 ;
  assign n9705 = ~n4228 & n9704 ;
  assign n9706 = n2049 | n9705 ;
  assign n9707 = n7826 ^ n7688 ^ 1'b0 ;
  assign n9708 = n9707 ^ n7053 ^ n1631 ;
  assign n9709 = n2116 & ~n7940 ;
  assign n9710 = ~n5778 & n9709 ;
  assign n9711 = n6369 ^ n5836 ^ 1'b0 ;
  assign n9712 = ~n324 & n9711 ;
  assign n9713 = n9712 ^ n4240 ^ 1'b0 ;
  assign n9714 = ~n5766 & n9713 ;
  assign n9715 = n5015 ^ n2827 ^ n2587 ;
  assign n9716 = n5537 & n9715 ;
  assign n9717 = x69 & ~n5810 ;
  assign n9718 = n9420 ^ n5351 ^ n4729 ;
  assign n9719 = n3505 | n5514 ;
  assign n9720 = n4547 & ~n9719 ;
  assign n9721 = n9385 ^ n7882 ^ n6427 ;
  assign n9725 = n175 | n3078 ;
  assign n9722 = x76 & n3489 ;
  assign n9723 = n9722 ^ n4340 ^ 1'b0 ;
  assign n9724 = n1865 | n9723 ;
  assign n9726 = n9725 ^ n9724 ^ 1'b0 ;
  assign n9727 = n9721 & n9726 ;
  assign n9728 = n4449 ^ n2779 ^ 1'b0 ;
  assign n9729 = n3872 | n9728 ;
  assign n9730 = x50 & ~n1708 ;
  assign n9731 = n6779 & n9730 ;
  assign n9732 = n9731 ^ n7877 ^ n7388 ;
  assign n9733 = ~n9729 & n9732 ;
  assign n9734 = n4527 & n8407 ;
  assign n9747 = n3289 ^ n1165 ^ 1'b0 ;
  assign n9748 = n2416 & ~n9747 ;
  assign n9749 = n3601 & ~n5822 ;
  assign n9750 = n9748 & n9749 ;
  assign n9751 = ~n9748 & n9750 ;
  assign n9735 = ~n414 & n585 ;
  assign n9736 = ~n585 & n9735 ;
  assign n9737 = n2605 & ~n8183 ;
  assign n9738 = ~n2605 & n9737 ;
  assign n9739 = n4737 | n9738 ;
  assign n9740 = n9738 & ~n9739 ;
  assign n9741 = n2993 | n3601 ;
  assign n9742 = n2993 & ~n9741 ;
  assign n9743 = n4456 & ~n9742 ;
  assign n9744 = ~n2313 & n9743 ;
  assign n9745 = n9740 & n9744 ;
  assign n9746 = n9736 | n9745 ;
  assign n9752 = n9751 ^ n9746 ^ 1'b0 ;
  assign n9753 = n801 & ~n7549 ;
  assign n9754 = n9413 | n9753 ;
  assign n9755 = ~n391 & n9754 ;
  assign n9758 = n2603 ^ n679 ^ 1'b0 ;
  assign n9756 = n4747 ^ n580 ^ 1'b0 ;
  assign n9757 = ~n3488 & n9756 ;
  assign n9759 = n9758 ^ n9757 ^ 1'b0 ;
  assign n9760 = n6800 & n9396 ;
  assign n9761 = n8816 ^ n801 ^ 1'b0 ;
  assign n9762 = n7018 & ~n9761 ;
  assign n9763 = n9760 & n9762 ;
  assign n9764 = n1620 & n2696 ;
  assign n9765 = n9764 ^ n5316 ^ 1'b0 ;
  assign n9766 = n9649 ^ n327 ^ 1'b0 ;
  assign n9767 = n1943 ^ n166 ^ 1'b0 ;
  assign n9768 = n2872 | n9767 ;
  assign n9769 = n901 & ~n9768 ;
  assign n9770 = n9769 ^ n278 ^ 1'b0 ;
  assign n9771 = n1079 | n9770 ;
  assign n9772 = n2234 & ~n2638 ;
  assign n9773 = n9772 ^ n6238 ^ 1'b0 ;
  assign n9774 = n9770 ^ n1507 ^ 1'b0 ;
  assign n9775 = n3420 | n6674 ;
  assign n9776 = n2831 | n9164 ;
  assign n9778 = n2192 & ~n2794 ;
  assign n9777 = ~n3200 & n9571 ;
  assign n9779 = n9778 ^ n9777 ^ 1'b0 ;
  assign n9780 = ( ~n1703 & n4051 ) | ( ~n1703 & n7350 ) | ( n4051 & n7350 ) ;
  assign n9781 = n5917 ^ n615 ^ 1'b0 ;
  assign n9782 = n4419 & ~n9781 ;
  assign n9783 = n9782 ^ n9160 ^ 1'b0 ;
  assign n9784 = n2597 ^ n2402 ^ 1'b0 ;
  assign n9785 = n9784 ^ n560 ^ 1'b0 ;
  assign n9786 = n1562 & ~n9785 ;
  assign n9787 = n6764 ^ n4498 ^ 1'b0 ;
  assign n9788 = n1157 & ~n9787 ;
  assign n9789 = n1478 & n9788 ;
  assign n9790 = n1439 ^ n577 ^ 1'b0 ;
  assign n9791 = n2382 ^ n530 ^ 1'b0 ;
  assign n9792 = ~n7358 & n9791 ;
  assign n9793 = ( ~n9100 & n9790 ) | ( ~n9100 & n9792 ) | ( n9790 & n9792 ) ;
  assign n9794 = n8386 ^ n3245 ^ n1617 ;
  assign n9795 = n9794 ^ n7655 ^ n2479 ;
  assign n9796 = n692 & ~n5590 ;
  assign n9797 = n4450 & ~n9796 ;
  assign n9799 = ( n386 & n2185 ) | ( n386 & n2869 ) | ( n2185 & n2869 ) ;
  assign n9800 = ~n7615 & n9799 ;
  assign n9798 = n915 & ~n3342 ;
  assign n9801 = n9800 ^ n9798 ^ n3431 ;
  assign n9802 = n5699 ^ n2769 ^ 1'b0 ;
  assign n9803 = n3936 | n8553 ;
  assign n9804 = n2318 | n6281 ;
  assign n9805 = n3418 & n9804 ;
  assign n9806 = ~n9803 & n9805 ;
  assign n9807 = n9806 ^ n7521 ^ 1'b0 ;
  assign n9808 = n2128 ^ n2028 ^ 1'b0 ;
  assign n9810 = ( n2372 & n4200 ) | ( n2372 & n5156 ) | ( n4200 & n5156 ) ;
  assign n9809 = n879 & n2782 ;
  assign n9811 = n9810 ^ n9809 ^ 1'b0 ;
  assign n9812 = n9655 ^ n272 ^ 1'b0 ;
  assign n9813 = n4386 ^ n3844 ^ n844 ;
  assign n9814 = n1770 | n8071 ;
  assign n9815 = n9813 | n9814 ;
  assign n9816 = n3174 & ~n4553 ;
  assign n9817 = n9816 ^ n4737 ^ 1'b0 ;
  assign n9818 = ~n7617 & n9817 ;
  assign n9819 = n8415 & n9818 ;
  assign n9820 = n1812 & ~n8280 ;
  assign n9821 = ~n2423 & n6222 ;
  assign n9823 = ~n2361 & n6147 ;
  assign n9822 = n5451 | n7128 ;
  assign n9824 = n9823 ^ n9822 ^ 1'b0 ;
  assign n9825 = n4468 ^ n861 ^ 1'b0 ;
  assign n9826 = n2158 & n9825 ;
  assign n9827 = ~n3280 & n9826 ;
  assign n9828 = x54 & n9827 ;
  assign n9829 = n9828 ^ n1761 ^ 1'b0 ;
  assign n9831 = n8817 & n9422 ;
  assign n9830 = n3288 & ~n5654 ;
  assign n9832 = n9831 ^ n9830 ^ 1'b0 ;
  assign n9833 = ( x82 & n2990 ) | ( x82 & n3865 ) | ( n2990 & n3865 ) ;
  assign n9834 = ( n5676 & n8577 ) | ( n5676 & ~n9833 ) | ( n8577 & ~n9833 ) ;
  assign n9836 = n3420 & n5132 ;
  assign n9837 = ~n3730 & n9836 ;
  assign n9838 = n9634 & n9837 ;
  assign n9839 = n1438 & n9838 ;
  assign n9840 = n3013 & n3124 ;
  assign n9841 = n9839 & n9840 ;
  assign n9835 = ~n4430 & n4578 ;
  assign n9842 = n9841 ^ n9835 ^ 1'b0 ;
  assign n9843 = n5647 ^ n3322 ^ 1'b0 ;
  assign n9846 = n3820 ^ n2378 ^ n2203 ;
  assign n9844 = n1182 & ~n5457 ;
  assign n9845 = n9844 ^ n1881 ^ 1'b0 ;
  assign n9847 = n9846 ^ n9845 ^ n2582 ;
  assign n9848 = n9847 ^ n4683 ^ 1'b0 ;
  assign n9850 = n4633 ^ n3247 ^ 1'b0 ;
  assign n9849 = n2380 & ~n9698 ;
  assign n9851 = n9850 ^ n9849 ^ 1'b0 ;
  assign n9852 = n2262 ^ n308 ^ 1'b0 ;
  assign n9853 = n6187 & ~n9130 ;
  assign n9854 = ~n9852 & n9853 ;
  assign n9855 = ~n4035 & n9854 ;
  assign n9859 = n1088 & n2003 ;
  assign n9860 = ~n2003 & n9859 ;
  assign n9856 = n4802 ^ n2765 ^ 1'b0 ;
  assign n9857 = n9856 ^ n2542 ^ 1'b0 ;
  assign n9858 = x124 & ~n9857 ;
  assign n9861 = n9860 ^ n9858 ^ n7968 ;
  assign n9862 = n829 & ~n1689 ;
  assign n9863 = ( ~n180 & n2769 ) | ( ~n180 & n9862 ) | ( n2769 & n9862 ) ;
  assign n9864 = n9863 ^ n4745 ^ 1'b0 ;
  assign n9865 = n6061 ^ n2794 ^ n2416 ;
  assign n9866 = x6 | n9865 ;
  assign n9867 = n1605 & ~n9866 ;
  assign n9868 = n2769 & ~n8852 ;
  assign n9872 = n8061 ^ n7688 ^ n7355 ;
  assign n9870 = ~n2537 & n2793 ;
  assign n9871 = n4314 & n9870 ;
  assign n9869 = n8074 ^ n7143 ^ 1'b0 ;
  assign n9873 = n9872 ^ n9871 ^ n9869 ;
  assign n9874 = ( n357 & n2937 ) | ( n357 & n7404 ) | ( n2937 & n7404 ) ;
  assign n9875 = n2248 & ~n3437 ;
  assign n9876 = n9875 ^ n7581 ^ 1'b0 ;
  assign n9877 = n5241 & ~n9876 ;
  assign n9878 = ~n5652 & n9877 ;
  assign n9879 = ~n303 & n1390 ;
  assign n9880 = ( ~n1638 & n5136 ) | ( ~n1638 & n7510 ) | ( n5136 & n7510 ) ;
  assign n9881 = n2833 & ~n7936 ;
  assign n9882 = n9880 & n9881 ;
  assign n9883 = n965 & n3169 ;
  assign n9884 = n1113 & n9883 ;
  assign n9885 = ( n362 & ~n7849 ) | ( n362 & n9146 ) | ( ~n7849 & n9146 ) ;
  assign n9886 = n9885 ^ n792 ^ 1'b0 ;
  assign n9890 = ~n1343 & n6232 ;
  assign n9887 = n5466 ^ n2955 ^ 1'b0 ;
  assign n9888 = n5635 & ~n9887 ;
  assign n9889 = n2243 & ~n9888 ;
  assign n9891 = n9890 ^ n9889 ^ 1'b0 ;
  assign n9892 = ~n1732 & n4564 ;
  assign n9893 = ~n999 & n5243 ;
  assign n9894 = ~n5356 & n9893 ;
  assign n9895 = n9894 ^ n8475 ^ 1'b0 ;
  assign n9896 = n5669 & ~n7488 ;
  assign n9897 = n9896 ^ n2288 ^ 1'b0 ;
  assign n9898 = n5992 ^ n4857 ^ 1'b0 ;
  assign n9899 = n6506 & n9898 ;
  assign n9900 = n9899 ^ x37 ^ 1'b0 ;
  assign n9901 = ~n9897 & n9900 ;
  assign n9902 = n437 & ~n1213 ;
  assign n9903 = n4263 ^ x84 ^ 1'b0 ;
  assign n9904 = n7234 | n9903 ;
  assign n9905 = ~n9089 & n9729 ;
  assign n9906 = n9904 & ~n9905 ;
  assign n9907 = ~n1999 & n4957 ;
  assign n9908 = n9907 ^ n5981 ^ 1'b0 ;
  assign n9909 = ~n2204 & n7468 ;
  assign n9910 = n2374 | n5669 ;
  assign n9911 = x22 & n3354 ;
  assign n9912 = n9910 & ~n9911 ;
  assign n9913 = n9912 ^ n4773 ^ 1'b0 ;
  assign n9914 = n3180 ^ n2648 ^ 1'b0 ;
  assign n9915 = n6894 | n9914 ;
  assign n9916 = n9013 & ~n9915 ;
  assign n9917 = ~n8452 & n9916 ;
  assign n9918 = ~n3806 & n4132 ;
  assign n9919 = ~n1929 & n9918 ;
  assign n9920 = n1639 | n6946 ;
  assign n9922 = n8292 ^ n2193 ^ 1'b0 ;
  assign n9923 = x69 & n9922 ;
  assign n9924 = n174 | n2829 ;
  assign n9925 = n9924 ^ n7057 ^ 1'b0 ;
  assign n9926 = n9923 & ~n9925 ;
  assign n9921 = n332 & ~n8308 ;
  assign n9927 = n9926 ^ n9921 ^ 1'b0 ;
  assign n9934 = ~n973 & n5574 ;
  assign n9932 = n3414 ^ n3004 ^ 1'b0 ;
  assign n9933 = n2828 & n9932 ;
  assign n9935 = n9934 ^ n9933 ^ 1'b0 ;
  assign n9928 = n7621 & ~n9410 ;
  assign n9929 = n9928 ^ n728 ^ 1'b0 ;
  assign n9930 = n2344 | n9929 ;
  assign n9931 = ( n8315 & ~n8786 ) | ( n8315 & n9930 ) | ( ~n8786 & n9930 ) ;
  assign n9936 = n9935 ^ n9931 ^ 1'b0 ;
  assign n9937 = n4526 | n9936 ;
  assign n9938 = n2937 ^ n220 ^ 1'b0 ;
  assign n9939 = n904 & n9938 ;
  assign n9940 = n8824 ^ n573 ^ 1'b0 ;
  assign n9941 = ( n4887 & n9939 ) | ( n4887 & ~n9940 ) | ( n9939 & ~n9940 ) ;
  assign n9942 = ~n1254 & n4292 ;
  assign n9943 = n3914 | n8906 ;
  assign n9944 = n9943 ^ n1893 ^ 1'b0 ;
  assign n9945 = n1248 | n2339 ;
  assign n9946 = n9945 ^ n5323 ^ 1'b0 ;
  assign n9947 = n7100 ^ x66 ^ 1'b0 ;
  assign n9955 = n458 & n3209 ;
  assign n9956 = n1047 & n9955 ;
  assign n9957 = ~n2545 & n9956 ;
  assign n9952 = ~n704 & n4452 ;
  assign n9953 = ~n2589 & n9952 ;
  assign n9954 = n5021 | n9953 ;
  assign n9958 = n9957 ^ n9954 ^ 1'b0 ;
  assign n9959 = ( x94 & n3768 ) | ( x94 & ~n9958 ) | ( n3768 & ~n9958 ) ;
  assign n9960 = ( n8945 & n9601 ) | ( n8945 & ~n9959 ) | ( n9601 & ~n9959 ) ;
  assign n9948 = n1791 | n3188 ;
  assign n9949 = n9948 ^ n3764 ^ 1'b0 ;
  assign n9950 = n9949 ^ n5062 ^ 1'b0 ;
  assign n9951 = n6131 & ~n9950 ;
  assign n9961 = n9960 ^ n9951 ^ 1'b0 ;
  assign n9962 = n3806 & n6384 ;
  assign n9963 = n5547 ^ n1770 ^ 1'b0 ;
  assign n9964 = n768 & n9963 ;
  assign n9965 = ~n5503 & n9964 ;
  assign n9966 = ~n9962 & n9965 ;
  assign n9967 = n9597 ^ n8124 ^ 1'b0 ;
  assign n9968 = n6120 | n9028 ;
  assign n9969 = n9968 ^ n4324 ^ 1'b0 ;
  assign n9970 = n8106 ^ n456 ^ 1'b0 ;
  assign n9971 = n9010 & n9970 ;
  assign n9972 = n5613 & ~n9971 ;
  assign n9973 = n2319 & n2517 ;
  assign n9974 = n4104 ^ n2829 ^ 1'b0 ;
  assign n9975 = ~n1876 & n9974 ;
  assign n9976 = n4708 & n9975 ;
  assign n9977 = n9976 ^ n1688 ^ 1'b0 ;
  assign n9978 = ~n6644 & n7213 ;
  assign n9979 = n2561 & ~n6132 ;
  assign n9980 = n9979 ^ n6821 ^ 1'b0 ;
  assign n9981 = n525 & ~n8304 ;
  assign n9982 = n9934 & n9981 ;
  assign n9983 = ~n1893 & n2228 ;
  assign n9984 = n9983 ^ n3755 ^ 1'b0 ;
  assign n9985 = n9984 ^ n3773 ^ 1'b0 ;
  assign n9986 = n9982 | n9985 ;
  assign n9987 = ~n1420 & n5615 ;
  assign n9988 = n2039 ^ x34 ^ 1'b0 ;
  assign n9989 = n2659 & ~n5448 ;
  assign n9990 = ~n9988 & n9989 ;
  assign n9991 = n9987 | n9990 ;
  assign n9992 = n9991 ^ n4281 ^ 1'b0 ;
  assign n9993 = n1174 & n6181 ;
  assign n9994 = n6610 & n9993 ;
  assign n9995 = n9994 ^ n2605 ^ 1'b0 ;
  assign n9996 = n2382 ^ n1585 ^ 1'b0 ;
  assign n9997 = n9996 ^ n1645 ^ 1'b0 ;
  assign n9998 = x25 & x81 ;
  assign n9999 = n9998 ^ n1560 ^ 1'b0 ;
  assign n10000 = n5181 & ~n5227 ;
  assign n10001 = n10000 ^ n481 ^ 1'b0 ;
  assign n10002 = n9107 & n10001 ;
  assign n10003 = ~n2435 & n10002 ;
  assign n10005 = n6206 ^ n3058 ^ 1'b0 ;
  assign n10006 = n8738 | n10005 ;
  assign n10004 = n2240 | n8938 ;
  assign n10007 = n10006 ^ n10004 ^ 1'b0 ;
  assign n10008 = ( ~x17 & n3830 ) | ( ~x17 & n6137 ) | ( n3830 & n6137 ) ;
  assign n10009 = n505 & n10008 ;
  assign n10010 = n10009 ^ n2877 ^ 1'b0 ;
  assign n10011 = ~n2654 & n3637 ;
  assign n10012 = n10011 ^ n5531 ^ 1'b0 ;
  assign n10013 = ( n3835 & n4264 ) | ( n3835 & ~n10012 ) | ( n4264 & ~n10012 ) ;
  assign n10021 = n6972 ^ n687 ^ 1'b0 ;
  assign n10014 = n2994 ^ n722 ^ 1'b0 ;
  assign n10015 = n888 & ~n7017 ;
  assign n10016 = n2188 | n10015 ;
  assign n10017 = n10016 ^ n3827 ^ 1'b0 ;
  assign n10018 = n10017 ^ n632 ^ 1'b0 ;
  assign n10019 = n10014 | n10018 ;
  assign n10020 = n985 & ~n10019 ;
  assign n10022 = n10021 ^ n10020 ^ 1'b0 ;
  assign n10025 = n3279 & n3492 ;
  assign n10026 = ~n391 & n10025 ;
  assign n10023 = n2188 ^ n742 ^ 1'b0 ;
  assign n10024 = n6531 & ~n10023 ;
  assign n10027 = n10026 ^ n10024 ^ n639 ;
  assign n10028 = ~n666 & n5971 ;
  assign n10029 = n10028 ^ n2103 ^ 1'b0 ;
  assign n10030 = n667 & n2985 ;
  assign n10031 = n8911 & n10030 ;
  assign n10032 = n10031 ^ n8294 ^ 1'b0 ;
  assign n10033 = n5574 | n10032 ;
  assign n10034 = n1342 ^ n150 ^ 1'b0 ;
  assign n10035 = n2819 | n10034 ;
  assign n10036 = n5836 | n8246 ;
  assign n10037 = n147 & ~n8840 ;
  assign n10038 = ~n1094 & n10037 ;
  assign n10039 = ~n1888 & n10038 ;
  assign n10040 = ~n3376 & n10039 ;
  assign n10041 = n678 & n7858 ;
  assign n10042 = n3381 | n8490 ;
  assign n10043 = n530 | n10042 ;
  assign n10044 = n2483 ^ n203 ^ 1'b0 ;
  assign n10045 = n6781 | n10044 ;
  assign n10046 = n10045 ^ n9504 ^ n719 ;
  assign n10047 = n911 & ~n10001 ;
  assign n10048 = n7674 ^ n4224 ^ 1'b0 ;
  assign n10049 = n9143 | n10048 ;
  assign n10050 = n261 & n5347 ;
  assign n10051 = n6712 & n10050 ;
  assign n10052 = n3734 ^ n366 ^ 1'b0 ;
  assign n10053 = ~n5662 & n10052 ;
  assign n10054 = n8704 ^ n3662 ^ n3413 ;
  assign n10055 = ( n4514 & n10053 ) | ( n4514 & ~n10054 ) | ( n10053 & ~n10054 ) ;
  assign n10056 = n3115 & ~n3981 ;
  assign n10057 = n10056 ^ n6561 ^ 1'b0 ;
  assign n10058 = n1418 | n8348 ;
  assign n10059 = n10058 ^ n902 ^ 1'b0 ;
  assign n10060 = n722 & n10059 ;
  assign n10061 = n5389 & n10060 ;
  assign n10062 = n2206 | n10061 ;
  assign n10063 = n10062 ^ n3100 ^ 1'b0 ;
  assign n10064 = n10063 ^ n2396 ^ 1'b0 ;
  assign n10065 = n8712 | n10064 ;
  assign n10066 = n4348 | n10065 ;
  assign n10067 = ~n2569 & n4510 ;
  assign n10068 = n3015 & ~n5082 ;
  assign n10069 = ~n10067 & n10068 ;
  assign n10070 = n7984 ^ n4743 ^ 1'b0 ;
  assign n10071 = ~n943 & n5246 ;
  assign n10072 = n4681 & n10071 ;
  assign n10073 = ~n976 & n10072 ;
  assign n10074 = n1254 | n5161 ;
  assign n10075 = n3535 & ~n10074 ;
  assign n10076 = n2715 & ~n4259 ;
  assign n10077 = n3907 & n10076 ;
  assign n10078 = n6544 ^ n3182 ^ n787 ;
  assign n10079 = n10078 ^ n9616 ^ n1990 ;
  assign n10080 = ~n593 & n657 ;
  assign n10081 = n10080 ^ n2782 ^ 1'b0 ;
  assign n10082 = ~n2558 & n10081 ;
  assign n10083 = n3752 & n10082 ;
  assign n10084 = n10083 ^ n6348 ^ 1'b0 ;
  assign n10086 = n4255 ^ n335 ^ 1'b0 ;
  assign n10085 = n1881 & ~n7004 ;
  assign n10087 = n10086 ^ n10085 ^ 1'b0 ;
  assign n10088 = n2240 ^ n1587 ^ x37 ;
  assign n10089 = n9272 | n10088 ;
  assign n10090 = n3348 ^ n770 ^ 1'b0 ;
  assign n10092 = n6297 ^ n730 ^ 1'b0 ;
  assign n10093 = ~n3346 & n9504 ;
  assign n10094 = ~n10092 & n10093 ;
  assign n10095 = ( n2280 & ~n9385 ) | ( n2280 & n10094 ) | ( ~n9385 & n10094 ) ;
  assign n10091 = n7250 ^ n3601 ^ 1'b0 ;
  assign n10096 = n10095 ^ n10091 ^ n832 ;
  assign n10097 = n1889 & n9302 ;
  assign n10098 = ~n1394 & n10097 ;
  assign n10099 = n6291 ^ x76 ^ 1'b0 ;
  assign n10100 = n2635 & ~n10099 ;
  assign n10101 = n1017 & ~n10100 ;
  assign n10105 = n6295 ^ n2054 ^ n1401 ;
  assign n10103 = n2303 | n5260 ;
  assign n10104 = n464 & ~n10103 ;
  assign n10106 = n10105 ^ n10104 ^ n496 ;
  assign n10107 = n10106 ^ n8482 ^ n6882 ;
  assign n10102 = ~n177 & n2009 ;
  assign n10108 = n10107 ^ n10102 ^ 1'b0 ;
  assign n10109 = n1174 & ~n4650 ;
  assign n10110 = n10109 ^ n10055 ^ 1'b0 ;
  assign n10111 = n6046 & n9303 ;
  assign n10112 = n10111 ^ n6027 ^ 1'b0 ;
  assign n10113 = n3547 & n4482 ;
  assign n10114 = n10113 ^ n5157 ^ 1'b0 ;
  assign n10115 = ( n8061 & ~n8722 ) | ( n8061 & n10114 ) | ( ~n8722 & n10114 ) ;
  assign n10116 = n3987 ^ n1623 ^ 1'b0 ;
  assign n10117 = n5435 ^ n4514 ^ 1'b0 ;
  assign n10118 = n4082 & n10117 ;
  assign n10119 = ~n5647 & n7654 ;
  assign n10120 = n7881 & n10119 ;
  assign n10122 = n8341 ^ n5839 ^ 1'b0 ;
  assign n10123 = ~n5176 & n10122 ;
  assign n10121 = n163 & n9946 ;
  assign n10124 = n10123 ^ n10121 ^ 1'b0 ;
  assign n10125 = n5547 ^ n4348 ^ 1'b0 ;
  assign n10126 = n308 & ~n412 ;
  assign n10127 = n4798 & n10126 ;
  assign n10128 = n10127 ^ n2455 ^ 1'b0 ;
  assign n10129 = x43 | n10128 ;
  assign n10130 = ~n5974 & n8122 ;
  assign n10131 = n1625 | n10130 ;
  assign n10132 = n4443 & n6207 ;
  assign n10133 = n7518 ^ n4452 ^ 1'b0 ;
  assign n10134 = n6092 ^ n3493 ^ 1'b0 ;
  assign n10135 = n4387 ^ n1250 ^ 1'b0 ;
  assign n10136 = n3610 & n10135 ;
  assign n10137 = n4345 | n5481 ;
  assign n10138 = n10136 | n10137 ;
  assign n10139 = n8854 ^ n1439 ^ 1'b0 ;
  assign n10140 = ~n3295 & n10139 ;
  assign n10141 = ~n2088 & n8643 ;
  assign n10142 = n10141 ^ n9270 ^ 1'b0 ;
  assign n10143 = n8383 & ~n10142 ;
  assign n10144 = ~n10140 & n10143 ;
  assign n10145 = n6396 & n10144 ;
  assign n10146 = ~n3485 & n10145 ;
  assign n10148 = n1242 ^ n556 ^ x17 ;
  assign n10149 = n10148 ^ n8210 ^ 1'b0 ;
  assign n10147 = n1572 | n3834 ;
  assign n10150 = n10149 ^ n10147 ^ 1'b0 ;
  assign n10154 = ( ~n2559 & n3701 ) | ( ~n2559 & n8183 ) | ( n3701 & n8183 ) ;
  assign n10155 = n7822 ^ n3246 ^ 1'b0 ;
  assign n10156 = n10154 & n10155 ;
  assign n10151 = n916 | n3935 ;
  assign n10152 = n10151 ^ n9778 ^ 1'b0 ;
  assign n10153 = ~n4468 & n10152 ;
  assign n10157 = n10156 ^ n10153 ^ 1'b0 ;
  assign n10158 = n4686 & n8005 ;
  assign n10159 = ~n9942 & n10158 ;
  assign n10160 = n925 & n1507 ;
  assign n10161 = n10160 ^ n1906 ^ 1'b0 ;
  assign n10162 = n10161 ^ n1732 ^ 1'b0 ;
  assign n10163 = n2229 ^ n2176 ^ 1'b0 ;
  assign n10164 = n10163 ^ x43 ^ 1'b0 ;
  assign n10165 = n1711 | n10164 ;
  assign n10166 = n5365 ^ n1056 ^ 1'b0 ;
  assign n10167 = n4204 & ~n5011 ;
  assign n10168 = n10167 ^ n9197 ^ 1'b0 ;
  assign n10169 = n8803 | n10168 ;
  assign n10170 = n2431 | n3140 ;
  assign n10171 = n10170 ^ n4505 ^ 1'b0 ;
  assign n10172 = n1245 ^ n907 ^ 1'b0 ;
  assign n10173 = n10171 & n10172 ;
  assign n10174 = n10173 ^ n7861 ^ 1'b0 ;
  assign n10175 = n4513 & n9009 ;
  assign n10176 = n10175 ^ n4616 ^ 1'b0 ;
  assign n10177 = n4581 & n10176 ;
  assign n10178 = ~n695 & n10177 ;
  assign n10179 = n5787 ^ n4722 ^ 1'b0 ;
  assign n10180 = n8580 ^ n7164 ^ n2517 ;
  assign n10181 = n7577 ^ n6131 ^ 1'b0 ;
  assign n10182 = n4447 & n10181 ;
  assign n10183 = n9110 ^ n292 ^ 1'b0 ;
  assign n10184 = n5995 & ~n10183 ;
  assign n10185 = ~n3825 & n10184 ;
  assign n10186 = ~n4568 & n5044 ;
  assign n10187 = ~n4033 & n10186 ;
  assign n10188 = x119 & n934 ;
  assign n10189 = n10188 ^ n729 ^ 1'b0 ;
  assign n10190 = ~n8460 & n10189 ;
  assign n10191 = n10190 ^ n9998 ^ n3883 ;
  assign n10192 = n10191 ^ n3523 ^ 1'b0 ;
  assign n10193 = n1481 & n2912 ;
  assign n10194 = n1416 & ~n3222 ;
  assign n10195 = n10193 | n10194 ;
  assign n10196 = n10195 ^ n8545 ^ 1'b0 ;
  assign n10197 = n3475 & n6491 ;
  assign n10198 = n10197 ^ n1334 ^ 1'b0 ;
  assign n10199 = n10198 ^ n4843 ^ n2333 ;
  assign n10200 = n1145 & n8816 ;
  assign n10201 = ~n4441 & n5643 ;
  assign n10202 = ( n401 & n941 ) | ( n401 & n4622 ) | ( n941 & n4622 ) ;
  assign n10203 = ( ~n2231 & n3825 ) | ( ~n2231 & n3890 ) | ( n3825 & n3890 ) ;
  assign n10204 = n2931 ^ n388 ^ 1'b0 ;
  assign n10205 = ~n4182 & n10204 ;
  assign n10206 = ~n692 & n10205 ;
  assign n10207 = n243 & n10206 ;
  assign n10208 = ~n3938 & n5634 ;
  assign n10209 = ( n2945 & n5756 ) | ( n2945 & ~n5812 ) | ( n5756 & ~n5812 ) ;
  assign n10210 = n4305 | n10209 ;
  assign n10211 = n10210 ^ n4556 ^ 1'b0 ;
  assign n10212 = n3259 | n5494 ;
  assign n10213 = n10212 ^ n7189 ^ 1'b0 ;
  assign n10214 = n6634 ^ n3504 ^ 1'b0 ;
  assign n10215 = n540 & n934 ;
  assign n10216 = n10215 ^ x18 ^ 1'b0 ;
  assign n10217 = ~n9473 & n10216 ;
  assign n10218 = n10217 ^ n2583 ^ 1'b0 ;
  assign n10219 = ~n10214 & n10218 ;
  assign n10220 = n4354 & ~n6114 ;
  assign n10221 = n4434 | n6473 ;
  assign n10222 = n10221 ^ n1532 ^ 1'b0 ;
  assign n10223 = ~n4123 & n10222 ;
  assign n10224 = n10223 ^ n2142 ^ 1'b0 ;
  assign n10225 = n5945 ^ n4522 ^ n3562 ;
  assign n10226 = ~n1229 & n10225 ;
  assign n10227 = n2994 ^ n1803 ^ n204 ;
  assign n10228 = n10227 ^ n5234 ^ 1'b0 ;
  assign n10229 = n4250 & ~n10228 ;
  assign n10231 = n2903 & n3424 ;
  assign n10232 = ~n3770 & n10231 ;
  assign n10230 = n269 & ~n9267 ;
  assign n10233 = n10232 ^ n10230 ^ 1'b0 ;
  assign n10234 = n1440 | n1523 ;
  assign n10235 = n7880 & ~n10234 ;
  assign n10236 = ~n5544 & n6310 ;
  assign n10237 = ( ~n1167 & n3795 ) | ( ~n1167 & n10236 ) | ( n3795 & n10236 ) ;
  assign n10238 = n4452 & ~n6967 ;
  assign n10239 = n10238 ^ n2233 ^ 1'b0 ;
  assign n10240 = n3848 | n10239 ;
  assign n10241 = n7584 & ~n10240 ;
  assign n10242 = n6012 ^ n854 ^ 1'b0 ;
  assign n10243 = ~n7199 & n10242 ;
  assign n10244 = n10243 ^ n4143 ^ 1'b0 ;
  assign n10246 = n4295 ^ n3336 ^ 1'b0 ;
  assign n10247 = n10246 ^ n1576 ^ 1'b0 ;
  assign n10248 = n8987 | n10247 ;
  assign n10245 = n1745 & n2103 ;
  assign n10249 = n10248 ^ n10245 ^ 1'b0 ;
  assign n10250 = ( n2684 & n3385 ) | ( n2684 & n10249 ) | ( n3385 & n10249 ) ;
  assign n10251 = n1476 | n9311 ;
  assign n10252 = x37 & ~n8700 ;
  assign n10253 = n4115 ^ n2412 ^ n437 ;
  assign n10254 = n1017 & n10253 ;
  assign n10255 = x24 | n4769 ;
  assign n10256 = n10255 ^ n8335 ^ 1'b0 ;
  assign n10257 = n6667 & ~n10256 ;
  assign n10258 = n3625 | n6167 ;
  assign n10259 = n852 & n10258 ;
  assign n10260 = n6392 ^ n398 ^ 1'b0 ;
  assign n10261 = n2174 ^ n787 ^ 1'b0 ;
  assign n10262 = n10253 & n10261 ;
  assign n10264 = ~n368 & n3240 ;
  assign n10265 = ~n1728 & n10264 ;
  assign n10266 = n10265 ^ n2838 ^ 1'b0 ;
  assign n10267 = ~n999 & n10266 ;
  assign n10263 = ~n8075 & n8399 ;
  assign n10268 = n10267 ^ n10263 ^ n9987 ;
  assign n10269 = n6401 | n9909 ;
  assign n10270 = ~n1863 & n5850 ;
  assign n10271 = n1750 ^ x69 ^ 1'b0 ;
  assign n10273 = n6474 ^ n3102 ^ 1'b0 ;
  assign n10274 = ~n2914 & n10273 ;
  assign n10272 = ~n1611 & n5265 ;
  assign n10275 = n10274 ^ n10272 ^ 1'b0 ;
  assign n10276 = n2935 & ~n3834 ;
  assign n10277 = n1970 & ~n2575 ;
  assign n10278 = ~n814 & n10277 ;
  assign n10279 = n10278 ^ x38 ^ 1'b0 ;
  assign n10280 = n10276 | n10279 ;
  assign n10281 = n9410 ^ n1804 ^ 1'b0 ;
  assign n10282 = n10281 ^ n8314 ^ 1'b0 ;
  assign n10283 = n8343 & ~n10282 ;
  assign n10284 = ~n2131 & n10283 ;
  assign n10285 = ~n4613 & n10284 ;
  assign n10286 = n10285 ^ n3231 ^ 1'b0 ;
  assign n10287 = n1862 & ~n10286 ;
  assign n10288 = n5357 | n9465 ;
  assign n10289 = n632 & n7646 ;
  assign n10290 = n10289 ^ n3804 ^ 1'b0 ;
  assign n10291 = n4474 ^ n855 ^ 1'b0 ;
  assign n10292 = n2663 & n10291 ;
  assign n10293 = ( n1675 & n2062 ) | ( n1675 & n10292 ) | ( n2062 & n10292 ) ;
  assign n10295 = n3996 & ~n5426 ;
  assign n10294 = n6936 & ~n7944 ;
  assign n10296 = n10295 ^ n10294 ^ 1'b0 ;
  assign n10298 = n4917 & n5077 ;
  assign n10297 = n3023 | n10224 ;
  assign n10299 = n10298 ^ n10297 ^ 1'b0 ;
  assign n10300 = n5707 ^ n4277 ^ n3896 ;
  assign n10301 = n6611 ^ n6526 ^ 1'b0 ;
  assign n10302 = n4578 & ~n5685 ;
  assign n10303 = ~n4810 & n7678 ;
  assign n10304 = n10303 ^ x103 ^ 1'b0 ;
  assign n10305 = n10302 & n10304 ;
  assign n10306 = ~n1476 & n10305 ;
  assign n10307 = ~n10301 & n10306 ;
  assign n10313 = n9382 ^ n6681 ^ 1'b0 ;
  assign n10314 = ~n2627 & n10313 ;
  assign n10312 = n1716 & ~n3784 ;
  assign n10315 = n10314 ^ n10312 ^ 1'b0 ;
  assign n10308 = n8918 ^ n1515 ^ 1'b0 ;
  assign n10309 = n6049 ^ n1070 ^ 1'b0 ;
  assign n10310 = ~n7521 & n10309 ;
  assign n10311 = n10308 & n10310 ;
  assign n10316 = n10315 ^ n10311 ^ 1'b0 ;
  assign n10317 = ~n1495 & n10316 ;
  assign n10319 = ~n2170 & n2462 ;
  assign n10320 = n10319 ^ n2593 ^ 1'b0 ;
  assign n10321 = n10320 ^ n5563 ^ n2911 ;
  assign n10318 = n747 & ~n994 ;
  assign n10322 = n10321 ^ n10318 ^ 1'b0 ;
  assign n10323 = n1124 & ~n2206 ;
  assign n10324 = n3344 & n8129 ;
  assign n10325 = ~n4814 & n10324 ;
  assign n10326 = n7553 | n10325 ;
  assign n10327 = n10326 ^ n8942 ^ 1'b0 ;
  assign n10328 = ( x71 & n2222 ) | ( x71 & n3278 ) | ( n2222 & n3278 ) ;
  assign n10329 = n1370 & n4041 ;
  assign n10330 = n10329 ^ n2128 ^ 1'b0 ;
  assign n10331 = n7319 & ~n7416 ;
  assign n10332 = n10330 & ~n10331 ;
  assign n10333 = ~n442 & n2627 ;
  assign n10334 = n2988 & ~n8971 ;
  assign n10335 = n10334 ^ n2654 ^ 1'b0 ;
  assign n10336 = ~n10333 & n10335 ;
  assign n10338 = n543 & n2218 ;
  assign n10339 = ~n509 & n10338 ;
  assign n10337 = n6877 & n6997 ;
  assign n10340 = n10339 ^ n10337 ^ 1'b0 ;
  assign n10341 = n2265 & n3476 ;
  assign n10342 = ~n2477 & n10341 ;
  assign n10343 = n1522 & ~n2399 ;
  assign n10344 = n10342 & n10343 ;
  assign n10345 = n10344 ^ n3604 ^ n577 ;
  assign n10346 = n10345 ^ n4330 ^ 1'b0 ;
  assign n10347 = n4558 ^ n2992 ^ 1'b0 ;
  assign n10348 = n10347 ^ n10295 ^ 1'b0 ;
  assign n10349 = n1163 & ~n6187 ;
  assign n10350 = ~n1463 & n10349 ;
  assign n10351 = n10350 ^ n8646 ^ 1'b0 ;
  assign n10352 = n2178 & n4678 ;
  assign n10353 = ~n4192 & n8165 ;
  assign n10354 = n10353 ^ n7866 ^ 1'b0 ;
  assign n10355 = n10352 & ~n10354 ;
  assign n10362 = n6125 ^ n5977 ^ 1'b0 ;
  assign n10356 = n1084 & ~n1633 ;
  assign n10357 = n2298 & n10356 ;
  assign n10360 = ( n2399 & n5427 ) | ( n2399 & n10357 ) | ( n5427 & n10357 ) ;
  assign n10361 = n10360 ^ n7383 ^ 1'b0 ;
  assign n10358 = n10357 ^ n2956 ^ 1'b0 ;
  assign n10359 = n357 & ~n10358 ;
  assign n10363 = n10362 ^ n10361 ^ n10359 ;
  assign n10364 = n4168 ^ n3530 ^ n2113 ;
  assign n10365 = n2353 & ~n10364 ;
  assign n10366 = n8210 ^ n1495 ^ 1'b0 ;
  assign n10367 = n2679 ^ n303 ^ 1'b0 ;
  assign n10368 = n3086 | n10367 ;
  assign n10369 = n10368 ^ n8164 ^ 1'b0 ;
  assign n10370 = ~n10263 & n10369 ;
  assign n10371 = n8195 ^ n5805 ^ 1'b0 ;
  assign n10372 = n8278 ^ n7975 ^ 1'b0 ;
  assign n10373 = n5148 ^ n278 ^ 1'b0 ;
  assign n10374 = n4806 & ~n9382 ;
  assign n10375 = n10374 ^ n6773 ^ 1'b0 ;
  assign n10376 = n1137 & ~n3910 ;
  assign n10377 = n10376 ^ n1370 ^ 1'b0 ;
  assign n10378 = n10377 ^ n5511 ^ 1'b0 ;
  assign n10379 = ~n2308 & n10378 ;
  assign n10380 = n10379 ^ n4614 ^ 1'b0 ;
  assign n10381 = n3592 | n10380 ;
  assign n10382 = n1975 ^ n246 ^ 1'b0 ;
  assign n10383 = n10382 ^ n6498 ^ 1'b0 ;
  assign n10384 = n5901 & n10383 ;
  assign n10385 = ~n6050 & n6478 ;
  assign n10386 = ~n10384 & n10385 ;
  assign n10387 = n257 & ~n9080 ;
  assign n10388 = n1556 ^ n240 ^ 1'b0 ;
  assign n10389 = n7110 ^ n2654 ^ n1225 ;
  assign n10390 = ~n4458 & n7470 ;
  assign n10391 = n10390 ^ n1899 ^ 1'b0 ;
  assign n10392 = n10389 & n10391 ;
  assign n10393 = n2622 | n8206 ;
  assign n10394 = n2324 | n10393 ;
  assign n10395 = n10201 ^ n1079 ^ 1'b0 ;
  assign n10396 = n2332 ^ n1270 ^ 1'b0 ;
  assign n10397 = n2461 & n10396 ;
  assign n10398 = n9628 | n10397 ;
  assign n10399 = n1188 & n2667 ;
  assign n10400 = n3815 & ~n10399 ;
  assign n10401 = n10400 ^ n9154 ^ 1'b0 ;
  assign n10402 = n281 & ~n1560 ;
  assign n10403 = n3990 ^ n577 ^ 1'b0 ;
  assign n10404 = n4418 & n10403 ;
  assign n10405 = n10404 ^ n6159 ^ n5136 ;
  assign n10406 = n10405 ^ n7112 ^ 1'b0 ;
  assign n10407 = n1431 & ~n10406 ;
  assign n10408 = n5073 ^ n2830 ^ 1'b0 ;
  assign n10409 = n10408 ^ n9389 ^ n3557 ;
  assign n10410 = ~n4975 & n10409 ;
  assign n10411 = n10410 ^ n2492 ^ 1'b0 ;
  assign n10412 = ~n4808 & n10008 ;
  assign n10413 = n10412 ^ n3789 ^ 1'b0 ;
  assign n10414 = n4438 | n10331 ;
  assign n10415 = n5840 ^ n3940 ^ 1'b0 ;
  assign n10416 = ( n1163 & ~n1670 ) | ( n1163 & n10333 ) | ( ~n1670 & n10333 ) ;
  assign n10417 = n10416 ^ n7558 ^ n2694 ;
  assign n10418 = n6914 & ~n10417 ;
  assign n10419 = n10418 ^ n1623 ^ 1'b0 ;
  assign n10420 = n1821 & ~n10419 ;
  assign n10421 = n4413 & ~n10332 ;
  assign n10422 = ~x94 & n10421 ;
  assign n10423 = n2087 | n5578 ;
  assign n10424 = n3276 & ~n10423 ;
  assign n10425 = n1867 & n2689 ;
  assign n10426 = n1509 ^ n1327 ^ 1'b0 ;
  assign n10427 = n10426 ^ n6778 ^ n2470 ;
  assign n10428 = n4947 ^ n4345 ^ 1'b0 ;
  assign n10429 = n4562 & ~n10428 ;
  assign n10430 = ~n3408 & n6485 ;
  assign n10431 = ~n10429 & n10430 ;
  assign n10432 = n3148 ^ n1237 ^ 1'b0 ;
  assign n10433 = n6093 & n10432 ;
  assign n10434 = n1895 ^ n369 ^ 1'b0 ;
  assign n10435 = n9392 & n10434 ;
  assign n10436 = ~n1211 & n2807 ;
  assign n10437 = n2537 & n10436 ;
  assign n10438 = n1995 & ~n10437 ;
  assign n10439 = n10437 & n10438 ;
  assign n10440 = n6734 & ~n10439 ;
  assign n10441 = n10440 ^ n4618 ^ 1'b0 ;
  assign n10442 = n297 & ~n5315 ;
  assign n10443 = n7006 & n10442 ;
  assign n10444 = n2639 ^ n1383 ^ 1'b0 ;
  assign n10445 = ( ~n2922 & n4159 ) | ( ~n2922 & n7855 ) | ( n4159 & n7855 ) ;
  assign n10446 = n8534 ^ n3818 ^ 1'b0 ;
  assign n10447 = ~n10445 & n10446 ;
  assign n10448 = ~n1927 & n9138 ;
  assign n10449 = n1283 | n8430 ;
  assign n10450 = n10449 ^ n2894 ^ 1'b0 ;
  assign n10451 = ~n456 & n10450 ;
  assign n10452 = n10451 ^ n3552 ^ 1'b0 ;
  assign n10453 = ( n829 & n4203 ) | ( n829 & n9955 ) | ( n4203 & n9955 ) ;
  assign n10454 = n6087 & n9323 ;
  assign n10455 = n10454 ^ n3065 ^ 1'b0 ;
  assign n10456 = n6569 ^ n6561 ^ 1'b0 ;
  assign n10457 = n10455 & ~n10456 ;
  assign n10458 = n8654 | n9454 ;
  assign n10459 = n10458 ^ n9471 ^ 1'b0 ;
  assign n10460 = n4324 & ~n8809 ;
  assign n10461 = n6695 ^ n1410 ^ 1'b0 ;
  assign n10462 = n10416 & ~n10461 ;
  assign n10463 = n5974 ^ n1741 ^ 1'b0 ;
  assign n10464 = n2481 & ~n6111 ;
  assign n10465 = n833 & n10464 ;
  assign n10466 = n10463 & n10465 ;
  assign n10469 = n2462 & ~n4418 ;
  assign n10467 = n646 & ~n1452 ;
  assign n10468 = n10467 ^ n3603 ^ 1'b0 ;
  assign n10470 = n10469 ^ n10468 ^ n4162 ;
  assign n10471 = n10470 ^ n1199 ^ 1'b0 ;
  assign n10472 = n241 & ~n5482 ;
  assign n10473 = n7793 ^ n4395 ^ 1'b0 ;
  assign n10474 = ~n6472 & n10473 ;
  assign n10475 = n10472 & n10474 ;
  assign n10476 = x50 & n10475 ;
  assign n10477 = n3550 ^ n152 ^ 1'b0 ;
  assign n10478 = n4657 | n9858 ;
  assign n10479 = n1588 | n3517 ;
  assign n10480 = n1439 & ~n10479 ;
  assign n10481 = ~n1871 & n10480 ;
  assign n10484 = n143 & ~n3601 ;
  assign n10485 = n10484 ^ n729 ^ 1'b0 ;
  assign n10483 = n1051 | n6151 ;
  assign n10486 = n10485 ^ n10483 ^ 1'b0 ;
  assign n10487 = n998 & n3781 ;
  assign n10488 = n10487 ^ n4335 ^ 1'b0 ;
  assign n10489 = n10486 | n10488 ;
  assign n10482 = ~n2105 & n3217 ;
  assign n10490 = n10489 ^ n10482 ^ 1'b0 ;
  assign n10491 = n8855 & ~n10490 ;
  assign n10492 = ~n254 & n2735 ;
  assign n10493 = n569 & ~n609 ;
  assign n10494 = ~n4731 & n10493 ;
  assign n10495 = n1198 & ~n9431 ;
  assign n10496 = ~n628 & n10495 ;
  assign n10497 = ~n8598 & n8832 ;
  assign n10498 = n3605 ^ n607 ^ 1'b0 ;
  assign n10499 = ~n272 & n10498 ;
  assign n10500 = ~n5696 & n10499 ;
  assign n10501 = ~n9826 & n10500 ;
  assign n10502 = n10501 ^ n1679 ^ x17 ;
  assign n10503 = n10502 ^ n3641 ^ 1'b0 ;
  assign n10504 = n4265 & ~n5741 ;
  assign n10505 = n2603 ^ n1225 ^ 1'b0 ;
  assign n10506 = n3511 & ~n10505 ;
  assign n10507 = n10506 ^ n5431 ^ 1'b0 ;
  assign n10508 = n1993 ^ n262 ^ 1'b0 ;
  assign n10509 = n10507 & n10508 ;
  assign n10513 = n675 & ~n5159 ;
  assign n10514 = ~n5909 & n10513 ;
  assign n10510 = n2521 & n2670 ;
  assign n10511 = ~n2113 & n10510 ;
  assign n10512 = ~n7991 & n10511 ;
  assign n10515 = n10514 ^ n10512 ^ 1'b0 ;
  assign n10516 = n1340 & n2144 ;
  assign n10517 = n10516 ^ n4981 ^ n159 ;
  assign n10518 = n7948 & ~n8856 ;
  assign n10519 = n10518 ^ n8425 ^ 1'b0 ;
  assign n10520 = n1766 ^ n767 ^ 1'b0 ;
  assign n10521 = n7595 ^ n1450 ^ 1'b0 ;
  assign n10522 = n8475 & n10521 ;
  assign n10523 = n6352 & n10522 ;
  assign n10524 = n5348 ^ n1309 ^ 1'b0 ;
  assign n10525 = ~n3054 & n10524 ;
  assign n10526 = n10001 ^ n7264 ^ 1'b0 ;
  assign n10527 = ~x67 & n8541 ;
  assign n10528 = ~n10526 & n10527 ;
  assign n10529 = n2982 | n10528 ;
  assign n10530 = n6111 ^ n3651 ^ 1'b0 ;
  assign n10531 = n10530 ^ n9817 ^ 1'b0 ;
  assign n10532 = n2028 | n10531 ;
  assign n10533 = n656 & ~n8608 ;
  assign n10534 = n10533 ^ n4243 ^ 1'b0 ;
  assign n10535 = n9380 & ~n10534 ;
  assign n10536 = n6025 ^ n5882 ^ 1'b0 ;
  assign n10537 = n4632 ^ n2413 ^ 1'b0 ;
  assign n10538 = n9441 & ~n10537 ;
  assign n10539 = n7401 ^ n163 ^ 1'b0 ;
  assign n10540 = n9408 & n10539 ;
  assign n10541 = n3517 & n10540 ;
  assign n10542 = ~n509 & n1832 ;
  assign n10543 = n3773 & ~n8415 ;
  assign n10544 = n10543 ^ n9923 ^ 1'b0 ;
  assign n10545 = n4100 ^ n1177 ^ n453 ;
  assign n10546 = n6270 & n10545 ;
  assign n10547 = n4922 & n10546 ;
  assign n10553 = n4264 | n8558 ;
  assign n10550 = n4257 ^ n2146 ^ n820 ;
  assign n10551 = ( n3226 & n7052 ) | ( n3226 & n10550 ) | ( n7052 & n10550 ) ;
  assign n10548 = n2046 & n4510 ;
  assign n10549 = n7666 & n10548 ;
  assign n10552 = n10551 ^ n10549 ^ 1'b0 ;
  assign n10554 = n10553 ^ n10552 ^ n6786 ;
  assign n10555 = n4662 & n7442 ;
  assign n10556 = ~n909 & n9868 ;
  assign n10557 = n10556 ^ n6663 ^ 1'b0 ;
  assign n10560 = n5000 | n9703 ;
  assign n10561 = n1913 & ~n10560 ;
  assign n10558 = n6455 & ~n7946 ;
  assign n10559 = n4048 | n10558 ;
  assign n10562 = n10561 ^ n10559 ^ 1'b0 ;
  assign n10563 = n809 ^ x53 ^ 1'b0 ;
  assign n10564 = ~n2947 & n10563 ;
  assign n10565 = n4348 ^ n1136 ^ 1'b0 ;
  assign n10566 = n10564 | n10565 ;
  assign n10567 = n6423 ^ n249 ^ 1'b0 ;
  assign n10568 = ~n9640 & n10567 ;
  assign n10569 = n2317 ^ x98 ^ 1'b0 ;
  assign n10570 = n8500 & ~n10569 ;
  assign n10571 = n10570 ^ n1999 ^ 1'b0 ;
  assign n10572 = n468 & n3632 ;
  assign n10573 = ( n3437 & n5530 ) | ( n3437 & n10572 ) | ( n5530 & n10572 ) ;
  assign n10574 = n10573 ^ n7932 ^ n2910 ;
  assign n10575 = ~n2130 & n10574 ;
  assign n10576 = n6974 ^ n4840 ^ 1'b0 ;
  assign n10577 = x67 & n10576 ;
  assign n10578 = n3590 | n10577 ;
  assign n10579 = ~n8688 & n10578 ;
  assign n10580 = n6757 | n10579 ;
  assign n10581 = ~n2012 & n3726 ;
  assign n10582 = ~n1241 & n3274 ;
  assign n10583 = n444 | n6957 ;
  assign n10584 = ~n3832 & n4630 ;
  assign n10585 = n10584 ^ n5424 ^ 1'b0 ;
  assign n10586 = n4950 & n10585 ;
  assign n10587 = n5345 & n8862 ;
  assign n10588 = n3373 | n10587 ;
  assign n10589 = n10588 ^ n10120 ^ 1'b0 ;
  assign n10590 = n7392 ^ n4179 ^ 1'b0 ;
  assign n10591 = ~n4009 & n10590 ;
  assign n10592 = ~n10204 & n10591 ;
  assign n10594 = n4657 ^ x79 ^ 1'b0 ;
  assign n10593 = n3164 & ~n3365 ;
  assign n10595 = n10594 ^ n10593 ^ 1'b0 ;
  assign n10596 = n7644 & ~n10595 ;
  assign n10597 = n236 | n3746 ;
  assign n10598 = n404 | n10597 ;
  assign n10599 = n969 & n9988 ;
  assign n10600 = n10599 ^ n8301 ^ n852 ;
  assign n10601 = n2633 | n3175 ;
  assign n10602 = n5815 | n10601 ;
  assign n10603 = x22 & n1865 ;
  assign n10605 = ( n2949 & ~n3465 ) | ( n2949 & n8247 ) | ( ~n3465 & n8247 ) ;
  assign n10606 = n10605 ^ n4359 ^ 1'b0 ;
  assign n10604 = n4776 & n10551 ;
  assign n10607 = n10606 ^ n10604 ^ 1'b0 ;
  assign n10608 = n10607 ^ n8395 ^ n1834 ;
  assign n10609 = n10608 ^ n417 ^ 1'b0 ;
  assign n10610 = n2731 & n10346 ;
  assign n10611 = ~n2078 & n7399 ;
  assign n10612 = n1953 & n10611 ;
  assign n10613 = n6020 ^ n4614 ^ 1'b0 ;
  assign n10614 = n10612 | n10613 ;
  assign n10615 = n3274 ^ n2543 ^ 1'b0 ;
  assign n10616 = n10615 ^ n8124 ^ 1'b0 ;
  assign n10617 = n6898 & ~n10516 ;
  assign n10618 = n10617 ^ n1698 ^ 1'b0 ;
  assign n10619 = n1193 | n10618 ;
  assign n10620 = n2838 | n5262 ;
  assign n10621 = n2838 & ~n10620 ;
  assign n10622 = n3657 | n10621 ;
  assign n10623 = n5870 & ~n10622 ;
  assign n10624 = n2022 & ~n10623 ;
  assign n10625 = n10624 ^ n2546 ^ 1'b0 ;
  assign n10626 = n2359 & ~n10625 ;
  assign n10627 = ~n719 & n10626 ;
  assign n10628 = n3240 & n8322 ;
  assign n10629 = n9959 ^ n3054 ^ 1'b0 ;
  assign n10630 = n3935 & ~n10629 ;
  assign n10631 = n9620 ^ n3576 ^ 1'b0 ;
  assign n10632 = ~n10398 & n10631 ;
  assign n10633 = n4708 ^ n4157 ^ 1'b0 ;
  assign n10634 = n10633 ^ n10453 ^ 1'b0 ;
  assign n10635 = n7321 ^ n7250 ^ 1'b0 ;
  assign n10636 = n7023 ^ n6212 ^ 1'b0 ;
  assign n10637 = x18 & n10636 ;
  assign n10638 = n9725 & ~n9850 ;
  assign n10639 = n171 | n3892 ;
  assign n10640 = n3558 & ~n10639 ;
  assign n10641 = n2579 & ~n3666 ;
  assign n10642 = ~n10640 & n10641 ;
  assign n10643 = n1089 & n10642 ;
  assign n10644 = n8804 | n10643 ;
  assign n10645 = n3431 ^ n2235 ^ 1'b0 ;
  assign n10646 = n4740 ^ n681 ^ 1'b0 ;
  assign n10647 = ~n2491 & n10646 ;
  assign n10648 = n2322 & n3262 ;
  assign n10649 = n9303 & n10648 ;
  assign n10650 = n5764 | n10649 ;
  assign n10651 = n6501 & n8273 ;
  assign n10652 = ~n3968 & n10651 ;
  assign n10653 = n973 | n10652 ;
  assign n10654 = n6836 | n10653 ;
  assign n10655 = n2293 ^ n2221 ^ 1'b0 ;
  assign n10656 = n2418 & n10655 ;
  assign n10657 = ~n4139 & n10656 ;
  assign n10658 = n1001 | n10657 ;
  assign n10659 = n10654 | n10658 ;
  assign n10660 = n5647 ^ n1084 ^ 1'b0 ;
  assign n10661 = n4564 & ~n4727 ;
  assign n10662 = n363 & n10661 ;
  assign n10663 = n2927 & ~n10662 ;
  assign n10664 = n3102 & n10663 ;
  assign n10665 = n10664 ^ n4538 ^ 1'b0 ;
  assign n10667 = n591 & ~n6230 ;
  assign n10668 = n1176 & n10667 ;
  assign n10666 = n8436 & n10024 ;
  assign n10669 = n10668 ^ n10666 ^ 1'b0 ;
  assign n10670 = n4053 ^ n3467 ^ n1271 ;
  assign n10671 = n10670 ^ n2088 ^ 1'b0 ;
  assign n10673 = x37 & ~n6794 ;
  assign n10672 = n1337 & n8415 ;
  assign n10674 = n10673 ^ n10672 ^ 1'b0 ;
  assign n10675 = n6655 ^ n600 ^ 1'b0 ;
  assign n10676 = n5029 ^ n1959 ^ 1'b0 ;
  assign n10677 = ~n9606 & n10676 ;
  assign n10678 = n5043 & n8957 ;
  assign n10679 = n180 | n8443 ;
  assign n10680 = n4222 & n4472 ;
  assign n10681 = n10680 ^ n7640 ^ 1'b0 ;
  assign n10682 = n4924 | n8817 ;
  assign n10683 = n10682 ^ n9141 ^ 1'b0 ;
  assign n10684 = n10683 ^ n6082 ^ 1'b0 ;
  assign n10685 = ~n3442 & n10684 ;
  assign n10686 = n5935 ^ n5891 ^ n3313 ;
  assign n10689 = n2417 ^ n555 ^ 1'b0 ;
  assign n10687 = n1632 & n6663 ;
  assign n10688 = ~n9973 & n10687 ;
  assign n10690 = n10689 ^ n10688 ^ 1'b0 ;
  assign n10691 = n7865 ^ n4736 ^ 1'b0 ;
  assign n10692 = n431 & n3450 ;
  assign n10693 = n4987 | n10692 ;
  assign n10694 = n10693 ^ n5899 ^ 1'b0 ;
  assign n10695 = n3755 & ~n4516 ;
  assign n10696 = n4347 & ~n4585 ;
  assign n10697 = n10696 ^ n9715 ^ 1'b0 ;
  assign n10698 = n3274 | n10697 ;
  assign n10699 = n10695 & ~n10698 ;
  assign n10700 = ( n7426 & n10694 ) | ( n7426 & ~n10699 ) | ( n10694 & ~n10699 ) ;
  assign n10701 = n4686 & ~n8268 ;
  assign n10702 = n2303 | n10701 ;
  assign n10703 = ~n1545 & n6744 ;
  assign n10704 = n4942 & ~n7879 ;
  assign n10705 = n5016 & ~n7631 ;
  assign n10706 = n2758 & ~n2788 ;
  assign n10707 = n3070 & n10706 ;
  assign n10708 = n3653 & n10707 ;
  assign n10709 = n10708 ^ x58 ^ 1'b0 ;
  assign n10710 = n2010 | n3699 ;
  assign n10711 = n5905 & ~n9228 ;
  assign n10712 = n1582 & n10711 ;
  assign n10713 = n8323 | n10712 ;
  assign n10714 = n10713 ^ n3633 ^ 1'b0 ;
  assign n10715 = ~n770 & n9182 ;
  assign n10716 = n10715 ^ n8337 ^ 1'b0 ;
  assign n10719 = n813 | n2809 ;
  assign n10720 = n10719 ^ n3564 ^ 1'b0 ;
  assign n10717 = ~n3869 & n6821 ;
  assign n10718 = n5962 & n10717 ;
  assign n10721 = n10720 ^ n10718 ^ n2945 ;
  assign n10722 = n3411 & n9909 ;
  assign n10723 = n8344 ^ n4765 ^ n939 ;
  assign n10724 = n8294 & ~n10723 ;
  assign n10725 = ~n7336 & n10724 ;
  assign n10726 = n1057 | n4769 ;
  assign n10727 = n5944 & n7036 ;
  assign n10728 = n2380 ^ n2018 ^ 1'b0 ;
  assign n10729 = n10728 ^ n4139 ^ 1'b0 ;
  assign n10730 = n3700 ^ n475 ^ 1'b0 ;
  assign n10731 = ~n5036 & n10730 ;
  assign n10732 = n10729 & n10731 ;
  assign n10733 = n2496 | n6266 ;
  assign n10734 = n10733 ^ n2428 ^ 1'b0 ;
  assign n10735 = n3061 ^ n326 ^ 1'b0 ;
  assign n10736 = n10734 & n10735 ;
  assign n10737 = n208 | n10061 ;
  assign n10738 = ~n5311 & n5819 ;
  assign n10739 = n10738 ^ n9050 ^ 1'b0 ;
  assign n10742 = n4675 | n7534 ;
  assign n10743 = n10742 ^ n1563 ^ 1'b0 ;
  assign n10740 = n2182 ^ n1891 ^ 1'b0 ;
  assign n10741 = n8227 & n10740 ;
  assign n10744 = n10743 ^ n10741 ^ 1'b0 ;
  assign n10745 = n7600 ^ n6225 ^ 1'b0 ;
  assign n10746 = n7245 ^ n1485 ^ 1'b0 ;
  assign n10747 = ~n10745 & n10746 ;
  assign n10748 = ~n6052 & n10747 ;
  assign n10749 = n3648 & ~n4838 ;
  assign n10750 = ~n10748 & n10749 ;
  assign n10751 = ~n2932 & n7854 ;
  assign n10752 = n3733 & ~n4395 ;
  assign n10753 = n10752 ^ n7984 ^ 1'b0 ;
  assign n10754 = ~n10715 & n10753 ;
  assign n10755 = ~n1825 & n7688 ;
  assign n10756 = ~n381 & n1157 ;
  assign n10757 = n10756 ^ n1888 ^ 1'b0 ;
  assign n10758 = n7083 ^ n1590 ^ n719 ;
  assign n10759 = n3072 & n10758 ;
  assign n10760 = n4983 & ~n6681 ;
  assign n10761 = ~n3122 & n10760 ;
  assign n10762 = n8457 ^ n632 ^ 1'b0 ;
  assign n10763 = n10761 | n10762 ;
  assign n10764 = n10763 ^ n6442 ^ 1'b0 ;
  assign n10765 = n10759 & n10764 ;
  assign n10766 = n6523 ^ n6107 ^ 1'b0 ;
  assign n10767 = ~n3999 & n10766 ;
  assign n10768 = n8248 | n10767 ;
  assign n10769 = n9008 ^ n7012 ^ 1'b0 ;
  assign n10770 = n1774 & ~n3533 ;
  assign n10771 = n10770 ^ n163 ^ 1'b0 ;
  assign n10772 = n10769 & ~n10771 ;
  assign n10773 = n10768 & n10772 ;
  assign n10774 = n890 | n1250 ;
  assign n10775 = n9763 ^ n643 ^ 1'b0 ;
  assign n10776 = n10775 ^ n4781 ^ 1'b0 ;
  assign n10777 = n10720 & n10776 ;
  assign n10778 = ~n6568 & n6584 ;
  assign n10779 = n6044 & n10778 ;
  assign n10780 = n9590 & n10779 ;
  assign n10781 = ~n6469 & n8601 ;
  assign n10782 = n10781 ^ n3328 ^ 1'b0 ;
  assign n10783 = ( ~x48 & n4765 ) | ( ~x48 & n10782 ) | ( n4765 & n10782 ) ;
  assign n10784 = n2477 & ~n3124 ;
  assign n10788 = n1804 | n5164 ;
  assign n10789 = n8403 | n10788 ;
  assign n10785 = x119 & n3982 ;
  assign n10786 = n3411 & n10785 ;
  assign n10787 = n8749 | n10786 ;
  assign n10790 = n10789 ^ n10787 ^ 1'b0 ;
  assign n10791 = n10784 & n10790 ;
  assign n10792 = n3550 ^ n762 ^ 1'b0 ;
  assign n10793 = n10791 & n10792 ;
  assign n10794 = n1391 | n1718 ;
  assign n10795 = n4301 | n10794 ;
  assign n10796 = n10795 ^ n9924 ^ 1'b0 ;
  assign n10798 = n397 | n10695 ;
  assign n10797 = n3226 & n6540 ;
  assign n10799 = n10798 ^ n10797 ^ 1'b0 ;
  assign n10800 = n3013 & ~n10799 ;
  assign n10801 = n10796 & n10800 ;
  assign n10802 = n2798 & n10343 ;
  assign n10803 = n10802 ^ n8841 ^ 1'b0 ;
  assign n10804 = n5561 ^ n4994 ^ n1295 ;
  assign n10805 = n2265 & n10804 ;
  assign n10806 = ( n1017 & n1259 ) | ( n1017 & n1909 ) | ( n1259 & n1909 ) ;
  assign n10807 = n2466 ^ n755 ^ 1'b0 ;
  assign n10808 = n243 | n10807 ;
  assign n10809 = n10806 & ~n10808 ;
  assign n10810 = ~n2113 & n3565 ;
  assign n10811 = n10809 & n10810 ;
  assign n10812 = n10811 ^ n1975 ^ n180 ;
  assign n10813 = ~n1076 & n7629 ;
  assign n10814 = ~n2965 & n10813 ;
  assign n10815 = n10814 ^ n4590 ^ 1'b0 ;
  assign n10816 = n10815 ^ n3951 ^ 1'b0 ;
  assign n10817 = n6055 ^ n4733 ^ 1'b0 ;
  assign n10818 = n7207 ^ n2953 ^ n597 ;
  assign n10819 = ~n5594 & n10670 ;
  assign n10824 = n2128 ^ n1535 ^ 1'b0 ;
  assign n10825 = n1488 | n10824 ;
  assign n10821 = ~n4502 & n6168 ;
  assign n10822 = n10821 ^ n7319 ^ 1'b0 ;
  assign n10823 = ~n7723 & n10822 ;
  assign n10820 = x40 | n529 ;
  assign n10826 = n10825 ^ n10823 ^ n10820 ;
  assign n10827 = n5163 | n5262 ;
  assign n10828 = n2084 | n10827 ;
  assign n10829 = n6195 ^ n1893 ^ 1'b0 ;
  assign n10830 = n334 & n2862 ;
  assign n10831 = n10830 ^ n3041 ^ 1'b0 ;
  assign n10832 = n7080 & ~n10831 ;
  assign n10833 = n10832 ^ n3687 ^ 1'b0 ;
  assign n10834 = ~n3547 & n4336 ;
  assign n10835 = n10834 ^ n2131 ^ 1'b0 ;
  assign n10836 = n143 & ~n344 ;
  assign n10837 = n8116 ^ n1705 ^ 1'b0 ;
  assign n10838 = ~n2925 & n3135 ;
  assign n10839 = ( n471 & n10837 ) | ( n471 & ~n10838 ) | ( n10837 & ~n10838 ) ;
  assign n10840 = x102 | n8286 ;
  assign n10842 = n3465 & ~n4089 ;
  assign n10841 = ~n3724 & n5958 ;
  assign n10843 = n10842 ^ n10841 ^ 1'b0 ;
  assign n10844 = ~n10840 & n10843 ;
  assign n10845 = ~n9823 & n10283 ;
  assign n10846 = n157 & n6646 ;
  assign n10847 = ~n530 & n10846 ;
  assign n10848 = n2946 ^ n456 ^ 1'b0 ;
  assign n10849 = n10453 ^ n8643 ^ 1'b0 ;
  assign n10850 = n7170 ^ n5157 ^ 1'b0 ;
  assign n10851 = n10850 ^ n6449 ^ 1'b0 ;
  assign n10852 = n10851 ^ n10368 ^ 1'b0 ;
  assign n10853 = n5763 ^ n5277 ^ 1'b0 ;
  assign n10854 = n4213 | n10853 ;
  assign n10855 = n1258 | n3270 ;
  assign n10856 = n3391 & ~n10855 ;
  assign n10857 = ~n1031 & n5035 ;
  assign n10858 = ( ~n3311 & n10856 ) | ( ~n3311 & n10857 ) | ( n10856 & n10857 ) ;
  assign n10859 = n4289 ^ n3021 ^ 1'b0 ;
  assign n10860 = n9517 | n10707 ;
  assign n10861 = n10860 ^ n2632 ^ 1'b0 ;
  assign n10862 = ~n7419 & n8810 ;
  assign n10863 = n7512 & n10862 ;
  assign n10864 = ~n2603 & n10863 ;
  assign n10865 = n143 & n1811 ;
  assign n10866 = n10865 ^ n7371 ^ n7023 ;
  assign n10867 = n6493 ^ n577 ^ 1'b0 ;
  assign n10868 = ~n4001 & n6416 ;
  assign n10869 = n188 & n5783 ;
  assign n10870 = n3386 & n9686 ;
  assign n10871 = n10869 & n10870 ;
  assign n10872 = n1888 & ~n7293 ;
  assign n10873 = n3646 | n9625 ;
  assign n10874 = n1147 & ~n10873 ;
  assign n10875 = ~n4478 & n10874 ;
  assign n10876 = n4877 ^ n2080 ^ 1'b0 ;
  assign n10877 = n10876 ^ n381 ^ 1'b0 ;
  assign n10878 = n3618 ^ n3214 ^ n1150 ;
  assign n10879 = n5230 | n10878 ;
  assign n10880 = x6 | n10879 ;
  assign n10881 = n10880 ^ n1804 ^ 1'b0 ;
  assign n10882 = n10522 & n10881 ;
  assign n10883 = n10882 ^ n7931 ^ 1'b0 ;
  assign n10884 = n5952 | n10883 ;
  assign n10885 = n4566 ^ n1576 ^ 1'b0 ;
  assign n10886 = n10885 ^ n7305 ^ 1'b0 ;
  assign n10887 = ~n7078 & n10886 ;
  assign n10888 = n10887 ^ n7534 ^ 1'b0 ;
  assign n10889 = n10888 ^ n10592 ^ 1'b0 ;
  assign n10890 = n8061 & ~n8897 ;
  assign n10891 = ~n1355 & n10890 ;
  assign n10892 = n9345 | n10891 ;
  assign n10893 = ~n145 & n6991 ;
  assign n10894 = n10893 ^ n4036 ^ 1'b0 ;
  assign n10895 = n5220 ^ n4287 ^ 1'b0 ;
  assign n10896 = n1033 & ~n9075 ;
  assign n10897 = ~n2987 & n5124 ;
  assign n10898 = n5442 & ~n8648 ;
  assign n10899 = ~n10897 & n10898 ;
  assign n10900 = n9071 ^ x98 ^ 1'b0 ;
  assign n10901 = ( n973 & n8262 ) | ( n973 & ~n10900 ) | ( n8262 & ~n10900 ) ;
  assign n10902 = n10615 ^ n1479 ^ 1'b0 ;
  assign n10903 = n8747 & ~n10902 ;
  assign n10904 = n3820 ^ n1695 ^ n273 ;
  assign n10905 = ~n3171 & n6145 ;
  assign n10906 = ~n10904 & n10905 ;
  assign n10907 = ~n1582 & n2462 ;
  assign n10908 = ~n4630 & n10907 ;
  assign n10909 = ~n4345 & n10908 ;
  assign n10910 = n10909 ^ n10330 ^ 1'b0 ;
  assign n10911 = ~n1666 & n10910 ;
  assign n10912 = n10911 ^ n8946 ^ 1'b0 ;
  assign n10913 = n4368 | n10912 ;
  assign n10914 = n4933 ^ n1481 ^ 1'b0 ;
  assign n10915 = n10054 & ~n10914 ;
  assign n10916 = ~n695 & n10915 ;
  assign n10917 = n3167 | n4661 ;
  assign n10918 = n10917 ^ n8491 ^ 1'b0 ;
  assign n10919 = ~n2782 & n3681 ;
  assign n10920 = n10919 ^ n5311 ^ 1'b0 ;
  assign n10921 = x52 & ~n927 ;
  assign n10922 = n10697 ^ n1015 ^ 1'b0 ;
  assign n10923 = ~n3119 & n10922 ;
  assign n10924 = n10322 | n10923 ;
  assign n10925 = ~n4268 & n10571 ;
  assign n10926 = n4125 & ~n4931 ;
  assign n10927 = n10926 ^ n2376 ^ 1'b0 ;
  assign n10928 = ~n4045 & n10927 ;
  assign n10929 = n1113 & ~n7337 ;
  assign n10930 = n3037 & ~n9410 ;
  assign n10931 = n10930 ^ n4264 ^ 1'b0 ;
  assign n10932 = n1394 ^ n1133 ^ 1'b0 ;
  assign n10933 = n690 | n1935 ;
  assign n10934 = n2634 & ~n10933 ;
  assign n10935 = n10934 ^ n725 ^ 1'b0 ;
  assign n10936 = n6837 & ~n8628 ;
  assign n10937 = n3140 ^ n1392 ^ 1'b0 ;
  assign n10938 = n4206 & ~n6411 ;
  assign n10939 = n10937 & n10938 ;
  assign n10940 = n5015 ^ n645 ^ 1'b0 ;
  assign n10941 = n6700 ^ n1740 ^ 1'b0 ;
  assign n10942 = n10941 ^ n5385 ^ 1'b0 ;
  assign n10943 = n7273 & ~n10942 ;
  assign n10944 = n10943 ^ n1910 ^ 1'b0 ;
  assign n10945 = n3214 ^ n1907 ^ 1'b0 ;
  assign n10946 = ~n4875 & n10945 ;
  assign n10947 = n2235 & ~n3963 ;
  assign n10948 = n10946 & n10947 ;
  assign n10951 = n4664 ^ n3294 ^ 1'b0 ;
  assign n10949 = x38 | n6628 ;
  assign n10950 = n536 | n10949 ;
  assign n10952 = n10951 ^ n10950 ^ 1'b0 ;
  assign n10953 = n217 & ~n8443 ;
  assign n10954 = n7350 & n10953 ;
  assign n10955 = n4098 & ~n10954 ;
  assign n10956 = n10955 ^ n8732 ^ 1'b0 ;
  assign n10957 = ( n2435 & n4831 ) | ( n2435 & n10956 ) | ( n4831 & n10956 ) ;
  assign n10958 = ( n4612 & n5119 ) | ( n4612 & ~n10281 ) | ( n5119 & ~n10281 ) ;
  assign n10959 = n3455 & ~n7396 ;
  assign n10960 = n3253 & n10959 ;
  assign n10961 = ( n1129 & n2969 ) | ( n1129 & n4477 ) | ( n2969 & n4477 ) ;
  assign n10962 = n1052 & n10961 ;
  assign n10963 = n4416 & n10962 ;
  assign n10964 = n2134 | n10963 ;
  assign n10965 = n10964 ^ n8452 ^ 1'b0 ;
  assign n10966 = ~n10583 & n10965 ;
  assign n10967 = n2315 ^ n240 ^ x67 ;
  assign n10968 = n2458 | n2733 ;
  assign n10969 = n10968 ^ n7241 ^ 1'b0 ;
  assign n10970 = n4973 ^ n901 ^ 1'b0 ;
  assign n10971 = ~n4334 & n6607 ;
  assign n10972 = n7459 & n9010 ;
  assign n10973 = n10971 & n10972 ;
  assign n10974 = n3386 ^ n2126 ^ 1'b0 ;
  assign n10976 = n5967 ^ n3738 ^ 1'b0 ;
  assign n10977 = ~n7871 & n10976 ;
  assign n10978 = ~n5026 & n10977 ;
  assign n10975 = n1877 | n4287 ;
  assign n10979 = n10978 ^ n10975 ^ 1'b0 ;
  assign n10980 = n3391 ^ n3110 ^ 1'b0 ;
  assign n10981 = n809 & n1350 ;
  assign n10982 = ~n4482 & n10981 ;
  assign n10983 = n10982 ^ n6478 ^ 1'b0 ;
  assign n10984 = n10983 ^ n10533 ^ 1'b0 ;
  assign n10988 = x74 & n2240 ;
  assign n10985 = n5764 ^ n2776 ^ 1'b0 ;
  assign n10986 = n673 & n10985 ;
  assign n10987 = n10986 ^ n1344 ^ 1'b0 ;
  assign n10989 = n10988 ^ n10987 ^ n2028 ;
  assign n10990 = ~n2414 & n3037 ;
  assign n10991 = n3035 & ~n3365 ;
  assign n10992 = n5086 ^ n775 ^ 1'b0 ;
  assign n10993 = ~n3479 & n10992 ;
  assign n10994 = n4252 | n5850 ;
  assign n10995 = ( n4972 & ~n6696 ) | ( n4972 & n8502 ) | ( ~n6696 & n8502 ) ;
  assign n10996 = n4903 ^ n4210 ^ 1'b0 ;
  assign n10997 = n10995 & ~n10996 ;
  assign n10998 = n4192 ^ n788 ^ 1'b0 ;
  assign n10999 = n8849 & ~n10998 ;
  assign n11000 = n1693 ^ x95 ^ 1'b0 ;
  assign n11001 = n3212 & ~n8056 ;
  assign n11002 = n1629 & n3318 ;
  assign n11003 = ~n10730 & n11002 ;
  assign n11004 = n7437 ^ n5004 ^ 1'b0 ;
  assign n11005 = ~n5930 & n11004 ;
  assign n11006 = ~n209 & n11005 ;
  assign n11011 = n600 | n7662 ;
  assign n11012 = n11011 ^ n4806 ^ n2331 ;
  assign n11009 = n722 & ~n2312 ;
  assign n11010 = n11009 ^ n577 ^ 1'b0 ;
  assign n11007 = n959 | n6857 ;
  assign n11008 = n11007 ^ n4686 ^ 1'b0 ;
  assign n11013 = n11012 ^ n11010 ^ n11008 ;
  assign n11014 = n1235 & n9258 ;
  assign n11015 = n11014 ^ n2364 ^ 1'b0 ;
  assign n11016 = n4798 ^ n4251 ^ 1'b0 ;
  assign n11017 = n1790 & ~n11016 ;
  assign n11018 = n11017 ^ n4380 ^ 1'b0 ;
  assign n11019 = n11018 ^ n867 ^ 1'b0 ;
  assign n11020 = x100 & n1353 ;
  assign n11021 = n9131 & n11020 ;
  assign n11022 = n1842 ^ n728 ^ 1'b0 ;
  assign n11023 = n7128 | n11022 ;
  assign n11024 = ~n2344 & n8776 ;
  assign n11025 = n5826 & n11024 ;
  assign n11026 = n4019 | n10045 ;
  assign n11027 = ~n3314 & n11026 ;
  assign n11028 = n2226 & n6392 ;
  assign n11029 = n381 & n11028 ;
  assign n11030 = n3408 | n8706 ;
  assign n11031 = x46 | n11030 ;
  assign n11032 = n11031 ^ n6032 ^ 1'b0 ;
  assign n11033 = n4543 | n11032 ;
  assign n11035 = n971 | n1623 ;
  assign n11036 = n3097 & ~n11035 ;
  assign n11034 = ( ~n347 & n2140 ) | ( ~n347 & n5397 ) | ( n2140 & n5397 ) ;
  assign n11037 = n11036 ^ n11034 ^ 1'b0 ;
  assign n11038 = n293 & ~n8844 ;
  assign n11039 = n11038 ^ n2481 ^ 1'b0 ;
  assign n11040 = n11037 & ~n11039 ;
  assign n11042 = ~n687 & n1350 ;
  assign n11041 = n3672 & ~n4898 ;
  assign n11043 = n11042 ^ n11041 ^ 1'b0 ;
  assign n11044 = n747 & n4661 ;
  assign n11045 = n3119 | n8869 ;
  assign n11046 = n8845 & ~n11045 ;
  assign n11049 = n4683 & ~n8385 ;
  assign n11050 = ~n894 & n10528 ;
  assign n11051 = n11050 ^ n9092 ^ 1'b0 ;
  assign n11052 = ~n11049 & n11051 ;
  assign n11053 = n6511 & n11052 ;
  assign n11047 = n1586 & ~n9435 ;
  assign n11048 = n8158 & n11047 ;
  assign n11054 = n11053 ^ n11048 ^ n7558 ;
  assign n11055 = n518 & ~n5662 ;
  assign n11056 = n11055 ^ n2356 ^ 1'b0 ;
  assign n11057 = n500 & ~n3209 ;
  assign n11058 = ~n500 & n11057 ;
  assign n11059 = ~n1325 & n11058 ;
  assign n11060 = n11059 ^ n4162 ^ 1'b0 ;
  assign n11061 = n11060 ^ n9490 ^ 1'b0 ;
  assign n11062 = n3441 ^ n2427 ^ 1'b0 ;
  assign n11063 = ~n7735 & n11062 ;
  assign n11064 = ~n10368 & n11063 ;
  assign n11065 = n9195 ^ n5426 ^ 1'b0 ;
  assign n11066 = ~n2613 & n5635 ;
  assign n11067 = n2424 ^ n2326 ^ n578 ;
  assign n11068 = n406 & ~n11067 ;
  assign n11069 = n11068 ^ n3384 ^ 1'b0 ;
  assign n11070 = n1077 ^ n339 ^ 1'b0 ;
  assign n11071 = n1911 & ~n11070 ;
  assign n11072 = n11071 ^ n10937 ^ 1'b0 ;
  assign n11073 = n11072 ^ n5358 ^ 1'b0 ;
  assign n11074 = n1670 | n11073 ;
  assign n11075 = n3324 & n3927 ;
  assign n11076 = n11075 ^ n6314 ^ 1'b0 ;
  assign n11078 = n3582 & ~n7042 ;
  assign n11077 = n10350 ^ n6354 ^ 1'b0 ;
  assign n11079 = n11078 ^ n11077 ^ n2717 ;
  assign n11081 = n2912 ^ n2165 ^ 1'b0 ;
  assign n11082 = n1919 & ~n7173 ;
  assign n11083 = ~x70 & n11082 ;
  assign n11084 = n11081 & n11083 ;
  assign n11080 = n722 & n5281 ;
  assign n11085 = n11084 ^ n11080 ^ 1'b0 ;
  assign n11086 = n3478 ^ n1600 ^ 1'b0 ;
  assign n11087 = ~n6715 & n11086 ;
  assign n11088 = n3431 ^ n588 ^ 1'b0 ;
  assign n11089 = n11087 & n11088 ;
  assign n11090 = ( n1206 & n2121 ) | ( n1206 & ~n10123 ) | ( n2121 & ~n10123 ) ;
  assign n11091 = n4085 & n10615 ;
  assign n11092 = n11091 ^ n10163 ^ 1'b0 ;
  assign n11093 = n900 & n4302 ;
  assign n11094 = ~n11092 & n11093 ;
  assign n11095 = n9884 ^ n8697 ^ 1'b0 ;
  assign n11096 = n8219 & ~n11095 ;
  assign n11097 = ~n3162 & n11096 ;
  assign n11098 = n11097 ^ x56 ^ 1'b0 ;
  assign n11099 = ~n157 & n7338 ;
  assign n11100 = n11099 ^ n11056 ^ 1'b0 ;
  assign n11101 = x106 & ~n7368 ;
  assign n11102 = n11101 ^ n2319 ^ 1'b0 ;
  assign n11103 = n8121 | n9344 ;
  assign n11104 = n4918 ^ n1057 ^ 1'b0 ;
  assign n11105 = n2546 & ~n11104 ;
  assign n11106 = n11105 ^ n2252 ^ 1'b0 ;
  assign n11107 = n10152 ^ n8568 ^ 1'b0 ;
  assign n11108 = n1268 | n7783 ;
  assign n11109 = n7848 ^ n574 ^ 1'b0 ;
  assign n11110 = n11108 | n11109 ;
  assign n11111 = n2627 & ~n6082 ;
  assign n11112 = n9779 ^ n351 ^ 1'b0 ;
  assign n11113 = n11111 | n11112 ;
  assign n11114 = n11113 ^ n6754 ^ 1'b0 ;
  assign n11115 = n3636 | n5896 ;
  assign n11116 = n5094 ^ n959 ^ 1'b0 ;
  assign n11117 = ~n1099 & n11116 ;
  assign n11118 = n11117 ^ n1412 ^ x116 ;
  assign n11119 = n11118 ^ n6066 ^ 1'b0 ;
  assign n11120 = n6259 ^ n2754 ^ 1'b0 ;
  assign n11121 = n8559 & ~n11120 ;
  assign n11122 = n10409 & n11121 ;
  assign n11123 = n2044 & n11122 ;
  assign n11124 = n2348 & n11031 ;
  assign n11125 = n11124 ^ n1691 ^ 1'b0 ;
  assign n11126 = n852 & ~n11125 ;
  assign n11127 = ~n1304 & n9731 ;
  assign n11128 = n11127 ^ n2539 ^ 1'b0 ;
  assign n11129 = ~n1346 & n1510 ;
  assign n11130 = n9643 & n11129 ;
  assign n11131 = ( n1550 & n8641 ) | ( n1550 & ~n11130 ) | ( n8641 & ~n11130 ) ;
  assign n11132 = n1325 ^ n607 ^ 1'b0 ;
  assign n11133 = n1898 & n11132 ;
  assign n11139 = ~n680 & n3300 ;
  assign n11140 = n2621 & n11139 ;
  assign n11141 = n11140 ^ n3405 ^ 1'b0 ;
  assign n11134 = n1470 & n8520 ;
  assign n11135 = n11134 ^ n1209 ^ 1'b0 ;
  assign n11136 = n9894 & ~n11135 ;
  assign n11137 = n903 & n7640 ;
  assign n11138 = n11136 & ~n11137 ;
  assign n11142 = n11141 ^ n11138 ^ 1'b0 ;
  assign n11143 = n3119 ^ n2206 ^ 1'b0 ;
  assign n11144 = n11143 ^ n1134 ^ 1'b0 ;
  assign n11145 = n1071 & ~n6846 ;
  assign n11146 = ~n2654 & n11145 ;
  assign n11147 = n11146 ^ n808 ^ 1'b0 ;
  assign n11148 = ~n9437 & n10001 ;
  assign n11149 = ~n311 & n11148 ;
  assign n11150 = ~n3236 & n10447 ;
  assign n11152 = n2084 & ~n8179 ;
  assign n11153 = n8796 & n11152 ;
  assign n11151 = n1813 & n8572 ;
  assign n11154 = n11153 ^ n11151 ^ 1'b0 ;
  assign n11155 = x43 & ~n7332 ;
  assign n11156 = n11155 ^ n5408 ^ 1'b0 ;
  assign n11157 = ( n2395 & n9115 ) | ( n2395 & n11156 ) | ( n9115 & n11156 ) ;
  assign n11158 = n11154 | n11157 ;
  assign n11159 = n927 ^ n137 ^ 1'b0 ;
  assign n11160 = n4566 | n11159 ;
  assign n11161 = n143 & n4748 ;
  assign n11162 = ~n1890 & n11161 ;
  assign n11163 = n11160 | n11162 ;
  assign n11164 = n3601 | n8337 ;
  assign n11165 = n9876 & ~n11164 ;
  assign n11166 = n7582 ^ n3189 ^ 1'b0 ;
  assign n11167 = n3346 | n11166 ;
  assign n11169 = x30 & ~n335 ;
  assign n11170 = ~x30 & n11169 ;
  assign n11171 = n994 | n11170 ;
  assign n11172 = n11170 & ~n11171 ;
  assign n11173 = n11172 ^ n7713 ^ 1'b0 ;
  assign n11168 = n8695 | n10386 ;
  assign n11174 = n11173 ^ n11168 ^ 1'b0 ;
  assign n11175 = n4025 & ~n9992 ;
  assign n11176 = n3636 | n7047 ;
  assign n11177 = n2435 & n3395 ;
  assign n11178 = n11177 ^ n973 ^ 1'b0 ;
  assign n11179 = n3192 & ~n11178 ;
  assign n11180 = n11176 & n11179 ;
  assign n11181 = ~n774 & n8408 ;
  assign n11182 = n2011 | n11181 ;
  assign n11183 = n11182 ^ n2737 ^ 1'b0 ;
  assign n11184 = x55 & ~n11183 ;
  assign n11185 = ~n9797 & n11184 ;
  assign n11186 = n3288 & n7244 ;
  assign n11187 = ~n4843 & n11186 ;
  assign n11188 = n2054 | n3324 ;
  assign n11189 = n6195 ^ n3135 ^ 1'b0 ;
  assign n11190 = n11188 & ~n11189 ;
  assign n11191 = n11190 ^ n5693 ^ n2370 ;
  assign n11192 = n10359 ^ n8025 ^ 1'b0 ;
  assign n11193 = n8556 ^ n7354 ^ 1'b0 ;
  assign n11194 = n666 | n11193 ;
  assign n11195 = n2543 & ~n10838 ;
  assign n11196 = ~n4933 & n11195 ;
  assign n11197 = n11196 ^ n1052 ^ 1'b0 ;
  assign n11199 = n2231 & n6852 ;
  assign n11198 = n1074 & n10497 ;
  assign n11200 = n11199 ^ n11198 ^ n1689 ;
  assign n11201 = ~n3880 & n4452 ;
  assign n11202 = n9012 & n11201 ;
  assign n11203 = n9959 & ~n11202 ;
  assign n11204 = n8770 & n11203 ;
  assign n11205 = ~n2070 & n7485 ;
  assign n11206 = n11205 ^ n10253 ^ 1'b0 ;
  assign n11207 = n7916 & ~n11206 ;
  assign n11208 = n2568 ^ n2319 ^ 1'b0 ;
  assign n11209 = n1252 | n11208 ;
  assign n11210 = n10482 ^ n6345 ^ 1'b0 ;
  assign n11211 = n11209 & n11210 ;
  assign n11212 = ~n2319 & n8116 ;
  assign n11213 = n5416 & ~n11212 ;
  assign n11214 = ~n2704 & n3367 ;
  assign n11215 = n11214 ^ n3202 ^ 1'b0 ;
  assign n11216 = ( n2802 & n7959 ) | ( n2802 & n11215 ) | ( n7959 & n11215 ) ;
  assign n11217 = n9314 | n11216 ;
  assign n11218 = n468 | n5159 ;
  assign n11219 = n639 & ~n11218 ;
  assign n11220 = n2987 & n5112 ;
  assign n11221 = n6621 & ~n11220 ;
  assign n11222 = n791 & ~n3666 ;
  assign n11223 = ~n9570 & n11222 ;
  assign n11224 = n3100 & n11223 ;
  assign n11225 = ~n1634 & n3269 ;
  assign n11226 = ( n992 & n6741 ) | ( n992 & ~n11225 ) | ( n6741 & ~n11225 ) ;
  assign n11227 = n11224 | n11226 ;
  assign n11228 = n11227 ^ n1560 ^ 1'b0 ;
  assign n11229 = n10364 | n11228 ;
  assign n11230 = n2679 ^ n1526 ^ 1'b0 ;
  assign n11231 = n4507 & ~n11230 ;
  assign n11233 = n2246 | n2542 ;
  assign n11234 = n11233 ^ n5005 ^ 1'b0 ;
  assign n11232 = ~n2697 & n2780 ;
  assign n11235 = n11234 ^ n11232 ^ 1'b0 ;
  assign n11236 = n11235 ^ n9012 ^ 1'b0 ;
  assign n11237 = n163 & n11236 ;
  assign n11238 = ~n8073 & n11237 ;
  assign n11239 = ~n11231 & n11238 ;
  assign n11240 = n660 | n6879 ;
  assign n11241 = n2412 & ~n11240 ;
  assign n11242 = n172 | n11241 ;
  assign n11243 = n11242 ^ n2655 ^ 1'b0 ;
  assign n11244 = n3352 ^ n2824 ^ 1'b0 ;
  assign n11245 = n11244 ^ n1674 ^ 1'b0 ;
  assign n11246 = n1058 & ~n11245 ;
  assign n11247 = ~n2840 & n11246 ;
  assign n11248 = n11247 ^ n1816 ^ 1'b0 ;
  assign n11249 = n722 & n866 ;
  assign n11250 = ~n897 & n11249 ;
  assign n11251 = n852 | n3671 ;
  assign n11252 = n3962 | n11251 ;
  assign n11253 = n11250 | n11252 ;
  assign n11254 = n5586 & ~n9132 ;
  assign n11255 = x94 & n699 ;
  assign n11256 = n7368 | n11255 ;
  assign n11257 = x85 & n5716 ;
  assign n11258 = n11257 ^ n9045 ^ 1'b0 ;
  assign n11259 = n773 & n980 ;
  assign n11260 = n489 & ~n11259 ;
  assign n11261 = ~n2450 & n3784 ;
  assign n11262 = n11261 ^ n4216 ^ 1'b0 ;
  assign n11263 = n8938 ^ n6972 ^ 1'b0 ;
  assign n11264 = n6551 ^ n5606 ^ 1'b0 ;
  assign n11265 = n1056 & n5972 ;
  assign n11272 = n3587 ^ n791 ^ n630 ;
  assign n11273 = n11272 ^ n913 ^ 1'b0 ;
  assign n11274 = n666 | n11273 ;
  assign n11275 = n3122 & ~n11274 ;
  assign n11267 = n3527 & ~n5285 ;
  assign n11268 = n2452 & n11267 ;
  assign n11269 = n11268 ^ n3517 ^ 1'b0 ;
  assign n11266 = n3270 | n9350 ;
  assign n11270 = n11269 ^ n11266 ^ 1'b0 ;
  assign n11271 = n10845 & n11270 ;
  assign n11276 = n11275 ^ n11271 ^ 1'b0 ;
  assign n11277 = n759 & ~n1308 ;
  assign n11278 = n11277 ^ n5112 ^ 1'b0 ;
  assign n11283 = n2302 & n6350 ;
  assign n11284 = n11283 ^ n9890 ^ 1'b0 ;
  assign n11279 = n4253 ^ n2421 ^ 1'b0 ;
  assign n11280 = n2969 | n11279 ;
  assign n11281 = n4644 & ~n11280 ;
  assign n11282 = ~n2479 & n11281 ;
  assign n11285 = n11284 ^ n11282 ^ 1'b0 ;
  assign n11286 = n3996 & n11285 ;
  assign n11287 = n8175 ^ n5661 ^ 1'b0 ;
  assign n11288 = n3556 & ~n11287 ;
  assign n11289 = n11288 ^ n2402 ^ 1'b0 ;
  assign n11290 = n4844 ^ n4548 ^ 1'b0 ;
  assign n11291 = ~n853 & n11290 ;
  assign n11292 = ~n1028 & n11291 ;
  assign n11293 = n10797 & ~n11292 ;
  assign n11294 = n7538 ^ x1 ^ 1'b0 ;
  assign n11295 = n6396 & ~n6813 ;
  assign n11296 = ~n1552 & n1664 ;
  assign n11297 = n11296 ^ n2387 ^ 1'b0 ;
  assign n11298 = n5164 | n7175 ;
  assign n11299 = n6555 ^ n771 ^ 1'b0 ;
  assign n11300 = n5980 & ~n11299 ;
  assign n11301 = ~n8584 & n11300 ;
  assign n11302 = n11301 ^ n2103 ^ 1'b0 ;
  assign n11303 = n4912 & n5855 ;
  assign n11304 = n11303 ^ n9121 ^ 1'b0 ;
  assign n11308 = n2084 & n4126 ;
  assign n11309 = n11308 ^ n2514 ^ 1'b0 ;
  assign n11305 = n404 & n5837 ;
  assign n11306 = n11305 ^ n3762 ^ 1'b0 ;
  assign n11307 = ~n5073 & n11306 ;
  assign n11310 = n11309 ^ n11307 ^ 1'b0 ;
  assign n11311 = n7225 ^ n1720 ^ 1'b0 ;
  assign n11312 = n1590 & ~n8858 ;
  assign n11313 = ~n833 & n11312 ;
  assign n11314 = n2660 ^ x103 ^ 1'b0 ;
  assign n11315 = n4644 & n11314 ;
  assign n11316 = n8916 ^ n8199 ^ 1'b0 ;
  assign n11317 = n1581 | n11181 ;
  assign n11318 = n11317 ^ n6075 ^ 1'b0 ;
  assign n11319 = n11318 ^ n1435 ^ 1'b0 ;
  assign n11320 = ~n1150 & n11319 ;
  assign n11321 = n8688 ^ n5506 ^ 1'b0 ;
  assign n11322 = n8403 & ~n11321 ;
  assign n11323 = ~n363 & n3579 ;
  assign n11324 = n11323 ^ n779 ^ 1'b0 ;
  assign n11325 = n11324 ^ n2075 ^ 1'b0 ;
  assign n11326 = n7035 ^ n2739 ^ 1'b0 ;
  assign n11327 = n7629 & n11326 ;
  assign n11328 = n2027 ^ x4 ^ 1'b0 ;
  assign n11329 = n11327 & n11328 ;
  assign n11330 = n11325 | n11329 ;
  assign n11331 = n3699 | n5345 ;
  assign n11332 = n4370 ^ n1977 ^ n281 ;
  assign n11333 = ~n1933 & n11332 ;
  assign n11334 = ( n6046 & n6905 ) | ( n6046 & ~n11333 ) | ( n6905 & ~n11333 ) ;
  assign n11335 = n4903 ^ n4076 ^ 1'b0 ;
  assign n11336 = n4357 | n11335 ;
  assign n11337 = n11334 & n11336 ;
  assign n11338 = ~n3084 & n4966 ;
  assign n11339 = n11338 ^ n3224 ^ 1'b0 ;
  assign n11340 = n11337 | n11339 ;
  assign n11341 = n5945 ^ n5367 ^ 1'b0 ;
  assign n11342 = n3675 | n4566 ;
  assign n11343 = n180 | n11342 ;
  assign n11344 = ~n1150 & n11343 ;
  assign n11345 = n10193 & n11344 ;
  assign n11346 = n3237 & ~n3605 ;
  assign n11347 = n11345 & n11346 ;
  assign n11348 = n1861 | n11347 ;
  assign n11349 = n7876 | n9322 ;
  assign n11350 = ~n8730 & n11349 ;
  assign n11351 = n6893 ^ n6811 ^ 1'b0 ;
  assign n11352 = ~n9689 & n11351 ;
  assign n11353 = n11352 ^ n640 ^ 1'b0 ;
  assign n11355 = n5096 | n7408 ;
  assign n11356 = n11355 ^ n1514 ^ 1'b0 ;
  assign n11354 = n9110 ^ n4705 ^ 1'b0 ;
  assign n11357 = n11356 ^ n11354 ^ 1'b0 ;
  assign n11358 = n8341 ^ n7331 ^ n1383 ;
  assign n11359 = n5304 ^ n1649 ^ 1'b0 ;
  assign n11360 = n874 & n11359 ;
  assign n11361 = ~n1641 & n11360 ;
  assign n11362 = n2441 & ~n4739 ;
  assign n11363 = n11362 ^ n7016 ^ 1'b0 ;
  assign n11364 = n665 & n11363 ;
  assign n11365 = n1039 | n9091 ;
  assign n11366 = n9190 ^ n6174 ^ 1'b0 ;
  assign n11367 = ~n5809 & n11366 ;
  assign n11368 = ( n7289 & n7430 ) | ( n7289 & n11367 ) | ( n7430 & n11367 ) ;
  assign n11369 = n716 & ~n2955 ;
  assign n11370 = n11369 ^ n10973 ^ 1'b0 ;
  assign n11371 = n6992 & ~n11370 ;
  assign n11373 = n3441 ^ n1612 ^ 1'b0 ;
  assign n11374 = ~n5450 & n11373 ;
  assign n11372 = ~n243 & n3799 ;
  assign n11375 = n11374 ^ n11372 ^ 1'b0 ;
  assign n11377 = n2790 & n5093 ;
  assign n11378 = n1769 & n11377 ;
  assign n11379 = ( n1689 & n2610 ) | ( n1689 & ~n4716 ) | ( n2610 & ~n4716 ) ;
  assign n11380 = ( n9068 & n11378 ) | ( n9068 & ~n11379 ) | ( n11378 & ~n11379 ) ;
  assign n11376 = n2153 | n10207 ;
  assign n11381 = n11380 ^ n11376 ^ 1'b0 ;
  assign n11382 = ( n1062 & n6099 ) | ( n1062 & n11381 ) | ( n6099 & n11381 ) ;
  assign n11383 = n7433 ^ n6183 ^ 1'b0 ;
  assign n11384 = ~n569 & n11383 ;
  assign n11385 = n9596 ^ n6759 ^ n3674 ;
  assign n11386 = n2160 | n11385 ;
  assign n11387 = n9077 | n11386 ;
  assign n11390 = ~n6377 & n7271 ;
  assign n11391 = ~n2639 & n11390 ;
  assign n11388 = n1975 & ~n7828 ;
  assign n11389 = n11388 ^ n8703 ^ 1'b0 ;
  assign n11392 = n11391 ^ n11389 ^ 1'b0 ;
  assign n11393 = x35 & n11392 ;
  assign n11394 = n2405 ^ n2233 ^ 1'b0 ;
  assign n11395 = ~n7155 & n11394 ;
  assign n11396 = n11395 ^ n11176 ^ n3192 ;
  assign n11397 = n8632 ^ n2924 ^ 1'b0 ;
  assign n11398 = n2224 | n11397 ;
  assign n11399 = n11398 ^ n2859 ^ n2376 ;
  assign n11400 = n7094 | n9212 ;
  assign n11402 = n7099 ^ n3000 ^ 1'b0 ;
  assign n11403 = n10822 & ~n11402 ;
  assign n11401 = n4903 ^ n2546 ^ 1'b0 ;
  assign n11404 = n11403 ^ n11401 ^ 1'b0 ;
  assign n11405 = n1967 & n5195 ;
  assign n11406 = n461 & n11405 ;
  assign n11407 = n9764 ^ n2124 ^ 1'b0 ;
  assign n11408 = n11406 | n11407 ;
  assign n11409 = n494 & n597 ;
  assign n11410 = n11409 ^ n742 ^ 1'b0 ;
  assign n11411 = ~n1791 & n9027 ;
  assign n11412 = n3327 & n8911 ;
  assign n11413 = n2675 & n3853 ;
  assign n11414 = n11413 ^ n9823 ^ n6490 ;
  assign n11415 = n11414 ^ n10590 ^ n2289 ;
  assign n11416 = n2712 & ~n3210 ;
  assign n11417 = n2845 | n11416 ;
  assign n11418 = n4259 ^ n1790 ^ 1'b0 ;
  assign n11419 = n11417 | n11418 ;
  assign n11420 = n9691 ^ n5981 ^ 1'b0 ;
  assign n11421 = n4917 & ~n11420 ;
  assign n11422 = n11421 ^ n6759 ^ 1'b0 ;
  assign n11423 = n1943 | n7619 ;
  assign n11424 = n3961 | n8650 ;
  assign n11425 = n5635 & n8235 ;
  assign n11426 = n2353 & n11425 ;
  assign n11427 = n8613 | n11426 ;
  assign n11428 = n9207 & ~n11427 ;
  assign n11429 = n232 | n7245 ;
  assign n11436 = ~n1301 & n5281 ;
  assign n11437 = ~n7839 & n11436 ;
  assign n11430 = n1396 | n6434 ;
  assign n11431 = n11430 ^ n8638 ^ 1'b0 ;
  assign n11432 = n7041 ^ n533 ^ 1'b0 ;
  assign n11433 = ~n4551 & n11432 ;
  assign n11434 = n11209 & n11433 ;
  assign n11435 = ~n11431 & n11434 ;
  assign n11438 = n11437 ^ n11435 ^ n11420 ;
  assign n11439 = n2344 | n3047 ;
  assign n11440 = n1327 & ~n11439 ;
  assign n11441 = n6895 ^ n6684 ^ 1'b0 ;
  assign n11442 = n9376 | n11441 ;
  assign n11443 = n1834 & n6409 ;
  assign n11444 = n11443 ^ n9373 ^ 1'b0 ;
  assign n11445 = n437 & ~n4733 ;
  assign n11446 = n11445 ^ n3212 ^ 1'b0 ;
  assign n11447 = n9863 ^ n2248 ^ 1'b0 ;
  assign n11448 = x69 & n4013 ;
  assign n11449 = n11447 & n11448 ;
  assign n11450 = n11446 & ~n11449 ;
  assign n11451 = n11450 ^ n521 ^ 1'b0 ;
  assign n11452 = n278 | n11451 ;
  assign n11453 = n523 & n7231 ;
  assign n11454 = n4305 | n4411 ;
  assign n11455 = n2978 & ~n11454 ;
  assign n11456 = ~n729 & n2062 ;
  assign n11457 = n11455 | n11456 ;
  assign n11463 = n824 & n3481 ;
  assign n11464 = ~n824 & n11463 ;
  assign n11465 = n11464 ^ n3784 ^ 1'b0 ;
  assign n11459 = n194 | n6610 ;
  assign n11460 = n6610 & ~n11459 ;
  assign n11461 = n816 | n11460 ;
  assign n11462 = n11460 & ~n11461 ;
  assign n11458 = ~n1780 & n4043 ;
  assign n11466 = n11465 ^ n11462 ^ n11458 ;
  assign n11467 = n4191 ^ n2170 ^ 1'b0 ;
  assign n11468 = n240 & n4213 ;
  assign n11469 = ~n4958 & n11468 ;
  assign n11470 = n11469 ^ n10740 ^ 1'b0 ;
  assign n11471 = n11467 & ~n11470 ;
  assign n11472 = n11471 ^ n5203 ^ 1'b0 ;
  assign n11473 = n2010 & n2132 ;
  assign n11474 = n355 | n6168 ;
  assign n11475 = n11473 & n11474 ;
  assign n11476 = n7690 ^ n3991 ^ 1'b0 ;
  assign n11477 = ~n11475 & n11476 ;
  assign n11478 = n11477 ^ n4906 ^ 1'b0 ;
  assign n11479 = n3806 ^ n468 ^ 1'b0 ;
  assign n11480 = n6667 ^ n5808 ^ 1'b0 ;
  assign n11481 = ~n4089 & n11480 ;
  assign n11482 = ~n1058 & n11481 ;
  assign n11483 = ~n988 & n3880 ;
  assign n11484 = n4851 ^ n3842 ^ 1'b0 ;
  assign n11485 = n4553 ^ n959 ^ n791 ;
  assign n11486 = n6810 & ~n7368 ;
  assign n11487 = n11486 ^ n3758 ^ 1'b0 ;
  assign n11488 = n1765 & n9630 ;
  assign n11489 = n1708 | n2957 ;
  assign n11490 = n11489 ^ n9871 ^ 1'b0 ;
  assign n11491 = n7105 & n11490 ;
  assign n11492 = n3386 & n4090 ;
  assign n11493 = n11492 ^ n2423 ^ 1'b0 ;
  assign n11494 = n11493 ^ n677 ^ 1'b0 ;
  assign n11495 = n11494 ^ n9503 ^ n7764 ;
  assign n11496 = n3672 ^ n3215 ^ 1'b0 ;
  assign n11497 = n4774 ^ n2101 ^ 1'b0 ;
  assign n11498 = n11497 ^ n6135 ^ 1'b0 ;
  assign n11499 = n7039 ^ n4935 ^ 1'b0 ;
  assign n11500 = n9037 | n11499 ;
  assign n11501 = n6716 ^ n3121 ^ n2156 ;
  assign n11502 = ( n2474 & ~n8212 ) | ( n2474 & n11501 ) | ( ~n8212 & n11501 ) ;
  assign n11503 = ~n362 & n4463 ;
  assign n11504 = n11503 ^ n1623 ^ 1'b0 ;
  assign n11505 = n10986 ^ n167 ^ 1'b0 ;
  assign n11506 = n4612 & n11027 ;
  assign n11507 = ~n1502 & n5798 ;
  assign n11508 = n11507 ^ n3334 ^ n1134 ;
  assign n11509 = n3916 | n11508 ;
  assign n11510 = n7203 & ~n11509 ;
  assign n11511 = n2328 | n2640 ;
  assign n11512 = n11511 ^ n2164 ^ n1346 ;
  assign n11513 = n9598 ^ n7838 ^ 1'b0 ;
  assign n11514 = n8943 & n11513 ;
  assign n11515 = n379 & n5086 ;
  assign n11516 = n303 & n11515 ;
  assign n11517 = n11122 & ~n11516 ;
  assign n11518 = n11517 ^ n3162 ^ 1'b0 ;
  assign n11521 = n10189 ^ n1001 ^ 1'b0 ;
  assign n11522 = ( ~n905 & n2123 ) | ( ~n905 & n11521 ) | ( n2123 & n11521 ) ;
  assign n11523 = n2813 | n11522 ;
  assign n11524 = n768 | n11523 ;
  assign n11525 = n11524 ^ n6958 ^ 1'b0 ;
  assign n11519 = ~n4727 & n7951 ;
  assign n11520 = ~n5317 & n11519 ;
  assign n11526 = n11525 ^ n11520 ^ 1'b0 ;
  assign n11527 = n1761 & n7170 ;
  assign n11528 = n3147 | n6197 ;
  assign n11529 = ~n3119 & n7416 ;
  assign n11530 = n2724 & n11529 ;
  assign n11531 = n11530 ^ n2615 ^ 1'b0 ;
  assign n11532 = ( n1337 & n9853 ) | ( n1337 & ~n11531 ) | ( n9853 & ~n11531 ) ;
  assign n11533 = n3514 | n9072 ;
  assign n11534 = n4203 | n11533 ;
  assign n11536 = n3483 ^ n2961 ^ 1'b0 ;
  assign n11537 = n6686 & n11536 ;
  assign n11538 = n6404 & n11537 ;
  assign n11535 = ~n829 & n4849 ;
  assign n11539 = n11538 ^ n11535 ^ 1'b0 ;
  assign n11540 = n6748 & n11334 ;
  assign n11541 = n11540 ^ n2870 ^ 1'b0 ;
  assign n11542 = n1184 & ~n7805 ;
  assign n11543 = n7558 & ~n11512 ;
  assign n11544 = ~n7022 & n11543 ;
  assign n11545 = n3770 ^ n901 ^ 1'b0 ;
  assign n11546 = n1824 ^ n1790 ^ 1'b0 ;
  assign n11547 = n11546 ^ n5000 ^ n4359 ;
  assign n11548 = n11547 ^ n9928 ^ 1'b0 ;
  assign n11549 = n4405 & n6532 ;
  assign n11550 = n4064 & n11549 ;
  assign n11551 = n210 & n11550 ;
  assign n11552 = ~n5613 & n11551 ;
  assign n11560 = n4335 ^ n2328 ^ 1'b0 ;
  assign n11553 = n391 | n10697 ;
  assign n11554 = n8853 & ~n11553 ;
  assign n11555 = n1642 & ~n11215 ;
  assign n11556 = n3879 | n11555 ;
  assign n11557 = n6187 | n11556 ;
  assign n11558 = ~n11554 & n11557 ;
  assign n11559 = n11558 ^ n3722 ^ 1'b0 ;
  assign n11561 = n11560 ^ n11559 ^ n6814 ;
  assign n11562 = n791 & ~n8370 ;
  assign n11563 = n11562 ^ x102 ^ 1'b0 ;
  assign n11564 = n1009 | n4903 ;
  assign n11565 = n11564 ^ n477 ^ 1'b0 ;
  assign n11566 = n6326 & n11565 ;
  assign n11567 = n9166 ^ n2221 ^ 1'b0 ;
  assign n11568 = n969 ^ n530 ^ 1'b0 ;
  assign n11569 = n11568 ^ x24 ^ 1'b0 ;
  assign n11570 = n11567 & n11569 ;
  assign n11571 = ~n4808 & n5766 ;
  assign n11572 = n11570 | n11571 ;
  assign n11574 = n4330 & ~n5457 ;
  assign n11573 = n175 & n2553 ;
  assign n11575 = n11574 ^ n11573 ^ 1'b0 ;
  assign n11576 = n1491 & ~n11575 ;
  assign n11577 = ~n9246 & n11576 ;
  assign n11578 = n7422 & n8420 ;
  assign n11579 = n4093 & ~n11578 ;
  assign n11580 = n1197 & n11579 ;
  assign n11581 = ~n5840 & n8184 ;
  assign n11582 = ~n3850 & n11581 ;
  assign n11583 = n8768 ^ n3564 ^ 1'b0 ;
  assign n11584 = n8948 | n11583 ;
  assign n11585 = n8116 ^ n6409 ^ 1'b0 ;
  assign n11586 = n2226 & n6926 ;
  assign n11587 = n3350 | n3666 ;
  assign n11588 = n11587 ^ n4779 ^ 1'b0 ;
  assign n11589 = n10236 ^ n7649 ^ 1'b0 ;
  assign n11590 = n6193 ^ n2224 ^ 1'b0 ;
  assign n11591 = n2494 & ~n10826 ;
  assign n11592 = n6861 & ~n11350 ;
  assign n11593 = n3188 & n8793 ;
  assign n11594 = n11593 ^ n11354 ^ 1'b0 ;
  assign n11595 = n7038 & n11594 ;
  assign n11596 = n1044 & ~n7392 ;
  assign n11597 = n10950 ^ n1710 ^ 1'b0 ;
  assign n11598 = n2156 & ~n11597 ;
  assign n11599 = n11099 ^ n987 ^ 1'b0 ;
  assign n11600 = n11598 & n11599 ;
  assign n11601 = n11600 ^ n808 ^ 1'b0 ;
  assign n11602 = ~n1588 & n7540 ;
  assign n11603 = ~n4200 & n8810 ;
  assign n11604 = n2517 & n11603 ;
  assign n11605 = n7790 & n11604 ;
  assign n11606 = n3552 ^ n1421 ^ 1'b0 ;
  assign n11607 = n11606 ^ n726 ^ n534 ;
  assign n11608 = n2543 & ~n11607 ;
  assign n11609 = ~n6181 & n11608 ;
  assign n11610 = n4445 ^ n1350 ^ 1'b0 ;
  assign n11611 = n3991 ^ n2262 ^ 1'b0 ;
  assign n11612 = n462 & ~n588 ;
  assign n11613 = ~n11477 & n11612 ;
  assign n11617 = ~n4898 & n5256 ;
  assign n11614 = x42 & ~n411 ;
  assign n11615 = n11614 ^ n844 ^ 1'b0 ;
  assign n11616 = n6689 & ~n11615 ;
  assign n11618 = n11617 ^ n11616 ^ 1'b0 ;
  assign n11619 = n1047 & n4884 ;
  assign n11620 = n10971 & n11619 ;
  assign n11621 = n6716 & n11620 ;
  assign n11622 = ( n489 & ~n9863 ) | ( n489 & n11305 ) | ( ~n9863 & n11305 ) ;
  assign n11626 = n244 & ~n293 ;
  assign n11627 = ~n244 & n11626 ;
  assign n11628 = n2220 & n11627 ;
  assign n11623 = n5662 | n8386 ;
  assign n11624 = n8386 & ~n11623 ;
  assign n11625 = n2107 & ~n11624 ;
  assign n11629 = n11628 ^ n11625 ^ 1'b0 ;
  assign n11630 = x6 & n3085 ;
  assign n11631 = n545 | n11630 ;
  assign n11632 = n2564 & ~n11631 ;
  assign n11633 = n11629 & ~n11632 ;
  assign n11634 = n11633 ^ n6595 ^ 1'b0 ;
  assign n11635 = ( n1308 & n1549 ) | ( n1308 & ~n4814 ) | ( n1549 & ~n4814 ) ;
  assign n11636 = n3815 & ~n11635 ;
  assign n11637 = n11636 ^ n157 ^ 1'b0 ;
  assign n11638 = n11637 ^ n742 ^ 1'b0 ;
  assign n11639 = n11638 ^ n2476 ^ 1'b0 ;
  assign n11640 = n2529 & n11639 ;
  assign n11641 = n5657 & n8602 ;
  assign n11642 = ~n4556 & n11641 ;
  assign n11643 = n11642 ^ n1723 ^ 1'b0 ;
  assign n11644 = n8932 & n11643 ;
  assign n11645 = n2172 & n11644 ;
  assign n11646 = n1880 | n3011 ;
  assign n11647 = n11646 ^ n335 ^ 1'b0 ;
  assign n11648 = n4866 ^ n1939 ^ 1'b0 ;
  assign n11649 = n11647 | n11648 ;
  assign n11650 = n11649 ^ n1661 ^ 1'b0 ;
  assign n11651 = n11650 ^ n5670 ^ 1'b0 ;
  assign n11652 = n9923 & n11651 ;
  assign n11653 = n9576 ^ n1666 ^ 1'b0 ;
  assign n11654 = n7022 ^ n1019 ^ 1'b0 ;
  assign n11655 = ~n11506 & n11654 ;
  assign n11656 = n293 | n7319 ;
  assign n11657 = n11656 ^ n6935 ^ 1'b0 ;
  assign n11658 = ~n4619 & n8218 ;
  assign n11659 = ( n1817 & ~n4186 ) | ( n1817 & n11658 ) | ( ~n4186 & n11658 ) ;
  assign n11662 = n3269 & ~n3918 ;
  assign n11663 = n11662 ^ n577 ^ 1'b0 ;
  assign n11664 = n11663 ^ n3751 ^ 1'b0 ;
  assign n11660 = n618 ^ n612 ^ 1'b0 ;
  assign n11661 = n3503 & ~n11660 ;
  assign n11665 = n11664 ^ n11661 ^ 1'b0 ;
  assign n11666 = n11665 ^ n645 ^ 1'b0 ;
  assign n11667 = n3465 | n11666 ;
  assign n11668 = n1880 & ~n7155 ;
  assign n11669 = n3289 | n5519 ;
  assign n11670 = n11669 ^ n4776 ^ 1'b0 ;
  assign n11671 = n1550 ^ n468 ^ 1'b0 ;
  assign n11672 = ~n9481 & n11671 ;
  assign n11673 = n8429 & ~n11401 ;
  assign n11674 = n10246 ^ n6126 ^ n340 ;
  assign n11675 = ~n10969 & n11674 ;
  assign n11676 = n6323 & ~n7673 ;
  assign n11677 = ~n4450 & n11676 ;
  assign n11678 = n4474 & ~n11677 ;
  assign n11679 = n11678 ^ n623 ^ 1'b0 ;
  assign n11680 = n7888 ^ n7729 ^ 1'b0 ;
  assign n11681 = n11680 ^ n2132 ^ 1'b0 ;
  assign n11682 = n1338 & n7025 ;
  assign n11685 = n4283 ^ n4217 ^ 1'b0 ;
  assign n11686 = n5308 & ~n11685 ;
  assign n11683 = ~n468 & n3815 ;
  assign n11684 = n11683 ^ n3489 ^ 1'b0 ;
  assign n11687 = n11686 ^ n11684 ^ n3126 ;
  assign n11688 = n3310 & n11687 ;
  assign n11689 = ~n11682 & n11688 ;
  assign n11692 = n5678 ^ n4773 ^ 1'b0 ;
  assign n11693 = n11692 ^ n3584 ^ 1'b0 ;
  assign n11690 = n9394 ^ n6790 ^ n417 ;
  assign n11691 = n1013 | n11690 ;
  assign n11694 = n11693 ^ n11691 ^ 1'b0 ;
  assign n11697 = n3547 ^ n2640 ^ n851 ;
  assign n11695 = n1517 ^ n1128 ^ 1'b0 ;
  assign n11696 = n10173 & ~n11695 ;
  assign n11698 = n11697 ^ n11696 ^ 1'b0 ;
  assign n11699 = n10905 ^ n7324 ^ 1'b0 ;
  assign n11700 = n6559 ^ n2392 ^ 1'b0 ;
  assign n11701 = n3632 | n5365 ;
  assign n11702 = n11701 ^ n2370 ^ 1'b0 ;
  assign n11703 = n11700 | n11702 ;
  assign n11704 = n2953 & ~n9763 ;
  assign n11705 = ~n2787 & n3968 ;
  assign n11706 = n2845 & n11705 ;
  assign n11707 = n5916 ^ n2947 ^ 1'b0 ;
  assign n11708 = n4640 | n11707 ;
  assign n11709 = n7137 & ~n11708 ;
  assign n11710 = n11709 ^ n6323 ^ n1882 ;
  assign n11711 = n9904 ^ n4833 ^ 1'b0 ;
  assign n11712 = n8379 ^ n6973 ^ 1'b0 ;
  assign n11713 = n11711 | n11712 ;
  assign n11714 = n6225 & ~n10418 ;
  assign n11715 = n2640 | n6529 ;
  assign n11716 = ( n131 & n627 ) | ( n131 & ~n6799 ) | ( n627 & ~n6799 ) ;
  assign n11717 = n7702 | n11716 ;
  assign n11718 = n8876 | n11717 ;
  assign n11719 = n11715 | n11718 ;
  assign n11720 = n8699 ^ n838 ^ 1'b0 ;
  assign n11721 = n4703 & n10708 ;
  assign n11722 = n11721 ^ n2506 ^ 1'b0 ;
  assign n11723 = n7221 ^ n709 ^ 1'b0 ;
  assign n11724 = ( n6573 & n11722 ) | ( n6573 & n11723 ) | ( n11722 & n11723 ) ;
  assign n11725 = n11724 ^ n7680 ^ n7538 ;
  assign n11726 = n2165 & n7425 ;
  assign n11727 = n3247 & n11726 ;
  assign n11728 = n1186 & n8077 ;
  assign n11729 = n10920 & ~n11728 ;
  assign n11730 = ( n4426 & n11727 ) | ( n4426 & n11729 ) | ( n11727 & n11729 ) ;
  assign n11731 = n2798 ^ n1094 ^ 1'b0 ;
  assign n11732 = n2844 & ~n11731 ;
  assign n11733 = n4697 & n11732 ;
  assign n11734 = n11733 ^ n5208 ^ 1'b0 ;
  assign n11735 = n1469 | n11734 ;
  assign n11736 = n4006 | n11735 ;
  assign n11737 = n5745 & n11519 ;
  assign n11738 = n11736 & n11737 ;
  assign n11739 = n3006 ^ n1916 ^ 1'b0 ;
  assign n11740 = n1231 & ~n6506 ;
  assign n11741 = n10242 ^ n9620 ^ n1683 ;
  assign n11742 = n4851 ^ n3209 ^ 1'b0 ;
  assign n11743 = n3933 & ~n11742 ;
  assign n11744 = n6079 | n11743 ;
  assign n11745 = ~n1432 & n11744 ;
  assign n11746 = n1556 & ~n7388 ;
  assign n11747 = n11746 ^ n8418 ^ n1404 ;
  assign n11748 = n533 & n4182 ;
  assign n11749 = ~n3894 & n11748 ;
  assign n11750 = ~n2410 & n11749 ;
  assign n11751 = n10644 ^ x25 ^ 1'b0 ;
  assign n11752 = x1 & n1886 ;
  assign n11753 = ~n8296 & n11752 ;
  assign n11754 = n11753 ^ n5431 ^ 1'b0 ;
  assign n11755 = ~n1370 & n11754 ;
  assign n11756 = n2187 ^ n1252 ^ n1083 ;
  assign n11757 = n5667 & ~n9171 ;
  assign n11758 = n11757 ^ n2451 ^ 1'b0 ;
  assign n11759 = n1353 & ~n2893 ;
  assign n11760 = ~n256 & n11759 ;
  assign n11761 = ~n7866 & n11760 ;
  assign n11762 = n6473 & n11761 ;
  assign n11763 = n5723 & ~n11762 ;
  assign n11764 = n6665 & n11763 ;
  assign n11765 = ( n4571 & n6724 ) | ( n4571 & n9382 ) | ( n6724 & n9382 ) ;
  assign n11766 = n6020 & n11765 ;
  assign n11767 = n2985 & ~n5702 ;
  assign n11768 = ~n5347 & n11767 ;
  assign n11769 = n8908 ^ n8247 ^ 1'b0 ;
  assign n11770 = n11768 | n11769 ;
  assign n11771 = ~n468 & n1681 ;
  assign n11772 = n11771 ^ n3709 ^ 1'b0 ;
  assign n11773 = ~n1909 & n8165 ;
  assign n11774 = n150 | n5703 ;
  assign n11782 = n4922 & n8449 ;
  assign n11775 = n2429 ^ n1919 ^ 1'b0 ;
  assign n11776 = x7 & ~n2328 ;
  assign n11777 = ~n11775 & n11776 ;
  assign n11778 = n5248 & n8342 ;
  assign n11779 = n11777 | n11778 ;
  assign n11780 = n11779 ^ n3190 ^ 1'b0 ;
  assign n11781 = n5080 & ~n11780 ;
  assign n11783 = n11782 ^ n11781 ^ 1'b0 ;
  assign n11784 = n2302 | n10368 ;
  assign n11785 = n2462 ^ n147 ^ 1'b0 ;
  assign n11786 = n5916 & ~n11785 ;
  assign n11787 = n6503 ^ n2931 ^ 1'b0 ;
  assign n11788 = ~n8960 & n10470 ;
  assign n11789 = n11788 ^ n3010 ^ 1'b0 ;
  assign n11790 = n11789 ^ n9329 ^ 1'b0 ;
  assign n11791 = n1847 & n2228 ;
  assign n11792 = ~n3069 & n11791 ;
  assign n11793 = n10169 & ~n11792 ;
  assign n11794 = n1313 & ~n2628 ;
  assign n11795 = n1079 & n11794 ;
  assign n11796 = n789 & ~n11795 ;
  assign n11797 = ( ~n174 & n1732 ) | ( ~n174 & n2529 ) | ( n1732 & n2529 ) ;
  assign n11798 = n11797 ^ n351 ^ 1'b0 ;
  assign n11799 = n4292 ^ n425 ^ 1'b0 ;
  assign n11800 = n11798 & n11799 ;
  assign n11801 = ~x6 & n6151 ;
  assign n11802 = n3532 & n8343 ;
  assign n11803 = n9467 & n11802 ;
  assign n11804 = n3274 & ~n10202 ;
  assign n11805 = n2886 & n11804 ;
  assign n11806 = n7514 | n10261 ;
  assign n11807 = n2293 | n11806 ;
  assign n11808 = n5206 & n11000 ;
  assign n11809 = n9961 ^ n7440 ^ 1'b0 ;
  assign n11810 = n7391 ^ n1761 ^ 1'b0 ;
  assign n11811 = n11759 & n11810 ;
  assign n11812 = n3327 & ~n11811 ;
  assign n11813 = ~n4428 & n11812 ;
  assign n11814 = n6639 & ~n11813 ;
  assign n11815 = n2972 & n11814 ;
  assign n11817 = n553 & ~n5473 ;
  assign n11816 = ~n1632 & n5967 ;
  assign n11818 = n11817 ^ n11816 ^ n5159 ;
  assign n11819 = n4972 ^ n3045 ^ 1'b0 ;
  assign n11820 = n10952 & n11819 ;
  assign n11821 = n2746 & ~n5399 ;
  assign n11822 = n11821 ^ n5803 ^ 1'b0 ;
  assign n11823 = n8092 ^ n6923 ^ 1'b0 ;
  assign n11824 = n9923 & ~n11823 ;
  assign n11825 = x84 & n8689 ;
  assign n11826 = n11825 ^ n10356 ^ 1'b0 ;
  assign n11827 = n3350 | n3984 ;
  assign n11828 = n8352 | n11827 ;
  assign n11829 = n11826 & n11828 ;
  assign n11830 = n3547 ^ n1120 ^ 1'b0 ;
  assign n11831 = n5756 & n11830 ;
  assign n11832 = n5611 & n11831 ;
  assign n11833 = n3884 & n11832 ;
  assign n11834 = n11833 ^ n7221 ^ n7088 ;
  assign n11835 = n9327 & n11834 ;
  assign n11836 = n3098 ^ n521 ^ 1'b0 ;
  assign n11837 = n1975 & ~n11836 ;
  assign n11838 = ~n196 & n11837 ;
  assign n11839 = n9663 & n11838 ;
  assign n11840 = ( ~n517 & n9004 ) | ( ~n517 & n11839 ) | ( n9004 & n11839 ) ;
  assign n11841 = n3048 & ~n8824 ;
  assign n11842 = n11841 ^ n4019 ^ 1'b0 ;
  assign n11843 = n11549 ^ n1079 ^ 1'b0 ;
  assign n11844 = n9525 | n11843 ;
  assign n11845 = n4398 ^ n3855 ^ n779 ;
  assign n11846 = n7080 ^ n2622 ^ 1'b0 ;
  assign n11847 = n11845 & ~n11846 ;
  assign n11848 = n1412 & n11847 ;
  assign n11849 = n2596 & ~n11241 ;
  assign n11850 = ~n4344 & n5419 ;
  assign n11851 = ~n7377 & n11850 ;
  assign n11852 = n10219 ^ n5713 ^ 1'b0 ;
  assign n11853 = n218 | n11852 ;
  assign n11854 = n826 & n8916 ;
  assign n11855 = n6681 & n11854 ;
  assign n11856 = n789 | n2039 ;
  assign n11857 = n2938 | n11856 ;
  assign n11865 = n4976 ^ n3066 ^ 1'b0 ;
  assign n11858 = n7141 & ~n7504 ;
  assign n11859 = n11858 ^ n5443 ^ 1'b0 ;
  assign n11860 = n3636 & n11859 ;
  assign n11861 = n11860 ^ n6036 ^ 1'b0 ;
  assign n11862 = n4316 | n8680 ;
  assign n11863 = n11861 & n11862 ;
  assign n11864 = n3979 & n11863 ;
  assign n11866 = n11865 ^ n11864 ^ 1'b0 ;
  assign n11867 = n9015 ^ n3130 ^ 1'b0 ;
  assign n11868 = n11351 ^ n5518 ^ n2691 ;
  assign n11869 = ~n6879 & n11868 ;
  assign n11870 = ~n11867 & n11869 ;
  assign n11871 = n11870 ^ n8833 ^ 1'b0 ;
  assign n11872 = n9331 | n11871 ;
  assign n11873 = n8987 ^ n1485 ^ 1'b0 ;
  assign n11874 = n11542 ^ n7604 ^ 1'b0 ;
  assign n11875 = ~n3655 & n11874 ;
  assign n11876 = n224 & ~n6775 ;
  assign n11881 = n1005 ^ n371 ^ 1'b0 ;
  assign n11882 = n6455 | n11881 ;
  assign n11877 = n3987 | n7571 ;
  assign n11878 = n10072 ^ n611 ^ 1'b0 ;
  assign n11879 = n11877 & ~n11878 ;
  assign n11880 = n1851 & ~n11879 ;
  assign n11883 = n11882 ^ n11880 ^ n6237 ;
  assign n11884 = n11876 & ~n11883 ;
  assign n11885 = n1237 & n1720 ;
  assign n11887 = n4666 ^ n1797 ^ 1'b0 ;
  assign n11888 = ~n2564 & n11887 ;
  assign n11886 = ~n607 & n3973 ;
  assign n11889 = n11888 ^ n11886 ^ 1'b0 ;
  assign n11890 = ~n2593 & n3188 ;
  assign n11891 = n8226 | n11890 ;
  assign n11892 = ~n1298 & n8353 ;
  assign n11893 = ( n11349 & n11891 ) | ( n11349 & n11892 ) | ( n11891 & n11892 ) ;
  assign n11897 = ~n1353 & n6227 ;
  assign n11898 = n1353 & n11897 ;
  assign n11899 = n9406 & ~n11898 ;
  assign n11900 = ~n6667 & n11899 ;
  assign n11894 = n374 & n2298 ;
  assign n11895 = n2567 & n11894 ;
  assign n11896 = n2957 & n11895 ;
  assign n11901 = n11900 ^ n11896 ^ n11413 ;
  assign n11902 = ~n3842 & n7852 ;
  assign n11903 = n11902 ^ n5539 ^ 1'b0 ;
  assign n11904 = ~n11901 & n11903 ;
  assign n11905 = ~n7753 & n11369 ;
  assign n11906 = n11905 ^ n6607 ^ 1'b0 ;
  assign n11907 = n1823 ^ x6 ^ 1'b0 ;
  assign n11908 = n808 & n1850 ;
  assign n11909 = n2248 & ~n5017 ;
  assign n11910 = ~n11908 & n11909 ;
  assign n11911 = n11910 ^ n3574 ^ 1'b0 ;
  assign n11912 = n11907 & ~n11911 ;
  assign n11913 = n11912 ^ n956 ^ 1'b0 ;
  assign n11914 = ~n5605 & n11913 ;
  assign n11915 = ~n11216 & n11914 ;
  assign n11916 = n7705 ^ n3389 ^ 1'b0 ;
  assign n11917 = n6335 ^ n1664 ^ 1'b0 ;
  assign n11918 = n4568 ^ n2207 ^ 1'b0 ;
  assign n11919 = n11917 | n11918 ;
  assign n11923 = n5416 & ~n8623 ;
  assign n11920 = n1192 | n3633 ;
  assign n11921 = n3272 & ~n5837 ;
  assign n11922 = n11920 | n11921 ;
  assign n11924 = n11923 ^ n11922 ^ 1'b0 ;
  assign n11925 = n9458 & ~n10547 ;
  assign n11926 = n5086 & ~n9408 ;
  assign n11927 = n11926 ^ n1605 ^ n279 ;
  assign n11928 = n8931 ^ n1285 ^ 1'b0 ;
  assign n11929 = n7137 ^ n2250 ^ 1'b0 ;
  assign n11930 = n3405 | n11929 ;
  assign n11931 = ( n340 & n628 ) | ( n340 & ~n2948 ) | ( n628 & ~n2948 ) ;
  assign n11932 = n11930 | n11931 ;
  assign n11933 = n5091 & n11334 ;
  assign n11934 = n9013 & n11933 ;
  assign n11935 = n11934 ^ n2679 ^ 1'b0 ;
  assign n11936 = n10967 ^ n9392 ^ n7528 ;
  assign n11937 = n4662 ^ n2188 ^ 1'b0 ;
  assign n11938 = ~n7436 & n11042 ;
  assign n11939 = n1714 & n5855 ;
  assign n11940 = n3021 & ~n11939 ;
  assign n11941 = ~n11938 & n11940 ;
  assign n11942 = n6901 ^ n209 ^ 1'b0 ;
  assign n11943 = n6392 | n11942 ;
  assign n11944 = ( ~n4301 & n10352 ) | ( ~n4301 & n11943 ) | ( n10352 & n11943 ) ;
  assign n11945 = ~n920 & n1991 ;
  assign n11946 = n1487 & n2164 ;
  assign n11947 = ~n692 & n11946 ;
  assign n11948 = ( n1458 & ~n4597 ) | ( n1458 & n9699 ) | ( ~n4597 & n9699 ) ;
  assign n11949 = n11948 ^ n8106 ^ 1'b0 ;
  assign n11950 = n1195 & ~n11949 ;
  assign n11951 = n11950 ^ n3947 ^ 1'b0 ;
  assign n11952 = n6972 | n11467 ;
  assign n11953 = x1 | n11952 ;
  assign n11954 = n7004 ^ n3073 ^ 1'b0 ;
  assign n11955 = n1993 & ~n11954 ;
  assign n11956 = ~x102 & n7585 ;
  assign n11957 = ~n1239 & n11956 ;
  assign n11958 = n3711 | n11957 ;
  assign n11959 = n9243 ^ n4824 ^ 1'b0 ;
  assign n11960 = n2668 ^ n556 ^ 1'b0 ;
  assign n11961 = n2008 & n11960 ;
  assign n11962 = n4066 ^ n2075 ^ 1'b0 ;
  assign n11963 = ~n3033 & n11332 ;
  assign n11964 = n9997 ^ n6275 ^ 1'b0 ;
  assign n11965 = n3442 ^ n2476 ^ n2195 ;
  assign n11966 = ( ~n2892 & n3648 ) | ( ~n2892 & n11965 ) | ( n3648 & n11965 ) ;
  assign n11967 = n718 | n11966 ;
  assign n11968 = n738 | n11967 ;
  assign n11969 = n11484 ^ n3447 ^ n276 ;
  assign n11970 = n5715 ^ n2091 ^ 1'b0 ;
  assign n11971 = ( n220 & n2084 ) | ( n220 & ~n4366 ) | ( n2084 & ~n4366 ) ;
  assign n11972 = n11971 ^ x98 ^ 1'b0 ;
  assign n11973 = n7697 & ~n9996 ;
  assign n11974 = n3389 & ~n8633 ;
  assign n11976 = n10961 ^ n1200 ^ 1'b0 ;
  assign n11975 = n1044 | n11165 ;
  assign n11977 = n11976 ^ n11975 ^ 1'b0 ;
  assign n11978 = n180 | n2530 ;
  assign n11979 = n11978 ^ n3445 ^ 1'b0 ;
  assign n11980 = n11979 ^ n1500 ^ 1'b0 ;
  assign n11981 = n4216 & ~n11980 ;
  assign n11982 = n3505 ^ n3189 ^ 1'b0 ;
  assign n11983 = n11981 & ~n11982 ;
  assign n11984 = n7930 & ~n9141 ;
  assign n11985 = ~n8736 & n11984 ;
  assign n11986 = n3145 | n11985 ;
  assign n11987 = n832 | n11986 ;
  assign n11988 = ~n4334 & n5358 ;
  assign n11989 = n3565 & ~n5351 ;
  assign n11990 = ~n6561 & n11989 ;
  assign n11991 = n11988 & n11990 ;
  assign n11992 = n11991 ^ x24 ^ 1'b0 ;
  assign n11993 = n11987 & ~n11992 ;
  assign n11994 = n2760 | n6716 ;
  assign n11995 = n3327 ^ n1876 ^ 1'b0 ;
  assign n11996 = n2012 & ~n11995 ;
  assign n11997 = n10692 ^ n10527 ^ 1'b0 ;
  assign n11998 = x30 & ~n11997 ;
  assign n11999 = n10034 ^ n6754 ^ 1'b0 ;
  assign n12000 = ~n9448 & n11999 ;
  assign n12001 = ~n431 & n843 ;
  assign n12002 = n431 & n12001 ;
  assign n12003 = n12002 ^ n8959 ^ 1'b0 ;
  assign n12004 = ~n1469 & n12003 ;
  assign n12005 = ~n12003 & n12004 ;
  assign n12006 = n12005 ^ n8442 ^ n5176 ;
  assign n12007 = ~n1842 & n3280 ;
  assign n12008 = n12007 ^ n4860 ^ 1'b0 ;
  assign n12009 = n4280 & ~n12008 ;
  assign n12010 = n591 & ~n5547 ;
  assign n12011 = n12010 ^ x20 ^ 1'b0 ;
  assign n12012 = n12011 ^ n6631 ^ 1'b0 ;
  assign n12013 = n6843 | n12012 ;
  assign n12014 = n8689 | n12013 ;
  assign n12015 = n12014 ^ n11888 ^ 1'b0 ;
  assign n12016 = ~n9037 & n12015 ;
  assign n12017 = n1979 & n3595 ;
  assign n12018 = n1603 & ~n12017 ;
  assign n12019 = ~n999 & n7222 ;
  assign n12020 = n12019 ^ n11759 ^ 1'b0 ;
  assign n12021 = ~n3444 & n12020 ;
  assign n12026 = n1166 & ~n8116 ;
  assign n12027 = n12026 ^ n2398 ^ 1'b0 ;
  assign n12022 = n2632 ^ n2346 ^ 1'b0 ;
  assign n12023 = n4987 & n12022 ;
  assign n12024 = n12023 ^ n3110 ^ 1'b0 ;
  assign n12025 = n4128 | n12024 ;
  assign n12028 = n12027 ^ n12025 ^ 1'b0 ;
  assign n12029 = n4394 ^ n2652 ^ 1'b0 ;
  assign n12030 = n2673 & n12029 ;
  assign n12031 = ~n8246 & n12030 ;
  assign n12032 = n12031 ^ n8435 ^ 1'b0 ;
  assign n12033 = n7385 | n8863 ;
  assign n12034 = n4905 & ~n12033 ;
  assign n12035 = n4329 | n12034 ;
  assign n12037 = n8760 ^ n5635 ^ n805 ;
  assign n12036 = n4441 & n8737 ;
  assign n12038 = n12037 ^ n12036 ^ 1'b0 ;
  assign n12039 = ~n3547 & n6984 ;
  assign n12040 = ( n1008 & ~n7122 ) | ( n1008 & n12039 ) | ( ~n7122 & n12039 ) ;
  assign n12041 = n6907 & ~n12040 ;
  assign n12042 = n1287 | n10344 ;
  assign n12043 = n147 | n12042 ;
  assign n12044 = n2292 ^ n476 ^ 1'b0 ;
  assign n12045 = ~n5907 & n12044 ;
  assign n12046 = n12045 ^ n8687 ^ n3572 ;
  assign n12047 = n12046 ^ n5207 ^ 1'b0 ;
  assign n12048 = n4531 ^ n1079 ^ 1'b0 ;
  assign n12049 = n8373 & n12048 ;
  assign n12050 = n7986 | n12049 ;
  assign n12051 = n12050 ^ n6921 ^ 1'b0 ;
  assign n12052 = n9865 | n12051 ;
  assign n12053 = n5911 | n12052 ;
  assign n12054 = n12053 ^ n143 ^ 1'b0 ;
  assign n12055 = ~n6202 & n8645 ;
  assign n12056 = n12055 ^ n6315 ^ 1'b0 ;
  assign n12057 = n2062 & n5462 ;
  assign n12058 = n12056 | n12057 ;
  assign n12059 = n12058 ^ n8730 ^ 1'b0 ;
  assign n12060 = ~n5457 & n7648 ;
  assign n12061 = n12060 ^ n1574 ^ 1'b0 ;
  assign n12062 = ~n6542 & n10359 ;
  assign n12063 = n1136 | n5157 ;
  assign n12064 = n5427 & ~n9267 ;
  assign n12065 = n4953 & n10779 ;
  assign n12066 = n12065 ^ n6049 ^ 1'b0 ;
  assign n12067 = x62 | n163 ;
  assign n12068 = n937 & ~n9192 ;
  assign n12069 = n12068 ^ n3741 ^ 1'b0 ;
  assign n12070 = ~n683 & n12069 ;
  assign n12071 = n4688 & n12070 ;
  assign n12072 = n6827 & n12071 ;
  assign n12073 = ~n10861 & n10906 ;
  assign n12074 = ~x39 & n12073 ;
  assign n12075 = n3924 ^ n2445 ^ 1'b0 ;
  assign n12076 = n5176 | n12075 ;
  assign n12077 = n869 & ~n1276 ;
  assign n12078 = n3112 & n11433 ;
  assign n12079 = n8961 & n12078 ;
  assign n12080 = n6397 ^ n5260 ^ 1'b0 ;
  assign n12081 = n4251 & n10530 ;
  assign n12082 = n11498 ^ n10838 ^ 1'b0 ;
  assign n12083 = n1107 & n12082 ;
  assign n12084 = n8856 | n11944 ;
  assign n12086 = ~n3109 & n4703 ;
  assign n12085 = ~n1502 & n7403 ;
  assign n12087 = n12086 ^ n12085 ^ 1'b0 ;
  assign n12088 = n1224 & n6020 ;
  assign n12089 = n1973 | n12088 ;
  assign n12090 = n12089 ^ n2460 ^ 1'b0 ;
  assign n12091 = ( n240 & n1714 ) | ( n240 & n12090 ) | ( n1714 & n12090 ) ;
  assign n12092 = n11177 ^ n5127 ^ n4683 ;
  assign n12093 = ( x24 & ~n1231 ) | ( x24 & n8543 ) | ( ~n1231 & n8543 ) ;
  assign n12094 = n12093 ^ n257 ^ 1'b0 ;
  assign n12095 = ~n1147 & n5081 ;
  assign n12096 = n2693 & ~n12095 ;
  assign n12097 = ~n5935 & n12096 ;
  assign n12098 = n7574 & n8659 ;
  assign n12099 = n3982 & n5075 ;
  assign n12100 = n12099 ^ n3613 ^ 1'b0 ;
  assign n12101 = ( ~n2556 & n2756 ) | ( ~n2556 & n6730 ) | ( n2756 & n6730 ) ;
  assign n12102 = n10323 & n12101 ;
  assign n12103 = ~n260 & n546 ;
  assign n12104 = ~n546 & n12103 ;
  assign n12105 = ~n920 & n12104 ;
  assign n12106 = n2805 & ~n12105 ;
  assign n12107 = ~n637 & n716 ;
  assign n12108 = ~n716 & n12107 ;
  assign n12109 = ~x121 & n12108 ;
  assign n12110 = n460 & n12109 ;
  assign n12111 = ~n1212 & n12110 ;
  assign n12112 = n3813 & n12111 ;
  assign n12113 = n515 & n5635 ;
  assign n12114 = n12112 & n12113 ;
  assign n12115 = n977 | n12114 ;
  assign n12116 = n12114 & ~n12115 ;
  assign n12117 = n679 & ~n2655 ;
  assign n12118 = n2655 & n12117 ;
  assign n12119 = n12118 ^ n10216 ^ 1'b0 ;
  assign n12120 = n11053 | n12119 ;
  assign n12121 = n12116 & ~n12120 ;
  assign n12122 = n12106 & ~n12121 ;
  assign n12123 = n2134 & n12122 ;
  assign n12124 = ( n1410 & n3073 ) | ( n1410 & n9258 ) | ( n3073 & n9258 ) ;
  assign n12125 = n3700 | n12124 ;
  assign n12126 = n12125 ^ n2049 ^ 1'b0 ;
  assign n12127 = n1898 & n12126 ;
  assign n12128 = ( n3207 & n8006 ) | ( n3207 & ~n12127 ) | ( n8006 & ~n12127 ) ;
  assign n12129 = n5206 ^ x75 ^ 1'b0 ;
  assign n12130 = n1748 & n9107 ;
  assign n12131 = n12130 ^ n3066 ^ 1'b0 ;
  assign n12132 = n1295 & n3827 ;
  assign n12133 = n9348 ^ n857 ^ 1'b0 ;
  assign n12134 = n6742 & ~n12133 ;
  assign n12135 = ~n3503 & n5268 ;
  assign n12137 = x75 & n8768 ;
  assign n12138 = n5556 & n12137 ;
  assign n12139 = n4745 & ~n12138 ;
  assign n12140 = ~n4396 & n12139 ;
  assign n12136 = ~n3527 & n9433 ;
  assign n12141 = n12140 ^ n12136 ^ 1'b0 ;
  assign n12142 = n7928 | n12141 ;
  assign n12143 = n11976 ^ n297 ^ 1'b0 ;
  assign n12144 = ~n1708 & n3210 ;
  assign n12145 = ~n1884 & n12144 ;
  assign n12146 = n12145 ^ n10357 ^ 1'b0 ;
  assign n12147 = n646 & n12146 ;
  assign n12148 = ~n9010 & n12147 ;
  assign n12149 = n9918 ^ n437 ^ 1'b0 ;
  assign n12150 = n11557 & ~n12041 ;
  assign n12151 = n4686 ^ n267 ^ 1'b0 ;
  assign n12152 = n2248 & n12151 ;
  assign n12153 = n4249 | n12152 ;
  assign n12154 = n4182 & ~n12153 ;
  assign n12155 = n11764 ^ n11575 ^ 1'b0 ;
  assign n12156 = ~n11410 & n12155 ;
  assign n12157 = n2632 & ~n7250 ;
  assign n12158 = n1585 & ~n6534 ;
  assign n12159 = ~n8073 & n12158 ;
  assign n12160 = n12159 ^ n6214 ^ 1'b0 ;
  assign n12161 = n459 | n1522 ;
  assign n12162 = n12161 ^ n11895 ^ x23 ;
  assign n12163 = n5294 ^ n4602 ^ 1'b0 ;
  assign n12164 = n3664 & n12163 ;
  assign n12165 = n12162 & ~n12164 ;
  assign n12166 = n3388 | n8129 ;
  assign n12167 = n12166 ^ n7584 ^ n3773 ;
  assign n12168 = ~n2187 & n2303 ;
  assign n12169 = x83 & n5312 ;
  assign n12170 = ~n1431 & n12169 ;
  assign n12171 = n2832 & ~n12170 ;
  assign n12172 = n1792 & ~n12171 ;
  assign n12173 = n9331 ^ n3957 ^ 1'b0 ;
  assign n12174 = n12173 ^ n7408 ^ 1'b0 ;
  assign n12175 = n11208 | n12174 ;
  assign n12176 = n8371 | n8993 ;
  assign n12177 = ( n1078 & n7600 ) | ( n1078 & ~n12176 ) | ( n7600 & ~n12176 ) ;
  assign n12178 = n3478 & n9022 ;
  assign n12179 = ~n12177 & n12178 ;
  assign n12180 = n3091 & ~n12179 ;
  assign n12181 = n12180 ^ n11246 ^ 1'b0 ;
  assign n12182 = n7475 ^ n4596 ^ n3687 ;
  assign n12183 = ( n1107 & ~n1680 ) | ( n1107 & n12182 ) | ( ~n1680 & n12182 ) ;
  assign n12184 = n1996 | n7077 ;
  assign n12185 = n6355 & ~n12184 ;
  assign n12186 = n4576 & ~n12185 ;
  assign n12187 = n7587 ^ n3170 ^ 1'b0 ;
  assign n12188 = n11724 & ~n12187 ;
  assign n12189 = n1552 | n7417 ;
  assign n12190 = n3700 ^ n450 ^ 1'b0 ;
  assign n12191 = n7971 | n12190 ;
  assign n12192 = n12191 ^ n2048 ^ 1'b0 ;
  assign n12193 = ~n6300 & n12192 ;
  assign n12194 = n10695 & n12193 ;
  assign n12195 = ~n1157 & n7548 ;
  assign n12196 = n12195 ^ n5511 ^ 1'b0 ;
  assign n12197 = ~n12194 & n12196 ;
  assign n12198 = ~n12189 & n12197 ;
  assign n12199 = n609 & n12198 ;
  assign n12200 = ( ~n2011 & n3892 ) | ( ~n2011 & n5080 ) | ( n3892 & n5080 ) ;
  assign n12202 = n540 & ~n639 ;
  assign n12201 = n4159 & n4956 ;
  assign n12203 = n12202 ^ n12201 ^ 1'b0 ;
  assign n12204 = n1898 ^ n225 ^ 1'b0 ;
  assign n12205 = n1720 & ~n12204 ;
  assign n12206 = n12205 ^ n302 ^ 1'b0 ;
  assign n12207 = n4683 | n5148 ;
  assign n12208 = n5807 & ~n12207 ;
  assign n12209 = n12208 ^ n5811 ^ 1'b0 ;
  assign n12210 = n12013 | n12209 ;
  assign n12213 = ~x38 & n9214 ;
  assign n12212 = ~n2082 & n7535 ;
  assign n12214 = n12213 ^ n12212 ^ 1'b0 ;
  assign n12211 = n6059 & n7094 ;
  assign n12215 = n12214 ^ n12211 ^ 1'b0 ;
  assign n12216 = n9097 & n12215 ;
  assign n12217 = n5315 ^ n2754 ^ 1'b0 ;
  assign n12218 = n8656 | n8671 ;
  assign n12219 = x122 & n12218 ;
  assign n12220 = n12219 ^ n5635 ^ n462 ;
  assign n12221 = n3333 & ~n3636 ;
  assign n12222 = n2289 | n10578 ;
  assign n12223 = n12221 | n12222 ;
  assign n12224 = n10815 | n12223 ;
  assign n12225 = n742 & n2828 ;
  assign n12226 = ~n6295 & n12225 ;
  assign n12227 = n12226 ^ n874 ^ 1'b0 ;
  assign n12228 = n2193 ^ n556 ^ 1'b0 ;
  assign n12229 = n12227 & ~n12228 ;
  assign n12230 = n10275 ^ n5772 ^ 1'b0 ;
  assign n12231 = n1695 | n12230 ;
  assign n12232 = n11387 ^ n2024 ^ n1570 ;
  assign n12233 = n4671 | n7925 ;
  assign n12234 = n2067 & ~n9549 ;
  assign n12235 = n12234 ^ n722 ^ 1'b0 ;
  assign n12236 = ( ~n515 & n8862 ) | ( ~n515 & n12235 ) | ( n8862 & n12235 ) ;
  assign n12237 = n8244 | n12236 ;
  assign n12238 = n12237 ^ n11665 ^ 1'b0 ;
  assign n12239 = n6478 ^ n6007 ^ 1'b0 ;
  assign n12240 = ~n865 & n4315 ;
  assign n12241 = n12240 ^ n10114 ^ 1'b0 ;
  assign n12242 = n11231 & n12241 ;
  assign n12243 = n2746 & n3764 ;
  assign n12244 = n1722 ^ n634 ^ 1'b0 ;
  assign n12245 = n3481 | n12244 ;
  assign n12246 = ( n488 & n11140 ) | ( n488 & ~n12245 ) | ( n11140 & ~n12245 ) ;
  assign n12247 = n753 & ~n1124 ;
  assign n12248 = n12247 ^ n7006 ^ 1'b0 ;
  assign n12249 = n3456 ^ n2036 ^ 1'b0 ;
  assign n12250 = n12249 ^ n2248 ^ 1'b0 ;
  assign n12251 = ( x107 & ~n12248 ) | ( x107 & n12250 ) | ( ~n12248 & n12250 ) ;
  assign n12252 = n1552 | n2332 ;
  assign n12253 = n6167 | n12252 ;
  assign n12254 = n625 | n8909 ;
  assign n12255 = n12253 | n12254 ;
  assign n12256 = ( ~n10325 & n11890 ) | ( ~n10325 & n12255 ) | ( n11890 & n12255 ) ;
  assign n12257 = n392 & n8429 ;
  assign n12260 = n5563 ^ n4601 ^ 1'b0 ;
  assign n12261 = n12260 ^ n8396 ^ 1'b0 ;
  assign n12262 = n12261 ^ n6704 ^ n6539 ;
  assign n12258 = n433 & n4909 ;
  assign n12259 = n5287 & n12258 ;
  assign n12263 = n12262 ^ n12259 ^ 1'b0 ;
  assign n12264 = n3266 & ~n7415 ;
  assign n12265 = n6171 ^ n308 ^ 1'b0 ;
  assign n12266 = n10053 & n12265 ;
  assign n12267 = n6116 & ~n11014 ;
  assign n12268 = n12267 ^ n8432 ^ 1'b0 ;
  assign n12269 = n4247 ^ n4116 ^ 1'b0 ;
  assign n12270 = ~x2 & n8391 ;
  assign n12271 = n4221 & n12270 ;
  assign n12272 = n4216 ^ n2170 ^ 1'b0 ;
  assign n12273 = n11988 ^ n1481 ^ 1'b0 ;
  assign n12274 = x109 | n7199 ;
  assign n12275 = ~n1402 & n7678 ;
  assign n12276 = n1497 & n12275 ;
  assign n12277 = n6040 ^ n1912 ^ 1'b0 ;
  assign n12278 = ~n7673 & n12277 ;
  assign n12279 = n2889 ^ n2593 ^ 1'b0 ;
  assign n12280 = n12278 & ~n12279 ;
  assign n12281 = n12280 ^ n8943 ^ 1'b0 ;
  assign n12282 = n2654 & ~n5168 ;
  assign n12283 = ~n7315 & n12282 ;
  assign n12284 = n6828 ^ n1588 ^ 1'b0 ;
  assign n12285 = n527 & ~n754 ;
  assign n12286 = n12285 ^ n7828 ^ 1'b0 ;
  assign n12287 = n5486 | n9529 ;
  assign n12288 = ~n2218 & n12287 ;
  assign n12289 = ( n3903 & n12286 ) | ( n3903 & ~n12288 ) | ( n12286 & ~n12288 ) ;
  assign n12290 = n11188 ^ n5240 ^ 1'b0 ;
  assign n12291 = n12290 ^ n5342 ^ n1535 ;
  assign n12292 = n10605 ^ n2628 ^ 1'b0 ;
  assign n12293 = ( n2989 & n5649 ) | ( n2989 & ~n5853 ) | ( n5649 & ~n5853 ) ;
  assign n12294 = n10656 & n12293 ;
  assign n12295 = n437 & ~n3558 ;
  assign n12296 = n12295 ^ n1710 ^ 1'b0 ;
  assign n12297 = ~n12294 & n12296 ;
  assign n12298 = n1414 | n3602 ;
  assign n12299 = n12298 ^ n1763 ^ 1'b0 ;
  assign n12303 = n6381 & ~n10426 ;
  assign n12300 = n9166 ^ n3120 ^ 1'b0 ;
  assign n12301 = n10055 ^ n742 ^ 1'b0 ;
  assign n12302 = ~n12300 & n12301 ;
  assign n12304 = n12303 ^ n12302 ^ n4759 ;
  assign n12305 = n5083 | n5279 ;
  assign n12306 = n6467 | n12305 ;
  assign n12307 = n2750 & ~n4102 ;
  assign n12308 = n4379 ^ n471 ^ 1'b0 ;
  assign n12309 = n1354 & n7028 ;
  assign n12310 = ~n10357 & n12309 ;
  assign n12311 = n186 & ~n9623 ;
  assign n12312 = n4068 ^ n1291 ^ 1'b0 ;
  assign n12313 = ~n12311 & n12312 ;
  assign n12314 = n12313 ^ n9077 ^ 1'b0 ;
  assign n12315 = n4726 | n12314 ;
  assign n12316 = n12315 ^ n11329 ^ 1'b0 ;
  assign n12317 = n3681 | n12316 ;
  assign n12318 = x12 & ~n931 ;
  assign n12319 = n931 & n12318 ;
  assign n12320 = n12319 ^ n2513 ^ 1'b0 ;
  assign n12321 = ~n894 & n2484 ;
  assign n12322 = ~n2484 & n12321 ;
  assign n12323 = n884 & ~n12322 ;
  assign n12324 = ~n884 & n12323 ;
  assign n12325 = n803 | n1298 ;
  assign n12326 = n1298 & ~n12325 ;
  assign n12327 = n4293 | n12326 ;
  assign n12328 = n12324 & ~n12327 ;
  assign n12329 = n5667 | n12328 ;
  assign n12330 = n12320 | n12329 ;
  assign n12331 = n9041 | n9331 ;
  assign n12332 = n12331 ^ n1418 ^ 1'b0 ;
  assign n12333 = ( ~n615 & n3527 ) | ( ~n615 & n4249 ) | ( n3527 & n4249 ) ;
  assign n12334 = n12333 ^ n8415 ^ 1'b0 ;
  assign n12335 = n12334 ^ n7039 ^ 1'b0 ;
  assign n12336 = n4836 & ~n12335 ;
  assign n12337 = ( n12330 & ~n12332 ) | ( n12330 & n12336 ) | ( ~n12332 & n12336 ) ;
  assign n12338 = n4323 | n8174 ;
  assign n12339 = n5693 ^ n3140 ^ 1'b0 ;
  assign n12340 = n8205 ^ n7949 ^ n1791 ;
  assign n12341 = n1947 ^ n581 ^ 1'b0 ;
  assign n12342 = x123 & ~n12341 ;
  assign n12343 = ~n6544 & n12342 ;
  assign n12344 = ~n1473 & n12343 ;
  assign n12345 = n4389 ^ n3278 ^ n3074 ;
  assign n12347 = n9610 ^ n3582 ^ 1'b0 ;
  assign n12348 = n7797 ^ n1898 ^ 1'b0 ;
  assign n12349 = n12347 & n12348 ;
  assign n12346 = ~n1832 & n2738 ;
  assign n12350 = n12349 ^ n12346 ^ 1'b0 ;
  assign n12351 = n12350 ^ n10107 ^ 1'b0 ;
  assign n12352 = n12345 | n12351 ;
  assign n12353 = n12352 ^ n6534 ^ 1'b0 ;
  assign n12354 = n5106 ^ n3319 ^ 1'b0 ;
  assign n12355 = ~n973 & n12354 ;
  assign n12356 = n163 & ~n2868 ;
  assign n12357 = n12355 & n12356 ;
  assign n12358 = n9388 ^ n4453 ^ 1'b0 ;
  assign n12359 = n11658 ^ n2518 ^ 1'b0 ;
  assign n12360 = n12359 ^ n9774 ^ 1'b0 ;
  assign n12361 = n12358 & ~n12360 ;
  assign n12362 = n9032 ^ n7775 ^ 1'b0 ;
  assign n12363 = n1052 & ~n6376 ;
  assign n12364 = ~n1414 & n2220 ;
  assign n12365 = n6756 & n12364 ;
  assign n12366 = n11928 ^ n2098 ^ 1'b0 ;
  assign n12367 = n8342 & ~n12366 ;
  assign n12368 = n3690 ^ n2067 ^ 1'b0 ;
  assign n12369 = n8641 & ~n12368 ;
  assign n12370 = n7525 ^ n519 ^ 1'b0 ;
  assign n12371 = n4429 & ~n12370 ;
  assign n12372 = n12371 ^ n5243 ^ 1'b0 ;
  assign n12373 = ~n3046 & n5958 ;
  assign n12374 = ~n6226 & n12373 ;
  assign n12375 = n959 | n6368 ;
  assign n12376 = n3099 & ~n12375 ;
  assign n12377 = ( n1484 & n12374 ) | ( n1484 & ~n12376 ) | ( n12374 & ~n12376 ) ;
  assign n12378 = n1588 | n11055 ;
  assign n12379 = n3594 ^ n2119 ^ 1'b0 ;
  assign n12380 = ~n12378 & n12379 ;
  assign n12381 = n4048 ^ n1192 ^ 1'b0 ;
  assign n12382 = n12381 ^ n1657 ^ 1'b0 ;
  assign n12383 = n7501 & ~n12382 ;
  assign n12384 = n5062 & ~n7102 ;
  assign n12385 = n12384 ^ n2777 ^ 1'b0 ;
  assign n12386 = n12385 ^ n1957 ^ 1'b0 ;
  assign n12387 = n9350 ^ n6396 ^ 1'b0 ;
  assign n12388 = n198 & n6074 ;
  assign n12389 = n12388 ^ n628 ^ 1'b0 ;
  assign n12390 = n12389 ^ n9445 ^ 1'b0 ;
  assign n12391 = n9662 ^ n2378 ^ 1'b0 ;
  assign n12392 = n1473 & ~n2059 ;
  assign n12393 = ~n8850 & n12392 ;
  assign n12394 = ~n5918 & n12393 ;
  assign n12395 = n12027 & n12394 ;
  assign n12396 = ( n1031 & ~n1898 ) | ( n1031 & n4010 ) | ( ~n1898 & n4010 ) ;
  assign n12397 = n2487 ^ n882 ^ 1'b0 ;
  assign n12398 = n3511 & ~n5315 ;
  assign n12399 = ~n1429 & n12398 ;
  assign n12400 = n2116 ^ n1992 ^ 1'b0 ;
  assign n12401 = n1189 ^ n397 ^ 1'b0 ;
  assign n12402 = ~n12400 & n12401 ;
  assign n12403 = x16 & ~n10448 ;
  assign n12404 = n12403 ^ n7715 ^ n4041 ;
  assign n12405 = x117 & n10129 ;
  assign n12406 = n4394 | n5829 ;
  assign n12407 = ~n11937 & n12309 ;
  assign n12408 = n5816 & n12407 ;
  assign n12411 = n2788 & ~n2884 ;
  assign n12412 = x65 | n12411 ;
  assign n12413 = n3704 & ~n12412 ;
  assign n12409 = ( n404 & n718 ) | ( n404 & n6628 ) | ( n718 & n6628 ) ;
  assign n12410 = n12409 ^ n1962 ^ 1'b0 ;
  assign n12414 = n12413 ^ n12410 ^ 1'b0 ;
  assign n12415 = n5281 & ~n10226 ;
  assign n12416 = n12415 ^ n4008 ^ 1'b0 ;
  assign n12417 = x75 | n8297 ;
  assign n12418 = n2071 & ~n3511 ;
  assign n12419 = n5356 ^ n1081 ^ 1'b0 ;
  assign n12420 = n12418 | n12419 ;
  assign n12421 = n12420 ^ n4715 ^ 1'b0 ;
  assign n12422 = n7012 & ~n7875 ;
  assign n12423 = n12422 ^ n11209 ^ n2639 ;
  assign n12424 = n1629 | n7483 ;
  assign n12425 = n2380 | n6416 ;
  assign n12426 = n404 | n12425 ;
  assign n12427 = n12426 ^ n8332 ^ 1'b0 ;
  assign n12428 = ( n1933 & ~n2858 ) | ( n1933 & n7325 ) | ( ~n2858 & n7325 ) ;
  assign n12429 = n8232 ^ n5834 ^ 1'b0 ;
  assign n12430 = n8119 | n12429 ;
  assign n12431 = n12430 ^ n10927 ^ 1'b0 ;
  assign n12432 = n6512 & ~n12431 ;
  assign n12433 = ( n1388 & n3335 ) | ( n1388 & n9336 ) | ( n3335 & n9336 ) ;
  assign n12434 = n12433 ^ n4604 ^ 1'b0 ;
  assign n12435 = n8297 ^ x7 ^ 1'b0 ;
  assign n12436 = n4010 & n12435 ;
  assign n12437 = ~n3251 & n4652 ;
  assign n12438 = ~n12436 & n12437 ;
  assign n12439 = ~n2087 & n4345 ;
  assign n12440 = ~n2924 & n3343 ;
  assign n12441 = ~n9068 & n10929 ;
  assign n12442 = n12441 ^ n2470 ^ 1'b0 ;
  assign n12443 = n6227 ^ n4122 ^ 1'b0 ;
  assign n12444 = n11837 & n12443 ;
  assign n12445 = n10573 ^ n7396 ^ 1'b0 ;
  assign n12446 = n1176 | n12445 ;
  assign n12447 = n6942 ^ n2617 ^ 1'b0 ;
  assign n12448 = n393 & ~n12447 ;
  assign n12449 = n2349 | n5933 ;
  assign n12450 = n1176 & ~n12449 ;
  assign n12451 = n8718 | n12450 ;
  assign n12452 = n12448 | n12451 ;
  assign n12453 = n285 | n3177 ;
  assign n12454 = ~n754 & n8986 ;
  assign n12455 = n12453 & n12454 ;
  assign n12456 = n1884 | n12455 ;
  assign n12457 = n12456 ^ n2330 ^ 1'b0 ;
  assign n12458 = n8762 ^ n4777 ^ 1'b0 ;
  assign n12463 = n1853 ^ n1639 ^ 1'b0 ;
  assign n12462 = n398 & n4596 ;
  assign n12464 = n12463 ^ n12462 ^ 1'b0 ;
  assign n12459 = n4645 | n9799 ;
  assign n12460 = n4000 & ~n12459 ;
  assign n12461 = n7347 & ~n12460 ;
  assign n12465 = n12464 ^ n12461 ^ 1'b0 ;
  assign n12466 = n1741 & n11797 ;
  assign n12467 = ~n7347 & n12466 ;
  assign n12468 = n12467 ^ n4005 ^ n2338 ;
  assign n12469 = n6225 ^ n4477 ^ 1'b0 ;
  assign n12470 = n8165 & n12469 ;
  assign n12471 = n2204 & n5592 ;
  assign n12472 = n692 | n7358 ;
  assign n12473 = n3839 | n12472 ;
  assign n12474 = n2512 & ~n5457 ;
  assign n12475 = ~n7512 & n12474 ;
  assign n12476 = n5167 | n12475 ;
  assign n12477 = n12476 ^ n5397 ^ 1'b0 ;
  assign n12478 = n12473 & ~n12477 ;
  assign n12479 = ~n12471 & n12478 ;
  assign n12480 = n3287 & ~n6649 ;
  assign n12481 = n12480 ^ n293 ^ 1'b0 ;
  assign n12482 = ~n3814 & n12481 ;
  assign n12483 = n5179 & n12482 ;
  assign n12484 = n5285 ^ n1664 ^ 1'b0 ;
  assign n12485 = n791 & ~n12484 ;
  assign n12486 = n5360 & n9444 ;
  assign n12487 = n8405 & ~n11743 ;
  assign n12489 = n2580 ^ n1152 ^ 1'b0 ;
  assign n12490 = n9481 | n12489 ;
  assign n12488 = ~n1231 & n5829 ;
  assign n12491 = n12490 ^ n12488 ^ 1'b0 ;
  assign n12498 = ~n2639 & n7007 ;
  assign n12499 = n760 & n12498 ;
  assign n12492 = x3 & ~n998 ;
  assign n12493 = n12492 ^ n2096 ^ 1'b0 ;
  assign n12494 = n12493 ^ n6750 ^ n1399 ;
  assign n12495 = n12494 ^ n4105 ^ 1'b0 ;
  assign n12496 = n8645 & ~n12495 ;
  assign n12497 = ~n254 & n12496 ;
  assign n12500 = n12499 ^ n12497 ^ 1'b0 ;
  assign n12501 = n9481 ^ n5544 ^ 1'b0 ;
  assign n12502 = n5684 ^ n2176 ^ 1'b0 ;
  assign n12503 = n12502 ^ n9258 ^ n347 ;
  assign n12504 = n6965 ^ n952 ^ 1'b0 ;
  assign n12505 = n4538 | n10849 ;
  assign n12506 = n3344 & n12505 ;
  assign n12507 = ~n3880 & n12506 ;
  assign n12508 = n10905 ^ n3319 ^ 1'b0 ;
  assign n12509 = n10736 & n12508 ;
  assign n12510 = n12509 ^ n11680 ^ 1'b0 ;
  assign n12511 = n2874 & ~n12510 ;
  assign n12512 = n3477 & n7781 ;
  assign n12513 = n12512 ^ n5561 ^ n2949 ;
  assign n12514 = n1452 | n7508 ;
  assign n12515 = n4174 | n12514 ;
  assign n12516 = n9382 ^ n1933 ^ 1'b0 ;
  assign n12517 = n1005 | n12516 ;
  assign n12518 = ( ~n4833 & n12515 ) | ( ~n4833 & n12517 ) | ( n12515 & n12517 ) ;
  assign n12519 = n5277 ^ n4390 ^ 1'b0 ;
  assign n12520 = n1342 & ~n12519 ;
  assign n12521 = n269 & n12192 ;
  assign n12522 = ~n12520 & n12521 ;
  assign n12523 = n7877 & n10474 ;
  assign n12524 = n12523 ^ n4307 ^ 1'b0 ;
  assign n12525 = n12308 ^ n1698 ^ 1'b0 ;
  assign n12526 = n8472 ^ n5592 ^ 1'b0 ;
  assign n12527 = n6252 & ~n12526 ;
  assign n12528 = n3328 & n11467 ;
  assign n12529 = n243 | n2876 ;
  assign n12530 = n12528 | n12529 ;
  assign n12531 = n1600 & ~n1778 ;
  assign n12532 = n12531 ^ n639 ^ 1'b0 ;
  assign n12533 = n3811 | n5537 ;
  assign n12534 = n1602 & ~n12533 ;
  assign n12535 = n6579 & ~n7779 ;
  assign n12536 = n4622 & ~n4876 ;
  assign n12537 = ~n7170 & n12536 ;
  assign n12538 = ( ~n3908 & n8310 ) | ( ~n3908 & n12537 ) | ( n8310 & n12537 ) ;
  assign n12539 = n1517 & n5647 ;
  assign n12540 = n900 & n6446 ;
  assign n12541 = n12540 ^ n8425 ^ 1'b0 ;
  assign n12542 = n12541 ^ n3744 ^ 1'b0 ;
  assign n12543 = n10379 & n12542 ;
  assign n12544 = n11051 ^ n5392 ^ 1'b0 ;
  assign n12545 = n6879 | n12544 ;
  assign n12546 = n3251 ^ n3145 ^ 1'b0 ;
  assign n12547 = n10579 | n10612 ;
  assign n12548 = n6563 & n12547 ;
  assign n12549 = n6563 & n11988 ;
  assign n12550 = n10241 ^ n6075 ^ 1'b0 ;
  assign n12551 = n12549 & n12550 ;
  assign n12552 = n6378 | n8736 ;
  assign n12553 = ~n673 & n809 ;
  assign n12554 = ~n12552 & n12553 ;
  assign n12555 = n1823 & n2207 ;
  assign n12556 = n6575 | n12555 ;
  assign n12557 = n3788 & n8885 ;
  assign n12558 = n12557 ^ x14 ^ 1'b0 ;
  assign n12559 = n5275 & ~n8293 ;
  assign n12560 = n2413 & n4987 ;
  assign n12561 = ~n987 & n12560 ;
  assign n12562 = ~n729 & n1886 ;
  assign n12563 = ~n2412 & n12562 ;
  assign n12564 = ~n3953 & n12563 ;
  assign n12565 = n12561 | n12564 ;
  assign n12566 = n578 & ~n1578 ;
  assign n12567 = ( n2192 & n8500 ) | ( n2192 & n10850 ) | ( n8500 & n10850 ) ;
  assign n12568 = n5915 ^ n1510 ^ 1'b0 ;
  assign n12569 = n5352 & ~n12568 ;
  assign n12570 = n11181 | n12569 ;
  assign n12571 = n12570 ^ n3964 ^ n900 ;
  assign n12572 = n2510 ^ n1275 ^ 1'b0 ;
  assign n12573 = n3359 & ~n12572 ;
  assign n12579 = n258 & ~n8108 ;
  assign n12580 = ~n3140 & n12579 ;
  assign n12577 = n1558 ^ n1511 ^ 1'b0 ;
  assign n12578 = n3896 & ~n12577 ;
  assign n12581 = n12580 ^ n12578 ^ 1'b0 ;
  assign n12574 = n8277 ^ n4113 ^ 1'b0 ;
  assign n12575 = n12574 ^ n5253 ^ x26 ;
  assign n12576 = n12575 ^ n159 ^ 1'b0 ;
  assign n12582 = n12581 ^ n12576 ^ 1'b0 ;
  assign n12586 = n5277 & ~n12138 ;
  assign n12583 = n6713 ^ n6473 ^ 1'b0 ;
  assign n12584 = n12583 ^ n433 ^ 1'b0 ;
  assign n12585 = n5981 & ~n12584 ;
  assign n12587 = n12586 ^ n12585 ^ 1'b0 ;
  assign n12588 = n3744 & n6661 ;
  assign n12589 = ~n5521 & n12588 ;
  assign n12590 = n10836 ^ n1603 ^ 1'b0 ;
  assign n12591 = n1338 ^ x33 ^ 1'b0 ;
  assign n12592 = n8151 ^ n1013 ^ 1'b0 ;
  assign n12593 = n10798 & n12592 ;
  assign n12594 = n10189 ^ n7542 ^ n208 ;
  assign n12595 = n12532 ^ n6734 ^ 1'b0 ;
  assign n12596 = x88 & ~n6526 ;
  assign n12597 = n12596 ^ n6712 ^ 1'b0 ;
  assign n12598 = n11188 & n12597 ;
  assign n12599 = n12598 ^ n11895 ^ 1'b0 ;
  assign n12600 = ~n673 & n1751 ;
  assign n12601 = n12600 ^ n1425 ^ 1'b0 ;
  assign n12602 = n11893 & n12601 ;
  assign n12603 = n5434 | n9055 ;
  assign n12604 = n12603 ^ n6501 ^ n404 ;
  assign n12605 = n3572 | n7797 ;
  assign n12606 = n3116 & n3274 ;
  assign n12607 = ~n163 & n556 ;
  assign n12608 = n12199 ^ n2596 ^ 1'b0 ;
  assign n12609 = n12607 & ~n12608 ;
  assign n12610 = n4474 & ~n8436 ;
  assign n12611 = n2603 & ~n11883 ;
  assign n12612 = n12611 ^ n1962 ^ 1'b0 ;
  assign n12613 = n5817 ^ n2611 ^ n2083 ;
  assign n12614 = n391 | n7697 ;
  assign n12615 = ~n11128 & n12614 ;
  assign n12616 = ~n5069 & n12615 ;
  assign n12617 = n4664 ^ n679 ^ 1'b0 ;
  assign n12618 = n2153 & n12617 ;
  assign n12619 = n1741 & n12287 ;
  assign n12620 = n12619 ^ n5035 ^ 1'b0 ;
  assign n12621 = n8333 ^ n4528 ^ 1'b0 ;
  assign n12622 = n8595 ^ n2969 ^ n2491 ;
  assign n12623 = n12622 ^ n4180 ^ 1'b0 ;
  assign n12624 = n12623 ^ n8444 ^ n7662 ;
  assign n12625 = n3100 ^ n1247 ^ 1'b0 ;
  assign n12626 = n2675 ^ n1103 ^ 1'b0 ;
  assign n12627 = ~n3357 & n12626 ;
  assign n12628 = ( n511 & n539 ) | ( n511 & n1386 ) | ( n539 & n1386 ) ;
  assign n12629 = n1518 | n4007 ;
  assign n12630 = n12628 & ~n12629 ;
  assign n12633 = n5614 ^ n2028 ^ 1'b0 ;
  assign n12634 = ~n6022 & n12633 ;
  assign n12631 = n6579 ^ n2127 ^ n1597 ;
  assign n12632 = n10999 & ~n12631 ;
  assign n12635 = n12634 ^ n12632 ^ 1'b0 ;
  assign n12636 = ~n1703 & n6852 ;
  assign n12637 = n5273 & n12636 ;
  assign n12638 = x29 | n815 ;
  assign n12639 = ~n709 & n12638 ;
  assign n12640 = ~n1897 & n12639 ;
  assign n12641 = n1937 & n12640 ;
  assign n12642 = n3809 & ~n4386 ;
  assign n12643 = n3874 & n4814 ;
  assign n12644 = n3666 & n12643 ;
  assign n12645 = ( n1556 & n12642 ) | ( n1556 & ~n12644 ) | ( n12642 & ~n12644 ) ;
  assign n12646 = n2228 & n4708 ;
  assign n12647 = ~n6813 & n12646 ;
  assign n12648 = n530 | n3027 ;
  assign n12649 = n8490 & ~n12648 ;
  assign n12650 = n2030 | n5235 ;
  assign n12651 = n6283 | n12650 ;
  assign n12652 = n4776 & n12651 ;
  assign n12653 = n12652 ^ n9574 ^ 1'b0 ;
  assign n12654 = n362 & n10055 ;
  assign n12655 = n3433 & ~n5805 ;
  assign n12656 = n2105 & n12655 ;
  assign n12657 = n3908 ^ n3475 ^ 1'b0 ;
  assign n12658 = n12657 ^ n10252 ^ 1'b0 ;
  assign n12662 = n8099 ^ n3540 ^ 1'b0 ;
  assign n12663 = n3498 ^ n2656 ^ 1'b0 ;
  assign n12664 = n12662 & ~n12663 ;
  assign n12665 = n11591 & n12664 ;
  assign n12666 = n12665 ^ n2998 ^ 1'b0 ;
  assign n12659 = n331 & n7967 ;
  assign n12660 = n12659 ^ n10938 ^ 1'b0 ;
  assign n12661 = n3792 & ~n12660 ;
  assign n12667 = n12666 ^ n12661 ^ 1'b0 ;
  assign n12668 = n6969 ^ n2697 ^ 1'b0 ;
  assign n12669 = n1367 & ~n7964 ;
  assign n12670 = n10708 ^ n4791 ^ 1'b0 ;
  assign n12671 = ( n867 & n2144 ) | ( n867 & ~n4423 ) | ( n2144 & ~n4423 ) ;
  assign n12672 = n3986 ^ n3841 ^ 1'b0 ;
  assign n12673 = n12671 | n12672 ;
  assign n12674 = n12673 ^ n3074 ^ 1'b0 ;
  assign n12675 = n8551 ^ n5624 ^ 1'b0 ;
  assign n12676 = n7054 & n12675 ;
  assign n12677 = n8554 & ~n10657 ;
  assign n12678 = n7280 ^ n351 ^ 1'b0 ;
  assign n12679 = n7146 & ~n11030 ;
  assign n12680 = n3567 | n7615 ;
  assign n12681 = n2629 & n10784 ;
  assign n12682 = n7955 ^ n3861 ^ 1'b0 ;
  assign n12683 = n799 & n3073 ;
  assign n12684 = n12683 ^ n3093 ^ 1'b0 ;
  assign n12685 = n177 | n4219 ;
  assign n12686 = n12685 ^ n8401 ^ 1'b0 ;
  assign n12687 = n2106 | n5731 ;
  assign n12688 = n12686 & ~n12687 ;
  assign n12689 = ~n1372 & n1788 ;
  assign n12690 = n2823 & n12689 ;
  assign n12691 = n642 & ~n4737 ;
  assign n12692 = n12691 ^ n9473 ^ 1'b0 ;
  assign n12693 = n12692 ^ n2108 ^ 1'b0 ;
  assign n12694 = ~n533 & n12693 ;
  assign n12695 = n12694 ^ n9337 ^ 1'b0 ;
  assign n12702 = n3225 & ~n6132 ;
  assign n12699 = ~n347 & n1237 ;
  assign n12700 = ~n4002 & n6044 ;
  assign n12701 = n12699 & n12700 ;
  assign n12703 = n12702 ^ n12701 ^ 1'b0 ;
  assign n12696 = n5721 & n10992 ;
  assign n12697 = ~n620 & n12696 ;
  assign n12698 = n6257 | n12697 ;
  assign n12704 = n12703 ^ n12698 ^ 1'b0 ;
  assign n12705 = n3704 ^ n3266 ^ 1'b0 ;
  assign n12706 = ~n10088 & n12705 ;
  assign n12707 = n12706 ^ n6844 ^ 1'b0 ;
  assign n12708 = n12707 ^ n10014 ^ 1'b0 ;
  assign n12709 = n12704 & n12708 ;
  assign n12710 = n4898 | n6594 ;
  assign n12711 = ~n1947 & n3809 ;
  assign n12712 = ~n1642 & n12711 ;
  assign n12713 = n2431 | n12712 ;
  assign n12714 = n10954 & ~n12713 ;
  assign n12715 = n12714 ^ n9372 ^ 1'b0 ;
  assign n12716 = n4712 & ~n12715 ;
  assign n12717 = n3064 ^ n2048 ^ n1755 ;
  assign n12718 = n7250 ^ n2898 ^ 1'b0 ;
  assign n12719 = ~n12717 & n12718 ;
  assign n12720 = n5825 ^ n180 ^ 1'b0 ;
  assign n12721 = ~n11593 & n12720 ;
  assign n12722 = n12625 ^ n11668 ^ 1'b0 ;
  assign n12723 = n12721 & ~n12722 ;
  assign n12724 = ~n6114 & n7514 ;
  assign n12725 = n12724 ^ n6035 ^ 1'b0 ;
  assign n12726 = n9114 ^ n3587 ^ 1'b0 ;
  assign n12727 = n7822 & ~n12726 ;
  assign n12728 = n2602 ^ n1121 ^ 1'b0 ;
  assign n12729 = ~n521 & n3665 ;
  assign n12730 = n2395 & n12729 ;
  assign n12731 = n12730 ^ n765 ^ 1'b0 ;
  assign n12732 = n12728 & n12731 ;
  assign n12733 = n9295 & n12732 ;
  assign n12734 = ~n1197 & n1266 ;
  assign n12735 = n12734 ^ n3559 ^ x6 ;
  assign n12736 = ( n1867 & n4861 ) | ( n1867 & ~n8286 ) | ( n4861 & ~n8286 ) ;
  assign n12737 = n5519 | n12736 ;
  assign n12738 = n12737 ^ n11084 ^ 1'b0 ;
  assign n12739 = n8036 | n12738 ;
  assign n12740 = ( n7848 & ~n12735 ) | ( n7848 & n12739 ) | ( ~n12735 & n12739 ) ;
  assign n12741 = n6225 & n9186 ;
  assign n12742 = n12741 ^ n3735 ^ 1'b0 ;
  assign n12743 = n6563 ^ n2989 ^ 1'b0 ;
  assign n12744 = ~n1211 & n4673 ;
  assign n12745 = n5455 ^ n3764 ^ n2746 ;
  assign n12746 = n2062 | n2288 ;
  assign n12747 = n12253 & ~n12746 ;
  assign n12748 = ~n12745 & n12747 ;
  assign n12749 = n12744 & n12748 ;
  assign n12750 = n12749 ^ n1747 ^ 1'b0 ;
  assign n12752 = ( n1001 & ~n4350 ) | ( n1001 & n5157 ) | ( ~n4350 & n5157 ) ;
  assign n12753 = n12752 ^ n11607 ^ 1'b0 ;
  assign n12751 = ~n5203 & n8747 ;
  assign n12754 = n12753 ^ n12751 ^ 1'b0 ;
  assign n12755 = n10453 ^ n4350 ^ 1'b0 ;
  assign n12756 = n4888 & n7106 ;
  assign n12762 = n2452 & n4979 ;
  assign n12757 = ~n3033 & n3709 ;
  assign n12758 = n1327 & n12757 ;
  assign n12759 = n11988 | n12758 ;
  assign n12760 = n2464 & n12759 ;
  assign n12761 = n5434 & n12760 ;
  assign n12763 = n12762 ^ n12761 ^ n8235 ;
  assign n12764 = n2412 ^ n2028 ^ 1'b0 ;
  assign n12765 = n1825 | n5800 ;
  assign n12766 = n12765 ^ n11923 ^ 1'b0 ;
  assign n12767 = n6415 & n12766 ;
  assign n12768 = x99 | n8317 ;
  assign n12769 = n5445 ^ n1121 ^ 1'b0 ;
  assign n12770 = n3808 & ~n12769 ;
  assign n12771 = n7619 ^ n6754 ^ n4212 ;
  assign n12772 = n5645 ^ n1742 ^ 1'b0 ;
  assign n12773 = x1 | n12772 ;
  assign n12774 = n12773 ^ n8902 ^ 1'b0 ;
  assign n12775 = n2156 | n12774 ;
  assign n12776 = n12771 & ~n12775 ;
  assign n12777 = n994 & ~n7666 ;
  assign n12778 = n1031 & n1079 ;
  assign n12779 = n658 | n12778 ;
  assign n12780 = n5664 ^ n4310 ^ 1'b0 ;
  assign n12781 = n11188 ^ n9295 ^ 1'b0 ;
  assign n12782 = ~n12780 & n12781 ;
  assign n12783 = n7928 | n12782 ;
  assign n12784 = n8803 ^ n1118 ^ 1'b0 ;
  assign n12785 = n12783 | n12784 ;
  assign n12786 = n1805 & ~n2218 ;
  assign n12787 = n6796 ^ n1189 ^ 1'b0 ;
  assign n12788 = n12786 | n12787 ;
  assign n12789 = ~n4708 & n9205 ;
  assign n12790 = n2302 & ~n3869 ;
  assign n12791 = ~n6242 & n12790 ;
  assign n12792 = n12791 ^ n150 ^ 1'b0 ;
  assign n12793 = n3015 ^ n2355 ^ n435 ;
  assign n12794 = n12792 & n12793 ;
  assign n12795 = n490 & n12794 ;
  assign n12796 = n11038 ^ n3536 ^ 1'b0 ;
  assign n12797 = n10031 ^ n9382 ^ n3567 ;
  assign n12798 = n12797 ^ n2952 ^ 1'b0 ;
  assign n12799 = n12796 | n12798 ;
  assign n12800 = n12799 ^ x63 ^ 1'b0 ;
  assign n12801 = n8309 ^ n7905 ^ 1'b0 ;
  assign n12802 = ~n10014 & n12801 ;
  assign n12803 = n12802 ^ n12249 ^ n2445 ;
  assign n12804 = n5985 & ~n10894 ;
  assign n12805 = n12804 ^ n4571 ^ 1'b0 ;
  assign n12806 = n10352 ^ n3156 ^ 1'b0 ;
  assign n12807 = ~n1424 & n5887 ;
  assign n12808 = n12807 ^ n4271 ^ 1'b0 ;
  assign n12809 = ~n10692 & n12808 ;
  assign n12810 = n12806 & n12809 ;
  assign n12820 = n3139 ^ n1710 ^ 1'b0 ;
  assign n12821 = n5779 & ~n12820 ;
  assign n12814 = ( n456 & n1611 ) | ( n456 & n2226 ) | ( n1611 & n2226 ) ;
  assign n12815 = n476 | n1689 ;
  assign n12816 = n12814 & ~n12815 ;
  assign n12811 = n4806 ^ n3804 ^ 1'b0 ;
  assign n12812 = n699 | n12811 ;
  assign n12813 = n12812 ^ n8541 ^ 1'b0 ;
  assign n12817 = n12816 ^ n12813 ^ n7678 ;
  assign n12818 = n12249 ^ n10474 ^ 1'b0 ;
  assign n12819 = ~n12817 & n12818 ;
  assign n12822 = n12821 ^ n12819 ^ 1'b0 ;
  assign n12823 = n2984 ^ n250 ^ x21 ;
  assign n12826 = n5901 ^ n2622 ^ 1'b0 ;
  assign n12827 = n5725 & ~n12826 ;
  assign n12824 = n4200 ^ n774 ^ 1'b0 ;
  assign n12825 = n856 | n12824 ;
  assign n12828 = n12827 ^ n12825 ^ n450 ;
  assign n12829 = n11374 ^ n6841 ^ 1'b0 ;
  assign n12830 = ~n12828 & n12829 ;
  assign n12831 = n12830 ^ n4179 ^ n695 ;
  assign n12832 = n12831 ^ n531 ^ 1'b0 ;
  assign n12833 = n12823 & ~n12832 ;
  assign n12834 = n3997 & n6482 ;
  assign n12835 = n5872 & n12834 ;
  assign n12836 = n5392 & n12835 ;
  assign n12837 = n4036 | n5599 ;
  assign n12838 = n12837 ^ n11322 ^ n4440 ;
  assign n12839 = ~n749 & n4482 ;
  assign n12840 = n12839 ^ n10941 ^ 1'b0 ;
  assign n12841 = ~n4204 & n10270 ;
  assign n12842 = n12841 ^ n5815 ^ 1'b0 ;
  assign n12843 = n12505 ^ n11417 ^ 1'b0 ;
  assign n12844 = ~n5844 & n9728 ;
  assign n12845 = ~n5374 & n11985 ;
  assign n12846 = n1985 & n9638 ;
  assign n12847 = n7417 ^ n3535 ^ 1'b0 ;
  assign n12848 = ~n7163 & n12847 ;
  assign n12849 = n8244 & n12848 ;
  assign n12850 = n12846 & n12849 ;
  assign n12851 = ~n1391 & n1568 ;
  assign n12852 = n3458 | n4073 ;
  assign n12853 = n12851 | n12852 ;
  assign n12854 = n2827 ^ n1853 ^ 1'b0 ;
  assign n12855 = n787 & ~n973 ;
  assign n12856 = ( n3615 & ~n10876 ) | ( n3615 & n12855 ) | ( ~n10876 & n12855 ) ;
  assign n12857 = ~n5872 & n12856 ;
  assign n12858 = ~n4104 & n12857 ;
  assign n12859 = n208 & n4840 ;
  assign n12860 = n12859 ^ n5977 ^ 1'b0 ;
  assign n12861 = n8451 & n12860 ;
  assign n12862 = n12861 ^ n4125 ^ 1'b0 ;
  assign n12863 = ~n4416 & n11923 ;
  assign n12864 = n1529 & n4064 ;
  assign n12866 = n6167 ^ n5857 ^ n1184 ;
  assign n12865 = n5398 & ~n6159 ;
  assign n12867 = n12866 ^ n12865 ^ n2626 ;
  assign n12868 = n6037 | n9722 ;
  assign n12869 = n11385 & ~n12868 ;
  assign n12870 = n6204 ^ n3988 ^ 1'b0 ;
  assign n12871 = ~n5015 & n12870 ;
  assign n12872 = n9259 ^ n2204 ^ 1'b0 ;
  assign n12873 = n12871 & ~n12872 ;
  assign n12875 = n2597 & n6310 ;
  assign n12874 = n1232 & n1429 ;
  assign n12876 = n12875 ^ n12874 ^ 1'b0 ;
  assign n12877 = n6569 & ~n6783 ;
  assign n12878 = n12877 ^ n4621 ^ 1'b0 ;
  assign n12879 = n334 | n5952 ;
  assign n12880 = n5684 & n11031 ;
  assign n12881 = ~n5240 & n12880 ;
  assign n12882 = ~n2142 & n12881 ;
  assign n12883 = n7782 ^ n1406 ^ 1'b0 ;
  assign n12884 = ~n10270 & n12883 ;
  assign n12885 = n12882 & n12884 ;
  assign n12886 = ( n5513 & n6172 ) | ( n5513 & ~n8774 ) | ( n6172 & ~n8774 ) ;
  assign n12888 = n3552 & ~n4159 ;
  assign n12889 = n12888 ^ n6678 ^ 1'b0 ;
  assign n12887 = n986 & ~n3589 ;
  assign n12890 = n12889 ^ n12887 ^ n3993 ;
  assign n12891 = ~n12886 & n12890 ;
  assign n12892 = ~n9177 & n12891 ;
  assign n12893 = n462 | n12892 ;
  assign n12894 = n3524 | n12440 ;
  assign n12895 = n12440 & ~n12894 ;
  assign n12896 = n8164 | n9888 ;
  assign n12897 = n5551 & ~n7195 ;
  assign n12898 = n12897 ^ n11703 ^ n8796 ;
  assign n12899 = n5133 ^ n3128 ^ 1'b0 ;
  assign n12900 = n6792 ^ n3604 ^ n2327 ;
  assign n12901 = n3335 | n12900 ;
  assign n12902 = n5710 & ~n12901 ;
  assign n12903 = n1810 | n2201 ;
  assign n12904 = n8106 ^ n939 ^ 1'b0 ;
  assign n12905 = n12903 & n12904 ;
  assign n12906 = n5627 | n12905 ;
  assign n12907 = n1066 & ~n5090 ;
  assign n12908 = n12906 & n12907 ;
  assign n12909 = n6493 ^ n803 ^ 1'b0 ;
  assign n12910 = n225 & ~n1057 ;
  assign n12911 = n3582 ^ n2312 ^ 1'b0 ;
  assign n12912 = n5018 ^ n2410 ^ 1'b0 ;
  assign n12913 = n12912 ^ n7856 ^ n4386 ;
  assign n12914 = ~n10209 & n12913 ;
  assign n12915 = n7380 & n12914 ;
  assign n12916 = x38 & ~n1651 ;
  assign n12917 = n3278 & n12916 ;
  assign n12918 = n5251 ^ n2458 ^ 1'b0 ;
  assign n12919 = n12917 & ~n12918 ;
  assign n12920 = ~n4403 & n12919 ;
  assign n12921 = n12920 ^ n4828 ^ 1'b0 ;
  assign n12922 = n11617 | n12921 ;
  assign n12923 = ( n4895 & ~n5358 ) | ( n4895 & n9058 ) | ( ~n5358 & n9058 ) ;
  assign n12924 = n9853 ^ n5420 ^ 1'b0 ;
  assign n12925 = n6571 & n8931 ;
  assign n12926 = ~n3479 & n8339 ;
  assign n12927 = ~n472 & n2908 ;
  assign n12928 = n472 & n12927 ;
  assign n12929 = n11019 & ~n12928 ;
  assign n12930 = ~n12926 & n12929 ;
  assign n12931 = n12926 & n12930 ;
  assign n12932 = n954 & n9392 ;
  assign n12933 = n208 & n12932 ;
  assign n12936 = n11795 ^ n6330 ^ n1754 ;
  assign n12934 = n244 & n4182 ;
  assign n12935 = n12934 ^ n759 ^ 1'b0 ;
  assign n12937 = n12936 ^ n12935 ^ 1'b0 ;
  assign n12938 = n2405 ^ n2192 ^ 1'b0 ;
  assign n12939 = n5857 & n10554 ;
  assign n12940 = n3973 ^ n927 ^ 1'b0 ;
  assign n12941 = n12940 ^ n7787 ^ n2126 ;
  assign n12946 = n4033 & ~n8342 ;
  assign n12942 = n2961 ^ n2769 ^ 1'b0 ;
  assign n12943 = n543 & ~n2756 ;
  assign n12944 = n12943 ^ n11209 ^ 1'b0 ;
  assign n12945 = n12942 | n12944 ;
  assign n12947 = n12946 ^ n12945 ^ n6841 ;
  assign n12948 = n2370 ^ n1791 ^ 1'b0 ;
  assign n12949 = n10944 ^ n840 ^ 1'b0 ;
  assign n12950 = n9597 & ~n12949 ;
  assign n12951 = n6509 | n8119 ;
  assign n12952 = n5694 ^ n718 ^ 1'b0 ;
  assign n12953 = n10948 ^ x70 ^ 1'b0 ;
  assign n12954 = n1213 | n1422 ;
  assign n12955 = n12953 & ~n12954 ;
  assign n12956 = n10463 ^ n6591 ^ 1'b0 ;
  assign n12957 = n9826 & ~n12956 ;
  assign n12958 = ~x45 & n12957 ;
  assign n12959 = n6717 | n9768 ;
  assign n12960 = n5997 ^ n2912 ^ 1'b0 ;
  assign n12961 = n6352 | n12960 ;
  assign n12962 = ( n3938 & n4703 ) | ( n3938 & ~n8410 ) | ( n4703 & ~n8410 ) ;
  assign n12963 = n4251 | n12962 ;
  assign n12964 = n5841 | n6719 ;
  assign n12965 = n9856 ^ n7649 ^ n2121 ;
  assign n12966 = n7749 ^ n4611 ^ n499 ;
  assign n12967 = n12966 ^ n9240 ^ 1'b0 ;
  assign n12968 = n587 | n5566 ;
  assign n12969 = n12968 ^ n2192 ^ 1'b0 ;
  assign n12970 = n12000 ^ n8428 ^ 1'b0 ;
  assign n12971 = n12970 ^ n5244 ^ 1'b0 ;
  assign n12972 = n12969 | n12971 ;
  assign n12973 = n1376 & n6786 ;
  assign n12974 = n12973 ^ n5308 ^ 1'b0 ;
  assign n12975 = n3903 | n11690 ;
  assign n12976 = n12975 ^ n8648 ^ 1'b0 ;
  assign n12977 = ( n6197 & ~n7504 ) | ( n6197 & n12976 ) | ( ~n7504 & n12976 ) ;
  assign n12978 = n10633 ^ n9585 ^ 1'b0 ;
  assign n12979 = n2034 & ~n2278 ;
  assign n12980 = n6331 ^ n1295 ^ 1'b0 ;
  assign n12981 = n12979 & n12980 ;
  assign n12982 = n12981 ^ n2164 ^ 1'b0 ;
  assign n12983 = n1627 & ~n11564 ;
  assign n12984 = n11965 ^ n7051 ^ 1'b0 ;
  assign n12985 = ~n8174 & n11399 ;
  assign n12986 = n3865 & n12985 ;
  assign n12987 = n4856 ^ n3550 ^ 1'b0 ;
  assign n12988 = x24 & n2057 ;
  assign n12989 = ~n2057 & n12988 ;
  assign n12990 = ( n3869 & ~n5649 ) | ( n3869 & n9884 ) | ( ~n5649 & n9884 ) ;
  assign n12991 = n236 | n12778 ;
  assign n12992 = n2113 | n12991 ;
  assign n12993 = n6187 ^ x47 ^ 1'b0 ;
  assign n12994 = n12993 ^ x6 ^ 1'b0 ;
  assign n12995 = n2303 | n8894 ;
  assign n12996 = n12995 ^ n5412 ^ 1'b0 ;
  assign n12997 = n3501 ^ n1248 ^ 1'b0 ;
  assign n12998 = ( n853 & ~n3866 ) | ( n853 & n6714 ) | ( ~n3866 & n6714 ) ;
  assign n12999 = n7920 & n12998 ;
  assign n13000 = n12999 ^ n12041 ^ 1'b0 ;
  assign n13001 = ~n10780 & n13000 ;
  assign n13002 = n1056 | n3395 ;
  assign n13003 = ~n10905 & n13002 ;
  assign n13004 = n13003 ^ n2554 ^ 1'b0 ;
  assign n13005 = n2223 ^ n2170 ^ 1'b0 ;
  assign n13006 = ( n5962 & n9351 ) | ( n5962 & n13005 ) | ( n9351 & n13005 ) ;
  assign n13007 = n2482 | n9656 ;
  assign n13008 = n13007 ^ n6577 ^ 1'b0 ;
  assign n13009 = ~n13006 & n13008 ;
  assign n13010 = n8280 & n12957 ;
  assign n13011 = n2064 | n13010 ;
  assign n13012 = n13011 ^ n853 ^ 1'b0 ;
  assign n13013 = n11389 ^ n10276 ^ 1'b0 ;
  assign n13014 = n8102 | n13013 ;
  assign n13015 = ( n1907 & n4624 ) | ( n1907 & ~n10672 ) | ( n4624 & ~n10672 ) ;
  assign n13016 = n4477 & n6428 ;
  assign n13017 = n8276 & n13016 ;
  assign n13018 = n6781 ^ n2958 ^ 1'b0 ;
  assign n13019 = ~n13017 & n13018 ;
  assign n13020 = n10395 & n13019 ;
  assign n13021 = n13020 ^ n2419 ^ 1'b0 ;
  assign n13022 = n7828 ^ n7529 ^ 1'b0 ;
  assign n13023 = n489 & n11188 ;
  assign n13024 = ~n1062 & n13023 ;
  assign n13025 = n1556 & n10665 ;
  assign n13026 = n7050 | n7076 ;
  assign n13027 = ( n999 & n3467 ) | ( n999 & ~n13026 ) | ( n3467 & ~n13026 ) ;
  assign n13028 = n13027 ^ n1111 ^ 1'b0 ;
  assign n13029 = n13025 & n13028 ;
  assign n13030 = ( n1616 & n11054 ) | ( n1616 & ~n13029 ) | ( n11054 & ~n13029 ) ;
  assign n13031 = ( n1361 & n1631 ) | ( n1361 & n6055 ) | ( n1631 & n6055 ) ;
  assign n13032 = n11391 ^ n4972 ^ n2224 ;
  assign n13033 = n13031 & n13032 ;
  assign n13034 = n13033 ^ n2893 ^ 1'b0 ;
  assign n13035 = n13034 ^ n9192 ^ 1'b0 ;
  assign n13036 = ~x45 & n2858 ;
  assign n13037 = n4285 | n13036 ;
  assign n13038 = n8916 & ~n13037 ;
  assign n13039 = n6773 ^ n3816 ^ 1'b0 ;
  assign n13040 = n6126 | n13039 ;
  assign n13041 = ~n569 & n2243 ;
  assign n13042 = n13041 ^ n9365 ^ 1'b0 ;
  assign n13043 = n13042 ^ n1973 ^ 1'b0 ;
  assign n13044 = n7824 ^ n1392 ^ 1'b0 ;
  assign n13045 = ~n1965 & n9166 ;
  assign n13046 = n3899 & n13045 ;
  assign n13047 = ( ~n3364 & n3544 ) | ( ~n3364 & n13046 ) | ( n3544 & n13046 ) ;
  assign n13048 = n7203 ^ n1899 ^ n1895 ;
  assign n13049 = n10417 & ~n13048 ;
  assign n13050 = ~n13047 & n13049 ;
  assign n13051 = n8950 | n13050 ;
  assign n13052 = n1121 | n13051 ;
  assign n13054 = ( x99 & n400 ) | ( x99 & ~n8443 ) | ( n400 & ~n8443 ) ;
  assign n13053 = n2724 & ~n3343 ;
  assign n13055 = n13054 ^ n13053 ^ 1'b0 ;
  assign n13056 = n13055 ^ n11334 ^ 1'b0 ;
  assign n13057 = n5855 ^ n4522 ^ 1'b0 ;
  assign n13058 = n1408 ^ n1276 ^ 1'b0 ;
  assign n13059 = n8199 | n11449 ;
  assign n13060 = n10573 & ~n13059 ;
  assign n13061 = ~n3467 & n10616 ;
  assign n13062 = n5786 & n13061 ;
  assign n13068 = n6062 ^ n5443 ^ 1'b0 ;
  assign n13063 = n10152 ^ n8794 ^ 1'b0 ;
  assign n13064 = ~n1039 & n13063 ;
  assign n13065 = n2802 ^ n2652 ^ 1'b0 ;
  assign n13066 = n13064 & ~n13065 ;
  assign n13067 = ~n12564 & n13066 ;
  assign n13069 = n13068 ^ n13067 ^ 1'b0 ;
  assign n13070 = ~n1599 & n3773 ;
  assign n13071 = n9696 & n13070 ;
  assign n13072 = n13071 ^ n986 ^ 1'b0 ;
  assign n13073 = ~n2670 & n3546 ;
  assign n13074 = n13073 ^ n3830 ^ 1'b0 ;
  assign n13075 = n12839 & n13074 ;
  assign n13076 = n2945 & ~n8597 ;
  assign n13077 = n3135 & ~n13076 ;
  assign n13078 = n3107 & n13077 ;
  assign n13079 = ~n746 & n1026 ;
  assign n13080 = n13079 ^ n232 ^ 1'b0 ;
  assign n13081 = n2683 & ~n13080 ;
  assign n13082 = ~n501 & n13081 ;
  assign n13083 = n1716 & n13082 ;
  assign n13084 = n13083 ^ n3452 ^ 1'b0 ;
  assign n13085 = n9909 & n13084 ;
  assign n13086 = n7002 & n7683 ;
  assign n13087 = n13086 ^ n8302 ^ 1'b0 ;
  assign n13088 = n13087 ^ n796 ^ 1'b0 ;
  assign n13089 = n1204 & ~n5312 ;
  assign n13090 = n13089 ^ n12300 ^ 1'b0 ;
  assign n13091 = n10031 ^ n4082 ^ 1'b0 ;
  assign n13092 = n10786 | n13091 ;
  assign n13093 = n8961 | n13092 ;
  assign n13094 = n13090 | n13093 ;
  assign n13095 = n4189 & ~n13094 ;
  assign n13097 = n4126 & n5086 ;
  assign n13098 = n13097 ^ n815 ^ 1'b0 ;
  assign n13099 = n13098 ^ n10968 ^ 1'b0 ;
  assign n13096 = n494 & ~n3848 ;
  assign n13100 = n13099 ^ n13096 ^ 1'b0 ;
  assign n13101 = n3482 ^ n1549 ^ 1'b0 ;
  assign n13102 = n13100 | n13101 ;
  assign n13103 = ~n10075 & n11968 ;
  assign n13104 = ~n5014 & n13103 ;
  assign n13105 = n1469 | n7863 ;
  assign n13106 = n1649 & ~n13105 ;
  assign n13107 = n6446 & n7953 ;
  assign n13108 = n1517 ^ n620 ^ 1'b0 ;
  assign n13109 = ( n2699 & n6220 ) | ( n2699 & ~n7540 ) | ( n6220 & ~n7540 ) ;
  assign n13110 = n13108 | n13109 ;
  assign n13111 = n13110 ^ n7238 ^ 1'b0 ;
  assign n13112 = n10489 ^ n2733 ^ 1'b0 ;
  assign n13113 = n13112 ^ n5357 ^ 1'b0 ;
  assign n13114 = n1659 ^ n1354 ^ 1'b0 ;
  assign n13115 = n2126 & n4929 ;
  assign n13116 = ~n13114 & n13115 ;
  assign n13117 = n11607 | n13116 ;
  assign n13118 = n13117 ^ n6721 ^ 1'b0 ;
  assign n13119 = ~n4437 & n5815 ;
  assign n13120 = n10946 & n13119 ;
  assign n13121 = n4159 | n6809 ;
  assign n13122 = n8532 | n13121 ;
  assign n13123 = n4179 ^ n2182 ^ 1'b0 ;
  assign n13124 = n6266 | n13123 ;
  assign n13125 = n13122 | n13124 ;
  assign n13126 = n1245 & n4331 ;
  assign n13127 = n5306 ^ n363 ^ 1'b0 ;
  assign n13128 = n2388 & ~n13127 ;
  assign n13129 = n13128 ^ n10652 ^ 1'b0 ;
  assign n13130 = n2660 & ~n3331 ;
  assign n13131 = ~n7403 & n12508 ;
  assign n13132 = n11341 | n12866 ;
  assign n13133 = n12352 ^ n10157 ^ 1'b0 ;
  assign n13136 = n2938 & ~n5088 ;
  assign n13137 = n13136 ^ n4345 ^ 1'b0 ;
  assign n13134 = ~n509 & n8575 ;
  assign n13135 = n13134 ^ n2477 ^ 1'b0 ;
  assign n13138 = n13137 ^ n13135 ^ n1361 ;
  assign n13139 = n3594 & n9438 ;
  assign n13140 = n2445 & n13139 ;
  assign n13141 = n6994 & ~n7091 ;
  assign n13142 = n227 & n5302 ;
  assign n13143 = n13142 ^ n11391 ^ 1'b0 ;
  assign n13144 = ~n5467 & n13143 ;
  assign n13145 = n2090 & n13144 ;
  assign n13146 = ~n11414 & n13145 ;
  assign n13147 = n338 & n1933 ;
  assign n13148 = n4820 & ~n13147 ;
  assign n13149 = ~n1568 & n13148 ;
  assign n13150 = ~n5941 & n10072 ;
  assign n13151 = n12746 ^ n9463 ^ 1'b0 ;
  assign n13152 = n6844 & n13151 ;
  assign n13153 = n3895 & ~n7245 ;
  assign n13154 = n6277 ^ n1009 ^ 1'b0 ;
  assign n13155 = ~n2652 & n13154 ;
  assign n13156 = n13155 ^ n4566 ^ 1'b0 ;
  assign n13157 = n1300 & n6608 ;
  assign n13158 = ~n1195 & n13157 ;
  assign n13159 = n13158 ^ n1133 ^ 1'b0 ;
  assign n13160 = n7518 ^ n1484 ^ 1'b0 ;
  assign n13161 = ~n12226 & n13160 ;
  assign n13162 = n13161 ^ n1157 ^ 1'b0 ;
  assign n13163 = ~x96 & n13162 ;
  assign n13164 = n5062 ^ n152 ^ 1'b0 ;
  assign n13165 = ~n3529 & n7980 ;
  assign n13166 = n4686 & ~n13165 ;
  assign n13167 = ~n12313 & n13166 ;
  assign n13168 = n364 | n6419 ;
  assign n13169 = ~n5548 & n13031 ;
  assign n13170 = n13169 ^ n7729 ^ 1'b0 ;
  assign n13171 = n10239 ^ n7809 ^ 1'b0 ;
  assign n13172 = n6246 & n13171 ;
  assign n13173 = n5691 ^ n643 ^ 1'b0 ;
  assign n13174 = n13173 ^ n9327 ^ 1'b0 ;
  assign n13175 = n1524 & n1780 ;
  assign n13176 = n3300 & ~n13175 ;
  assign n13177 = n13176 ^ n10595 ^ n3505 ;
  assign n13178 = n10798 ^ n653 ^ 1'b0 ;
  assign n13179 = n12030 & ~n13178 ;
  assign n13180 = n1898 & n7625 ;
  assign n13181 = ~n4380 & n13180 ;
  assign n13182 = ~n5148 & n6813 ;
  assign n13183 = ~n5360 & n13182 ;
  assign n13184 = n13183 ^ n9810 ^ n1295 ;
  assign n13185 = n5963 ^ n5398 ^ 1'b0 ;
  assign n13186 = n2330 & ~n13185 ;
  assign n13187 = x34 | n5214 ;
  assign n13188 = ( n773 & n2564 ) | ( n773 & n4290 ) | ( n2564 & n4290 ) ;
  assign n13189 = n13188 ^ n8559 ^ n3203 ;
  assign n13190 = n13187 & ~n13189 ;
  assign n13191 = ~n13186 & n13190 ;
  assign n13192 = n2170 ^ x97 ^ 1'b0 ;
  assign n13193 = n11590 ^ n5644 ^ 1'b0 ;
  assign n13195 = n3706 ^ n817 ^ 1'b0 ;
  assign n13194 = ~n1860 & n12041 ;
  assign n13196 = n13195 ^ n13194 ^ 1'b0 ;
  assign n13197 = n10270 ^ n2785 ^ 1'b0 ;
  assign n13198 = n10152 & ~n10204 ;
  assign n13199 = n4897 & n6326 ;
  assign n13200 = n12969 & n13199 ;
  assign n13201 = n12807 ^ n12173 ^ 1'b0 ;
  assign n13202 = ~n2819 & n13201 ;
  assign n13203 = n6815 ^ n3561 ^ 1'b0 ;
  assign n13204 = n7428 & ~n13203 ;
  assign n13205 = n3745 | n10106 ;
  assign n13206 = n13204 | n13205 ;
  assign n13207 = n998 | n3113 ;
  assign n13208 = n3081 & ~n9990 ;
  assign n13209 = ~n801 & n13208 ;
  assign n13210 = n13209 ^ n7230 ^ n163 ;
  assign n13211 = n1150 & ~n8558 ;
  assign n13212 = ( ~n1748 & n13210 ) | ( ~n1748 & n13211 ) | ( n13210 & n13211 ) ;
  assign n13213 = n13207 & ~n13212 ;
  assign n13214 = ~n2486 & n5403 ;
  assign n13215 = n3875 & ~n11226 ;
  assign n13216 = ~n677 & n13215 ;
  assign n13217 = n3403 & n13216 ;
  assign n13218 = n11877 ^ n9258 ^ 1'b0 ;
  assign n13219 = ~n4155 & n12668 ;
  assign n13220 = n11444 ^ n2933 ^ n1792 ;
  assign n13230 = n2518 & ~n5069 ;
  assign n13231 = x39 | n1027 ;
  assign n13232 = n13230 & n13231 ;
  assign n13233 = ~n6348 & n12692 ;
  assign n13234 = ( ~n2514 & n13232 ) | ( ~n2514 & n13233 ) | ( n13232 & n13233 ) ;
  assign n13235 = n1088 & ~n13234 ;
  assign n13236 = ~n5699 & n13235 ;
  assign n13221 = n1627 ^ x22 ^ 1'b0 ;
  assign n13222 = n2433 & ~n13221 ;
  assign n13224 = n8109 ^ n257 ^ 1'b0 ;
  assign n13223 = ~n7432 & n8490 ;
  assign n13225 = n13224 ^ n13223 ^ 1'b0 ;
  assign n13226 = n13222 & ~n13225 ;
  assign n13227 = n13226 ^ n6005 ^ 1'b0 ;
  assign n13228 = n3806 & n9216 ;
  assign n13229 = n13227 & n13228 ;
  assign n13237 = n13236 ^ n13229 ^ n10687 ;
  assign n13238 = n1689 & n13237 ;
  assign n13239 = n5142 | n5227 ;
  assign n13240 = n3493 | n13239 ;
  assign n13241 = n13240 ^ n9826 ^ n4967 ;
  assign n13242 = n6048 ^ n4640 ^ 1'b0 ;
  assign n13243 = ~n1044 & n6569 ;
  assign n13244 = n13243 ^ n471 ^ 1'b0 ;
  assign n13245 = n2793 & n3378 ;
  assign n13246 = n3773 & ~n12821 ;
  assign n13247 = ~n12842 & n13246 ;
  assign n13248 = n13245 & n13247 ;
  assign n13249 = n3672 & ~n7332 ;
  assign n13250 = n13249 ^ n9094 ^ 1'b0 ;
  assign n13251 = ~n4701 & n9955 ;
  assign n13252 = n13251 ^ n6418 ^ 1'b0 ;
  assign n13253 = ~n2414 & n13252 ;
  assign n13254 = n13253 ^ n2044 ^ 1'b0 ;
  assign n13255 = n11531 & n12238 ;
  assign n13256 = n2042 & n5557 ;
  assign n13257 = n13256 ^ n11127 ^ 1'b0 ;
  assign n13258 = n6108 & ~n13257 ;
  assign n13259 = n13255 & ~n13258 ;
  assign n13260 = n1623 & ~n8613 ;
  assign n13261 = n10472 ^ n7263 ^ 1'b0 ;
  assign n13265 = n6864 ^ n4081 ^ 1'b0 ;
  assign n13263 = n7844 ^ n4250 ^ 1'b0 ;
  assign n13262 = ~n3419 & n5107 ;
  assign n13264 = n13263 ^ n13262 ^ 1'b0 ;
  assign n13266 = n13265 ^ n13264 ^ 1'b0 ;
  assign n13267 = x75 | n1941 ;
  assign n13268 = n8043 & ~n13267 ;
  assign n13269 = n1627 | n13268 ;
  assign n13270 = n13269 ^ n11723 ^ 1'b0 ;
  assign n13273 = n3918 ^ n2861 ^ 1'b0 ;
  assign n13274 = n13273 ^ n5109 ^ n3362 ;
  assign n13271 = ~n5234 & n6087 ;
  assign n13272 = n3697 & ~n13271 ;
  assign n13275 = n13274 ^ n13272 ^ 1'b0 ;
  assign n13276 = n2681 & ~n8991 ;
  assign n13277 = n4264 & n5723 ;
  assign n13278 = n1642 ^ n1582 ^ 1'b0 ;
  assign n13279 = n5012 & ~n13278 ;
  assign n13280 = ~n5248 & n13279 ;
  assign n13281 = n12418 ^ n8873 ^ n1077 ;
  assign n13282 = n11729 ^ n10831 ^ n5836 ;
  assign n13283 = n3528 | n8265 ;
  assign n13284 = n2318 & ~n13283 ;
  assign n13285 = ~n6142 & n13284 ;
  assign n13286 = n12397 & ~n13285 ;
  assign n13287 = n13286 ^ n9013 ^ 1'b0 ;
  assign n13288 = n3895 ^ n1879 ^ 1'b0 ;
  assign n13289 = n13005 & ~n13288 ;
  assign n13290 = n927 & n5320 ;
  assign n13291 = ~n3639 & n8657 ;
  assign n13292 = ~n6449 & n13291 ;
  assign n13293 = n13292 ^ n6410 ^ 1'b0 ;
  assign n13294 = n5274 & n9452 ;
  assign n13295 = ~n8368 & n8842 ;
  assign n13296 = n13295 ^ n2697 ^ 1'b0 ;
  assign n13297 = n5909 & n13296 ;
  assign n13298 = n2462 ^ x46 ^ 1'b0 ;
  assign n13299 = n942 ^ x66 ^ 1'b0 ;
  assign n13300 = n13298 & ~n13299 ;
  assign n13301 = n13300 ^ n8688 ^ 1'b0 ;
  assign n13302 = n13301 ^ n2936 ^ 1'b0 ;
  assign n13303 = n13297 & ~n13302 ;
  assign n13304 = n8339 & ~n10848 ;
  assign n13305 = n2286 & ~n8869 ;
  assign n13306 = n633 & n13305 ;
  assign n13307 = n7834 ^ n1899 ^ n733 ;
  assign n13308 = n2855 & ~n10404 ;
  assign n13309 = ~n1884 & n7437 ;
  assign n13310 = ~n13308 & n13309 ;
  assign n13311 = n3603 & ~n7320 ;
  assign n13312 = n13310 & n13311 ;
  assign n13313 = n12381 ^ n9101 ^ n6009 ;
  assign n13314 = n8335 ^ n7096 ^ n6792 ;
  assign n13315 = n2670 ^ n1250 ^ 1'b0 ;
  assign n13316 = n13315 ^ n12297 ^ 1'b0 ;
  assign n13317 = ~n9174 & n13316 ;
  assign n13318 = n1313 & ~n1776 ;
  assign n13319 = ( n11617 & n11928 ) | ( n11617 & ~n13318 ) | ( n11928 & ~n13318 ) ;
  assign n13322 = ~n1083 & n2546 ;
  assign n13323 = n13322 ^ n559 ^ 1'b0 ;
  assign n13324 = n2308 | n5075 ;
  assign n13325 = n13324 ^ n7353 ^ 1'b0 ;
  assign n13326 = ~n13323 & n13325 ;
  assign n13320 = n1393 | n12125 ;
  assign n13321 = n5569 | n13320 ;
  assign n13327 = n13326 ^ n13321 ^ 1'b0 ;
  assign n13328 = n1597 | n8183 ;
  assign n13329 = n4478 & n13328 ;
  assign n13330 = n3470 | n3751 ;
  assign n13331 = n5389 | n13330 ;
  assign n13332 = n13329 | n13331 ;
  assign n13333 = n6423 & n10901 ;
  assign n13334 = ~n3367 & n13333 ;
  assign n13336 = n1225 | n4514 ;
  assign n13335 = ~n1257 & n2673 ;
  assign n13337 = n13336 ^ n13335 ^ 1'b0 ;
  assign n13338 = n9992 ^ n3844 ^ 1'b0 ;
  assign n13341 = ( n867 & n5358 ) | ( n867 & ~n6636 ) | ( n5358 & ~n6636 ) ;
  assign n13339 = n3422 | n9192 ;
  assign n13340 = n13339 ^ n7934 ^ 1'b0 ;
  assign n13342 = n13341 ^ n13340 ^ 1'b0 ;
  assign n13343 = n1545 | n1662 ;
  assign n13344 = n13343 ^ n4808 ^ 1'b0 ;
  assign n13345 = n6631 & n13344 ;
  assign n13346 = n13345 ^ n9656 ^ 1'b0 ;
  assign n13347 = n2288 & n2512 ;
  assign n13348 = n13347 ^ n7097 ^ 1'b0 ;
  assign n13349 = n13348 ^ n2217 ^ 1'b0 ;
  assign n13350 = n13346 & ~n13349 ;
  assign n13351 = n7982 ^ n488 ^ 1'b0 ;
  assign n13352 = n7417 ^ n6259 ^ x121 ;
  assign n13353 = n5276 | n7148 ;
  assign n13354 = n1281 & ~n13353 ;
  assign n13355 = n6695 ^ n1769 ^ 1'b0 ;
  assign n13356 = x101 & ~n3410 ;
  assign n13357 = n5547 ^ n2288 ^ 1'b0 ;
  assign n13358 = n2085 | n13357 ;
  assign n13359 = n13358 ^ n4141 ^ n633 ;
  assign n13360 = ( ~n4831 & n4981 ) | ( ~n4831 & n6684 ) | ( n4981 & n6684 ) ;
  assign n13361 = n13360 ^ n1827 ^ 1'b0 ;
  assign n13362 = n9172 & n13361 ;
  assign n13363 = n6990 & n10072 ;
  assign n13364 = n11222 ^ n3604 ^ 1'b0 ;
  assign n13365 = ~n10295 & n13364 ;
  assign n13366 = n5247 & ~n12525 ;
  assign n13367 = n4865 ^ x24 ^ 1'b0 ;
  assign n13368 = n287 | n13367 ;
  assign n13369 = n9283 | n13368 ;
  assign n13370 = n13369 ^ n6700 ^ 1'b0 ;
  assign n13371 = n13370 ^ n8610 ^ n4368 ;
  assign n13372 = n3937 & ~n13371 ;
  assign n13373 = n6071 ^ n969 ^ 1'b0 ;
  assign n13374 = n13373 ^ n11280 ^ n4115 ;
  assign n13375 = ( ~n4944 & n8772 ) | ( ~n4944 & n11564 ) | ( n8772 & n11564 ) ;
  assign n13376 = n5600 ^ n985 ^ 1'b0 ;
  assign n13377 = n7519 & n13376 ;
  assign n13378 = n1450 ^ x72 ^ 1'b0 ;
  assign n13379 = n13074 & ~n13378 ;
  assign n13380 = n374 & ~n760 ;
  assign n13381 = ~n205 & n9500 ;
  assign n13382 = n884 ^ n446 ^ 1'b0 ;
  assign n13383 = ~n13381 & n13382 ;
  assign n13384 = ( n3006 & n3438 ) | ( n3006 & n8532 ) | ( n3438 & n8532 ) ;
  assign n13385 = n11142 | n13384 ;
  assign n13386 = ~n3676 & n9850 ;
  assign n13387 = n7130 ^ n1136 ^ 1'b0 ;
  assign n13388 = ~n13386 & n13387 ;
  assign n13389 = n4443 & n9706 ;
  assign n13390 = n13389 ^ n12476 ^ 1'b0 ;
  assign n13391 = n1552 | n8891 ;
  assign n13392 = n180 & ~n13391 ;
  assign n13393 = x116 & ~n13392 ;
  assign n13394 = ~n2062 & n13393 ;
  assign n13395 = ~n4566 & n7486 ;
  assign n13396 = n8548 ^ n7164 ^ 1'b0 ;
  assign n13397 = n2537 | n13396 ;
  assign n13398 = n10330 | n13397 ;
  assign n13399 = n9003 ^ n3124 ^ 1'b0 ;
  assign n13400 = ~n2130 & n2983 ;
  assign n13401 = n9351 & n13400 ;
  assign n13402 = n1469 ^ n925 ^ 1'b0 ;
  assign n13403 = n13402 ^ n11316 ^ 1'b0 ;
  assign n13404 = n1405 & n13403 ;
  assign n13405 = n5937 & ~n7510 ;
  assign n13406 = n12669 & n13405 ;
  assign n13407 = n1838 & n4262 ;
  assign n13408 = n13407 ^ n7737 ^ 1'b0 ;
  assign n13409 = n1512 & ~n13408 ;
  assign n13410 = n11873 & n13409 ;
  assign n13411 = n2849 & n3148 ;
  assign n13412 = n3308 & n13411 ;
  assign n13413 = n6700 & n13412 ;
  assign n13414 = n3251 | n13413 ;
  assign n13415 = ~n4666 & n13414 ;
  assign n13416 = ~n3381 & n12573 ;
  assign n13417 = n13416 ^ x93 ^ 1'b0 ;
  assign n13418 = n13417 ^ n9784 ^ 1'b0 ;
  assign n13419 = n7154 & n13418 ;
  assign n13420 = n13419 ^ n1599 ^ 1'b0 ;
  assign n13421 = ~n9041 & n13420 ;
  assign n13431 = n6893 & ~n9066 ;
  assign n13432 = n11736 & n13431 ;
  assign n13433 = ~n7741 & n13432 ;
  assign n13425 = n4719 ^ n4142 ^ n612 ;
  assign n13426 = n1195 & ~n13425 ;
  assign n13427 = x99 & n6636 ;
  assign n13428 = n5494 | n7130 ;
  assign n13429 = n13427 | n13428 ;
  assign n13430 = ( n1969 & ~n13426 ) | ( n1969 & n13429 ) | ( ~n13426 & n13429 ) ;
  assign n13423 = n3015 & n7049 ;
  assign n13422 = n2554 & ~n10732 ;
  assign n13424 = n13423 ^ n13422 ^ 1'b0 ;
  assign n13434 = n13433 ^ n13430 ^ n13424 ;
  assign n13435 = n3761 | n8832 ;
  assign n13436 = n2754 & n6876 ;
  assign n13439 = ( n820 & n2049 ) | ( n820 & n7829 ) | ( n2049 & n7829 ) ;
  assign n13437 = n4662 & ~n7301 ;
  assign n13438 = n1847 & ~n13437 ;
  assign n13440 = n13439 ^ n13438 ^ 1'b0 ;
  assign n13441 = ~n5945 & n13440 ;
  assign n13442 = n6277 ^ n3429 ^ 1'b0 ;
  assign n13443 = n2630 & ~n13442 ;
  assign n13444 = n11065 & n13443 ;
  assign n13445 = ~n1643 & n13444 ;
  assign n13446 = n6781 ^ n5953 ^ 1'b0 ;
  assign n13447 = ~n4705 & n5830 ;
  assign n13448 = n13447 ^ n4661 ^ 1'b0 ;
  assign n13449 = n4768 & n13448 ;
  assign n13450 = n13449 ^ n3116 ^ 1'b0 ;
  assign n13451 = n13450 ^ n8468 ^ n2476 ;
  assign n13452 = n7759 ^ n5283 ^ 1'b0 ;
  assign n13453 = n4879 ^ n1927 ^ 1'b0 ;
  assign n13454 = n1856 & n13453 ;
  assign n13455 = n371 | n10751 ;
  assign n13456 = n6245 ^ n2456 ^ 1'b0 ;
  assign n13457 = n13456 ^ n10857 ^ n883 ;
  assign n13458 = n7811 | n8651 ;
  assign n13459 = ~n290 & n13458 ;
  assign n13460 = n10334 ^ n620 ^ 1'b0 ;
  assign n13461 = n12166 & ~n13460 ;
  assign n13462 = n2042 & n4468 ;
  assign n13463 = n4299 & ~n6990 ;
  assign n13464 = n13463 ^ n8974 ^ 1'b0 ;
  assign n13465 = n9964 & n13464 ;
  assign n13466 = ( n12671 & ~n12705 ) | ( n12671 & n13465 ) | ( ~n12705 & n13465 ) ;
  assign n13467 = n4592 & n13466 ;
  assign n13468 = n8101 & n10968 ;
  assign n13469 = n8641 ^ n1538 ^ 1'b0 ;
  assign n13470 = n1535 & ~n13469 ;
  assign n13471 = n13470 ^ n6871 ^ 1'b0 ;
  assign n13472 = n2487 | n8314 ;
  assign n13473 = ~n13471 & n13472 ;
  assign n13474 = n499 | n4738 ;
  assign n13475 = n3336 & n13474 ;
  assign n13476 = ( ~n2428 & n3110 ) | ( ~n2428 & n11696 ) | ( n3110 & n11696 ) ;
  assign n13477 = ~n154 & n3726 ;
  assign n13478 = n778 & n2249 ;
  assign n13479 = ~n13477 & n13478 ;
  assign n13480 = n8040 & n8602 ;
  assign n13481 = ~n3951 & n13480 ;
  assign n13482 = n13481 ^ n11605 ^ 1'b0 ;
  assign n13483 = ~n13479 & n13482 ;
  assign n13484 = ( n12690 & ~n13476 ) | ( n12690 & n13483 ) | ( ~n13476 & n13483 ) ;
  assign n13485 = n6540 | n7337 ;
  assign n13486 = n393 & ~n13485 ;
  assign n13487 = n4301 ^ n575 ^ 1'b0 ;
  assign n13488 = n13487 ^ n3398 ^ 1'b0 ;
  assign n13489 = n205 & n11953 ;
  assign n13490 = ~n13488 & n13489 ;
  assign n13493 = n12703 ^ n4782 ^ 1'b0 ;
  assign n13494 = n4909 | n13493 ;
  assign n13491 = n1785 ^ x3 ^ 1'b0 ;
  assign n13492 = n3951 & ~n13491 ;
  assign n13495 = n13494 ^ n13492 ^ 1'b0 ;
  assign n13496 = n515 & n1376 ;
  assign n13497 = n1950 & n13496 ;
  assign n13498 = n2787 & ~n13497 ;
  assign n13499 = n13498 ^ n8712 ^ 1'b0 ;
  assign n13500 = ~n1503 & n13499 ;
  assign n13502 = n7942 ^ n4930 ^ 1'b0 ;
  assign n13501 = n3749 & ~n9344 ;
  assign n13503 = n13502 ^ n13501 ^ 1'b0 ;
  assign n13504 = ~n5965 & n8391 ;
  assign n13505 = n5747 & n13504 ;
  assign n13506 = n902 | n13505 ;
  assign n13507 = ~n1250 & n6907 ;
  assign n13508 = n9071 ^ n2433 ^ 1'b0 ;
  assign n13509 = n1708 & ~n2456 ;
  assign n13510 = n4643 | n6775 ;
  assign n13511 = n9587 & ~n13510 ;
  assign n13512 = ~n461 & n9677 ;
  assign n13513 = n13511 & n13512 ;
  assign n13514 = n1487 | n11944 ;
  assign n13515 = n8019 ^ n5634 ^ 1'b0 ;
  assign n13516 = n3439 | n13515 ;
  assign n13517 = n417 | n13516 ;
  assign n13518 = n3407 | n13517 ;
  assign n13519 = n13518 ^ n9039 ^ 1'b0 ;
  assign n13520 = n7102 ^ n3112 ^ 1'b0 ;
  assign n13521 = ( n9544 & n13235 ) | ( n9544 & n13520 ) | ( n13235 & n13520 ) ;
  assign n13522 = ~x1 & n13521 ;
  assign n13523 = n5674 ^ n3243 ^ 1'b0 ;
  assign n13524 = n737 | n4199 ;
  assign n13525 = n13523 | n13524 ;
  assign n13526 = n13525 ^ n7394 ^ 1'b0 ;
  assign n13527 = n2396 | n13526 ;
  assign n13528 = n11295 ^ n1675 ^ 1'b0 ;
  assign n13529 = n9338 ^ n2518 ^ 1'b0 ;
  assign n13530 = n13529 ^ n8571 ^ 1'b0 ;
  assign n13531 = n4338 & ~n6598 ;
  assign n13532 = n13531 ^ n10156 ^ 1'b0 ;
  assign n13533 = n9358 ^ n1338 ^ 1'b0 ;
  assign n13534 = ~n2426 & n13533 ;
  assign n13535 = n13534 ^ n1337 ^ 1'b0 ;
  assign n13536 = n2759 | n7344 ;
  assign n13537 = n7316 & ~n9524 ;
  assign n13538 = n3046 & n13537 ;
  assign n13539 = n1914 ^ n456 ^ 1'b0 ;
  assign n13540 = n5505 | n13539 ;
  assign n13541 = n12251 & ~n13540 ;
  assign n13542 = n9715 ^ n3952 ^ 1'b0 ;
  assign n13543 = n5223 & ~n13542 ;
  assign n13544 = n5574 ^ n2551 ^ 1'b0 ;
  assign n13545 = n5309 & ~n8469 ;
  assign n13552 = ~n1065 & n8431 ;
  assign n13553 = ~n4296 & n13552 ;
  assign n13547 = n1788 & n4555 ;
  assign n13548 = ~n13231 & n13547 ;
  assign n13549 = n13548 ^ n8559 ^ n7102 ;
  assign n13550 = n2593 & n13549 ;
  assign n13546 = n763 & n2154 ;
  assign n13551 = n13550 ^ n13546 ^ 1'b0 ;
  assign n13554 = n13553 ^ n13551 ^ 1'b0 ;
  assign n13555 = n7371 ^ n1599 ^ 1'b0 ;
  assign n13556 = n5034 ^ n3927 ^ 1'b0 ;
  assign n13557 = n479 & n13556 ;
  assign n13558 = n3249 | n3527 ;
  assign n13559 = n9486 | n13558 ;
  assign n13560 = n2908 | n13559 ;
  assign n13561 = ( n3514 & n9480 ) | ( n3514 & n11426 ) | ( n9480 & n11426 ) ;
  assign n13562 = n10342 | n13561 ;
  assign n13563 = n13562 ^ n7253 ^ 1'b0 ;
  assign n13564 = n464 | n11008 ;
  assign n13565 = n13564 ^ n144 ^ 1'b0 ;
  assign n13566 = ~n6148 & n13565 ;
  assign n13568 = ( x24 & n4588 ) | ( x24 & n6437 ) | ( n4588 & n6437 ) ;
  assign n13567 = n3642 & n10404 ;
  assign n13569 = n13568 ^ n13567 ^ 1'b0 ;
  assign n13570 = n2933 ^ n2890 ^ 1'b0 ;
  assign n13571 = ~n10803 & n13570 ;
  assign n13572 = n13569 | n13571 ;
  assign n13573 = ~n330 & n2494 ;
  assign n13574 = n1817 & n13573 ;
  assign n13575 = ~n5803 & n7577 ;
  assign n13576 = ~n5191 & n13575 ;
  assign n13577 = n1261 | n1485 ;
  assign n13578 = n13577 ^ n9498 ^ 1'b0 ;
  assign n13579 = n7734 | n13578 ;
  assign n13580 = n13083 ^ n11768 ^ n2146 ;
  assign n13581 = n5181 ^ n3528 ^ 1'b0 ;
  assign n13582 = n2356 & n13581 ;
  assign n13583 = n1686 & ~n6718 ;
  assign n13584 = n2735 & n10728 ;
  assign n13585 = n13583 & n13584 ;
  assign n13586 = n861 & ~n2397 ;
  assign n13587 = n7514 ^ n6151 ^ 1'b0 ;
  assign n13588 = ~n10574 & n13587 ;
  assign n13589 = n7848 ^ n3287 ^ n1555 ;
  assign n13590 = n9077 ^ n3981 ^ n3894 ;
  assign n13591 = n4793 & n11828 ;
  assign n13592 = n3603 & ~n6378 ;
  assign n13593 = n13592 ^ n2126 ^ 1'b0 ;
  assign n13594 = n5709 & ~n13593 ;
  assign n13595 = n8610 ^ x53 ^ 1'b0 ;
  assign n13596 = n1680 | n13595 ;
  assign n13597 = n13596 ^ n5224 ^ 1'b0 ;
  assign n13598 = n13594 | n13597 ;
  assign n13599 = ~n3136 & n11522 ;
  assign n13600 = n13599 ^ n1588 ^ 1'b0 ;
  assign n13601 = n3186 & n5828 ;
  assign n13602 = n4447 ^ n1742 ^ n388 ;
  assign n13603 = n3694 | n4365 ;
  assign n13604 = ~n13602 & n13603 ;
  assign n13605 = n3990 & n13604 ;
  assign n13606 = n12882 ^ n4989 ^ 1'b0 ;
  assign n13607 = n7854 | n13606 ;
  assign n13608 = ( n13601 & n13605 ) | ( n13601 & ~n13607 ) | ( n13605 & ~n13607 ) ;
  assign n13609 = n2627 ^ n816 ^ 1'b0 ;
  assign n13610 = n9165 & n10323 ;
  assign n13611 = n13469 ^ n1183 ^ 1'b0 ;
  assign n13617 = n278 | n820 ;
  assign n13618 = n278 & ~n13617 ;
  assign n13619 = ~n2109 & n13618 ;
  assign n13620 = n13619 ^ n8021 ^ 1'b0 ;
  assign n13621 = n2088 | n13620 ;
  assign n13616 = n302 | n2085 ;
  assign n13622 = n13621 ^ n13616 ^ 1'b0 ;
  assign n13612 = ~n1479 & n6279 ;
  assign n13613 = n13612 ^ n6323 ^ 1'b0 ;
  assign n13614 = n1586 & n13613 ;
  assign n13615 = ~n499 & n13614 ;
  assign n13623 = n13622 ^ n13615 ^ 1'b0 ;
  assign n13624 = n261 & n4275 ;
  assign n13625 = ~n1132 & n13624 ;
  assign n13626 = n8167 | n13625 ;
  assign n13627 = n13626 ^ n3290 ^ 1'b0 ;
  assign n13628 = n2783 | n13627 ;
  assign n13629 = n13628 ^ n13012 ^ 1'b0 ;
  assign n13630 = n2289 ^ n1355 ^ 1'b0 ;
  assign n13631 = n10198 & n11737 ;
  assign n13632 = n7790 ^ n6571 ^ 1'b0 ;
  assign n13633 = n2033 & ~n7846 ;
  assign n13634 = n3303 | n4566 ;
  assign n13635 = n3706 & n8719 ;
  assign n13636 = n10208 & n13635 ;
  assign n13637 = n5096 | n12831 ;
  assign n13638 = n13636 | n13637 ;
  assign n13639 = n13638 ^ n8872 ^ 1'b0 ;
  assign n13640 = n5277 & n10701 ;
  assign n13641 = n6657 | n11263 ;
  assign n13642 = n13641 ^ n7230 ^ 1'b0 ;
  assign n13643 = ( x24 & n6095 ) | ( x24 & ~n6684 ) | ( n6095 & ~n6684 ) ;
  assign n13644 = n12440 ^ n4773 ^ 1'b0 ;
  assign n13645 = n13643 & ~n13644 ;
  assign n13646 = ~n1863 & n7654 ;
  assign n13647 = ( ~n7505 & n9987 ) | ( ~n7505 & n13646 ) | ( n9987 & n13646 ) ;
  assign n13648 = ~n10017 & n10187 ;
  assign n13649 = n9023 & n13648 ;
  assign n13650 = n2563 & n13649 ;
  assign n13651 = n12640 ^ n8430 ^ n2222 ;
  assign n13652 = n4824 | n13651 ;
  assign n13653 = ( x119 & n5267 ) | ( x119 & n7578 ) | ( n5267 & n7578 ) ;
  assign n13654 = n2961 & n10540 ;
  assign n13655 = n5493 & ~n7527 ;
  assign n13656 = n13655 ^ n5365 ^ 1'b0 ;
  assign n13657 = n10333 ^ n7992 ^ 1'b0 ;
  assign n13658 = n6107 & n13657 ;
  assign n13659 = n13658 ^ n1446 ^ 1'b0 ;
  assign n13660 = n13656 & n13659 ;
  assign n13661 = n4018 ^ n901 ^ 1'b0 ;
  assign n13662 = n6667 & n12206 ;
  assign n13663 = ~n5709 & n7621 ;
  assign n13664 = ~n362 & n13663 ;
  assign n13665 = ~n922 & n2596 ;
  assign n13666 = n13665 ^ n3196 ^ 1'b0 ;
  assign n13667 = n6306 | n6695 ;
  assign n13668 = n12634 ^ n11487 ^ n1596 ;
  assign n13669 = n1625 ^ n1611 ^ 1'b0 ;
  assign n13670 = n10318 & ~n13669 ;
  assign n13671 = n5951 & n13670 ;
  assign n13672 = n13671 ^ n8959 ^ n7749 ;
  assign n13673 = ~n699 & n5302 ;
  assign n13674 = n13673 ^ n1353 ^ 1'b0 ;
  assign n13675 = ( ~n6273 & n6629 ) | ( ~n6273 & n13674 ) | ( n6629 & n13674 ) ;
  assign n13676 = n13675 ^ n3110 ^ 1'b0 ;
  assign n13677 = n3620 & n13676 ;
  assign n13678 = n11917 ^ n1037 ^ 1'b0 ;
  assign n13679 = x113 & ~n10545 ;
  assign n13680 = n13679 ^ n5885 ^ n4527 ;
  assign n13681 = n5050 & n10528 ;
  assign n13682 = n13681 ^ n1558 ^ 1'b0 ;
  assign n13683 = n7192 & ~n13682 ;
  assign n13684 = ~n9811 & n13683 ;
  assign n13685 = n13684 ^ n2615 ^ 1'b0 ;
  assign n13686 = n11144 | n13685 ;
  assign n13687 = ~n13680 & n13686 ;
  assign n13688 = n13687 ^ n5245 ^ 1'b0 ;
  assign n13689 = ~n1639 & n8946 ;
  assign n13690 = n8227 ^ n2872 ^ 1'b0 ;
  assign n13691 = n10140 & ~n13690 ;
  assign n13692 = n7818 ^ n3681 ^ 1'b0 ;
  assign n13693 = n13692 ^ n5694 ^ 1'b0 ;
  assign n13695 = n2364 ^ n363 ^ 1'b0 ;
  assign n13696 = n3595 & ~n13695 ;
  assign n13694 = n3733 & n11143 ;
  assign n13697 = n13696 ^ n13694 ^ 1'b0 ;
  assign n13698 = ~n2762 & n13697 ;
  assign n13699 = n6264 ^ n3165 ^ 1'b0 ;
  assign n13700 = n3655 ^ n3601 ^ 1'b0 ;
  assign n13701 = n2778 & n13700 ;
  assign n13702 = n13699 & n13701 ;
  assign n13703 = n8940 & ~n11783 ;
  assign n13704 = n1046 & n6103 ;
  assign n13705 = ~n12625 & n13704 ;
  assign n13706 = ~n3757 & n13705 ;
  assign n13709 = ~n884 & n1429 ;
  assign n13708 = ~n2201 & n8219 ;
  assign n13710 = n13709 ^ n13708 ^ 1'b0 ;
  assign n13711 = n363 | n13710 ;
  assign n13712 = n13711 ^ n6011 ^ 1'b0 ;
  assign n13713 = n13712 ^ n4348 ^ 1'b0 ;
  assign n13707 = x35 & n5219 ;
  assign n13714 = n13713 ^ n13707 ^ 1'b0 ;
  assign n13715 = n3793 & n13196 ;
  assign n13716 = ~n12998 & n13715 ;
  assign n13717 = n5857 ^ n614 ^ 1'b0 ;
  assign n13718 = n1337 & n13717 ;
  assign n13719 = ~n10144 & n13718 ;
  assign n13720 = n1898 ^ n1481 ^ 1'b0 ;
  assign n13721 = n13215 & n13720 ;
  assign n13722 = n3238 ^ n484 ^ 1'b0 ;
  assign n13723 = n180 | n5036 ;
  assign n13724 = n13723 ^ n580 ^ 1'b0 ;
  assign n13725 = n1874 & n13724 ;
  assign n13726 = n13725 ^ n12308 ^ 1'b0 ;
  assign n13727 = n13722 | n13726 ;
  assign n13728 = n13568 ^ n6135 ^ 1'b0 ;
  assign n13729 = n152 | n5365 ;
  assign n13730 = n4353 & n4765 ;
  assign n13731 = n13729 | n13730 ;
  assign n13733 = n1908 & n3630 ;
  assign n13734 = n13733 ^ n2603 ^ 1'b0 ;
  assign n13732 = n1285 | n4944 ;
  assign n13735 = n13734 ^ n13732 ^ 1'b0 ;
  assign n13736 = n4824 & ~n5191 ;
  assign n13737 = n6557 ^ n855 ^ 1'b0 ;
  assign n13738 = n8343 & n13737 ;
  assign n13739 = n13128 & ~n13738 ;
  assign n13740 = n2176 & n2679 ;
  assign n13741 = n13740 ^ n1037 ^ 1'b0 ;
  assign n13742 = n2140 & ~n12918 ;
  assign n13743 = ~n13741 & n13742 ;
  assign n13744 = n8746 ^ n4416 ^ n2000 ;
  assign n13745 = n2752 | n13744 ;
  assign n13746 = n1145 & n10683 ;
  assign n13747 = n13746 ^ n9176 ^ n7032 ;
  assign n13748 = n559 & ~n13747 ;
  assign n13749 = n857 & ~n3283 ;
  assign n13750 = n13749 ^ n13340 ^ 1'b0 ;
  assign n13751 = n4028 & ~n13750 ;
  assign n13752 = ~n3333 & n13751 ;
  assign n13753 = n5061 & ~n10330 ;
  assign n13754 = n13753 ^ n6181 ^ 1'b0 ;
  assign n13755 = n12887 ^ n8304 ^ n3802 ;
  assign n13756 = ( ~n8284 & n13754 ) | ( ~n8284 & n13755 ) | ( n13754 & n13755 ) ;
  assign n13757 = n4742 | n12308 ;
  assign n13758 = n799 & ~n956 ;
  assign n13759 = n3626 & ~n13758 ;
  assign n13760 = n13759 ^ n12974 ^ 1'b0 ;
  assign n13761 = n13757 | n13760 ;
  assign n13762 = n7002 & n12282 ;
  assign n13763 = ~n4836 & n13762 ;
  assign n13764 = n9525 ^ n6981 ^ 1'b0 ;
  assign n13765 = n2739 & n12500 ;
  assign n13766 = n12144 ^ n11910 ^ 1'b0 ;
  assign n13767 = ~n5494 & n13766 ;
  assign n13768 = n13767 ^ n11111 ^ 1'b0 ;
  assign n13769 = n13551 ^ n8335 ^ 1'b0 ;
  assign n13770 = n5319 ^ n3368 ^ 1'b0 ;
  assign n13771 = n4734 & n13770 ;
  assign n13772 = ( n569 & n9813 ) | ( n569 & ~n13771 ) | ( n9813 & ~n13771 ) ;
  assign n13773 = ~n3198 & n3758 ;
  assign n13774 = n12813 & n13773 ;
  assign n13775 = n4633 | n6071 ;
  assign n13776 = ~n852 & n13775 ;
  assign n13777 = n13776 ^ n4708 ^ 1'b0 ;
  assign n13778 = n2696 & n3058 ;
  assign n13779 = n13777 & n13778 ;
  assign n13780 = n9801 & ~n13779 ;
  assign n13781 = n1045 & ~n4817 ;
  assign n13782 = n6038 ^ n636 ^ 1'b0 ;
  assign n13783 = n11162 ^ n8365 ^ 1'b0 ;
  assign n13784 = n8720 ^ n5193 ^ 1'b0 ;
  assign n13785 = n13230 | n13784 ;
  assign n13786 = n13210 ^ n8916 ^ 1'b0 ;
  assign n13788 = n986 ^ n376 ^ 1'b0 ;
  assign n13789 = n7185 & n13788 ;
  assign n13790 = ~n4778 & n13789 ;
  assign n13791 = n4443 & n13790 ;
  assign n13787 = n4868 & ~n5683 ;
  assign n13792 = n13791 ^ n13787 ^ 1'b0 ;
  assign n13793 = n1172 & ~n3090 ;
  assign n13794 = n13793 ^ n5214 ^ 1'b0 ;
  assign n13795 = n13794 ^ n1985 ^ 1'b0 ;
  assign n13796 = n8693 ^ x35 ^ 1'b0 ;
  assign n13797 = n8654 ^ n1300 ^ n763 ;
  assign n13798 = n12221 ^ n7472 ^ 1'b0 ;
  assign n13799 = ( ~n7348 & n13797 ) | ( ~n7348 & n13798 ) | ( n13797 & n13798 ) ;
  assign n13800 = ( n2450 & n7971 ) | ( n2450 & n13799 ) | ( n7971 & n13799 ) ;
  assign n13801 = n2348 & n5871 ;
  assign n13802 = n13801 ^ x73 ^ 1'b0 ;
  assign n13803 = n13802 ^ n3528 ^ 1'b0 ;
  assign n13804 = n4212 & n13803 ;
  assign n13805 = n1026 | n12715 ;
  assign n13806 = n2093 & n5119 ;
  assign n13807 = n1505 & ~n13806 ;
  assign n13808 = n5643 & n13807 ;
  assign n13809 = n1205 | n5319 ;
  assign n13810 = n3751 | n7358 ;
  assign n13811 = n6604 & ~n11768 ;
  assign n13812 = n13811 ^ n713 ^ 1'b0 ;
  assign n13813 = n2086 & n13812 ;
  assign n13814 = n13813 ^ n3249 ^ 1'b0 ;
  assign n13815 = n13814 ^ n1914 ^ 1'b0 ;
  assign n13816 = n3811 & ~n3869 ;
  assign n13817 = n4765 & ~n11437 ;
  assign n13823 = n4230 & n6465 ;
  assign n13824 = ~x18 & n13823 ;
  assign n13818 = n2518 & ~n4075 ;
  assign n13819 = n13818 ^ n2856 ^ 1'b0 ;
  assign n13820 = n11272 & n13819 ;
  assign n13821 = n12601 ^ n3098 ^ 1'b0 ;
  assign n13822 = n13820 & n13821 ;
  assign n13825 = n13824 ^ n13822 ^ 1'b0 ;
  assign n13826 = n13825 ^ n9997 ^ 1'b0 ;
  assign n13827 = n7102 & ~n13826 ;
  assign n13828 = n5367 ^ n3433 ^ 1'b0 ;
  assign n13829 = n11160 & ~n13828 ;
  assign n13830 = n511 & n13829 ;
  assign n13831 = n1801 & ~n2827 ;
  assign n13832 = n13831 ^ n4548 ^ 1'b0 ;
  assign n13833 = n10362 & n13832 ;
  assign n13834 = n12295 ^ n8662 ^ 1'b0 ;
  assign n13835 = x57 & n11212 ;
  assign n13836 = n13835 ^ n1511 ^ 1'b0 ;
  assign n13837 = n9879 & ~n13836 ;
  assign n13838 = n13837 ^ n4973 ^ 1'b0 ;
  assign n13839 = n7033 & n13838 ;
  assign n13840 = ( n1737 & n2206 ) | ( n1737 & n3171 ) | ( n2206 & n3171 ) ;
  assign n13841 = ~n6294 & n11995 ;
  assign n13842 = n4476 | n7942 ;
  assign n13843 = n13119 ^ n2704 ^ 1'b0 ;
  assign n13844 = n13842 & n13843 ;
  assign n13845 = n9340 ^ n4084 ^ 1'b0 ;
  assign n13846 = ~n7419 & n13845 ;
  assign n13847 = n13846 ^ n5962 ^ 1'b0 ;
  assign n13848 = n8641 ^ n1532 ^ 1'b0 ;
  assign n13849 = n13847 | n13848 ;
  assign n13850 = ~n4872 & n8158 ;
  assign n13851 = ( n3840 & ~n13593 ) | ( n3840 & n13850 ) | ( ~n13593 & n13850 ) ;
  assign n13852 = n10882 ^ n7438 ^ 1'b0 ;
  assign n13853 = n4503 & n13852 ;
  assign n13854 = n3374 ^ n2484 ^ 1'b0 ;
  assign n13855 = n6949 | n13854 ;
  assign n13856 = n8976 ^ n3203 ^ 1'b0 ;
  assign n13857 = n2846 & ~n13856 ;
  assign n13858 = n5728 | n12420 ;
  assign n13859 = n13857 | n13858 ;
  assign n13860 = n9894 ^ n2866 ^ 1'b0 ;
  assign n13861 = n11822 & n13860 ;
  assign n13862 = ~n3750 & n8868 ;
  assign n13863 = n13862 ^ n4505 ^ 1'b0 ;
  assign n13864 = ~n362 & n2351 ;
  assign n13865 = n13864 ^ n1487 ^ 1'b0 ;
  assign n13866 = n3764 | n13865 ;
  assign n13867 = n13866 ^ n5403 ^ 1'b0 ;
  assign n13868 = n6079 ^ n4944 ^ 1'b0 ;
  assign n13869 = ~n3482 & n13868 ;
  assign n13870 = ~n13867 & n13869 ;
  assign n13871 = ~n674 & n2851 ;
  assign n13872 = n13871 ^ n3778 ^ 1'b0 ;
  assign n13873 = n13872 ^ n4002 ^ 1'b0 ;
  assign n13874 = ~n6335 & n13873 ;
  assign n13875 = ~n4605 & n10417 ;
  assign n13876 = n5111 & n13875 ;
  assign n13877 = ~n2794 & n3115 ;
  assign n13878 = n13877 ^ n2889 ^ 1'b0 ;
  assign n13879 = n13878 ^ n8910 ^ 1'b0 ;
  assign n13880 = n3930 & n13879 ;
  assign n13881 = n2308 & n11379 ;
  assign n13882 = n13881 ^ n484 ^ 1'b0 ;
  assign n13883 = n4888 & n13882 ;
  assign n13884 = n7948 & n13883 ;
  assign n13885 = n7992 ^ n7426 ^ n5915 ;
  assign n13886 = n10296 ^ n1473 ^ 1'b0 ;
  assign n13887 = n3039 & ~n13886 ;
  assign n13888 = n13887 ^ n4888 ^ 1'b0 ;
  assign n13889 = n8297 ^ n3119 ^ 1'b0 ;
  assign n13890 = n11598 & ~n13889 ;
  assign n13891 = n7542 ^ n3755 ^ 1'b0 ;
  assign n13892 = ~n11367 & n13891 ;
  assign n13893 = n224 & n3207 ;
  assign n13894 = n13893 ^ n916 ^ 1'b0 ;
  assign n13895 = n2696 ^ n1865 ^ 1'b0 ;
  assign n13896 = n10198 | n13895 ;
  assign n13897 = ~n1879 & n2046 ;
  assign n13898 = n1446 & n13897 ;
  assign n13899 = n3822 | n8945 ;
  assign n13900 = n8517 ^ n951 ^ 1'b0 ;
  assign n13901 = n904 & ~n2769 ;
  assign n13902 = n13901 ^ n8491 ^ 1'b0 ;
  assign n13903 = ~n4324 & n11507 ;
  assign n13904 = ( ~n1398 & n11475 ) | ( ~n1398 & n12017 ) | ( n11475 & n12017 ) ;
  assign n13905 = ( n8658 & ~n13903 ) | ( n8658 & n13904 ) | ( ~n13903 & n13904 ) ;
  assign n13907 = n7988 & n11554 ;
  assign n13906 = n3241 & n10527 ;
  assign n13908 = n13907 ^ n13906 ^ 1'b0 ;
  assign n13909 = n10001 ^ n6904 ^ 1'b0 ;
  assign n13910 = n7175 ^ n4498 ^ 1'b0 ;
  assign n13911 = n2330 | n2797 ;
  assign n13912 = n10252 ^ x56 ^ 1'b0 ;
  assign n13913 = n1828 | n2924 ;
  assign n13914 = n1662 & ~n13913 ;
  assign n13915 = n4553 ^ n1786 ^ 1'b0 ;
  assign n13916 = n1500 | n13915 ;
  assign n13917 = ~n637 & n9039 ;
  assign n13918 = n4014 & ~n8304 ;
  assign n13919 = n13918 ^ x18 ^ 1'b0 ;
  assign n13920 = n2234 & ~n13919 ;
  assign n13921 = ~n6985 & n13920 ;
  assign n13922 = n11379 & ~n13921 ;
  assign n13923 = ~n1740 & n6423 ;
  assign n13924 = n7416 & n13923 ;
  assign n13925 = n2293 | n5484 ;
  assign n13926 = n13925 ^ n8704 ^ 1'b0 ;
  assign n13927 = n1182 | n5134 ;
  assign n13928 = n1971 | n13927 ;
  assign n13929 = n13928 ^ n7324 ^ 1'b0 ;
  assign n13930 = n10157 ^ n835 ^ 1'b0 ;
  assign n13931 = n525 | n1469 ;
  assign n13932 = n3165 | n12677 ;
  assign n13933 = n826 ^ n351 ^ 1'b0 ;
  assign n13934 = n3481 & n13933 ;
  assign n13935 = n4182 | n9476 ;
  assign n13936 = ( n431 & ~n11265 ) | ( n431 & n13935 ) | ( ~n11265 & n13935 ) ;
  assign n13937 = n2306 ^ n2113 ^ 1'b0 ;
  assign n13938 = n13937 ^ n2905 ^ 1'b0 ;
  assign n13939 = n2433 & ~n13938 ;
  assign n13940 = n13939 ^ n9446 ^ 1'b0 ;
  assign n13941 = ~n7008 & n13940 ;
  assign n13942 = ~n4757 & n6244 ;
  assign n13943 = n13591 ^ n6364 ^ n1040 ;
  assign n13945 = n3403 | n5952 ;
  assign n13946 = n13945 ^ n11250 ^ 1'b0 ;
  assign n13944 = n879 & ~n7055 ;
  assign n13947 = n13946 ^ n13944 ^ 1'b0 ;
  assign n13948 = n2435 & n10008 ;
  assign n13949 = ~n4299 & n13948 ;
  assign n13950 = n4838 | n12310 ;
  assign n13951 = ( n3206 & n7536 ) | ( n3206 & n7946 ) | ( n7536 & n7946 ) ;
  assign n13952 = n1338 & n4983 ;
  assign n13953 = n1254 & n13952 ;
  assign n13954 = n10739 | n13953 ;
  assign n13955 = n13951 | n13954 ;
  assign n13956 = n1862 & ~n5424 ;
  assign n13957 = ~n7529 & n13956 ;
  assign n13958 = x93 & n3444 ;
  assign n13959 = n6628 | n13958 ;
  assign n13960 = n4619 ^ n4240 ^ 1'b0 ;
  assign n13961 = n4953 | n5133 ;
  assign n13962 = n6461 & n8448 ;
  assign n13963 = n2602 & n3974 ;
  assign n13964 = n978 & ~n2656 ;
  assign n13965 = n1888 ^ n574 ^ x81 ;
  assign n13966 = n13965 ^ n10090 ^ 1'b0 ;
  assign n13969 = ~n2170 & n3368 ;
  assign n13967 = n2228 & n8346 ;
  assign n13968 = n13967 ^ n3850 ^ 1'b0 ;
  assign n13970 = n13969 ^ n13968 ^ n6899 ;
  assign n13971 = n13775 & ~n13970 ;
  assign n13972 = n9189 ^ n5268 ^ n1754 ;
  assign n13973 = n269 & n13972 ;
  assign n13974 = n4206 & n5599 ;
  assign n13975 = ~n6408 & n13974 ;
  assign n13976 = n10225 ^ n8490 ^ 1'b0 ;
  assign n13978 = ~n742 & n3501 ;
  assign n13977 = n6523 & ~n11389 ;
  assign n13979 = n13978 ^ n13977 ^ 1'b0 ;
  assign n13980 = n9529 ^ n4942 ^ 1'b0 ;
  assign n13981 = ~n756 & n13980 ;
  assign n13982 = n13981 ^ n2933 ^ n1847 ;
  assign n13983 = n4527 ^ n928 ^ 1'b0 ;
  assign n13984 = ~n13982 & n13983 ;
  assign n13985 = n3799 ^ n2235 ^ 1'b0 ;
  assign n13986 = n13820 & ~n13985 ;
  assign n13987 = ( n3606 & ~n9012 ) | ( n3606 & n9827 ) | ( ~n9012 & n9827 ) ;
  assign n13988 = n1681 & n7465 ;
  assign n13992 = n4792 | n7828 ;
  assign n13993 = n13992 ^ n4895 ^ 1'b0 ;
  assign n13994 = n5874 & ~n13993 ;
  assign n13991 = n12448 & n13758 ;
  assign n13995 = n13994 ^ n13991 ^ n406 ;
  assign n13989 = n6961 ^ n3950 ^ 1'b0 ;
  assign n13990 = n12702 & ~n13989 ;
  assign n13996 = n13995 ^ n13990 ^ 1'b0 ;
  assign n13997 = n13996 ^ n2740 ^ 1'b0 ;
  assign n13998 = n236 | n5705 ;
  assign n13999 = n13998 ^ n760 ^ 1'b0 ;
  assign n14000 = n5161 & ~n13999 ;
  assign n14001 = ~n1793 & n14000 ;
  assign n14002 = n7951 & n14001 ;
  assign n14003 = n788 & ~n8298 ;
  assign n14004 = n14002 & n14003 ;
  assign n14005 = n9538 & n10586 ;
  assign n14006 = n14005 ^ n7609 ^ 1'b0 ;
  assign n14007 = n2020 | n7181 ;
  assign n14008 = n5592 & ~n7260 ;
  assign n14009 = n922 & n14008 ;
  assign n14010 = n14007 | n14009 ;
  assign n14011 = n6157 | n14010 ;
  assign n14012 = n4307 & ~n4661 ;
  assign n14013 = n2601 & n8013 ;
  assign n14014 = n4351 & n14013 ;
  assign n14015 = n3615 ^ n414 ^ 1'b0 ;
  assign n14016 = n6323 & ~n14015 ;
  assign n14017 = ~n4970 & n14016 ;
  assign n14018 = n14014 & n14017 ;
  assign n14019 = n695 & n11732 ;
  assign n14020 = n14018 | n14019 ;
  assign n14021 = n2694 ^ x75 ^ 1'b0 ;
  assign n14022 = n1206 & ~n14021 ;
  assign n14023 = n14022 ^ n6677 ^ 1'b0 ;
  assign n14024 = n1761 ^ x117 ^ 1'b0 ;
  assign n14025 = n3717 ^ n1011 ^ 1'b0 ;
  assign n14027 = ( n3626 & ~n6049 ) | ( n3626 & n7112 ) | ( ~n6049 & n7112 ) ;
  assign n14026 = n5417 | n9871 ;
  assign n14028 = n14027 ^ n14026 ^ 1'b0 ;
  assign n14029 = ( n1771 & n14025 ) | ( n1771 & n14028 ) | ( n14025 & n14028 ) ;
  assign n14030 = n9366 | n12842 ;
  assign n14031 = n14030 ^ n13599 ^ 1'b0 ;
  assign n14032 = ~n2958 & n12342 ;
  assign n14033 = n12283 & n14032 ;
  assign n14034 = ( ~n2450 & n3131 ) | ( ~n2450 & n4969 ) | ( n3131 & n4969 ) ;
  assign n14035 = n3673 ^ n1861 ^ 1'b0 ;
  assign n14036 = n1206 & ~n14035 ;
  assign n14037 = n3143 & n14036 ;
  assign n14038 = n14037 ^ n13979 ^ n7875 ;
  assign n14039 = n6972 ^ n5378 ^ 1'b0 ;
  assign n14040 = n11527 ^ n2679 ^ 1'b0 ;
  assign n14041 = n14040 ^ n4846 ^ 1'b0 ;
  assign n14042 = n4710 | n6655 ;
  assign n14043 = n14042 ^ n5514 ^ 1'b0 ;
  assign n14044 = n8314 ^ n7855 ^ 1'b0 ;
  assign n14045 = n4557 & ~n14044 ;
  assign n14046 = ~n14043 & n14045 ;
  assign n14047 = n8122 ^ n6630 ^ 1'b0 ;
  assign n14048 = n5316 & ~n14047 ;
  assign n14049 = n14048 ^ n6770 ^ n1114 ;
  assign n14050 = n9098 ^ n4678 ^ n3951 ;
  assign n14051 = n3993 | n9367 ;
  assign n14052 = n14050 & ~n14051 ;
  assign n14053 = n14049 & ~n14052 ;
  assign n14054 = n14053 ^ n8267 ^ 1'b0 ;
  assign n14055 = n12095 ^ x14 ^ 1'b0 ;
  assign n14056 = n5015 | n5165 ;
  assign n14057 = n14056 ^ n2458 ^ 1'b0 ;
  assign n14058 = n2464 & n4010 ;
  assign n14059 = n14058 ^ n7558 ^ 1'b0 ;
  assign n14060 = n2180 & n4731 ;
  assign n14061 = ~n688 & n14060 ;
  assign n14062 = n14061 ^ n1132 ^ 1'b0 ;
  assign n14063 = n8185 | n14062 ;
  assign n14064 = n2136 | n12852 ;
  assign n14065 = n4190 ^ n3442 ^ 1'b0 ;
  assign n14066 = ~n3437 & n14065 ;
  assign n14067 = n14066 ^ n2091 ^ 1'b0 ;
  assign n14068 = ~n14064 & n14067 ;
  assign n14069 = n6742 ^ n4089 ^ 1'b0 ;
  assign n14070 = n6508 | n14069 ;
  assign n14071 = ~n1913 & n11933 ;
  assign n14072 = n14070 & n14071 ;
  assign n14081 = n6938 ^ n1939 ^ 1'b0 ;
  assign n14073 = n7683 ^ n7527 ^ n458 ;
  assign n14074 = n6876 & ~n14073 ;
  assign n14075 = n14074 ^ n12235 ^ 1'b0 ;
  assign n14076 = n2492 | n10291 ;
  assign n14077 = n679 & ~n4068 ;
  assign n14078 = n14076 & ~n14077 ;
  assign n14079 = n14078 ^ n6401 ^ 1'b0 ;
  assign n14080 = n14075 & n14079 ;
  assign n14082 = n14081 ^ n14080 ^ 1'b0 ;
  assign n14083 = n7977 ^ n5268 ^ n860 ;
  assign n14084 = n14083 ^ n3415 ^ 1'b0 ;
  assign n14085 = x14 & ~n12267 ;
  assign n14086 = n11153 & ~n14085 ;
  assign n14087 = n7645 ^ n4260 ^ 1'b0 ;
  assign n14088 = n6050 & n14087 ;
  assign n14089 = ( n1076 & n3072 ) | ( n1076 & n8144 ) | ( n3072 & n8144 ) ;
  assign n14090 = n374 | n8317 ;
  assign n14091 = n14090 ^ n14040 ^ n2059 ;
  assign n14092 = n2313 | n14091 ;
  assign n14093 = n2057 | n3204 ;
  assign n14094 = n14093 ^ n13736 ^ n1438 ;
  assign n14095 = n11828 ^ n7505 ^ 1'b0 ;
  assign n14096 = n14094 & n14095 ;
  assign n14097 = n6550 ^ n2712 ^ n1361 ;
  assign n14098 = n5868 ^ n4355 ^ 1'b0 ;
  assign n14099 = n3907 | n14098 ;
  assign n14100 = n14099 ^ n7846 ^ 1'b0 ;
  assign n14101 = n12866 ^ n6775 ^ 1'b0 ;
  assign n14102 = ~n14100 & n14101 ;
  assign n14103 = n12309 ^ n7126 ^ 1'b0 ;
  assign n14104 = n8195 | n14103 ;
  assign n14105 = n2351 | n8643 ;
  assign n14106 = n7158 & n14105 ;
  assign n14107 = n11795 & n14106 ;
  assign n14108 = ( n2044 & n3719 ) | ( n2044 & ~n10105 ) | ( n3719 & ~n10105 ) ;
  assign n14109 = n14108 ^ n2130 ^ 1'b0 ;
  assign n14110 = ~n4881 & n9523 ;
  assign n14111 = n3334 & n4348 ;
  assign n14112 = n14111 ^ n4136 ^ 1'b0 ;
  assign n14113 = n8726 & ~n14112 ;
  assign n14114 = ~n8545 & n10161 ;
  assign n14115 = n14114 ^ n4536 ^ 1'b0 ;
  assign n14116 = ~n2295 & n13274 ;
  assign n14117 = ( n4018 & ~n9093 ) | ( n4018 & n13227 ) | ( ~n9093 & n13227 ) ;
  assign n14118 = n3222 | n5983 ;
  assign n14119 = n14118 ^ n5134 ^ 1'b0 ;
  assign n14120 = n14119 ^ n6523 ^ 1'b0 ;
  assign n14121 = n709 | n14120 ;
  assign n14125 = n6568 ^ n4676 ^ 1'b0 ;
  assign n14126 = n4640 & ~n14125 ;
  assign n14122 = n1464 & ~n11882 ;
  assign n14123 = n14122 ^ n5034 ^ 1'b0 ;
  assign n14124 = n8915 | n14123 ;
  assign n14127 = n14126 ^ n14124 ^ 1'b0 ;
  assign n14128 = n1083 & n6827 ;
  assign n14129 = n12505 & n14128 ;
  assign n14130 = n14127 & n14129 ;
  assign n14131 = n6374 ^ n4701 ^ 1'b0 ;
  assign n14132 = n3478 & n14131 ;
  assign n14133 = n14132 ^ n13518 ^ 1'b0 ;
  assign n14134 = n3875 & n14133 ;
  assign n14135 = n7982 ^ x109 ^ 1'b0 ;
  assign n14136 = ~n685 & n5855 ;
  assign n14137 = n14136 ^ n941 ^ 1'b0 ;
  assign n14138 = n13143 ^ n1024 ^ x6 ;
  assign n14139 = n14137 & ~n14138 ;
  assign n14140 = ~n12549 & n14139 ;
  assign n14141 = n13899 & ~n14140 ;
  assign n14142 = n5803 & n14141 ;
  assign n14143 = n2392 & ~n7481 ;
  assign n14144 = n3246 & ~n14143 ;
  assign n14147 = n4345 ^ n1948 ^ 1'b0 ;
  assign n14148 = n14147 ^ n6004 ^ n5415 ;
  assign n14149 = ( ~n546 & n2558 ) | ( ~n546 & n14148 ) | ( n2558 & n14148 ) ;
  assign n14145 = ~n749 & n6060 ;
  assign n14146 = ~n6114 & n14145 ;
  assign n14150 = n14149 ^ n14146 ^ 1'b0 ;
  assign n14151 = n2603 & ~n14150 ;
  assign n14152 = n9356 & ~n14151 ;
  assign n14153 = n8384 ^ n1479 ^ 1'b0 ;
  assign n14154 = ~n655 & n1211 ;
  assign n14155 = n742 ^ x8 ^ 1'b0 ;
  assign n14156 = n666 | n14155 ;
  assign n14157 = n1996 & ~n14156 ;
  assign n14158 = n10453 & ~n14157 ;
  assign n14159 = ~n14154 & n14158 ;
  assign n14160 = n14159 ^ n8710 ^ 1'b0 ;
  assign n14161 = ~n8155 & n9290 ;
  assign n14162 = n14161 ^ n2660 ^ 1'b0 ;
  assign n14163 = n4468 ^ n909 ^ 1'b0 ;
  assign n14164 = n10361 | n14163 ;
  assign n14165 = n2948 | n7221 ;
  assign n14166 = n5043 | n14165 ;
  assign n14167 = n2026 & n3069 ;
  assign n14168 = n14167 ^ n8384 ^ 1'b0 ;
  assign n14169 = n14166 & ~n14168 ;
  assign n14170 = n2659 | n9787 ;
  assign n14171 = n4877 | n13867 ;
  assign n14172 = n1458 & ~n5163 ;
  assign n14173 = x100 & n3384 ;
  assign n14174 = n5007 & ~n14173 ;
  assign n14175 = ~n14172 & n14174 ;
  assign n14176 = n3353 & ~n6707 ;
  assign n14177 = n3249 & n14176 ;
  assign n14178 = n6416 ^ x87 ^ 1'b0 ;
  assign n14179 = n2965 & n14178 ;
  assign n14180 = n10934 ^ n5277 ^ 1'b0 ;
  assign n14181 = n1931 & ~n14180 ;
  assign n14182 = n14181 ^ n12236 ^ 1'b0 ;
  assign n14183 = ~n324 & n14045 ;
  assign n14184 = n14183 ^ n10072 ^ 1'b0 ;
  assign n14185 = n3547 ^ n801 ^ 1'b0 ;
  assign n14186 = n14185 ^ n2412 ^ 1'b0 ;
  assign n14187 = n6854 | n14186 ;
  assign n14188 = n324 | n5059 ;
  assign n14189 = ~n9773 & n14188 ;
  assign n14190 = ~n14187 & n14189 ;
  assign n14191 = n7905 | n8006 ;
  assign n14192 = n6673 & ~n14191 ;
  assign n14193 = ~n6105 & n6508 ;
  assign n14194 = n11931 & n12062 ;
  assign n14195 = n14193 & n14194 ;
  assign n14197 = n3682 | n6378 ;
  assign n14198 = n4675 & ~n14197 ;
  assign n14199 = n1568 & ~n5865 ;
  assign n14200 = n14198 & n14199 ;
  assign n14196 = n12561 ^ n506 ^ 1'b0 ;
  assign n14201 = n14200 ^ n14196 ^ 1'b0 ;
  assign n14202 = n14201 ^ n9590 ^ 1'b0 ;
  assign n14203 = n11081 ^ n7575 ^ 1'b0 ;
  assign n14204 = n7927 | n14203 ;
  assign n14205 = n198 & ~n2751 ;
  assign n14206 = n9885 ^ n1819 ^ 1'b0 ;
  assign n14207 = n7277 ^ n3594 ^ n2265 ;
  assign n14208 = ( n4874 & ~n7008 ) | ( n4874 & n9010 ) | ( ~n7008 & n9010 ) ;
  assign n14209 = n876 & n14208 ;
  assign n14210 = ~n3027 & n12853 ;
  assign n14211 = n5156 & n14210 ;
  assign n14212 = ~n545 & n14211 ;
  assign n14213 = n7658 ^ n5102 ^ 1'b0 ;
  assign n14214 = ~n9567 & n14213 ;
  assign n14215 = n14214 ^ n486 ^ x57 ;
  assign n14217 = n6120 | n6385 ;
  assign n14218 = n5931 ^ n1661 ^ 1'b0 ;
  assign n14219 = n14217 | n14218 ;
  assign n14216 = n11912 & ~n12796 ;
  assign n14220 = n14219 ^ n14216 ^ 1'b0 ;
  assign n14221 = n506 | n8183 ;
  assign n14222 = n618 | n6515 ;
  assign n14223 = n1094 & ~n14222 ;
  assign n14224 = n14223 ^ n6099 ^ 1'b0 ;
  assign n14225 = n14224 ^ n4319 ^ n490 ;
  assign n14226 = ( x102 & n6061 ) | ( x102 & ~n12145 ) | ( n6061 & ~n12145 ) ;
  assign n14227 = n8414 | n10982 ;
  assign n14228 = n437 & n5494 ;
  assign n14229 = n14228 ^ n3606 ^ 1'b0 ;
  assign n14230 = n14229 ^ x6 ^ 1'b0 ;
  assign n14231 = n2150 & ~n11765 ;
  assign n14232 = n2438 ^ n1922 ^ 1'b0 ;
  assign n14233 = n688 & n14232 ;
  assign n14235 = ~n3126 & n3755 ;
  assign n14236 = n14235 ^ n7525 ^ 1'b0 ;
  assign n14234 = n941 | n1353 ;
  assign n14237 = n14236 ^ n14234 ^ 1'b0 ;
  assign n14238 = n14233 & n14237 ;
  assign n14239 = n14231 & n14238 ;
  assign n14240 = ( n3435 & n8189 ) | ( n3435 & ~n8650 ) | ( n8189 & ~n8650 ) ;
  assign n14241 = ~n7376 & n9561 ;
  assign n14242 = ~n14240 & n14241 ;
  assign n14243 = n536 & n2805 ;
  assign n14244 = n2084 & ~n11162 ;
  assign n14245 = n4906 ^ n3203 ^ 1'b0 ;
  assign n14246 = n14244 & ~n14245 ;
  assign n14247 = ~n5348 & n14246 ;
  assign n14248 = n14243 & n14247 ;
  assign n14249 = n5063 ^ n4561 ^ 1'b0 ;
  assign n14250 = n6118 ^ n1621 ^ 1'b0 ;
  assign n14251 = ( n7800 & ~n11195 ) | ( n7800 & n14250 ) | ( ~n11195 & n14250 ) ;
  assign n14252 = n5834 ^ n3459 ^ 1'b0 ;
  assign n14253 = n3489 & n8988 ;
  assign n14254 = n2900 | n3861 ;
  assign n14255 = n3860 & n10507 ;
  assign n14256 = n14255 ^ n9623 ^ 1'b0 ;
  assign n14257 = ~n14254 & n14256 ;
  assign n14258 = n14257 ^ n11275 ^ 1'b0 ;
  assign n14262 = n5240 ^ n859 ^ 1'b0 ;
  assign n14263 = n7968 | n14262 ;
  assign n14259 = n2074 | n4600 ;
  assign n14260 = n2288 | n14259 ;
  assign n14261 = n9279 & n14260 ;
  assign n14264 = n14263 ^ n14261 ^ 1'b0 ;
  assign n14265 = n12976 ^ n5837 ^ 1'b0 ;
  assign n14266 = ~n6043 & n14265 ;
  assign n14267 = n12176 | n12812 ;
  assign n14268 = n4292 & ~n5822 ;
  assign n14269 = ~n6345 & n14268 ;
  assign n14270 = n6529 ^ n4712 ^ 1'b0 ;
  assign n14271 = ~n7730 & n14270 ;
  assign n14272 = n2642 | n14271 ;
  assign n14273 = n14269 & ~n14272 ;
  assign n14274 = n11730 | n14273 ;
  assign n14275 = n5885 | n14274 ;
  assign n14276 = n14267 & n14275 ;
  assign n14277 = n14276 ^ n10132 ^ 1'b0 ;
  assign n14278 = n7839 & ~n13627 ;
  assign n14279 = n14278 ^ n12669 ^ 1'b0 ;
  assign n14280 = n14279 ^ n4768 ^ 1'b0 ;
  assign n14281 = n14280 ^ n1619 ^ 1'b0 ;
  assign n14282 = x77 & ~n14281 ;
  assign n14283 = n3678 & n7350 ;
  assign n14284 = ~n4588 & n14283 ;
  assign n14285 = n3676 & ~n8280 ;
  assign n14286 = ~n13646 & n14285 ;
  assign n14287 = n6935 | n14286 ;
  assign n14288 = n11617 ^ n8677 ^ 1'b0 ;
  assign n14289 = n9190 & n14288 ;
  assign n14290 = n14228 ^ n6671 ^ n625 ;
  assign n14291 = ( ~n1033 & n10694 ) | ( ~n1033 & n14290 ) | ( n10694 & n14290 ) ;
  assign n14292 = ~n2987 & n13047 ;
  assign n14293 = n14292 ^ n12658 ^ 1'b0 ;
  assign n14294 = n2154 & n5207 ;
  assign n14295 = n14294 ^ n5352 ^ 1'b0 ;
  assign n14296 = n988 & n3245 ;
  assign n14297 = n6702 | n14296 ;
  assign n14298 = n3027 ^ n1118 ^ 1'b0 ;
  assign n14299 = n5804 ^ n5605 ^ n307 ;
  assign n14300 = ~n775 & n14299 ;
  assign n14301 = n14300 ^ n3276 ^ 1'b0 ;
  assign n14302 = n5471 ^ n4429 ^ n2667 ;
  assign n14303 = ( n1919 & ~n9279 ) | ( n1919 & n14302 ) | ( ~n9279 & n14302 ) ;
  assign n14304 = n6238 ^ n6099 ^ 1'b0 ;
  assign n14305 = n1531 | n14304 ;
  assign n14306 = n13539 ^ n3064 ^ 1'b0 ;
  assign n14307 = n8942 & ~n14306 ;
  assign n14308 = n14307 ^ n12168 ^ 1'b0 ;
  assign n14309 = n7019 & n7055 ;
  assign n14310 = n14309 ^ n7888 ^ 1'b0 ;
  assign n14311 = ~n2991 & n14310 ;
  assign n14312 = n5594 | n5781 ;
  assign n14313 = n900 & ~n14312 ;
  assign n14314 = n13463 ^ n11379 ^ 1'b0 ;
  assign n14315 = n7474 ^ n2892 ^ 1'b0 ;
  assign n14316 = ~n1079 & n14315 ;
  assign n14317 = n4610 & n14316 ;
  assign n14318 = n8134 ^ n2028 ^ 1'b0 ;
  assign n14319 = n1737 | n2044 ;
  assign n14320 = n2330 | n12463 ;
  assign n14321 = ( n2413 & n14319 ) | ( n2413 & ~n14320 ) | ( n14319 & ~n14320 ) ;
  assign n14322 = n8462 ^ n518 ^ 1'b0 ;
  assign n14323 = n1206 & ~n6644 ;
  assign n14324 = ~n1948 & n14323 ;
  assign n14325 = n4716 | n11435 ;
  assign n14326 = n14325 ^ n5547 ^ 1'b0 ;
  assign n14327 = n11554 ^ n2925 ^ 1'b0 ;
  assign n14328 = ( n1943 & ~n3182 ) | ( n1943 & n6359 ) | ( ~n3182 & n6359 ) ;
  assign n14329 = ~n4491 & n14328 ;
  assign n14331 = ~n1483 & n7980 ;
  assign n14332 = n288 & n3641 ;
  assign n14333 = ~n7984 & n14332 ;
  assign n14334 = n1024 | n14333 ;
  assign n14335 = n14334 ^ n5285 ^ 1'b0 ;
  assign n14336 = n14335 ^ n11188 ^ n540 ;
  assign n14337 = ( n10670 & n14331 ) | ( n10670 & ~n14336 ) | ( n14331 & ~n14336 ) ;
  assign n14330 = n10861 | n13452 ;
  assign n14338 = n14337 ^ n14330 ^ 1'b0 ;
  assign n14339 = n1500 ^ n967 ^ 1'b0 ;
  assign n14340 = n14339 ^ n3631 ^ n2718 ;
  assign n14341 = ~n1088 & n14340 ;
  assign n14342 = n12293 ^ n4019 ^ n1897 ;
  assign n14343 = n13857 & ~n14342 ;
  assign n14344 = n14343 ^ n4381 ^ 1'b0 ;
  assign n14345 = n9053 ^ n8277 ^ n6043 ;
  assign n14346 = ~n3481 & n9939 ;
  assign n14347 = n2676 & n4739 ;
  assign n14348 = ~n14346 & n14347 ;
  assign n14349 = n12793 ^ n3342 ^ 1'b0 ;
  assign n14350 = n11307 ^ n10222 ^ 1'b0 ;
  assign n14351 = n3597 & n14350 ;
  assign n14352 = n6708 & n14351 ;
  assign n14353 = ~n13819 & n14352 ;
  assign n14354 = ( x93 & n4655 ) | ( x93 & n14353 ) | ( n4655 & n14353 ) ;
  assign n14355 = ( n1703 & n6759 ) | ( n1703 & n10415 ) | ( n6759 & n10415 ) ;
  assign n14356 = n10463 ^ n166 ^ 1'b0 ;
  assign n14357 = ~n9365 & n14356 ;
  assign n14358 = n5645 & ~n14357 ;
  assign n14359 = n942 & n4774 ;
  assign n14360 = ( ~n5439 & n13806 ) | ( ~n5439 & n14359 ) | ( n13806 & n14359 ) ;
  assign n14361 = n11337 & n14360 ;
  assign n14362 = ~n4424 & n6187 ;
  assign n14363 = n14362 ^ n13099 ^ 1'b0 ;
  assign n14364 = n2363 ^ n774 ^ 1'b0 ;
  assign n14365 = n14363 | n14364 ;
  assign n14366 = n14365 ^ n10612 ^ 1'b0 ;
  assign n14368 = n2298 ^ n709 ^ 1'b0 ;
  assign n14369 = n1908 & n14368 ;
  assign n14367 = n2412 & ~n10015 ;
  assign n14370 = n14369 ^ n14367 ^ 1'b0 ;
  assign n14371 = n277 & n3438 ;
  assign n14372 = ( ~n933 & n4186 ) | ( ~n933 & n7592 ) | ( n4186 & n7592 ) ;
  assign n14373 = n5243 ^ n1433 ^ 1'b0 ;
  assign n14374 = n4652 & n14373 ;
  assign n14375 = n14372 & n14374 ;
  assign n14376 = n1363 & ~n14375 ;
  assign n14377 = ~n14371 & n14376 ;
  assign n14378 = ( n2342 & n3153 ) | ( n2342 & n3740 ) | ( n3153 & n3740 ) ;
  assign n14379 = ~n1719 & n14378 ;
  assign n14380 = n7466 ^ n4285 ^ 1'b0 ;
  assign n14381 = n6877 & n14380 ;
  assign n14382 = ( x6 & ~n4141 ) | ( x6 & n14381 ) | ( ~n4141 & n14381 ) ;
  assign n14383 = n1672 | n14382 ;
  assign n14384 = n8532 | n14383 ;
  assign n14385 = n8921 & n14384 ;
  assign n14386 = n6792 ^ n2622 ^ 1'b0 ;
  assign n14387 = n4785 | n14386 ;
  assign n14390 = ~n222 & n5077 ;
  assign n14388 = n6735 ^ n5351 ^ 1'b0 ;
  assign n14389 = n8617 & ~n14388 ;
  assign n14391 = n14390 ^ n14389 ^ n11945 ;
  assign n14392 = ~n14387 & n14391 ;
  assign n14394 = ( n476 & n491 ) | ( n476 & n5681 ) | ( n491 & n5681 ) ;
  assign n14393 = n2814 & n11933 ;
  assign n14395 = n14394 ^ n14393 ^ 1'b0 ;
  assign n14396 = n14395 ^ n10533 ^ 1'b0 ;
  assign n14397 = n12706 | n14396 ;
  assign n14398 = n5443 | n14397 ;
  assign n14399 = n240 & ~n732 ;
  assign n14400 = n5962 & n6323 ;
  assign n14401 = n8986 & n14400 ;
  assign n14402 = n4318 ^ n2307 ^ 1'b0 ;
  assign n14405 = n257 | n1188 ;
  assign n14403 = n5522 ^ n4348 ^ 1'b0 ;
  assign n14404 = n11710 | n14403 ;
  assign n14406 = n14405 ^ n14404 ^ 1'b0 ;
  assign n14407 = n9452 ^ n5865 ^ 1'b0 ;
  assign n14408 = n3192 & ~n14407 ;
  assign n14409 = n2211 ^ n1691 ^ 1'b0 ;
  assign n14410 = n14409 ^ n13982 ^ n13472 ;
  assign n14412 = n7519 ^ n1189 ^ 1'b0 ;
  assign n14413 = ~n1383 & n14412 ;
  assign n14411 = n1586 | n5610 ;
  assign n14414 = n14413 ^ n14411 ^ 1'b0 ;
  assign n14415 = n14414 ^ n6299 ^ 1'b0 ;
  assign n14416 = n551 | n14415 ;
  assign n14417 = x72 & n3015 ;
  assign n14418 = ~n12903 & n14417 ;
  assign n14419 = ( n905 & n5816 ) | ( n905 & ~n14418 ) | ( n5816 & ~n14418 ) ;
  assign n14420 = n2976 & n14419 ;
  assign n14421 = n9448 | n14420 ;
  assign n14422 = n3010 | n6426 ;
  assign n14423 = n3010 & ~n14422 ;
  assign n14424 = n14423 ^ n7856 ^ 1'b0 ;
  assign n14425 = n9964 & ~n14424 ;
  assign n14427 = n2113 & n6384 ;
  assign n14428 = n14427 ^ n6864 ^ 1'b0 ;
  assign n14426 = n620 & ~n3120 ;
  assign n14429 = n14428 ^ n14426 ^ 1'b0 ;
  assign n14430 = n13806 ^ n6448 ^ 1'b0 ;
  assign n14431 = n5937 & ~n6972 ;
  assign n14432 = n14431 ^ n13950 ^ 1'b0 ;
  assign n14433 = n5832 ^ n5195 ^ 1'b0 ;
  assign n14434 = n7368 & n14433 ;
  assign n14435 = n14434 ^ n9445 ^ 1'b0 ;
  assign n14436 = n14208 & n14435 ;
  assign n14437 = ~n9039 & n9199 ;
  assign n14438 = n3041 & n14437 ;
  assign n14440 = ~n2579 & n3386 ;
  assign n14441 = n14440 ^ n6549 ^ 1'b0 ;
  assign n14442 = n4318 & n14441 ;
  assign n14439 = n2288 & n4244 ;
  assign n14443 = n14442 ^ n14439 ^ 1'b0 ;
  assign n14444 = n4257 | n12400 ;
  assign n14445 = n2794 | n14444 ;
  assign n14446 = n645 & n799 ;
  assign n14447 = n8736 & ~n10694 ;
  assign n14448 = ~n13437 & n14447 ;
  assign n14449 = n13231 & ~n14448 ;
  assign n14450 = ~n14446 & n14449 ;
  assign n14451 = n5737 & ~n14450 ;
  assign n14452 = ~n14445 & n14451 ;
  assign n14453 = n7221 ^ n6565 ^ 1'b0 ;
  assign n14454 = ( n4167 & n6461 ) | ( n4167 & ~n7426 ) | ( n6461 & ~n7426 ) ;
  assign n14459 = n5323 & n11329 ;
  assign n14460 = ~n7712 & n14459 ;
  assign n14455 = n3641 & n13109 ;
  assign n14456 = n7396 ^ n6631 ^ 1'b0 ;
  assign n14457 = n8063 & ~n14456 ;
  assign n14458 = n14455 & ~n14457 ;
  assign n14461 = n14460 ^ n14458 ^ 1'b0 ;
  assign n14462 = n5042 ^ n4549 ^ 1'b0 ;
  assign n14463 = n1737 & n14462 ;
  assign n14464 = n3687 ^ n2650 ^ n630 ;
  assign n14465 = n7001 | n14464 ;
  assign n14466 = n6458 & ~n6549 ;
  assign n14467 = ~n10284 & n14466 ;
  assign n14468 = ~n9856 & n10354 ;
  assign n14469 = n6258 ^ n5820 ^ n672 ;
  assign n14470 = n13223 & ~n14469 ;
  assign n14471 = n6613 ^ n324 ^ 1'b0 ;
  assign n14472 = ~n208 & n5836 ;
  assign n14473 = n6333 ^ n308 ^ 1'b0 ;
  assign n14474 = n3289 | n11632 ;
  assign n14475 = n8650 & ~n14474 ;
  assign n14476 = n3824 | n14475 ;
  assign n14477 = n14476 ^ n8074 ^ 1'b0 ;
  assign n14478 = n10755 ^ n2036 ^ 1'b0 ;
  assign n14479 = n3629 & n14478 ;
  assign n14480 = n6479 & ~n13443 ;
  assign n14481 = n14479 | n14480 ;
  assign n14482 = n7802 & ~n10158 ;
  assign n14483 = n13491 ^ n3832 ^ 1'b0 ;
  assign n14484 = ~n2837 & n5069 ;
  assign n14485 = n14484 ^ n3324 ^ 1'b0 ;
  assign n14486 = n2756 & n13817 ;
  assign n14487 = ~n4612 & n5345 ;
  assign n14488 = n6109 ^ n3326 ^ 1'b0 ;
  assign n14489 = ~n2137 & n14488 ;
  assign n14490 = n6930 & n14489 ;
  assign n14491 = n14490 ^ n327 ^ 1'b0 ;
  assign n14492 = n3883 | n14491 ;
  assign n14494 = n2397 ^ n2354 ^ 1'b0 ;
  assign n14495 = n5613 & n14494 ;
  assign n14496 = n2686 & n14495 ;
  assign n14497 = ~n4440 & n14496 ;
  assign n14493 = n9376 ^ n7185 ^ 1'b0 ;
  assign n14498 = n14497 ^ n14493 ^ 1'b0 ;
  assign n14499 = n2673 & n14498 ;
  assign n14500 = n1888 & n3294 ;
  assign n14501 = ~n652 & n14500 ;
  assign n14502 = n5886 ^ n1309 ^ 1'b0 ;
  assign n14503 = ~n14501 & n14502 ;
  assign n14504 = n11912 & ~n14503 ;
  assign n14505 = ~n369 & n1128 ;
  assign n14506 = n8431 & ~n14505 ;
  assign n14507 = n9537 & n14506 ;
  assign n14508 = n2395 & ~n14507 ;
  assign n14509 = n13098 ^ n353 ^ 1'b0 ;
  assign n14510 = n2712 & ~n14509 ;
  assign n14511 = ~n6449 & n14510 ;
  assign n14512 = n5573 ^ x103 ^ 1'b0 ;
  assign n14513 = n14512 ^ n8987 ^ n8938 ;
  assign n14514 = ( n1586 & ~n3518 ) | ( n1586 & n10190 ) | ( ~n3518 & n10190 ) ;
  assign n14515 = ~n1937 & n14514 ;
  assign n14516 = n14515 ^ n3343 ^ 1'b0 ;
  assign n14517 = ( n1531 & n3367 ) | ( n1531 & n7201 ) | ( n3367 & n7201 ) ;
  assign n14518 = ~n351 & n797 ;
  assign n14519 = n4778 & ~n11404 ;
  assign n14520 = n14519 ^ n9265 ^ 1'b0 ;
  assign n14521 = n667 & ~n14520 ;
  assign n14522 = ~n14518 & n14521 ;
  assign n14523 = ~n339 & n556 ;
  assign n14524 = n4682 ^ n1790 ^ n852 ;
  assign n14526 = x33 & ~n6439 ;
  assign n14525 = n7727 & n10935 ;
  assign n14527 = n14526 ^ n14525 ^ 1'b0 ;
  assign n14529 = n1801 & ~n2470 ;
  assign n14530 = n14529 ^ n13958 ^ 1'b0 ;
  assign n14531 = n2330 ^ n1295 ^ 1'b0 ;
  assign n14532 = n14530 & ~n14531 ;
  assign n14528 = ~n11437 & n12898 ;
  assign n14533 = n14532 ^ n14528 ^ 1'b0 ;
  assign n14534 = n3906 ^ n2477 ^ n323 ;
  assign n14535 = n14534 ^ n14019 ^ 1'b0 ;
  assign n14536 = n10573 | n14535 ;
  assign n14537 = n1981 & ~n3104 ;
  assign n14538 = n14537 ^ n1230 ^ 1'b0 ;
  assign n14539 = n13032 & ~n14538 ;
  assign n14540 = n533 & n14539 ;
  assign n14541 = n11630 | n14540 ;
  assign n14542 = n3334 & ~n8580 ;
  assign n14543 = n14542 ^ n156 ^ 1'b0 ;
  assign n14544 = ~n1380 & n3278 ;
  assign n14545 = n14544 ^ n3306 ^ 1'b0 ;
  assign n14546 = n7126 | n14545 ;
  assign n14547 = n5245 & ~n14546 ;
  assign n14548 = n471 | n2370 ;
  assign n14549 = n14548 ^ n2293 ^ 1'b0 ;
  assign n14550 = ( ~n4057 & n12059 ) | ( ~n4057 & n14549 ) | ( n12059 & n14549 ) ;
  assign n14551 = n4895 ^ n154 ^ 1'b0 ;
  assign n14552 = ~n13982 & n14551 ;
  assign n14553 = n14552 ^ n1496 ^ 1'b0 ;
  assign n14554 = n1920 & n10087 ;
  assign n14555 = n8268 ^ n3626 ^ 1'b0 ;
  assign n14556 = n9856 | n14555 ;
  assign n14557 = n10615 ^ n2667 ^ 1'b0 ;
  assign n14558 = n4797 ^ n3753 ^ 1'b0 ;
  assign n14559 = n14557 & ~n14558 ;
  assign n14560 = n3755 ^ n1097 ^ 1'b0 ;
  assign n14561 = n10216 ^ n4007 ^ 1'b0 ;
  assign n14562 = n11267 & n14561 ;
  assign n14563 = n14562 ^ n4505 ^ 1'b0 ;
  assign n14564 = n14563 ^ n7185 ^ 1'b0 ;
  assign n14565 = n6596 | n14564 ;
  assign n14566 = n3697 & ~n3789 ;
  assign n14567 = n14565 & n14566 ;
  assign n14568 = ( ~n3869 & n10017 ) | ( ~n3869 & n12030 ) | ( n10017 & n12030 ) ;
  assign n14569 = n3576 | n8158 ;
  assign n14570 = n2242 & ~n14569 ;
  assign n14571 = n2969 & ~n3167 ;
  assign n14572 = ~n11261 & n14571 ;
  assign n14576 = ( n1432 & ~n2086 ) | ( n1432 & n7029 ) | ( ~n2086 & n7029 ) ;
  assign n14574 = n1303 & ~n1390 ;
  assign n14575 = n14270 & n14574 ;
  assign n14573 = n2252 ^ n1854 ^ 1'b0 ;
  assign n14577 = n14576 ^ n14575 ^ n14573 ;
  assign n14578 = n3212 & ~n14577 ;
  assign n14579 = n14578 ^ n4793 ^ 1'b0 ;
  assign n14580 = n8323 ^ n3366 ^ x100 ;
  assign n14581 = n559 & ~n3498 ;
  assign n14582 = ~n10547 & n14581 ;
  assign n14584 = n3960 ^ x69 ^ 1'b0 ;
  assign n14585 = n2778 & n14584 ;
  assign n14586 = n517 | n14585 ;
  assign n14587 = ~n9852 & n14586 ;
  assign n14583 = n1450 & n12195 ;
  assign n14588 = n14587 ^ n14583 ^ 1'b0 ;
  assign n14589 = n1206 & ~n3401 ;
  assign n14590 = n1015 ^ x57 ^ 1'b0 ;
  assign n14591 = n14589 | n14590 ;
  assign n14592 = n14591 ^ n3237 ^ n695 ;
  assign n14593 = n1487 & ~n14592 ;
  assign n14594 = ~n1344 & n14593 ;
  assign n14595 = ~n3248 & n4840 ;
  assign n14596 = n5226 & n14595 ;
  assign n14597 = n1850 | n14596 ;
  assign n14598 = n4266 & ~n6940 ;
  assign n14599 = n8797 & n14598 ;
  assign n14600 = ( ~n10619 & n14597 ) | ( ~n10619 & n14599 ) | ( n14597 & n14599 ) ;
  assign n14601 = ~n3082 & n10099 ;
  assign n14606 = ~n9473 & n11431 ;
  assign n14607 = n14606 ^ n9439 ^ 1'b0 ;
  assign n14608 = ( n6263 & n9692 ) | ( n6263 & n14607 ) | ( n9692 & n14607 ) ;
  assign n14603 = n1897 & n2031 ;
  assign n14602 = n6813 & ~n7953 ;
  assign n14604 = n14603 ^ n14602 ^ 1'b0 ;
  assign n14605 = n6731 & ~n14604 ;
  assign n14609 = n14608 ^ n14605 ^ 1'b0 ;
  assign n14613 = n180 | n1635 ;
  assign n14614 = n147 | n14613 ;
  assign n14610 = n2481 & ~n3935 ;
  assign n14611 = n8911 | n14610 ;
  assign n14612 = n3093 & ~n14611 ;
  assign n14615 = n14614 ^ n14612 ^ n4940 ;
  assign n14616 = n11512 ^ n224 ^ 1'b0 ;
  assign n14617 = n8165 & n14616 ;
  assign n14622 = n8262 ^ n7467 ^ n5894 ;
  assign n14618 = n6035 & n6340 ;
  assign n14619 = n14618 ^ n7328 ^ 1'b0 ;
  assign n14620 = n3116 | n14619 ;
  assign n14621 = n14620 ^ n2213 ^ 1'b0 ;
  assign n14623 = n14622 ^ n14621 ^ 1'b0 ;
  assign n14624 = n12009 ^ n10455 ^ 1'b0 ;
  assign n14625 = n3863 & ~n14624 ;
  assign n14626 = n14625 ^ n3825 ^ 1'b0 ;
  assign n14627 = n8249 & n14626 ;
  assign n14628 = n459 & ~n12602 ;
  assign n14629 = n14628 ^ n1899 ^ 1'b0 ;
  assign n14630 = ~n3365 & n5492 ;
  assign n14631 = ~n1929 & n11527 ;
  assign n14632 = n6497 & n14631 ;
  assign n14633 = n8910 ^ n1277 ^ n1103 ;
  assign n14634 = n805 ^ n294 ^ 1'b0 ;
  assign n14635 = n11120 | n14634 ;
  assign n14636 = n14635 ^ x72 ^ 1'b0 ;
  assign n14637 = n4085 & ~n10772 ;
  assign n14638 = n6625 & n11107 ;
  assign n14639 = n3784 & n14638 ;
  assign n14640 = n3981 ^ n732 ^ 1'b0 ;
  assign n14641 = n1676 & ~n14640 ;
  assign n14642 = n14641 ^ n2783 ^ 1'b0 ;
  assign n14643 = n4319 & n11877 ;
  assign n14644 = n14643 ^ n4655 ^ 1'b0 ;
  assign n14645 = n3166 | n14644 ;
  assign n14646 = n12627 ^ n1145 ^ 1'b0 ;
  assign n14647 = ~n13919 & n14646 ;
  assign n14648 = ~n8365 & n10784 ;
  assign n14649 = n14648 ^ n6268 ^ 1'b0 ;
  assign n14650 = n10656 ^ n8181 ^ 1'b0 ;
  assign n14654 = ( n3099 & n5102 ) | ( n3099 & n6661 ) | ( n5102 & n6661 ) ;
  assign n14651 = n1329 ^ n586 ^ 1'b0 ;
  assign n14652 = n2170 & ~n14651 ;
  assign n14653 = ~n6348 & n14652 ;
  assign n14655 = n14654 ^ n14653 ^ 1'b0 ;
  assign n14656 = x90 & n1920 ;
  assign n14657 = ~n588 & n14656 ;
  assign n14658 = ~n14655 & n14657 ;
  assign n14661 = n3787 ^ n2699 ^ 1'b0 ;
  assign n14659 = n4430 & ~n6909 ;
  assign n14660 = n11380 & n14659 ;
  assign n14662 = n14661 ^ n14660 ^ n14363 ;
  assign n14663 = n2905 & ~n3869 ;
  assign n14664 = n551 & n14663 ;
  assign n14665 = n14664 ^ n8610 ^ 1'b0 ;
  assign n14666 = n3110 & n6166 ;
  assign n14667 = ~n5935 & n14666 ;
  assign n14668 = ~n3635 & n4775 ;
  assign n14669 = n2827 & n14668 ;
  assign n14670 = n1391 & n12008 ;
  assign n14671 = n6488 & n9060 ;
  assign n14672 = n14671 ^ n1483 ^ 1'b0 ;
  assign n14673 = ( n2998 & ~n3169 ) | ( n2998 & n7093 ) | ( ~n3169 & n7093 ) ;
  assign n14674 = ~x60 & n14673 ;
  assign n14675 = n2158 & ~n14674 ;
  assign n14676 = n1569 & n14675 ;
  assign n14677 = n14676 ^ n10091 ^ 1'b0 ;
  assign n14678 = n9071 & n10154 ;
  assign n14679 = n6628 ^ n1511 ^ 1'b0 ;
  assign n14680 = n10748 ^ n9758 ^ 1'b0 ;
  assign n14681 = n14680 ^ n6148 ^ 1'b0 ;
  assign n14682 = n5002 | n14681 ;
  assign n14683 = n2395 | n3118 ;
  assign n14684 = n468 | n5709 ;
  assign n14685 = n14684 ^ n2285 ^ 1'b0 ;
  assign n14686 = n11562 ^ n2131 ^ 1'b0 ;
  assign n14687 = n14685 & ~n14686 ;
  assign n14688 = n6557 ^ n1152 ^ 1'b0 ;
  assign n14689 = n1597 ^ n335 ^ 1'b0 ;
  assign n14690 = ~n12677 & n14689 ;
  assign n14691 = n14688 & n14690 ;
  assign n14692 = n5297 & ~n11552 ;
  assign n14694 = n6730 ^ n5492 ^ 1'b0 ;
  assign n14693 = n338 & ~n9382 ;
  assign n14695 = n14694 ^ n14693 ^ 1'b0 ;
  assign n14696 = n11018 & ~n12879 ;
  assign n14697 = n1899 & ~n14696 ;
  assign n14698 = n7422 & n14697 ;
  assign n14699 = n7048 ^ n2677 ^ 1'b0 ;
  assign n14700 = n7689 | n12269 ;
  assign n14701 = n14700 ^ n6259 ^ 1'b0 ;
  assign n14702 = n8800 & n10144 ;
  assign n14703 = n5092 ^ n738 ^ 1'b0 ;
  assign n14704 = n4922 & ~n14703 ;
  assign n14705 = ~n4769 & n12266 ;
  assign n14706 = ~n12823 & n14705 ;
  assign n14707 = n9803 ^ n7493 ^ 1'b0 ;
  assign n14708 = n172 & n14707 ;
  assign n14709 = n14708 ^ n4149 ^ 1'b0 ;
  assign n14710 = ~n5537 & n14709 ;
  assign n14711 = ~n4843 & n14710 ;
  assign n14712 = ~n4030 & n5942 ;
  assign n14713 = n14712 ^ n2561 ^ 1'b0 ;
  assign n14714 = n10640 & ~n14713 ;
  assign n14715 = n7569 ^ n6794 ^ 1'b0 ;
  assign n14716 = n5568 & n14715 ;
  assign n14717 = n10936 ^ n10453 ^ 1'b0 ;
  assign n14718 = ~n745 & n3048 ;
  assign n14719 = n6542 & n14718 ;
  assign n14720 = n5737 & n8273 ;
  assign n14721 = n5331 & n12790 ;
  assign n14722 = n14721 ^ n1411 ^ 1'b0 ;
  assign n14723 = n1880 & ~n8399 ;
  assign n14724 = n14723 ^ n5371 ^ 1'b0 ;
  assign n14725 = n9982 ^ n3630 ^ 1'b0 ;
  assign n14726 = n12839 & ~n14725 ;
  assign n14727 = n14726 ^ n486 ^ 1'b0 ;
  assign n14728 = n1103 & n14727 ;
  assign n14729 = n6532 & n14728 ;
  assign n14730 = n5408 ^ n1338 ^ 1'b0 ;
  assign n14731 = n14730 ^ n6928 ^ 1'b0 ;
  assign n14732 = n12759 ^ n7388 ^ 1'b0 ;
  assign n14733 = n3225 | n9784 ;
  assign n14734 = n14732 | n14733 ;
  assign n14735 = ~n2044 & n2758 ;
  assign n14736 = n14735 ^ n7258 ^ 1'b0 ;
  assign n14737 = n8800 | n14736 ;
  assign n14738 = n9132 ^ n1526 ^ 1'b0 ;
  assign n14739 = n14737 | n14738 ;
  assign n14740 = n4558 | n6950 ;
  assign n14741 = n11030 & ~n14740 ;
  assign n14742 = x78 & ~n6399 ;
  assign n14743 = n5458 & n14742 ;
  assign n14744 = ~n5458 & n14743 ;
  assign n14745 = x86 & ~n542 ;
  assign n14746 = ~x86 & n14745 ;
  assign n14747 = n14746 ^ n3727 ^ 1'b0 ;
  assign n14748 = x71 & x97 ;
  assign n14749 = ~x71 & n14748 ;
  assign n14750 = ~n937 & n7347 ;
  assign n14751 = n14749 & n14750 ;
  assign n14752 = n3300 & ~n14751 ;
  assign n14753 = n14747 & n14752 ;
  assign n14754 = n14744 & n14753 ;
  assign n14755 = n5197 & n12903 ;
  assign n14756 = ~n12903 & n14755 ;
  assign n14757 = n7928 | n14756 ;
  assign n14758 = n14754 & ~n14757 ;
  assign n14759 = n6074 & ~n9514 ;
  assign n14760 = ~n10602 & n14759 ;
  assign n14761 = n9508 | n12586 ;
  assign n14762 = n4408 & ~n10578 ;
  assign n14763 = n9176 ^ n5120 ^ n2428 ;
  assign n14764 = n14763 ^ n6177 ^ n2823 ;
  assign n14765 = ~n9994 & n14585 ;
  assign n14766 = ~n1119 & n14765 ;
  assign n14767 = n2635 | n14766 ;
  assign n14768 = n14767 ^ n11990 ^ n139 ;
  assign n14769 = n1578 | n8314 ;
  assign n14770 = n5811 ^ n2607 ^ 1'b0 ;
  assign n14771 = n14769 & ~n14770 ;
  assign n14772 = n14771 ^ n3873 ^ 1'b0 ;
  assign n14773 = n5357 ^ n3730 ^ 1'b0 ;
  assign n14774 = n1898 | n14773 ;
  assign n14775 = n4428 & n6991 ;
  assign n14776 = n14775 ^ n13008 ^ 1'b0 ;
  assign n14777 = n2965 ^ n875 ^ 1'b0 ;
  assign n14778 = n14777 ^ n10726 ^ 1'b0 ;
  assign n14779 = n2353 | n11298 ;
  assign n14780 = n14778 & ~n14779 ;
  assign n14781 = n376 & ~n935 ;
  assign n14782 = n868 & n14781 ;
  assign n14783 = n3540 & ~n4527 ;
  assign n14784 = n14783 ^ n11391 ^ 1'b0 ;
  assign n14785 = n6279 & n14784 ;
  assign n14786 = n7886 | n14785 ;
  assign n14787 = n11351 ^ n1140 ^ 1'b0 ;
  assign n14788 = n4115 | n12902 ;
  assign n14789 = n4973 | n14788 ;
  assign n14790 = n5727 & n7198 ;
  assign n14791 = n14790 ^ n1664 ^ n1342 ;
  assign n14792 = n266 | n14791 ;
  assign n14793 = n5350 & ~n8126 ;
  assign n14794 = ~n1337 & n14793 ;
  assign n14795 = n234 | n9121 ;
  assign n14796 = n9320 & n14795 ;
  assign n14797 = n14796 ^ n4315 ^ 1'b0 ;
  assign n14798 = n14797 ^ n4197 ^ 1'b0 ;
  assign n14799 = ~n14794 & n14798 ;
  assign n14800 = n12315 ^ n954 ^ x19 ;
  assign n14801 = n7753 ^ n1939 ^ 1'b0 ;
  assign n14802 = x70 & n10416 ;
  assign n14803 = ~n3933 & n14802 ;
  assign n14804 = n7879 | n14803 ;
  assign n14805 = n14801 & ~n14804 ;
  assign n14812 = n3179 & n9504 ;
  assign n14813 = ~n5544 & n14812 ;
  assign n14807 = x105 & n4895 ;
  assign n14808 = n14807 ^ n2810 ^ 1'b0 ;
  assign n14809 = ~n7130 & n14808 ;
  assign n14810 = ~n14428 & n14809 ;
  assign n14806 = ~n2470 & n14357 ;
  assign n14811 = n14810 ^ n14806 ^ 1'b0 ;
  assign n14814 = n14813 ^ n14811 ^ n9165 ;
  assign n14815 = n2948 ^ n2632 ^ 1'b0 ;
  assign n14816 = n8803 | n14815 ;
  assign n14817 = ~n1925 & n13459 ;
  assign n14818 = n14817 ^ n10507 ^ 1'b0 ;
  assign n14819 = n5437 | n9714 ;
  assign n14820 = n14819 ^ n5999 ^ n5951 ;
  assign n14821 = n7543 & n14820 ;
  assign n14822 = n2987 | n10146 ;
  assign n14823 = n14604 & ~n14822 ;
  assign n14824 = ( n1552 & ~n5852 ) | ( n1552 & n5973 ) | ( ~n5852 & n5973 ) ;
  assign n14825 = ( ~n6423 & n6655 ) | ( ~n6423 & n14824 ) | ( n6655 & n14824 ) ;
  assign n14826 = n9431 | n14825 ;
  assign n14827 = n14826 ^ n6770 ^ 1'b0 ;
  assign n14828 = n14827 ^ n1842 ^ 1'b0 ;
  assign n14829 = n6790 | n11768 ;
  assign n14830 = n3295 | n7371 ;
  assign n14831 = n14830 ^ n3866 ^ 1'b0 ;
  assign n14832 = ( n1646 & n3284 ) | ( n1646 & n14831 ) | ( n3284 & n14831 ) ;
  assign n14833 = n2961 & n6043 ;
  assign n14834 = n14833 ^ n2844 ^ 1'b0 ;
  assign n14835 = n14832 & ~n14834 ;
  assign n14836 = n14835 ^ n3140 ^ 1'b0 ;
  assign n14837 = n12091 & n14836 ;
  assign n14838 = n1880 & ~n4602 ;
  assign n14841 = ( n478 & ~n1854 ) | ( n478 & n5289 ) | ( ~n1854 & n5289 ) ;
  assign n14839 = ~n6064 & n7049 ;
  assign n14840 = ~n10679 & n14839 ;
  assign n14842 = n14841 ^ n14840 ^ 1'b0 ;
  assign n14843 = n14838 & ~n14842 ;
  assign n14844 = n7568 ^ n6158 ^ n3714 ;
  assign n14845 = n995 | n14844 ;
  assign n14846 = n3112 & n14845 ;
  assign n14847 = n14846 ^ n6132 ^ n3380 ;
  assign n14848 = n14847 ^ n4027 ^ 1'b0 ;
  assign n14849 = n6486 ^ n1817 ^ 1'b0 ;
  assign n14850 = n971 | n14849 ;
  assign n14851 = n3106 | n14850 ;
  assign n14852 = n14851 ^ n9610 ^ 1'b0 ;
  assign n14853 = n11867 ^ n10253 ^ 1'b0 ;
  assign n14854 = n13326 ^ n574 ^ 1'b0 ;
  assign n14855 = n7646 ^ n855 ^ 1'b0 ;
  assign n14856 = n971 | n14855 ;
  assign n14857 = n14856 ^ n11632 ^ 1'b0 ;
  assign n14858 = ~n14854 & n14857 ;
  assign n14859 = n9962 ^ n3935 ^ 1'b0 ;
  assign n14860 = n2673 & n3672 ;
  assign n14861 = n2884 & n14860 ;
  assign n14862 = n2564 ^ n1939 ^ 1'b0 ;
  assign n14863 = n14861 | n14862 ;
  assign n14864 = n1394 ^ n428 ^ 1'b0 ;
  assign n14865 = ~n1083 & n14864 ;
  assign n14866 = ~n4527 & n14865 ;
  assign n14867 = n2246 & n14866 ;
  assign n14868 = n487 & n3227 ;
  assign n14869 = n14868 ^ n7291 ^ 1'b0 ;
  assign n14870 = n14869 ^ n2723 ^ 1'b0 ;
  assign n14871 = n14870 ^ n5254 ^ 1'b0 ;
  assign n14872 = ~n9653 & n14871 ;
  assign n14873 = ~n1015 & n14872 ;
  assign n14874 = n14867 & n14873 ;
  assign n14875 = n4323 | n14874 ;
  assign n14877 = n517 ^ x21 ^ 1'b0 ;
  assign n14878 = n3403 | n14877 ;
  assign n14876 = n12066 & n14048 ;
  assign n14879 = n14878 ^ n14876 ^ 1'b0 ;
  assign n14880 = n840 | n1031 ;
  assign n14881 = n9473 ^ n5451 ^ 1'b0 ;
  assign n14882 = n3839 & n14881 ;
  assign n14883 = ( n1714 & ~n3272 ) | ( n1714 & n8601 ) | ( ~n3272 & n8601 ) ;
  assign n14884 = ~n1970 & n14883 ;
  assign n14885 = n14884 ^ n3179 ^ n1350 ;
  assign n14886 = ( n3618 & n4379 ) | ( n3618 & n14885 ) | ( n4379 & n14885 ) ;
  assign n14887 = n6802 | n11663 ;
  assign n14888 = n8584 | n11228 ;
  assign n14889 = n14888 ^ n4293 ^ 1'b0 ;
  assign n14890 = ~n9121 & n11191 ;
  assign n14891 = n14890 ^ n4119 ^ 1'b0 ;
  assign n14892 = n9469 ^ n2821 ^ 1'b0 ;
  assign n14893 = n14892 ^ n202 ^ 1'b0 ;
  assign n14894 = n4856 & ~n14893 ;
  assign n14895 = ~n9136 & n14460 ;
  assign n14896 = n458 & n3665 ;
  assign n14897 = n3614 ^ n3548 ^ 1'b0 ;
  assign n14898 = ~n3968 & n14897 ;
  assign n14900 = n2637 | n11882 ;
  assign n14901 = n2211 & ~n14900 ;
  assign n14899 = ~n755 & n1536 ;
  assign n14902 = n14901 ^ n14899 ^ 1'b0 ;
  assign n14903 = ~n9203 & n12297 ;
  assign n14904 = n2886 ^ n651 ^ 1'b0 ;
  assign n14905 = n14903 & ~n14904 ;
  assign n14906 = n12654 ^ n9928 ^ n3599 ;
  assign n14907 = n2425 & ~n9876 ;
  assign n14908 = n14907 ^ n12626 ^ 1'b0 ;
  assign n14909 = n14321 & ~n14908 ;
  assign n14910 = ~n14906 & n14909 ;
  assign n14912 = ~n5018 & n9327 ;
  assign n14913 = n14912 ^ n1155 ^ 1'b0 ;
  assign n14911 = n6549 | n6584 ;
  assign n14914 = n14913 ^ n14911 ^ 1'b0 ;
  assign n14915 = n2942 ^ n1221 ^ 1'b0 ;
  assign n14916 = n14914 | n14915 ;
  assign n14917 = n9319 ^ n3874 ^ 1'b0 ;
  assign n14918 = n14917 ^ n677 ^ 1'b0 ;
  assign n14919 = n336 & ~n8406 ;
  assign n14920 = n14919 ^ n2394 ^ 1'b0 ;
  assign n14921 = n14920 ^ n9961 ^ 1'b0 ;
  assign n14922 = n6315 & n14921 ;
  assign n14923 = n1093 | n7030 ;
  assign n14924 = n14923 ^ n11320 ^ 1'b0 ;
  assign n14925 = n4540 ^ n1578 ^ 1'b0 ;
  assign n14926 = n7713 & ~n14925 ;
  assign n14927 = n14926 ^ n6494 ^ 1'b0 ;
  assign n14928 = ~n907 & n4902 ;
  assign n14929 = n1197 & n14928 ;
  assign n14930 = n5468 | n11391 ;
  assign n14931 = n14930 ^ n6394 ^ 1'b0 ;
  assign n14932 = n14931 ^ n12856 ^ 1'b0 ;
  assign n14933 = n7806 ^ n7519 ^ 1'b0 ;
  assign n14934 = ~n9101 & n14933 ;
  assign n14935 = ( ~n141 & n7343 ) | ( ~n141 & n14934 ) | ( n7343 & n14934 ) ;
  assign n14936 = n11783 ^ n10344 ^ 1'b0 ;
  assign n14941 = n2412 & ~n11225 ;
  assign n14937 = ~n5493 & n11807 ;
  assign n14938 = n3781 ^ n3369 ^ 1'b0 ;
  assign n14939 = ~n2579 & n14938 ;
  assign n14940 = ~n14937 & n14939 ;
  assign n14942 = n14941 ^ n14940 ^ 1'b0 ;
  assign n14943 = n8760 | n10033 ;
  assign n14944 = n14943 ^ n7393 ^ 1'b0 ;
  assign n14945 = ( n2442 & ~n9621 ) | ( n2442 & n14944 ) | ( ~n9621 & n14944 ) ;
  assign n14946 = n5906 ^ n892 ^ 1'b0 ;
  assign n14947 = n12271 ^ n2364 ^ 1'b0 ;
  assign n14948 = n692 | n14947 ;
  assign n14949 = n4616 ^ n973 ^ 1'b0 ;
  assign n14950 = ~n13268 & n14949 ;
  assign n14951 = n7878 ^ n404 ^ 1'b0 ;
  assign n14952 = ~n12561 & n14951 ;
  assign n14953 = n14952 ^ n11040 ^ n4647 ;
  assign n14954 = n9894 ^ n2336 ^ 1'b0 ;
  assign n14955 = n699 ^ n250 ^ 1'b0 ;
  assign n14956 = ~n3143 & n14955 ;
  assign n14957 = n5855 ^ n3960 ^ 1'b0 ;
  assign n14958 = n14956 & ~n14957 ;
  assign n14959 = n14958 ^ n3603 ^ 1'b0 ;
  assign n14960 = ~n1992 & n5993 ;
  assign n14961 = n7574 & n14960 ;
  assign n14962 = n3405 | n9802 ;
  assign n14963 = n14962 ^ n630 ^ 1'b0 ;
  assign n14964 = n941 | n1402 ;
  assign n14965 = n14964 ^ n435 ^ 1'b0 ;
  assign n14966 = n989 & n5755 ;
  assign n14967 = n5264 | n7345 ;
  assign n14968 = n9690 ^ n4224 ^ 1'b0 ;
  assign n14969 = n308 & ~n3339 ;
  assign n14970 = n14969 ^ n309 ^ 1'b0 ;
  assign n14971 = n14968 | n14970 ;
  assign n14972 = ~n3708 & n14048 ;
  assign n14973 = n14972 ^ n10558 ^ 1'b0 ;
  assign n14974 = n675 & n10700 ;
  assign n14975 = ~n9899 & n14974 ;
  assign n14976 = n6110 & ~n8710 ;
  assign n14977 = n6359 & n14976 ;
  assign n14978 = n2250 & ~n3874 ;
  assign n14979 = n2330 | n7860 ;
  assign n14980 = n14979 ^ n10271 ^ 1'b0 ;
  assign n14981 = n14980 ^ n13602 ^ n4531 ;
  assign n14982 = ~n4748 & n5819 ;
  assign n14983 = n139 & ~n5678 ;
  assign n14984 = ~n5290 & n14983 ;
  assign n14985 = n14984 ^ n6025 ^ 1'b0 ;
  assign n14986 = n14985 ^ n4639 ^ 1'b0 ;
  assign n14987 = ~n8770 & n14986 ;
  assign n14988 = n8550 & n14987 ;
  assign n14989 = ~n4193 & n14293 ;
  assign n14990 = n14989 ^ n14395 ^ 1'b0 ;
  assign n14991 = n5647 ^ n3869 ^ 1'b0 ;
  assign n14992 = n14991 ^ n3727 ^ 1'b0 ;
  assign n14993 = n12957 ^ n6919 ^ 1'b0 ;
  assign n14994 = n1085 & ~n2687 ;
  assign n14995 = n14994 ^ n4769 ^ 1'b0 ;
  assign n14996 = n14995 ^ n14456 ^ n7428 ;
  assign n14997 = n6025 | n13802 ;
  assign n14998 = ( n859 & ~n3931 ) | ( n859 & n6800 ) | ( ~n3931 & n6800 ) ;
  assign n14999 = n3189 | n14998 ;
  assign n15000 = n2113 & n6270 ;
  assign n15001 = ~n10447 & n15000 ;
  assign n15002 = n6208 & ~n14884 ;
  assign n15003 = n3011 & ~n15002 ;
  assign n15004 = n3399 ^ n2733 ^ 1'b0 ;
  assign n15005 = ~n7348 & n15004 ;
  assign n15006 = n646 & ~n4175 ;
  assign n15007 = n15006 ^ n6848 ^ 1'b0 ;
  assign n15008 = n3092 & ~n15007 ;
  assign n15009 = ~n15005 & n15008 ;
  assign n15010 = ( ~n6169 & n10295 ) | ( ~n6169 & n15009 ) | ( n10295 & n15009 ) ;
  assign n15011 = n4037 ^ n2382 ^ 1'b0 ;
  assign n15012 = n4156 ^ n805 ^ 1'b0 ;
  assign n15013 = n15012 ^ n9068 ^ 1'b0 ;
  assign n15014 = n8482 | n15013 ;
  assign n15015 = ( n5891 & n6178 ) | ( n5891 & n8000 ) | ( n6178 & n8000 ) ;
  assign n15016 = n13962 ^ n3367 ^ 1'b0 ;
  assign n15017 = n15015 | n15016 ;
  assign n15018 = n5736 ^ n2156 ^ 1'b0 ;
  assign n15019 = n15018 ^ n225 ^ 1'b0 ;
  assign n15020 = n14844 | n15019 ;
  assign n15021 = n15020 ^ n7816 ^ 1'b0 ;
  assign n15022 = n5798 ^ n4370 ^ 1'b0 ;
  assign n15023 = n7627 & ~n15022 ;
  assign n15024 = ~n5350 & n15023 ;
  assign n15025 = n7000 ^ n4048 ^ 1'b0 ;
  assign n15026 = ~n10227 & n15025 ;
  assign n15030 = ~n2949 & n7177 ;
  assign n15031 = n2847 & n15030 ;
  assign n15027 = n2221 ^ x93 ^ 1'b0 ;
  assign n15028 = n7023 & n15027 ;
  assign n15029 = ( ~n2980 & n3290 ) | ( ~n2980 & n15028 ) | ( n3290 & n15028 ) ;
  assign n15032 = n15031 ^ n15029 ^ n14596 ;
  assign n15033 = ~n6136 & n6410 ;
  assign n15034 = n2823 & n15033 ;
  assign n15035 = n7228 | n15034 ;
  assign n15036 = n8080 ^ n3987 ^ 1'b0 ;
  assign n15037 = n10968 | n15036 ;
  assign n15038 = n15037 ^ n1027 ^ 1'b0 ;
  assign n15039 = ~n13108 & n15038 ;
  assign n15041 = n464 & n1351 ;
  assign n15042 = n15041 ^ n5329 ^ 1'b0 ;
  assign n15040 = n8722 & n9068 ;
  assign n15043 = n15042 ^ n15040 ^ 1'b0 ;
  assign n15044 = n15043 ^ n7306 ^ 1'b0 ;
  assign n15045 = n7437 & n15044 ;
  assign n15046 = n4721 & ~n7764 ;
  assign n15047 = ~n973 & n15046 ;
  assign n15048 = n2412 & n15047 ;
  assign n15049 = n4021 ^ n3515 ^ 1'b0 ;
  assign n15050 = n15049 ^ n10580 ^ 1'b0 ;
  assign n15051 = n13308 ^ n1761 ^ 1'b0 ;
  assign n15052 = n15051 ^ n4437 ^ n1035 ;
  assign n15053 = n14289 & n15052 ;
  assign n15054 = n15053 ^ n10574 ^ 1'b0 ;
  assign n15055 = ~n556 & n9085 ;
  assign n15056 = n1414 & n13308 ;
  assign n15057 = n2837 & ~n6681 ;
  assign n15058 = n8299 & n15057 ;
  assign n15059 = n2494 & ~n15058 ;
  assign n15060 = ~n11107 & n15059 ;
  assign n15061 = n14950 & ~n15060 ;
  assign n15062 = n15061 ^ n3413 ^ 1'b0 ;
  assign n15063 = n1821 & n9643 ;
  assign n15064 = n2904 & ~n15063 ;
  assign n15065 = n673 | n3415 ;
  assign n15066 = n13625 | n15065 ;
  assign n15067 = ~n5832 & n15066 ;
  assign n15068 = n10692 ^ n8436 ^ 1'b0 ;
  assign n15069 = n15068 ^ n5381 ^ n208 ;
  assign n15070 = n15067 & n15069 ;
  assign n15071 = n9162 & n9646 ;
  assign n15072 = ~n3143 & n4895 ;
  assign n15073 = n8353 ^ n6108 ^ 1'b0 ;
  assign n15074 = n1157 & n11603 ;
  assign n15075 = ~n15073 & n15074 ;
  assign n15076 = n3207 ^ n620 ^ 1'b0 ;
  assign n15077 = n15076 ^ n6174 ^ 1'b0 ;
  assign n15079 = n2098 ^ n1661 ^ 1'b0 ;
  assign n15080 = n1313 & ~n15079 ;
  assign n15078 = n2456 & ~n7594 ;
  assign n15081 = n15080 ^ n15078 ^ 1'b0 ;
  assign n15082 = n811 | n1880 ;
  assign n15083 = n10551 ^ n8906 ^ n3520 ;
  assign n15084 = ~n3343 & n3693 ;
  assign n15085 = ~n393 & n15084 ;
  assign n15086 = n15085 ^ n5061 ^ 1'b0 ;
  assign n15087 = ( n2206 & ~n10571 ) | ( n2206 & n15086 ) | ( ~n10571 & n15086 ) ;
  assign n15088 = n11008 ^ n2622 ^ 1'b0 ;
  assign n15089 = n9781 ^ n2014 ^ 1'b0 ;
  assign n15090 = n1147 & n15089 ;
  assign n15091 = ~n14987 & n15090 ;
  assign n15092 = n11269 ^ n192 ^ 1'b0 ;
  assign n15093 = n11143 ^ n7848 ^ 1'b0 ;
  assign n15094 = x21 & ~n15093 ;
  assign n15095 = n13046 ^ n3489 ^ 1'b0 ;
  assign n15097 = n4088 ^ n2958 ^ 1'b0 ;
  assign n15098 = n5559 & ~n15097 ;
  assign n15096 = ~n2448 & n9863 ;
  assign n15099 = n15098 ^ n15096 ^ 1'b0 ;
  assign n15100 = n15099 ^ n13104 ^ 1'b0 ;
  assign n15101 = n8832 ^ n5492 ^ 1'b0 ;
  assign n15102 = n5971 ^ n5238 ^ 1'b0 ;
  assign n15103 = ~n2497 & n15102 ;
  assign n15104 = n15103 ^ n8710 ^ 1'b0 ;
  assign n15112 = n2223 | n4519 ;
  assign n15107 = ~n1476 & n11521 ;
  assign n15108 = ~n11521 & n15107 ;
  assign n15109 = n1664 | n15108 ;
  assign n15105 = n3633 & ~n5096 ;
  assign n15106 = n15105 ^ n7431 ^ n3381 ;
  assign n15110 = n15109 ^ n15106 ^ 1'b0 ;
  assign n15111 = n5976 & ~n15110 ;
  assign n15113 = n15112 ^ n15111 ^ 1'b0 ;
  assign n15114 = n2915 ^ n1353 ^ 1'b0 ;
  assign n15115 = n740 & n5437 ;
  assign n15116 = n8317 & n15115 ;
  assign n15117 = n4950 | n15116 ;
  assign n15118 = n11607 & ~n15117 ;
  assign n15119 = n258 & ~n1176 ;
  assign n15120 = n11822 ^ n2395 ^ 1'b0 ;
  assign n15121 = n2758 & n9127 ;
  assign n15122 = n2827 | n7021 ;
  assign n15123 = ( ~n2886 & n10782 ) | ( ~n2886 & n14883 ) | ( n10782 & n14883 ) ;
  assign n15124 = n15123 ^ n7031 ^ 1'b0 ;
  assign n15126 = n12247 ^ n391 ^ 1'b0 ;
  assign n15125 = n6821 & ~n10558 ;
  assign n15127 = n15126 ^ n15125 ^ 1'b0 ;
  assign n15128 = n3844 | n6032 ;
  assign n15129 = n2794 ^ n719 ^ 1'b0 ;
  assign n15130 = n7120 & n15129 ;
  assign n15131 = n8571 ^ n4595 ^ 1'b0 ;
  assign n15132 = n4052 | n10733 ;
  assign n15133 = n2042 & ~n3599 ;
  assign n15134 = ( n1498 & n2848 ) | ( n1498 & ~n10382 ) | ( n2848 & ~n10382 ) ;
  assign n15135 = x38 & ~n15134 ;
  assign n15136 = ~n1691 & n15135 ;
  assign n15137 = n14641 & n15136 ;
  assign n15138 = n12697 ^ n981 ^ 1'b0 ;
  assign n15139 = n15137 | n15138 ;
  assign n15140 = n6663 ^ n5871 ^ n5628 ;
  assign n15141 = ~n4246 & n15140 ;
  assign n15142 = n10061 ^ n9286 ^ 1'b0 ;
  assign n15143 = ~n4638 & n15142 ;
  assign n15144 = n2134 | n4012 ;
  assign n15146 = x70 & n1012 ;
  assign n15147 = ~n2364 & n15146 ;
  assign n15145 = ~n1672 & n3976 ;
  assign n15148 = n15147 ^ n15145 ^ 1'b0 ;
  assign n15149 = n475 & ~n4549 ;
  assign n15150 = n2429 & n15149 ;
  assign n15151 = n15150 ^ n3083 ^ 1'b0 ;
  assign n15152 = ~n2274 & n5627 ;
  assign n15153 = n6640 | n15152 ;
  assign n15154 = n15153 ^ n14187 ^ 1'b0 ;
  assign n15155 = n4930 & n5942 ;
  assign n15156 = ~n9845 & n15155 ;
  assign n15157 = n15156 ^ n1361 ^ 1'b0 ;
  assign n15158 = n2840 | n15157 ;
  assign n15159 = n5535 ^ n5273 ^ 1'b0 ;
  assign n15160 = ~n15158 & n15159 ;
  assign n15161 = n15078 ^ n2064 ^ 1'b0 ;
  assign n15162 = n6153 ^ n3993 ^ 1'b0 ;
  assign n15163 = ~n939 & n3020 ;
  assign n15164 = ~n4362 & n15163 ;
  assign n15165 = n15162 & n15164 ;
  assign n15166 = ~n2217 & n15165 ;
  assign n15167 = n2948 | n10021 ;
  assign n15168 = n15167 ^ n2074 ^ 1'b0 ;
  assign n15169 = n10300 ^ n7018 ^ 1'b0 ;
  assign n15170 = n5277 & n15169 ;
  assign n15171 = n3681 ^ n3472 ^ 1'b0 ;
  assign n15172 = n3455 & ~n15171 ;
  assign n15173 = x69 & n3429 ;
  assign n15174 = ~n2170 & n15173 ;
  assign n15175 = n7526 | n15174 ;
  assign n15176 = n3130 & ~n15175 ;
  assign n15177 = ~n10951 & n15176 ;
  assign n15180 = n5293 & ~n12756 ;
  assign n15181 = n14766 & n15180 ;
  assign n15178 = ~n1422 & n11867 ;
  assign n15179 = n14225 | n15178 ;
  assign n15182 = n15181 ^ n15179 ^ 1'b0 ;
  assign n15183 = n6963 ^ n1794 ^ 1'b0 ;
  assign n15184 = n5896 & ~n15183 ;
  assign n15185 = n11923 ^ n3560 ^ 1'b0 ;
  assign n15186 = n1916 ^ n1742 ^ 1'b0 ;
  assign n15187 = n15185 & n15186 ;
  assign n15188 = n15187 ^ n13308 ^ 1'b0 ;
  assign n15189 = ~n4605 & n10983 ;
  assign n15193 = n6954 ^ n3524 ^ 1'b0 ;
  assign n15194 = n15193 ^ n7216 ^ 1'b0 ;
  assign n15195 = n2802 & ~n15194 ;
  assign n15190 = n11212 ^ n7837 ^ 1'b0 ;
  assign n15191 = n10743 | n15190 ;
  assign n15192 = n15191 ^ n2201 ^ 1'b0 ;
  assign n15196 = n15195 ^ n15192 ^ n14654 ;
  assign n15197 = n15196 ^ n9446 ^ 1'b0 ;
  assign n15198 = n8853 ^ n440 ^ 1'b0 ;
  assign n15199 = n5662 ^ n5457 ^ 1'b0 ;
  assign n15200 = ~n15034 & n15199 ;
  assign n15201 = n3284 ^ n3020 ^ n1102 ;
  assign n15202 = n6854 & ~n15201 ;
  assign n15203 = n15202 ^ n13514 ^ 1'b0 ;
  assign n15204 = ~n732 & n15203 ;
  assign n15205 = n15204 ^ n6809 ^ 1'b0 ;
  assign n15206 = n7260 ^ n6935 ^ n2636 ;
  assign n15207 = n15206 ^ n5628 ^ n2656 ;
  assign n15208 = n5188 | n14161 ;
  assign n15210 = x20 & n4848 ;
  assign n15211 = n15210 ^ n5036 ^ 1'b0 ;
  assign n15209 = n1920 & n6702 ;
  assign n15212 = n15211 ^ n15209 ^ 1'b0 ;
  assign n15213 = n3789 & n5921 ;
  assign n15214 = n5946 ^ n897 ^ 1'b0 ;
  assign n15215 = n3369 & n9472 ;
  assign n15216 = n1624 & n4849 ;
  assign n15217 = n14054 ^ n9458 ^ 1'b0 ;
  assign n15218 = n15187 ^ n14654 ^ 1'b0 ;
  assign n15219 = n9611 & n13231 ;
  assign n15220 = ( ~n5378 & n10516 ) | ( ~n5378 & n15219 ) | ( n10516 & n15219 ) ;
  assign n15221 = ~n6787 & n7765 ;
  assign n15222 = ~n6933 & n15221 ;
  assign n15223 = n758 & ~n3113 ;
  assign n15224 = ~n15222 & n15223 ;
  assign n15225 = n15224 ^ n6511 ^ 1'b0 ;
  assign n15226 = n11566 ^ n6458 ^ 1'b0 ;
  assign n15227 = n14642 ^ n9208 ^ 1'b0 ;
  assign n15228 = n12197 & n15227 ;
  assign n15229 = n4265 | n9474 ;
  assign n15230 = n9645 | n15229 ;
  assign n15231 = n15230 ^ n7175 ^ 1'b0 ;
  assign n15232 = n2948 ^ n1967 ^ 1'b0 ;
  assign n15233 = n1166 | n6445 ;
  assign n15234 = n15233 ^ n14229 ^ 1'b0 ;
  assign n15235 = ~n2189 & n3750 ;
  assign n15236 = x45 | n3082 ;
  assign n15237 = ~n1688 & n9071 ;
  assign n15238 = n12993 ^ n6299 ^ n2896 ;
  assign n15239 = n3458 | n15238 ;
  assign n15240 = n15239 ^ n3158 ^ 1'b0 ;
  assign n15241 = n1788 & n15240 ;
  assign n15242 = n1963 ^ n1219 ^ 1'b0 ;
  assign n15243 = ~n6400 & n15242 ;
  assign n15244 = n13667 ^ n1245 ^ 1'b0 ;
  assign n15245 = ~n4354 & n15244 ;
  assign n15246 = n2814 | n3601 ;
  assign n15247 = n8934 & n15246 ;
  assign n15248 = ~n1195 & n12481 ;
  assign n15249 = n15247 & n15248 ;
  assign n15250 = n5707 & n12861 ;
  assign n15251 = n15250 ^ n10843 ^ 1'b0 ;
  assign n15253 = n8224 ^ n998 ^ 1'b0 ;
  assign n15254 = n4032 | n15253 ;
  assign n15252 = ~n5159 & n8268 ;
  assign n15255 = n15254 ^ n15252 ^ 1'b0 ;
  assign n15256 = n3459 ^ x3 ^ 1'b0 ;
  assign n15257 = ~n7986 & n9487 ;
  assign n15258 = ~n7371 & n10568 ;
  assign n15259 = n15258 ^ n4564 ^ 1'b0 ;
  assign n15260 = n1629 ^ x121 ^ 1'b0 ;
  assign n15261 = n6317 ^ n2026 ^ 1'b0 ;
  assign n15262 = ~n15260 & n15261 ;
  assign n15263 = n9662 ^ n5203 ^ 1'b0 ;
  assign n15264 = n15262 & ~n15263 ;
  assign n15265 = n4470 & ~n9342 ;
  assign n15266 = n8921 ^ n658 ^ 1'b0 ;
  assign n15267 = n11143 & n15266 ;
  assign n15268 = ~n5362 & n15267 ;
  assign n15269 = x19 | n1247 ;
  assign n15270 = n8342 ^ n1510 ^ 1'b0 ;
  assign n15271 = ~n9812 & n15270 ;
  assign n15272 = n2696 | n7163 ;
  assign n15273 = n3602 & n15272 ;
  assign n15275 = ~n976 & n5211 ;
  assign n15276 = ~n7110 & n15275 ;
  assign n15274 = n5728 | n11699 ;
  assign n15277 = n15276 ^ n15274 ^ 1'b0 ;
  assign n15278 = n14333 ^ n8319 ^ 1'b0 ;
  assign n15284 = n1639 ^ n384 ^ 1'b0 ;
  assign n15279 = x114 & ~n1489 ;
  assign n15280 = n1801 ^ n456 ^ 1'b0 ;
  assign n15281 = n15279 | n15280 ;
  assign n15282 = n13978 ^ n5872 ^ 1'b0 ;
  assign n15283 = ( n9334 & n15281 ) | ( n9334 & n15282 ) | ( n15281 & n15282 ) ;
  assign n15285 = n15284 ^ n15283 ^ n556 ;
  assign n15286 = n4452 ^ n2134 ^ 1'b0 ;
  assign n15287 = n10536 & n15286 ;
  assign n15288 = n4917 & ~n13207 ;
  assign n15289 = ~n254 & n14596 ;
  assign n15290 = n931 & n2008 ;
  assign n15291 = n4152 & ~n5157 ;
  assign n15292 = n15290 & n15291 ;
  assign n15293 = n509 & ~n11768 ;
  assign n15294 = n2562 & n15293 ;
  assign n15295 = ~n14073 & n15294 ;
  assign n15297 = n4742 ^ n704 ^ 1'b0 ;
  assign n15298 = n1096 & ~n15297 ;
  assign n15296 = n1331 & ~n4162 ;
  assign n15299 = n15298 ^ n15296 ^ 1'b0 ;
  assign n15303 = n5631 ^ n5104 ^ 1'b0 ;
  assign n15300 = n7463 ^ n1096 ^ 1'b0 ;
  assign n15301 = n2126 & n15300 ;
  assign n15302 = ~n3564 & n15301 ;
  assign n15304 = n15303 ^ n15302 ^ 1'b0 ;
  assign n15305 = n2484 | n9307 ;
  assign n15306 = ( n421 & n3153 ) | ( n421 & n3818 ) | ( n3153 & n3818 ) ;
  assign n15307 = ( ~n6975 & n12634 ) | ( ~n6975 & n15306 ) | ( n12634 & n15306 ) ;
  assign n15308 = n9878 ^ n7995 ^ 1'b0 ;
  assign n15309 = n13187 & n15308 ;
  assign n15310 = n15309 ^ n15202 ^ n2567 ;
  assign n15311 = n4989 & n15310 ;
  assign n15312 = n7851 & n15311 ;
  assign n15313 = n1756 | n3478 ;
  assign n15314 = n273 & n10479 ;
  assign n15315 = n14312 | n15314 ;
  assign n15316 = n5762 & ~n15315 ;
  assign n15317 = n3903 & ~n15316 ;
  assign n15318 = n1424 & ~n1522 ;
  assign n15319 = n7554 & n15318 ;
  assign n15320 = n7980 | n9080 ;
  assign n15321 = n15320 ^ n179 ^ 1'b0 ;
  assign n15322 = n11920 | n13627 ;
  assign n15323 = n4553 & ~n15322 ;
  assign n15324 = n5996 ^ n5945 ^ 1'b0 ;
  assign n15325 = ~n2275 & n15324 ;
  assign n15326 = n2140 & ~n4345 ;
  assign n15327 = n2170 & n15326 ;
  assign n15328 = n1570 & n8124 ;
  assign n15329 = n2622 ^ n2113 ^ 1'b0 ;
  assign n15330 = n6078 & n15329 ;
  assign n15331 = n15330 ^ n3693 ^ 1'b0 ;
  assign n15332 = n15328 & n15331 ;
  assign n15333 = n11295 ^ n6179 ^ 1'b0 ;
  assign n15334 = n5830 & ~n9110 ;
  assign n15335 = n8982 ^ n6613 ^ 1'b0 ;
  assign n15336 = n15334 | n15335 ;
  assign n15337 = n15336 ^ n6930 ^ n749 ;
  assign n15338 = n5744 ^ n3110 ^ 1'b0 ;
  assign n15339 = ~n829 & n9447 ;
  assign n15340 = n15339 ^ n3965 ^ 1'b0 ;
  assign n15341 = n15338 & ~n15340 ;
  assign n15342 = n5413 ^ n2419 ^ 1'b0 ;
  assign n15343 = n4836 & ~n15342 ;
  assign n15344 = n15343 ^ n10558 ^ 1'b0 ;
  assign n15345 = ( n5853 & n6998 ) | ( n5853 & n15344 ) | ( n6998 & n15344 ) ;
  assign n15346 = n15341 & ~n15345 ;
  assign n15347 = ( n1052 & n1168 ) | ( n1052 & n2123 ) | ( n1168 & n2123 ) ;
  assign n15348 = n11519 & ~n15347 ;
  assign n15349 = n5674 | n7343 ;
  assign n15350 = n15349 ^ n4618 ^ 1'b0 ;
  assign n15351 = n13857 ^ n9813 ^ 1'b0 ;
  assign n15352 = ~n14198 & n15351 ;
  assign n15353 = n2146 & n6844 ;
  assign n15354 = ~n15352 & n15353 ;
  assign n15357 = n2234 & ~n2419 ;
  assign n15358 = n3590 & n15357 ;
  assign n15359 = n15358 ^ n7368 ^ 1'b0 ;
  assign n15355 = ~n3300 & n3386 ;
  assign n15356 = n15355 ^ n8446 ^ 1'b0 ;
  assign n15360 = n15359 ^ n15356 ^ 1'b0 ;
  assign n15361 = n5470 & ~n15360 ;
  assign n15362 = n4251 ^ n2751 ^ 1'b0 ;
  assign n15363 = n8286 & ~n15362 ;
  assign n15364 = n3944 & n15363 ;
  assign n15365 = ~n8543 & n15364 ;
  assign n15366 = n4616 | n13592 ;
  assign n15367 = n15241 ^ n1790 ^ 1'b0 ;
  assign n15368 = n5062 ^ n4576 ^ 1'b0 ;
  assign n15369 = n9115 & ~n11936 ;
  assign n15370 = ~n2211 & n15369 ;
  assign n15371 = n4707 & ~n5073 ;
  assign n15372 = n15371 ^ n8043 ^ 1'b0 ;
  assign n15373 = ~n7383 & n15372 ;
  assign n15374 = ~n1761 & n5569 ;
  assign n15375 = n5592 & n6187 ;
  assign n15376 = n4273 & n15375 ;
  assign n15377 = n6208 & ~n15376 ;
  assign n15378 = n12355 ^ n2107 ^ 1'b0 ;
  assign n15379 = ( ~n12673 & n14083 ) | ( ~n12673 & n15378 ) | ( n14083 & n15378 ) ;
  assign n15380 = n5385 ^ n4336 ^ 1'b0 ;
  assign n15381 = n5020 | n15081 ;
  assign n15383 = n4061 & n4700 ;
  assign n15382 = n2855 & n5569 ;
  assign n15384 = n15383 ^ n15382 ^ 1'b0 ;
  assign n15385 = n9729 ^ n7133 ^ 1'b0 ;
  assign n15386 = n13665 & n15385 ;
  assign n15387 = n1597 & ~n5220 ;
  assign n15388 = n5814 | n12778 ;
  assign n15389 = n4315 & ~n10794 ;
  assign n15390 = n14093 ^ n1111 ^ 1'b0 ;
  assign n15391 = ~n5258 & n15390 ;
  assign n15392 = n13099 ^ n978 ^ 1'b0 ;
  assign n15393 = n8797 ^ n5437 ^ 1'b0 ;
  assign n15394 = n1552 | n15393 ;
  assign n15395 = n15394 ^ n8700 ^ 1'b0 ;
  assign n15396 = n15392 & ~n15395 ;
  assign n15397 = n15022 ^ n13024 ^ n11000 ;
  assign n15399 = ( ~n799 & n4056 ) | ( ~n799 & n8194 ) | ( n4056 & n8194 ) ;
  assign n15398 = ~n8809 & n15045 ;
  assign n15400 = n15399 ^ n15398 ^ 1'b0 ;
  assign n15401 = n9561 ^ n5499 ^ n393 ;
  assign n15402 = ( ~n5374 & n14842 ) | ( ~n5374 & n15401 ) | ( n14842 & n15401 ) ;
  assign n15403 = n5206 ^ n3920 ^ 1'b0 ;
  assign n15404 = n3372 & ~n15403 ;
  assign n15405 = n15404 ^ n8249 ^ 1'b0 ;
  assign n15406 = n4950 ^ n353 ^ 1'b0 ;
  assign n15407 = n15406 ^ n2246 ^ 1'b0 ;
  assign n15408 = n1097 | n15407 ;
  assign n15409 = n15408 ^ n7157 ^ 1'b0 ;
  assign n15410 = n15409 ^ n4938 ^ 1'b0 ;
  assign n15411 = n2398 | n13602 ;
  assign n15412 = n15410 | n15411 ;
  assign n15413 = ~n10073 & n13215 ;
  assign n15414 = n1388 ^ n171 ^ 1'b0 ;
  assign n15415 = n559 & ~n15414 ;
  assign n15416 = n9098 & n15415 ;
  assign n15417 = ~n15413 & n15416 ;
  assign n15418 = n3511 & ~n3668 ;
  assign n15419 = ~n3450 & n15418 ;
  assign n15420 = n15419 ^ n3348 ^ 1'b0 ;
  assign n15421 = n15420 ^ n3951 ^ 1'b0 ;
  assign n15422 = n13592 ^ n2151 ^ 1'b0 ;
  assign n15423 = n143 & n15422 ;
  assign n15424 = n3458 ^ n3311 ^ n903 ;
  assign n15425 = n15423 & ~n15424 ;
  assign n15426 = ~n6216 & n7385 ;
  assign n15427 = n732 & n1133 ;
  assign n15428 = ~n11065 & n15427 ;
  assign n15430 = ~n3398 & n3546 ;
  assign n15429 = n1898 & n2662 ;
  assign n15431 = n15430 ^ n15429 ^ 1'b0 ;
  assign n15432 = ( n759 & n13325 ) | ( n759 & ~n15431 ) | ( n13325 & ~n15431 ) ;
  assign n15433 = n7029 & n11501 ;
  assign n15434 = n11216 & ~n15433 ;
  assign n15435 = n3844 & n15434 ;
  assign n15436 = n3615 & ~n10707 ;
  assign n15437 = ~n2444 & n15436 ;
  assign n15438 = n716 & ~n8914 ;
  assign n15439 = n4755 | n11250 ;
  assign n15440 = n15438 | n15439 ;
  assign n15441 = n11622 ^ n10402 ^ 1'b0 ;
  assign n15442 = n4066 | n15441 ;
  assign n15443 = n1143 & n12623 ;
  assign n15444 = n2460 & n14786 ;
  assign n15445 = n759 & ~n3182 ;
  assign n15446 = n15445 ^ n1586 ^ 1'b0 ;
  assign n15447 = ~n301 & n12161 ;
  assign n15448 = n15447 ^ n2483 ^ 1'b0 ;
  assign n15449 = n2866 ^ x89 ^ 1'b0 ;
  assign n15450 = n1737 & ~n15449 ;
  assign n15452 = n4561 | n13318 ;
  assign n15453 = ~n4808 & n15452 ;
  assign n15451 = n9864 | n15222 ;
  assign n15454 = n15453 ^ n15451 ^ 1'b0 ;
  assign n15455 = n3029 | n15454 ;
  assign n15456 = n15455 ^ n8747 ^ 1'b0 ;
  assign n15457 = n3691 | n15080 ;
  assign n15458 = n3708 | n10729 ;
  assign n15459 = n3601 & ~n15458 ;
  assign n15460 = n1805 | n4021 ;
  assign n15461 = n7542 & ~n14610 ;
  assign n15462 = n15461 ^ n224 ^ 1'b0 ;
  assign n15463 = n4844 | n9089 ;
  assign n15464 = n12202 & n12993 ;
  assign n15465 = n7775 ^ n7602 ^ 1'b0 ;
  assign n15466 = ~n745 & n1578 ;
  assign n15467 = ~n2948 & n15466 ;
  assign n15468 = n868 | n15467 ;
  assign n15469 = n15465 | n15468 ;
  assign n15470 = n5389 ^ n1354 ^ 1'b0 ;
  assign n15471 = n1372 & ~n15470 ;
  assign n15474 = n2763 & n2960 ;
  assign n15475 = n4436 | n15474 ;
  assign n15476 = n15475 ^ n14661 ^ 1'b0 ;
  assign n15472 = x46 & ~n3287 ;
  assign n15473 = ~n2560 & n15472 ;
  assign n15477 = n15476 ^ n15473 ^ n2722 ;
  assign n15478 = n10296 ^ n1635 ^ 1'b0 ;
  assign n15479 = n12851 & n15478 ;
  assign n15480 = n2543 & n15479 ;
  assign n15481 = ~n4556 & n15480 ;
  assign n15482 = n9053 | n14997 ;
  assign n15483 = n14128 ^ n13692 ^ 1'b0 ;
  assign n15484 = n6972 | n15483 ;
  assign n15485 = n9169 | n10934 ;
  assign n15486 = n2267 & ~n15485 ;
  assign n15487 = n3249 & ~n15486 ;
  assign n15488 = n15487 ^ n7960 ^ 1'b0 ;
  assign n15489 = ~n10677 & n15488 ;
  assign n15490 = n15095 ^ n1092 ^ 1'b0 ;
  assign n15491 = n4030 | n11740 ;
  assign n15492 = ( ~n5669 & n7755 ) | ( ~n5669 & n10216 ) | ( n7755 & n10216 ) ;
  assign n15493 = ( n3806 & ~n15491 ) | ( n3806 & n15492 ) | ( ~n15491 & n15492 ) ;
  assign n15494 = n8209 | n9729 ;
  assign n15495 = n15493 & ~n15494 ;
  assign n15498 = n5416 & n11775 ;
  assign n15499 = n15498 ^ n3318 ^ 1'b0 ;
  assign n15496 = n14877 ^ n1552 ^ 1'b0 ;
  assign n15497 = n4523 & ~n15496 ;
  assign n15500 = n15499 ^ n15497 ^ n6894 ;
  assign n15501 = n792 & ~n15500 ;
  assign n15502 = n5486 & n15501 ;
  assign n15503 = ~n3437 & n4567 ;
  assign n15504 = n810 & ~n6036 ;
  assign n15505 = ~n15503 & n15504 ;
  assign n15506 = n15505 ^ n1056 ^ 1'b0 ;
  assign n15507 = n8911 & n11315 ;
  assign n15508 = n9212 & ~n12179 ;
  assign n15509 = n13904 ^ n7547 ^ 1'b0 ;
  assign n15510 = ~n15508 & n15509 ;
  assign n15512 = n5784 ^ n3153 ^ 1'b0 ;
  assign n15513 = n4728 & ~n15512 ;
  assign n15511 = n9662 ^ n2357 ^ n430 ;
  assign n15514 = n15513 ^ n15511 ^ 1'b0 ;
  assign n15515 = n14846 ^ n12905 ^ 1'b0 ;
  assign n15516 = n12394 | n14612 ;
  assign n15517 = n1569 & ~n5296 ;
  assign n15518 = n9731 ^ n243 ^ 1'b0 ;
  assign n15519 = n14991 ^ n11692 ^ 1'b0 ;
  assign n15520 = n15518 & n15519 ;
  assign n15521 = n7813 ^ n4555 ^ 1'b0 ;
  assign n15522 = n2497 | n4315 ;
  assign n15524 = ~n488 & n1116 ;
  assign n15523 = n1567 & ~n14854 ;
  assign n15525 = n15524 ^ n15523 ^ 1'b0 ;
  assign n15526 = n3750 ^ n3350 ^ 1'b0 ;
  assign n15527 = ~n5090 & n15526 ;
  assign n15528 = n10409 ^ n283 ^ 1'b0 ;
  assign n15530 = n3297 & n8601 ;
  assign n15531 = ~n5253 & n15530 ;
  assign n15532 = n9323 & ~n15531 ;
  assign n15533 = ~n3937 & n15532 ;
  assign n15529 = n4521 & ~n5481 ;
  assign n15534 = n15533 ^ n15529 ^ 1'b0 ;
  assign n15535 = n14654 ^ n9966 ^ 1'b0 ;
  assign n15536 = x75 & n15535 ;
  assign n15537 = n400 | n15391 ;
  assign n15538 = n14109 ^ n10669 ^ 1'b0 ;
  assign n15539 = n4253 & ~n4777 ;
  assign n15540 = n1743 | n6415 ;
  assign n15541 = ~n5254 & n9213 ;
  assign n15542 = n15541 ^ n400 ^ 1'b0 ;
  assign n15544 = n461 | n6731 ;
  assign n15545 = n2985 & ~n4240 ;
  assign n15546 = n8601 ^ n4090 ^ 1'b0 ;
  assign n15547 = ~n15545 & n15546 ;
  assign n15548 = ~n15544 & n15547 ;
  assign n15543 = n479 & n10767 ;
  assign n15549 = n15548 ^ n15543 ^ 1'b0 ;
  assign n15550 = n12627 ^ n4010 ^ n1510 ;
  assign n15551 = n3964 & ~n15099 ;
  assign n15552 = n1392 & n15551 ;
  assign n15553 = ~n7936 & n13342 ;
  assign n15554 = n15553 ^ n6073 ^ 1'b0 ;
  assign n15555 = ~n9834 & n12192 ;
  assign n15556 = n15555 ^ n15078 ^ 1'b0 ;
  assign n15557 = n9784 & n13951 ;
  assign n15558 = n13154 & ~n15557 ;
  assign n15559 = ~n2168 & n4666 ;
  assign n15560 = n15042 & n15559 ;
  assign n15562 = ~n3459 & n7784 ;
  assign n15563 = n15562 ^ n4068 ^ 1'b0 ;
  assign n15561 = n12796 ^ n10673 ^ 1'b0 ;
  assign n15564 = n15563 ^ n15561 ^ n13483 ;
  assign n15565 = ~n2506 & n6291 ;
  assign n15566 = n15565 ^ n5193 ^ 1'b0 ;
  assign n15567 = n362 | n15566 ;
  assign n15568 = n15567 ^ n6718 ^ 1'b0 ;
  assign n15569 = n13356 ^ n6437 ^ 1'b0 ;
  assign n15570 = ~n3601 & n15569 ;
  assign n15571 = n10794 ^ n971 ^ 1'b0 ;
  assign n15572 = ~n9653 & n10214 ;
  assign n15573 = n3776 ^ n1606 ^ 1'b0 ;
  assign n15574 = ~n2935 & n15573 ;
  assign n15575 = n14585 & n15574 ;
  assign n15576 = n1784 & n15575 ;
  assign n15577 = n11595 & ~n15576 ;
  assign n15578 = n15576 & n15577 ;
  assign n15579 = n15578 ^ n7574 ^ n874 ;
  assign n15580 = n4458 ^ n4155 ^ 1'b0 ;
  assign n15581 = n741 & n15580 ;
  assign n15582 = n15581 ^ n1835 ^ 1'b0 ;
  assign n15583 = ~n2708 & n15582 ;
  assign n15584 = n13082 ^ n3135 ^ 1'b0 ;
  assign n15585 = n15584 ^ n5150 ^ n2913 ;
  assign n15586 = n1291 & n15585 ;
  assign n15587 = n8856 & n15586 ;
  assign n15591 = n3629 & ~n8151 ;
  assign n15589 = n4810 | n5486 ;
  assign n15590 = n15589 ^ n5834 ^ 1'b0 ;
  assign n15588 = n738 & ~n8231 ;
  assign n15592 = n15591 ^ n15590 ^ n15588 ;
  assign n15593 = n15078 ^ n13872 ^ 1'b0 ;
  assign n15594 = n10799 ^ n1491 ^ 1'b0 ;
  assign n15595 = n11381 ^ n10024 ^ 1'b0 ;
  assign n15599 = n4255 | n7953 ;
  assign n15596 = n9068 ^ n391 ^ 1'b0 ;
  assign n15597 = n3328 & n15596 ;
  assign n15598 = n1346 | n15597 ;
  assign n15600 = n15599 ^ n15598 ^ 1'b0 ;
  assign n15601 = n5811 ^ n3642 ^ 1'b0 ;
  assign n15602 = n6291 & n15601 ;
  assign n15603 = n15602 ^ n4048 ^ 1'b0 ;
  assign n15604 = n15603 ^ n6609 ^ 1'b0 ;
  assign n15605 = n13463 | n15604 ;
  assign n15606 = ~n4955 & n7767 ;
  assign n15607 = n15605 & n15606 ;
  assign n15608 = n11205 & ~n15607 ;
  assign n15609 = n6135 & ~n12866 ;
  assign n15610 = n11611 ^ n2330 ^ 1'b0 ;
  assign n15611 = n15609 & ~n15610 ;
  assign n15612 = ~n7073 & n15611 ;
  assign n15613 = ~n3704 & n7403 ;
  assign n15614 = n7649 & ~n15613 ;
  assign n15615 = n9691 ^ n7036 ^ 1'b0 ;
  assign n15616 = ~n4643 & n6863 ;
  assign n15617 = ~n10665 & n15616 ;
  assign n15618 = n666 & ~n3054 ;
  assign n15619 = ~n10699 & n15618 ;
  assign n15620 = n3241 ^ n1847 ^ 1'b0 ;
  assign n15621 = n15609 ^ n8153 ^ 1'b0 ;
  assign n15622 = ( n213 & n15620 ) | ( n213 & ~n15621 ) | ( n15620 & ~n15621 ) ;
  assign n15623 = ~n1526 & n8990 ;
  assign n15624 = n15623 ^ n2959 ^ 1'b0 ;
  assign n15625 = n13669 | n15624 ;
  assign n15626 = n6040 ^ n3485 ^ 1'b0 ;
  assign n15627 = ~n15625 & n15626 ;
  assign n15628 = n4639 & ~n6362 ;
  assign n15629 = n15628 ^ n371 ^ 1'b0 ;
  assign n15630 = n14293 & n15629 ;
  assign n15631 = n9812 & n15630 ;
  assign n15632 = n10982 ^ n1157 ^ 1'b0 ;
  assign n15633 = n7736 & n13284 ;
  assign n15634 = n2050 & ~n15633 ;
  assign n15635 = n15632 & n15634 ;
  assign n15636 = ~n6168 & n15635 ;
  assign n15637 = n4424 ^ n3389 ^ 1'b0 ;
  assign n15638 = n4844 & n15637 ;
  assign n15639 = n15638 ^ n11279 ^ 1'b0 ;
  assign n15640 = n208 | n4183 ;
  assign n15641 = ~n6779 & n13301 ;
  assign n15642 = ~n15640 & n15641 ;
  assign n15643 = n5598 | n15642 ;
  assign n15644 = n1862 | n9768 ;
  assign n15645 = n1787 & ~n15644 ;
  assign n15647 = n6669 ^ n4247 ^ 1'b0 ;
  assign n15646 = n13440 & n14205 ;
  assign n15648 = n15647 ^ n15646 ^ 1'b0 ;
  assign n15649 = n9236 ^ n5787 ^ 1'b0 ;
  assign n15650 = ~n4808 & n15649 ;
  assign n15651 = n5510 & n15650 ;
  assign n15652 = n13798 ^ n3613 ^ 1'b0 ;
  assign n15653 = n15652 ^ n5497 ^ 1'b0 ;
  assign n15654 = ~n2489 & n2492 ;
  assign n15655 = n11727 & n15654 ;
  assign n15656 = n15655 ^ n6839 ^ 1'b0 ;
  assign n15657 = n9139 & n15656 ;
  assign n15658 = ( n3459 & ~n10026 ) | ( n3459 & n15657 ) | ( ~n10026 & n15657 ) ;
  assign n15659 = n7548 ^ n4233 ^ 1'b0 ;
  assign n15660 = n15659 ^ n8430 ^ n3987 ;
  assign n15661 = n12238 ^ n10187 ^ 1'b0 ;
  assign n15662 = n5891 ^ n1147 ^ 1'b0 ;
  assign n15663 = n14121 | n15662 ;
  assign n15664 = n12684 | n15663 ;
  assign n15665 = n8568 & n15664 ;
  assign n15666 = n14641 & ~n15652 ;
  assign n15667 = n15666 ^ n2020 ^ 1'b0 ;
  assign n15668 = n15667 ^ n11435 ^ n2193 ;
  assign n15670 = n6385 | n9748 ;
  assign n15669 = ~n6472 & n8235 ;
  assign n15671 = n15670 ^ n15669 ^ 1'b0 ;
  assign n15672 = n6107 & n8737 ;
  assign n15673 = n15672 ^ n6295 ^ 1'b0 ;
  assign n15674 = n3172 | n14370 ;
  assign n15675 = n7809 & ~n15674 ;
  assign n15676 = n2127 | n4075 ;
  assign n15677 = n15598 ^ n4872 ^ 1'b0 ;
  assign n15678 = n15676 | n15677 ;
  assign n15679 = n15678 ^ n1186 ^ 1'b0 ;
  assign n15680 = n6437 ^ n6224 ^ 1'b0 ;
  assign n15681 = n5874 & n15680 ;
  assign n15682 = ~n2396 & n15681 ;
  assign n15686 = n5715 & ~n7248 ;
  assign n15687 = n15686 ^ n11019 ^ 1'b0 ;
  assign n15688 = ~n4683 & n15687 ;
  assign n15683 = n676 & n1382 ;
  assign n15684 = n833 & ~n12229 ;
  assign n15685 = n15683 | n15684 ;
  assign n15689 = n15688 ^ n15685 ^ 1'b0 ;
  assign n15690 = n10447 ^ n2126 ^ 1'b0 ;
  assign n15691 = ~n14596 & n15690 ;
  assign n15692 = ~n6467 & n7185 ;
  assign n15693 = n692 & ~n11201 ;
  assign n15694 = n4389 & n15693 ;
  assign n15695 = n12658 ^ n1295 ^ 1'b0 ;
  assign n15696 = n171 | n15695 ;
  assign n15697 = n7797 ^ n7002 ^ 1'b0 ;
  assign n15698 = n13709 & n15697 ;
  assign n15699 = n3354 & n15698 ;
  assign n15700 = n1406 & ~n6916 ;
  assign n15701 = n15700 ^ n12549 ^ 1'b0 ;
  assign n15702 = n2397 & n4495 ;
  assign n15703 = ~n169 & n7755 ;
  assign n15704 = n1860 & n15703 ;
  assign n15705 = n913 | n15704 ;
  assign n15706 = n7496 | n15705 ;
  assign n15707 = ~n1266 & n5193 ;
  assign n15708 = n2935 & n15707 ;
  assign n15709 = n4461 ^ n2381 ^ 1'b0 ;
  assign n15710 = ~n6426 & n15709 ;
  assign n15711 = ( ~n7038 & n9845 ) | ( ~n7038 & n15710 ) | ( n9845 & n15710 ) ;
  assign n15712 = n5181 & n15711 ;
  assign n15713 = ~n15708 & n15712 ;
  assign n15714 = ~n15706 & n15713 ;
  assign n15715 = n4778 & n6270 ;
  assign n15716 = n15715 ^ n767 ^ 1'b0 ;
  assign n15718 = n2924 ^ n1995 ^ 1'b0 ;
  assign n15719 = n5268 & ~n15718 ;
  assign n15717 = n2328 & n7531 ;
  assign n15720 = n15719 ^ n15717 ^ n4967 ;
  assign n15721 = n5662 & n6619 ;
  assign n15722 = n15720 & n15721 ;
  assign n15723 = ( ~n3287 & n11032 ) | ( ~n3287 & n15584 ) | ( n11032 & n15584 ) ;
  assign n15724 = n10873 & n15723 ;
  assign n15725 = n13271 | n13699 ;
  assign n15726 = n1773 & n4863 ;
  assign n15729 = n1030 & n11267 ;
  assign n15730 = n6529 & n15729 ;
  assign n15731 = n1038 & n15730 ;
  assign n15727 = n9207 ^ n1076 ^ 1'b0 ;
  assign n15728 = ~n4115 & n15727 ;
  assign n15732 = n15731 ^ n15728 ^ 1'b0 ;
  assign n15733 = n8530 ^ n3188 ^ 1'b0 ;
  assign n15734 = n1995 & n3148 ;
  assign n15735 = n8650 ^ n774 ^ 1'b0 ;
  assign n15736 = ~n6864 & n15735 ;
  assign n15737 = n4280 | n7662 ;
  assign n15738 = n15737 ^ n319 ^ 1'b0 ;
  assign n15739 = ~n15736 & n15738 ;
  assign n15740 = n1787 | n7145 ;
  assign n15741 = n15740 ^ n8508 ^ 1'b0 ;
  assign n15742 = n147 | n5102 ;
  assign n15743 = n548 & ~n15742 ;
  assign n15745 = n1066 & ~n3995 ;
  assign n15746 = ~n1422 & n15745 ;
  assign n15747 = n5069 & ~n15746 ;
  assign n15748 = n15747 ^ n11715 ^ 1'b0 ;
  assign n15744 = x86 & ~n1811 ;
  assign n15749 = n15748 ^ n15744 ^ 1'b0 ;
  assign n15750 = ~n2327 & n8653 ;
  assign n15751 = n15750 ^ n1625 ^ 1'b0 ;
  assign n15752 = n7011 & n15751 ;
  assign n15753 = n1448 | n15752 ;
  assign n15754 = n3320 & n6953 ;
  assign n15755 = ~n905 & n15754 ;
  assign n15756 = n15755 ^ n3822 ^ n1058 ;
  assign n15757 = n15756 ^ n12654 ^ 1'b0 ;
  assign n15758 = n5486 & ~n14880 ;
  assign n15759 = n11280 & n15758 ;
  assign n15760 = n267 | n855 ;
  assign n15761 = n9191 & ~n15760 ;
  assign n15762 = n15761 ^ n6969 ^ 1'b0 ;
  assign n15763 = n13726 | n15762 ;
  assign n15764 = ~n4766 & n9603 ;
  assign n15765 = ~n7332 & n11292 ;
  assign n15766 = n14138 ^ n13761 ^ n4011 ;
  assign n15767 = n4433 ^ n666 ^ 1'b0 ;
  assign n15768 = n6378 ^ n5090 ^ n1440 ;
  assign n15769 = ( ~n3344 & n4265 ) | ( ~n3344 & n15768 ) | ( n4265 & n15768 ) ;
  assign n15770 = n15769 ^ n2318 ^ 1'b0 ;
  assign n15771 = n9366 | n15770 ;
  assign n15772 = n14903 ^ n6540 ^ 1'b0 ;
  assign n15773 = n1199 | n4608 ;
  assign n15774 = n351 & ~n3146 ;
  assign n15775 = n1338 & ~n5977 ;
  assign n15776 = n15775 ^ n10346 ^ 1'b0 ;
  assign n15777 = n976 & ~n7680 ;
  assign n15778 = n4355 | n12610 ;
  assign n15779 = n8826 & n10322 ;
  assign n15780 = n8916 ^ n240 ^ 1'b0 ;
  assign n15781 = n4138 & n15780 ;
  assign n15782 = ~n9718 & n15781 ;
  assign n15783 = n4438 | n12129 ;
  assign n15784 = n15782 | n15783 ;
  assign n15786 = n6714 & n8012 ;
  assign n15787 = n15786 ^ n773 ^ 1'b0 ;
  assign n15785 = n2701 ^ n1867 ^ 1'b0 ;
  assign n15788 = n15787 ^ n15785 ^ n11978 ;
  assign n15789 = ~n2213 & n2723 ;
  assign n15790 = n15789 ^ x116 ^ 1'b0 ;
  assign n15791 = n3988 & ~n15790 ;
  assign n15792 = n4703 & n11759 ;
  assign n15793 = n15792 ^ n7695 ^ 1'b0 ;
  assign n15794 = n4379 | n15793 ;
  assign n15795 = n15794 ^ n5347 ^ 1'b0 ;
  assign n15796 = n3091 & ~n15795 ;
  assign n15797 = ~n13273 & n15796 ;
  assign n15798 = n2447 & ~n5599 ;
  assign n15799 = n15798 ^ n12758 ^ 1'b0 ;
  assign n15800 = ( n671 & ~n1537 ) | ( n671 & n1743 ) | ( ~n1537 & n1743 ) ;
  assign n15801 = n6652 & n15800 ;
  assign n15802 = n7008 & n15801 ;
  assign n15803 = n2886 & ~n15802 ;
  assign n15804 = n15803 ^ n13106 ^ 1'b0 ;
  assign n15805 = n14479 & n15804 ;
  assign n15806 = ~n15799 & n15805 ;
  assign n15807 = n2610 ^ n1977 ^ n1602 ;
  assign n15808 = ~n2697 & n15807 ;
  assign n15809 = ~n3986 & n15808 ;
  assign n15810 = n14390 ^ n591 ^ 1'b0 ;
  assign n15811 = n15809 | n15810 ;
  assign n15812 = n1005 & ~n3823 ;
  assign n15813 = ( n8910 & ~n15811 ) | ( n8910 & n15812 ) | ( ~n15811 & n15812 ) ;
  assign n15814 = n9653 & n14832 ;
  assign n15815 = n9805 ^ n4450 ^ n2802 ;
  assign n15816 = n2948 | n6476 ;
  assign n15817 = n15815 & ~n15816 ;
  assign n15818 = n293 | n1172 ;
  assign n15819 = n15818 ^ n2049 ^ 1'b0 ;
  assign n15820 = n8391 & ~n15819 ;
  assign n15821 = ~n4861 & n9495 ;
  assign n15822 = n12817 ^ n2477 ^ 1'b0 ;
  assign n15823 = n4044 | n4853 ;
  assign n15824 = n1497 & ~n15823 ;
  assign n15825 = n15824 ^ n9396 ^ 1'b0 ;
  assign n15826 = n3147 ^ n795 ^ 1'b0 ;
  assign n15827 = n5362 & ~n15826 ;
  assign n15828 = n2589 & n15827 ;
  assign n15830 = n12790 ^ n3240 ^ n1130 ;
  assign n15829 = ~n10067 & n12223 ;
  assign n15831 = n15830 ^ n15829 ^ 1'b0 ;
  assign n15832 = n1861 | n13886 ;
  assign n15833 = n7090 & ~n15832 ;
  assign n15834 = ~n351 & n4934 ;
  assign n15835 = n15834 ^ n8043 ^ 1'b0 ;
  assign n15836 = n15210 & n15835 ;
  assign n15837 = n12226 & n15836 ;
  assign n15838 = ~n699 & n2470 ;
  assign n15839 = n15837 & n15838 ;
  assign n15840 = n3746 & n4548 ;
  assign n15841 = n15840 ^ n3313 ^ 1'b0 ;
  assign n15842 = n11506 ^ n2289 ^ 1'b0 ;
  assign n15843 = ~n2349 & n15842 ;
  assign n15844 = n4094 & n7797 ;
  assign n15845 = ( n309 & n15843 ) | ( n309 & n15844 ) | ( n15843 & n15844 ) ;
  assign n15846 = n177 | n11378 ;
  assign n15847 = n15846 ^ n12642 ^ 1'b0 ;
  assign n15851 = n395 | n4909 ;
  assign n15852 = n2725 | n15851 ;
  assign n15848 = n556 & ~n3200 ;
  assign n15849 = n15848 ^ n9824 ^ 1'b0 ;
  assign n15850 = x69 & ~n15849 ;
  assign n15853 = n15852 ^ n15850 ^ 1'b0 ;
  assign n15854 = n2730 & ~n8590 ;
  assign n15855 = n5676 & n10475 ;
  assign n15856 = ~n5676 & n15855 ;
  assign n15857 = n15854 & ~n15856 ;
  assign n15858 = ~n15854 & n15857 ;
  assign n15859 = n7241 ^ n1606 ^ 1'b0 ;
  assign n15860 = n4558 & ~n15859 ;
  assign n15861 = ~n363 & n15860 ;
  assign n15862 = ~n4126 & n15861 ;
  assign n15863 = n9639 ^ n2785 ^ 1'b0 ;
  assign n15864 = ( n6799 & n10352 ) | ( n6799 & ~n15863 ) | ( n10352 & ~n15863 ) ;
  assign n15865 = n4342 & ~n11531 ;
  assign n15866 = n6340 & n11122 ;
  assign n15867 = ~n12552 & n15866 ;
  assign n15868 = ~n11705 & n15867 ;
  assign n15869 = n1495 | n15868 ;
  assign n15870 = n6054 ^ n4450 ^ 1'b0 ;
  assign n15871 = n2403 ^ n1454 ^ 1'b0 ;
  assign n15872 = n468 & ~n15871 ;
  assign n15873 = n995 & n15872 ;
  assign n15874 = ~n821 & n4036 ;
  assign n15875 = n675 & ~n3162 ;
  assign n15876 = ~n15874 & n15875 ;
  assign n15877 = n7854 & ~n9176 ;
  assign n15878 = ~n8352 & n15877 ;
  assign n15879 = n15564 ^ n1523 ^ 1'b0 ;
  assign n15880 = ~n15878 & n15879 ;
  assign n15881 = n11529 ^ n10014 ^ 1'b0 ;
  assign n15882 = n8099 ^ n4247 ^ 1'b0 ;
  assign n15883 = n12347 & n15882 ;
  assign n15884 = ( n4408 & ~n12494 ) | ( n4408 & n15883 ) | ( ~n12494 & n15883 ) ;
  assign n15885 = ( ~n593 & n3846 ) | ( ~n593 & n5350 ) | ( n3846 & n5350 ) ;
  assign n15886 = n12728 ^ n3156 ^ 1'b0 ;
  assign n15887 = n15886 ^ n12238 ^ 1'b0 ;
  assign n15888 = n5034 & n14511 ;
  assign n15889 = n3378 | n12753 ;
  assign n15890 = n3530 & ~n6301 ;
  assign n15891 = n11640 & ~n14813 ;
  assign n15898 = ( n240 & ~n241 ) | ( n240 & n252 ) | ( ~n241 & n252 ) ;
  assign n15899 = n14137 & ~n15898 ;
  assign n15895 = ~n12714 & n14585 ;
  assign n15896 = ~n200 & n15895 ;
  assign n15892 = n2438 & n3816 ;
  assign n15893 = ~n4073 & n15892 ;
  assign n15894 = n3870 | n15893 ;
  assign n15897 = n15896 ^ n15894 ^ 1'b0 ;
  assign n15900 = n15899 ^ n15897 ^ 1'b0 ;
  assign n15901 = n10990 ^ n7157 ^ 1'b0 ;
  assign n15903 = n5916 ^ n1873 ^ 1'b0 ;
  assign n15904 = n2546 & n15903 ;
  assign n15905 = ~n14742 & n15904 ;
  assign n15902 = n3687 | n10278 ;
  assign n15906 = n15905 ^ n15902 ^ 1'b0 ;
  assign n15907 = ~n15901 & n15906 ;
  assign n15908 = n1068 & n2611 ;
  assign n15909 = ~n7164 & n9132 ;
  assign n15910 = n15445 & ~n15909 ;
  assign n15913 = n7206 | n8503 ;
  assign n15914 = n14382 & ~n15913 ;
  assign n15911 = n7925 ^ n4601 ^ 1'b0 ;
  assign n15912 = ~n1556 & n15911 ;
  assign n15915 = n15914 ^ n15912 ^ n2297 ;
  assign n15916 = n9872 & n11690 ;
  assign n15917 = n3059 & ~n14123 ;
  assign n15918 = n7844 ^ n5092 ^ 1'b0 ;
  assign n15919 = n15917 & ~n15918 ;
  assign n15920 = ~n1012 & n2835 ;
  assign n15921 = n964 | n15920 ;
  assign n15922 = n10801 | n15921 ;
  assign n15923 = n279 & ~n8950 ;
  assign n15924 = n15923 ^ n1745 ^ 1'b0 ;
  assign n15925 = n2745 & n3761 ;
  assign n15926 = ~n13633 & n15925 ;
  assign n15927 = ~n15585 & n15926 ;
  assign n15928 = n7043 & ~n8895 ;
  assign n15929 = n1948 & ~n2053 ;
  assign n15930 = n15929 ^ n1270 ^ 1'b0 ;
  assign n15931 = n13497 ^ n5277 ^ n2328 ;
  assign n15932 = n358 | n2619 ;
  assign n15933 = n15932 ^ n9013 ^ 1'b0 ;
  assign n15934 = n15933 ^ n7820 ^ 1'b0 ;
  assign n15935 = n4027 ^ n3331 ^ 1'b0 ;
  assign n15936 = n1623 | n6220 ;
  assign n15937 = ~n1906 & n15936 ;
  assign n15938 = n15935 & n15937 ;
  assign n15939 = n4739 & n13477 ;
  assign n15940 = n15939 ^ n13013 ^ 1'b0 ;
  assign n15942 = ( n904 & n5472 ) | ( n904 & ~n8816 ) | ( n5472 & ~n8816 ) ;
  assign n15941 = ~n2717 & n3790 ;
  assign n15943 = n15942 ^ n15941 ^ 1'b0 ;
  assign n15944 = n14002 | n15943 ;
  assign n15945 = ~n5519 & n6730 ;
  assign n15946 = n15945 ^ n15893 ^ 1'b0 ;
  assign n15947 = ~n842 & n15946 ;
  assign n15948 = n3974 | n13393 ;
  assign n15949 = n12197 ^ n10569 ^ n8198 ;
  assign n15950 = ~n3354 & n15949 ;
  assign n15951 = n1046 & ~n13263 ;
  assign n15952 = n12664 & n13601 ;
  assign n15953 = n15952 ^ n10339 ^ 1'b0 ;
  assign n15954 = n3376 & ~n6991 ;
  assign n15955 = n8240 & ~n9330 ;
  assign n15956 = ~n4316 & n15903 ;
  assign n15957 = n9978 & n15956 ;
  assign n15958 = n5971 ^ n4592 ^ 1'b0 ;
  assign n15959 = ~n12239 & n13701 ;
  assign n15970 = ~n175 & n12164 ;
  assign n15960 = ~n6009 & n11904 ;
  assign n15961 = n2371 & n15960 ;
  assign n15962 = n279 | n3086 ;
  assign n15963 = n15962 ^ n6526 ^ 1'b0 ;
  assign n15964 = n8170 & ~n15963 ;
  assign n15965 = ~n1469 & n15964 ;
  assign n15966 = n256 & n15965 ;
  assign n15967 = n11292 | n15966 ;
  assign n15968 = n15961 & ~n15967 ;
  assign n15969 = n14869 & ~n15968 ;
  assign n15971 = n15970 ^ n15969 ^ 1'b0 ;
  assign n15972 = n1907 & n7238 ;
  assign n15973 = n6385 | n14372 ;
  assign n15974 = n15973 ^ n1027 ^ 1'b0 ;
  assign n15975 = n10944 & n14236 ;
  assign n15976 = n15974 & n15975 ;
  assign n15977 = n1079 | n8164 ;
  assign n15978 = n6060 | n15977 ;
  assign n15979 = n1201 & n15978 ;
  assign n15980 = ~n2508 & n14128 ;
  assign n15981 = ~n11600 & n15980 ;
  assign n15982 = n2445 & n14345 ;
  assign n15983 = n7050 & ~n15867 ;
  assign n15984 = n11225 ^ x28 ^ 1'b0 ;
  assign n15985 = n2924 & n3099 ;
  assign n15986 = ~n673 & n15985 ;
  assign n15987 = n1535 & n8543 ;
  assign n15988 = n15987 ^ n6449 ^ n611 ;
  assign n15989 = n12235 | n15988 ;
  assign n15990 = n6608 & n15989 ;
  assign n15991 = n240 & n15990 ;
  assign n15992 = ~n1337 & n10429 ;
  assign n15993 = n15992 ^ n8206 ^ 1'b0 ;
  assign n15994 = n15993 ^ n2670 ^ 1'b0 ;
  assign n15995 = ( ~n331 & n2502 ) | ( ~n331 & n2927 ) | ( n2502 & n2927 ) ;
  assign n15996 = n7767 & ~n13025 ;
  assign n15997 = ~n8736 & n15996 ;
  assign n15998 = ~n15995 & n15997 ;
  assign n15999 = n6263 ^ n2471 ^ n2380 ;
  assign n16000 = n5245 | n8803 ;
  assign n16001 = n12597 & ~n16000 ;
  assign n16002 = n7837 & n16001 ;
  assign n16003 = n16002 ^ n5179 ^ 1'b0 ;
  assign n16004 = n6472 ^ n3321 ^ 1'b0 ;
  assign n16005 = n10453 | n15378 ;
  assign n16006 = n2222 | n16005 ;
  assign n16007 = n15017 ^ n1572 ^ 1'b0 ;
  assign n16009 = n2953 & ~n5355 ;
  assign n16010 = n16009 ^ n4002 ^ 1'b0 ;
  assign n16011 = n11351 & ~n16010 ;
  assign n16008 = n471 & ~n5082 ;
  assign n16012 = n16011 ^ n16008 ^ 1'b0 ;
  assign n16013 = n513 & n13330 ;
  assign n16014 = n6715 ^ n971 ^ 1'b0 ;
  assign n16015 = n7711 ^ n4315 ^ 1'b0 ;
  assign n16016 = ~n16014 & n16015 ;
  assign n16017 = n7445 & n16016 ;
  assign n16018 = ( n7544 & n16013 ) | ( n7544 & n16017 ) | ( n16013 & n16017 ) ;
  assign n16019 = n8520 ^ n4426 ^ 1'b0 ;
  assign n16020 = n5539 & ~n16019 ;
  assign n16021 = n16020 ^ n1308 ^ 1'b0 ;
  assign n16022 = n1163 & n16021 ;
  assign n16023 = n2910 & ~n13138 ;
  assign n16024 = n3073 & ~n6545 ;
  assign n16025 = n2942 | n16024 ;
  assign n16026 = n1735 | n16025 ;
  assign n16029 = x25 & n8942 ;
  assign n16030 = ~n5569 & n16029 ;
  assign n16031 = ( ~n2665 & n4187 ) | ( ~n2665 & n16030 ) | ( n4187 & n16030 ) ;
  assign n16032 = n16031 ^ n3255 ^ 1'b0 ;
  assign n16033 = n5742 & n16032 ;
  assign n16034 = n16033 ^ n4200 ^ 1'b0 ;
  assign n16035 = n16034 ^ n5969 ^ 1'b0 ;
  assign n16027 = n2557 | n8887 ;
  assign n16028 = n15662 & ~n16027 ;
  assign n16036 = n16035 ^ n16028 ^ n9266 ;
  assign n16037 = n16036 ^ n2806 ^ 1'b0 ;
  assign n16038 = n16037 ^ n14142 ^ 1'b0 ;
  assign n16039 = n14549 | n16038 ;
  assign n16040 = n2067 & ~n12877 ;
  assign n16042 = n14339 ^ n6734 ^ 1'b0 ;
  assign n16043 = n6990 & n16042 ;
  assign n16041 = ~n765 & n2409 ;
  assign n16044 = n16043 ^ n16041 ^ 1'b0 ;
  assign n16045 = n799 & ~n4403 ;
  assign n16046 = n16045 ^ n5355 ^ 1'b0 ;
  assign n16047 = n3295 | n6948 ;
  assign n16048 = n16047 ^ n745 ^ 1'b0 ;
  assign n16049 = n2979 ^ n531 ^ 1'b0 ;
  assign n16050 = n6584 | n16049 ;
  assign n16051 = n16048 & ~n16050 ;
  assign n16052 = n15404 & ~n16051 ;
  assign n16053 = n6339 & n16052 ;
  assign n16054 = n15552 ^ n3601 ^ 1'b0 ;
  assign n16055 = n5440 | n9469 ;
  assign n16056 = n16055 ^ n675 ^ 1'b0 ;
  assign n16057 = n8295 & ~n16056 ;
  assign n16058 = ~n7971 & n8249 ;
  assign n16059 = n16058 ^ n6148 ^ 1'b0 ;
  assign n16062 = n10281 ^ n548 ^ 1'b0 ;
  assign n16063 = n8007 | n16062 ;
  assign n16064 = n2486 & ~n16063 ;
  assign n16060 = n2327 & ~n3402 ;
  assign n16061 = n14406 & n16060 ;
  assign n16065 = n16064 ^ n16061 ^ 1'b0 ;
  assign n16066 = ~n896 & n10123 ;
  assign n16067 = n16066 ^ n2503 ^ 1'b0 ;
  assign n16068 = n2438 & ~n16067 ;
  assign n16069 = n7170 & n16068 ;
  assign n16070 = n3762 | n7678 ;
  assign n16071 = n709 & n16070 ;
  assign n16072 = n6550 ^ n3944 ^ 1'b0 ;
  assign n16073 = ~n2483 & n16001 ;
  assign n16074 = n16073 ^ n13654 ^ 1'b0 ;
  assign n16075 = n3336 | n7524 ;
  assign n16076 = n16075 ^ n8849 ^ 1'b0 ;
  assign n16077 = n450 | n9051 ;
  assign n16078 = n11561 ^ n8606 ^ 1'b0 ;
  assign n16080 = n4183 | n11609 ;
  assign n16081 = n11609 & ~n16080 ;
  assign n16079 = n1166 | n7178 ;
  assign n16082 = n16081 ^ n16079 ^ 1'b0 ;
  assign n16083 = n5281 & n6421 ;
  assign n16084 = n12627 ^ n5608 ^ 1'b0 ;
  assign n16085 = ~n2341 & n12168 ;
  assign n16086 = ~n4696 & n16085 ;
  assign n16087 = n16086 ^ n4555 ^ 1'b0 ;
  assign n16088 = n6309 & n7237 ;
  assign n16089 = ~n7964 & n16088 ;
  assign n16090 = n16089 ^ n15581 ^ 1'b0 ;
  assign n16091 = n3097 & ~n16090 ;
  assign n16092 = n16091 ^ n1560 ^ 1'b0 ;
  assign n16093 = n14341 ^ n11923 ^ n6988 ;
  assign n16094 = n2938 ^ n442 ^ 1'b0 ;
  assign n16095 = n3749 & n16094 ;
  assign n16096 = n1912 & ~n10894 ;
  assign n16097 = n16096 ^ n13713 ^ 1'b0 ;
  assign n16098 = n2281 & ~n16097 ;
  assign n16099 = n16095 & ~n16098 ;
  assign n16100 = n2699 & ~n2996 ;
  assign n16101 = n15557 & ~n16100 ;
  assign n16102 = n16101 ^ n4411 ^ 1'b0 ;
  assign n16103 = n6029 & ~n6327 ;
  assign n16104 = ~n7300 & n16103 ;
  assign n16105 = n1527 | n9011 ;
  assign n16106 = n14557 & n16105 ;
  assign n16107 = ~n6591 & n16035 ;
  assign n16108 = n10761 ^ n5370 ^ 1'b0 ;
  assign n16109 = ~n6760 & n10880 ;
  assign n16110 = n16109 ^ x69 ^ 1'b0 ;
  assign n16111 = n16108 | n16110 ;
  assign n16112 = n2621 & ~n16111 ;
  assign n16113 = n4630 ^ n778 ^ x62 ;
  assign n16114 = n4389 ^ n3340 ^ 1'b0 ;
  assign n16115 = n11366 & n16114 ;
  assign n16116 = n13348 ^ n6469 ^ 1'b0 ;
  assign n16117 = n1914 ^ x110 ^ 1'b0 ;
  assign n16118 = n5537 | n16117 ;
  assign n16119 = n3477 & ~n14643 ;
  assign n16120 = n16119 ^ n2442 ^ 1'b0 ;
  assign n16121 = n16120 ^ n3431 ^ 1'b0 ;
  assign n16122 = n496 | n6916 ;
  assign n16123 = n16121 | n16122 ;
  assign n16124 = n12226 ^ n4430 ^ 1'b0 ;
  assign n16125 = x23 & ~n16124 ;
  assign n16127 = n8921 & ~n12135 ;
  assign n16128 = n16127 ^ n7977 ^ 1'b0 ;
  assign n16126 = ~n2138 & n5410 ;
  assign n16129 = n16128 ^ n16126 ^ 1'b0 ;
  assign n16130 = n7321 & ~n11378 ;
  assign n16131 = n4115 & ~n5227 ;
  assign n16132 = n1681 | n16131 ;
  assign n16133 = n7577 ^ n3691 ^ n1450 ;
  assign n16134 = ( ~n905 & n5948 ) | ( ~n905 & n16133 ) | ( n5948 & n16133 ) ;
  assign n16135 = n16134 ^ n4152 ^ 1'b0 ;
  assign n16136 = n15338 ^ n9764 ^ n9211 ;
  assign n16137 = n2103 & n5319 ;
  assign n16138 = ~n3648 & n16137 ;
  assign n16139 = n8008 | n16138 ;
  assign n16140 = n16136 & ~n16139 ;
  assign n16141 = n10512 ^ n10133 ^ 1'b0 ;
  assign n16142 = n2581 | n16141 ;
  assign n16143 = n1003 & n2451 ;
  assign n16144 = n16143 ^ n3403 ^ 1'b0 ;
  assign n16145 = n5052 & ~n13379 ;
  assign n16146 = ~n16144 & n16145 ;
  assign n16147 = n1570 & n15928 ;
  assign n16148 = n8077 ^ n3691 ^ 1'b0 ;
  assign n16149 = n4289 & ~n4658 ;
  assign n16150 = n2935 & n16149 ;
  assign n16151 = n16150 ^ n256 ^ 1'b0 ;
  assign n16152 = n1372 & n16151 ;
  assign n16153 = n16148 | n16152 ;
  assign n16154 = n2738 & n6403 ;
  assign n16155 = n7645 | n10008 ;
  assign n16156 = n16155 ^ n10459 ^ 1'b0 ;
  assign n16157 = n5973 ^ n3491 ^ 1'b0 ;
  assign n16158 = n11859 & ~n11883 ;
  assign n16159 = n8787 ^ n1700 ^ 1'b0 ;
  assign n16160 = n3455 & n16159 ;
  assign n16161 = x50 | n11872 ;
  assign n16162 = n16161 ^ n10526 ^ 1'b0 ;
  assign n16163 = n10960 ^ n3858 ^ 1'b0 ;
  assign n16164 = ~n3441 & n16163 ;
  assign n16165 = n13734 ^ n11868 ^ 1'b0 ;
  assign n16166 = ~n2189 & n4623 ;
  assign n16167 = ~n16165 & n16166 ;
  assign n16168 = ~n6403 & n16167 ;
  assign n16169 = n651 & n2233 ;
  assign n16170 = n6785 | n16169 ;
  assign n16171 = n14939 ^ n2822 ^ 1'b0 ;
  assign n16172 = ( x107 & n897 ) | ( x107 & ~n11948 ) | ( n897 & ~n11948 ) ;
  assign n16173 = ~n4073 & n16172 ;
  assign n16174 = ~n9392 & n16173 ;
  assign n16175 = ~n5928 & n15818 ;
  assign n16176 = ~n11889 & n16175 ;
  assign n16177 = n15598 ^ n9279 ^ 1'b0 ;
  assign n16182 = n8840 ^ n6159 ^ 1'b0 ;
  assign n16183 = n2796 & ~n16182 ;
  assign n16181 = n694 | n2014 ;
  assign n16178 = ~n499 & n1552 ;
  assign n16179 = n16178 ^ n8184 ^ 1'b0 ;
  assign n16180 = n16179 ^ n3641 ^ 1'b0 ;
  assign n16184 = n16183 ^ n16181 ^ n16180 ;
  assign n16185 = n1261 & n1385 ;
  assign n16186 = n8823 ^ n3461 ^ 1'b0 ;
  assign n16187 = ~n16185 & n16186 ;
  assign n16188 = ( n2270 & ~n2816 ) | ( n2270 & n5249 ) | ( ~n2816 & n5249 ) ;
  assign n16189 = n10755 ^ n386 ^ 1'b0 ;
  assign n16190 = ~n7346 & n16189 ;
  assign n16191 = n16188 & n16190 ;
  assign n16192 = n16191 ^ n8422 ^ 1'b0 ;
  assign n16193 = n7575 ^ n4068 ^ 1'b0 ;
  assign n16194 = n16192 | n16193 ;
  assign n16195 = n5681 & ~n10463 ;
  assign n16196 = n351 | n16195 ;
  assign n16197 = n16196 ^ n15818 ^ 1'b0 ;
  assign n16198 = n3382 | n4966 ;
  assign n16199 = n12809 ^ n881 ^ 1'b0 ;
  assign n16200 = n2752 & ~n13670 ;
  assign n16201 = n6776 & ~n14418 ;
  assign n16202 = n6273 & n11729 ;
  assign n16203 = ~n9322 & n16202 ;
  assign n16204 = ~n13636 & n16203 ;
  assign n16205 = n4726 ^ n3799 ^ 1'b0 ;
  assign n16206 = n5909 & n16205 ;
  assign n16207 = n13177 | n16206 ;
  assign n16208 = n5431 | n16207 ;
  assign n16209 = n3282 | n15928 ;
  assign n16210 = n16209 ^ n8776 ^ 1'b0 ;
  assign n16211 = n2192 | n12278 ;
  assign n16212 = n7103 & n10260 ;
  assign n16213 = ~n506 & n9236 ;
  assign n16214 = n1512 & ~n13754 ;
  assign n16215 = n16214 ^ n10761 ^ n10087 ;
  assign n16216 = n4408 | n5347 ;
  assign n16217 = n8249 | n16216 ;
  assign n16218 = n14511 | n16217 ;
  assign n16219 = n4204 ^ n1421 ^ 1'b0 ;
  assign n16220 = n13775 ^ n1738 ^ 1'b0 ;
  assign n16221 = ~n10468 & n16220 ;
  assign n16222 = n2426 & n3105 ;
  assign n16223 = n2053 & ~n11103 ;
  assign n16224 = n16222 & n16223 ;
  assign n16225 = ~n4162 & n16224 ;
  assign n16226 = n9650 & ~n15286 ;
  assign n16227 = n16226 ^ n143 ^ 1'b0 ;
  assign n16228 = x23 & n4940 ;
  assign n16229 = n2875 & ~n5634 ;
  assign n16230 = n16229 ^ n3370 ^ 1'b0 ;
  assign n16231 = n16230 ^ n1682 ^ 1'b0 ;
  assign n16232 = n660 & ~n4969 ;
  assign n16233 = ~n16231 & n16232 ;
  assign n16234 = ( ~n1959 & n2758 ) | ( ~n1959 & n3806 ) | ( n2758 & n3806 ) ;
  assign n16235 = n16234 ^ n3557 ^ 1'b0 ;
  assign n16236 = n3899 | n16235 ;
  assign n16237 = ~n3143 & n5592 ;
  assign n16238 = n4863 & n10321 ;
  assign n16239 = n13619 ^ n1258 ^ 1'b0 ;
  assign n16240 = n1713 & n16239 ;
  assign n16241 = ~n896 & n16240 ;
  assign n16242 = n16241 ^ n5574 ^ 1'b0 ;
  assign n16243 = n4182 & n6412 ;
  assign n16244 = ( n6970 & n8838 ) | ( n6970 & ~n15489 ) | ( n8838 & ~n15489 ) ;
  assign n16245 = n8581 ^ n7948 ^ 1'b0 ;
  assign n16246 = n692 & n7766 ;
  assign n16247 = n16246 ^ n8323 ^ 1'b0 ;
  assign n16248 = n8244 | n11818 ;
  assign n16249 = n16248 ^ n4657 ^ 1'b0 ;
  assign n16250 = n2986 & ~n16249 ;
  assign n16251 = n16250 ^ n2317 ^ 1'b0 ;
  assign n16252 = ~n2038 & n2810 ;
  assign n16253 = n4380 & n5557 ;
  assign n16254 = n16253 ^ n13798 ^ 1'b0 ;
  assign n16255 = n4531 | n16254 ;
  assign n16256 = n13147 ^ n12721 ^ 1'b0 ;
  assign n16257 = ~n9837 & n10547 ;
  assign n16258 = n16257 ^ n5927 ^ 1'b0 ;
  assign n16259 = n7252 ^ n2418 ^ 1'b0 ;
  assign n16260 = n9792 & ~n16259 ;
  assign n16261 = n14204 ^ n361 ^ 1'b0 ;
  assign n16262 = n13471 ^ n5953 ^ 1'b0 ;
  assign n16263 = ~n3350 & n4697 ;
  assign n16264 = ~n4766 & n16263 ;
  assign n16265 = ( n15452 & ~n16262 ) | ( n15452 & n16264 ) | ( ~n16262 & n16264 ) ;
  assign n16266 = n16150 ^ n4733 ^ 1'b0 ;
  assign n16267 = n12145 & n16266 ;
  assign n16268 = n1200 & n10499 ;
  assign n16269 = ~n16267 & n16268 ;
  assign n16270 = n13098 & n16269 ;
  assign n16271 = ( n2012 & n2153 ) | ( n2012 & n3641 ) | ( n2153 & n3641 ) ;
  assign n16272 = n16271 ^ n7305 ^ 1'b0 ;
  assign n16273 = n8723 | n12780 ;
  assign n16274 = n16273 ^ n4507 ^ 1'b0 ;
  assign n16275 = n13990 & ~n16274 ;
  assign n16276 = n4315 ^ n556 ^ 1'b0 ;
  assign n16277 = n2196 & n16276 ;
  assign n16278 = ~n15409 & n16277 ;
  assign n16279 = n11380 ^ n3533 ^ 1'b0 ;
  assign n16280 = n4759 & n16279 ;
  assign n16281 = n2501 & n13047 ;
  assign n16282 = n16281 ^ n10740 ^ 1'b0 ;
  assign n16283 = n10149 ^ n3543 ^ 1'b0 ;
  assign n16284 = n14819 ^ n1884 ^ n1176 ;
  assign n16285 = ~n16283 & n16284 ;
  assign n16286 = n8630 ^ n5889 ^ n1277 ;
  assign n16287 = n6811 & n6933 ;
  assign n16288 = n4960 | n16287 ;
  assign n16289 = n16286 | n16288 ;
  assign n16290 = n2346 | n11378 ;
  assign n16291 = n5756 & n16290 ;
  assign n16292 = n1239 & ~n10703 ;
  assign n16293 = n16291 & n16292 ;
  assign n16294 = ( x65 & n6017 ) | ( x65 & n6101 ) | ( n6017 & n6101 ) ;
  assign n16295 = n7662 ^ n2827 ^ 1'b0 ;
  assign n16296 = ~n14418 & n16295 ;
  assign n16297 = n16296 ^ n3029 ^ 1'b0 ;
  assign n16298 = n598 | n16297 ;
  assign n16299 = n14270 & ~n16298 ;
  assign n16300 = ~n14641 & n16299 ;
  assign n16301 = ~n6721 & n9408 ;
  assign n16302 = n9097 ^ n8233 ^ n4100 ;
  assign n16303 = n8352 ^ n8247 ^ 1'b0 ;
  assign n16304 = n1077 | n16303 ;
  assign n16305 = n9407 & ~n16304 ;
  assign n16306 = n2859 & n16305 ;
  assign n16307 = n2249 | n5638 ;
  assign n16308 = n6202 & ~n10763 ;
  assign n16309 = n3764 & n16308 ;
  assign n16310 = n722 & n2021 ;
  assign n16311 = n1623 & n10692 ;
  assign n16312 = n8559 ^ n4729 ^ 1'b0 ;
  assign n16316 = n4881 & ~n5206 ;
  assign n16317 = n16316 ^ n3413 ^ 1'b0 ;
  assign n16313 = ~n3764 & n5319 ;
  assign n16314 = n3251 & n16313 ;
  assign n16315 = n16314 ^ n3240 ^ 1'b0 ;
  assign n16318 = n16317 ^ n16315 ^ n3666 ;
  assign n16319 = n3968 & ~n13599 ;
  assign n16320 = n16319 ^ n5575 ^ 1'b0 ;
  assign n16321 = n1817 & ~n5379 ;
  assign n16322 = n16321 ^ n2948 ^ 1'b0 ;
  assign n16326 = n6746 | n8577 ;
  assign n16327 = n8577 & ~n16326 ;
  assign n16324 = n6323 ^ n2805 ^ 1'b0 ;
  assign n16325 = n3993 | n16324 ;
  assign n16323 = n9473 & n16095 ;
  assign n16328 = n16327 ^ n16325 ^ n16323 ;
  assign n16329 = ~n11333 & n16328 ;
  assign n16330 = n613 & ~n4019 ;
  assign n16331 = n16330 ^ n3888 ^ 1'b0 ;
  assign n16332 = n16331 ^ n10035 ^ 1'b0 ;
  assign n16333 = ~n14081 & n16332 ;
  assign n16334 = n16333 ^ n3729 ^ 1'b0 ;
  assign n16335 = n3085 & n16334 ;
  assign n16337 = n4029 & n11092 ;
  assign n16336 = n5692 & n7529 ;
  assign n16338 = n16337 ^ n16336 ^ 1'b0 ;
  assign n16342 = n4071 | n7360 ;
  assign n16343 = n6800 | n16342 ;
  assign n16339 = n5055 ^ n4467 ^ 1'b0 ;
  assign n16340 = n4319 | n7612 ;
  assign n16341 = n16339 & n16340 ;
  assign n16344 = n16343 ^ n16341 ^ 1'b0 ;
  assign n16345 = n476 | n16344 ;
  assign n16346 = n16345 ^ n1893 ^ 1'b0 ;
  assign n16347 = n8940 ^ n2036 ^ 1'b0 ;
  assign n16348 = n13936 ^ n4107 ^ 1'b0 ;
  assign n16349 = n4322 & n16348 ;
  assign n16350 = n5016 ^ n2370 ^ 1'b0 ;
  assign n16351 = n13431 ^ n4542 ^ 1'b0 ;
  assign n16352 = n5951 & n16351 ;
  assign n16353 = n1823 & ~n12740 ;
  assign n16354 = n8496 | n8946 ;
  assign n16355 = n13398 ^ n11123 ^ 1'b0 ;
  assign n16356 = n16354 & n16355 ;
  assign n16357 = n4623 ^ n4293 ^ n3709 ;
  assign n16358 = n1263 | n16357 ;
  assign n16359 = n16358 ^ n3321 ^ 1'b0 ;
  assign n16360 = n16359 ^ n8847 ^ 1'b0 ;
  assign n16361 = n7426 | n9376 ;
  assign n16362 = n4726 & ~n8341 ;
  assign n16363 = n9996 ^ n6187 ^ 1'b0 ;
  assign n16364 = n8282 & n16363 ;
  assign n16365 = n1256 & n16364 ;
  assign n16366 = n16362 & n16365 ;
  assign n16367 = n9522 ^ n8509 ^ 1'b0 ;
  assign n16368 = n12315 ^ n1241 ^ 1'b0 ;
  assign n16369 = n13950 ^ n5739 ^ 1'b0 ;
  assign n16370 = n477 & ~n2931 ;
  assign n16371 = n14229 & n16108 ;
  assign n16372 = n1483 & ~n15561 ;
  assign n16373 = n4918 ^ n3618 ^ 1'b0 ;
  assign n16374 = n4918 & ~n10640 ;
  assign n16375 = n16374 ^ n14312 ^ 1'b0 ;
  assign n16376 = n851 | n11242 ;
  assign n16377 = n8006 & ~n16376 ;
  assign n16378 = n16377 ^ n7839 ^ 1'b0 ;
  assign n16379 = ~n14326 & n15196 ;
  assign n16380 = n3342 & ~n4715 ;
  assign n16381 = n16380 ^ n147 ^ 1'b0 ;
  assign n16382 = n15912 ^ n10244 ^ 1'b0 ;
  assign n16383 = n11320 ^ n1212 ^ 1'b0 ;
  assign n16384 = n258 & n16383 ;
  assign n16385 = n16384 ^ n1005 ^ n666 ;
  assign n16386 = n13539 ^ n362 ^ 1'b0 ;
  assign n16387 = n4354 | n5124 ;
  assign n16388 = n16387 ^ n4329 ^ 1'b0 ;
  assign n16389 = n7737 & ~n9638 ;
  assign n16390 = n15164 & n16389 ;
  assign n16391 = n14303 ^ n11987 ^ n10356 ;
  assign n16392 = n9001 | n11357 ;
  assign n16393 = n7500 ^ n5897 ^ 1'b0 ;
  assign n16394 = n1283 & ~n11287 ;
  assign n16395 = ~n2374 & n2946 ;
  assign n16396 = n16395 ^ n15603 ^ 1'b0 ;
  assign n16397 = n2044 | n16396 ;
  assign n16398 = n5327 & n16397 ;
  assign n16399 = n16398 ^ n14608 ^ 1'b0 ;
  assign n16400 = ( n3573 & n11680 ) | ( n3573 & ~n14639 ) | ( n11680 & ~n14639 ) ;
  assign n16401 = n2440 ^ n1398 ^ 1'b0 ;
  assign n16402 = ~n466 & n6843 ;
  assign n16403 = n8653 ^ n2020 ^ 1'b0 ;
  assign n16404 = n15330 & ~n16403 ;
  assign n16405 = n10270 ^ n6148 ^ 1'b0 ;
  assign n16406 = ~n6398 & n12410 ;
  assign n16407 = n2234 & ~n16406 ;
  assign n16408 = n16407 ^ n9968 ^ 1'b0 ;
  assign n16409 = n2249 & n16408 ;
  assign n16410 = n16405 & n16409 ;
  assign n16413 = n4059 | n13320 ;
  assign n16411 = n11371 ^ n5991 ^ 1'b0 ;
  assign n16412 = n10665 & n16411 ;
  assign n16414 = n16413 ^ n16412 ^ 1'b0 ;
  assign n16416 = n2826 ^ n2567 ^ 1'b0 ;
  assign n16415 = x28 & n5107 ;
  assign n16417 = n16416 ^ n16415 ^ 1'b0 ;
  assign n16418 = n15170 ^ n685 ^ 1'b0 ;
  assign n16419 = n16026 ^ n9775 ^ 1'b0 ;
  assign n16420 = n14565 ^ n137 ^ 1'b0 ;
  assign n16421 = n4434 | n7505 ;
  assign n16422 = n1599 | n16421 ;
  assign n16423 = n16422 ^ n605 ^ 1'b0 ;
  assign n16424 = n12389 ^ n8276 ^ n2050 ;
  assign n16425 = n15502 | n16424 ;
  assign n16426 = n1844 & ~n9656 ;
  assign n16427 = n16426 ^ n10701 ^ 1'b0 ;
  assign n16428 = n3319 & ~n7594 ;
  assign n16429 = ( n6839 & ~n10707 ) | ( n6839 & n16271 ) | ( ~n10707 & n16271 ) ;
  assign n16430 = n7916 ^ n6199 ^ n3174 ;
  assign n16431 = n845 | n5431 ;
  assign n16432 = n13473 & ~n16431 ;
  assign n16433 = n959 & n16432 ;
  assign n16434 = n8296 ^ n6592 ^ 1'b0 ;
  assign n16435 = n1213 | n16434 ;
  assign n16436 = n16433 & ~n16435 ;
  assign n16437 = n11019 ^ n6268 ^ 1'b0 ;
  assign n16438 = n8003 & ~n15293 ;
  assign n16439 = n9454 ^ n9338 ^ 1'b0 ;
  assign n16440 = n9651 & ~n16439 ;
  assign n16441 = n10011 ^ n9418 ^ n1263 ;
  assign n16442 = n11034 ^ n5011 ^ x47 ;
  assign n16443 = n778 & n9760 ;
  assign n16444 = n2295 | n3576 ;
  assign n16445 = n16444 ^ n7861 ^ 1'b0 ;
  assign n16446 = n2554 & n10455 ;
  assign n16447 = ~n2131 & n16446 ;
  assign n16448 = n16447 ^ n12124 ^ 1'b0 ;
  assign n16449 = ~n16445 & n16448 ;
  assign n16450 = ~n8571 & n16449 ;
  assign n16451 = n16450 ^ n713 ^ 1'b0 ;
  assign n16452 = n2722 & ~n4175 ;
  assign n16453 = n16452 ^ n13645 ^ 1'b0 ;
  assign n16454 = n3651 ^ n3474 ^ 1'b0 ;
  assign n16455 = n1578 & ~n16454 ;
  assign n16456 = n14475 ^ x110 ^ 1'b0 ;
  assign n16457 = n15812 ^ n8711 ^ 1'b0 ;
  assign n16458 = n16457 ^ n14708 ^ 1'b0 ;
  assign n16459 = n10497 & ~n16458 ;
  assign n16460 = ~n16456 & n16459 ;
  assign n16462 = n4804 ^ n2482 ^ 1'b0 ;
  assign n16463 = n879 & ~n16462 ;
  assign n16461 = ~n5891 & n9127 ;
  assign n16464 = n16463 ^ n16461 ^ 1'b0 ;
  assign n16465 = n3761 & ~n7220 ;
  assign n16466 = n2705 ^ x117 ^ 1'b0 ;
  assign n16467 = ~n999 & n16466 ;
  assign n16468 = n13046 | n16467 ;
  assign n16469 = n730 & n4514 ;
  assign n16470 = ~n6437 & n16469 ;
  assign n16471 = n1212 | n16470 ;
  assign n16472 = n16468 & ~n16471 ;
  assign n16473 = n1767 | n4357 ;
  assign n16474 = n9447 | n16473 ;
  assign n16475 = n706 & ~n11336 ;
  assign n16476 = n4013 ^ n2170 ^ 1'b0 ;
  assign n16477 = n2780 & ~n16476 ;
  assign n16478 = n8877 & n16477 ;
  assign n16479 = n16478 ^ n8314 ^ 1'b0 ;
  assign n16480 = n16479 ^ n11487 ^ 1'b0 ;
  assign n16482 = ~n2685 & n4210 ;
  assign n16483 = n16482 ^ n1100 ^ 1'b0 ;
  assign n16481 = ~n3912 & n15935 ;
  assign n16484 = n16483 ^ n16481 ^ 1'b0 ;
  assign n16485 = x94 & n729 ;
  assign n16486 = ~n7510 & n16485 ;
  assign n16487 = n12418 & n16486 ;
  assign n16488 = n7674 & ~n7960 ;
  assign n16489 = n13027 ^ n987 ^ 1'b0 ;
  assign n16490 = n11348 ^ n577 ^ 1'b0 ;
  assign n16491 = n7219 ^ n3474 ^ 1'b0 ;
  assign n16492 = n5390 & n13734 ;
  assign n16494 = ~n1209 & n9833 ;
  assign n16495 = n992 | n16494 ;
  assign n16496 = n3383 & ~n16495 ;
  assign n16497 = ~n3391 & n16496 ;
  assign n16493 = n1145 & n10482 ;
  assign n16498 = n16497 ^ n16493 ^ 1'b0 ;
  assign n16499 = n14797 ^ n12622 ^ 1'b0 ;
  assign n16500 = n4065 & ~n6620 ;
  assign n16501 = n6327 & n16500 ;
  assign n16502 = ~n3899 & n5355 ;
  assign n16503 = ~n184 & n1959 ;
  assign n16504 = ~n5775 & n16503 ;
  assign n16505 = n7951 ^ n2969 ^ 1'b0 ;
  assign n16506 = ~n16504 & n16505 ;
  assign n16507 = n7463 ^ n1416 ^ 1'b0 ;
  assign n16508 = n6038 & ~n16507 ;
  assign n16509 = n7261 & ~n13299 ;
  assign n16510 = n7783 ^ n1635 ^ 1'b0 ;
  assign n16511 = ~n13469 & n16510 ;
  assign n16512 = n16511 ^ n6698 ^ 1'b0 ;
  assign n16513 = n7942 | n16512 ;
  assign n16514 = n1204 | n16513 ;
  assign n16515 = n2176 & ~n11519 ;
  assign n16516 = n371 & ~n16376 ;
  assign n16517 = n16516 ^ n6631 ^ 1'b0 ;
  assign n16518 = n351 & n1204 ;
  assign n16519 = n5779 | n16518 ;
  assign n16520 = n3196 & n5995 ;
  assign n16521 = n16520 ^ n2386 ^ 1'b0 ;
  assign n16522 = n555 & ~n15998 ;
  assign n16523 = ( ~n2300 & n15187 ) | ( ~n2300 & n16522 ) | ( n15187 & n16522 ) ;
  assign n16524 = ~n8244 & n9193 ;
  assign n16525 = n16524 ^ n13746 ^ 1'b0 ;
  assign n16526 = n16525 ^ n7353 ^ 1'b0 ;
  assign n16527 = n8580 ^ n2739 ^ n1250 ;
  assign n16528 = n12452 & n15753 ;
  assign n16529 = n8552 & n11213 ;
  assign n16530 = n2802 & n16529 ;
  assign n16531 = n3542 ^ n2479 ^ 1'b0 ;
  assign n16532 = n2235 | n16531 ;
  assign n16533 = n16532 ^ n12882 ^ 1'b0 ;
  assign n16534 = n2116 & n4382 ;
  assign n16535 = n16534 ^ n12026 ^ 1'b0 ;
  assign n16536 = n1611 | n13236 ;
  assign n16537 = n16535 & ~n16536 ;
  assign n16538 = ~n7485 & n13187 ;
  assign n16539 = n16538 ^ n5159 ^ 1'b0 ;
  assign n16540 = n16539 ^ n1200 ^ 1'b0 ;
  assign n16541 = n5231 | n16540 ;
  assign n16542 = n5345 ^ n4056 ^ 1'b0 ;
  assign n16543 = n14486 ^ n11979 ^ n11632 ;
  assign n16544 = n3789 | n14280 ;
  assign n16545 = ~n231 & n16544 ;
  assign n16546 = n5242 ^ n5085 ^ 1'b0 ;
  assign n16547 = n12362 & ~n16546 ;
  assign n16548 = n4793 & ~n6122 ;
  assign n16549 = n16548 ^ n13735 ^ 1'b0 ;
  assign n16550 = n12031 ^ n6235 ^ 1'b0 ;
  assign n16551 = n8548 ^ n131 ^ 1'b0 ;
  assign n16552 = n722 & n16551 ;
  assign n16553 = n16148 ^ n12854 ^ 1'b0 ;
  assign n16554 = n16552 & ~n16553 ;
  assign n16555 = n9753 ^ n7281 ^ 1'b0 ;
  assign n16556 = n5889 & ~n15797 ;
  assign n16557 = n16556 ^ n6545 ^ 1'b0 ;
  assign n16558 = n6054 & ~n6135 ;
  assign n16559 = n16558 ^ n551 ^ 1'b0 ;
  assign n16560 = n16559 ^ n3811 ^ 1'b0 ;
  assign n16561 = n8346 & ~n11316 ;
  assign n16562 = ~n13186 & n16561 ;
  assign n16563 = ( n5971 & n10657 ) | ( n5971 & n14198 ) | ( n10657 & n14198 ) ;
  assign n16564 = n5445 ^ n2905 ^ 1'b0 ;
  assign n16565 = ~n9121 & n16564 ;
  assign n16566 = n16565 ^ n7429 ^ 1'b0 ;
  assign n16567 = n16566 ^ n13686 ^ 1'b0 ;
  assign n16568 = n11552 ^ n3762 ^ 1'b0 ;
  assign n16569 = n8432 ^ n5262 ^ 1'b0 ;
  assign n16570 = ~n1913 & n11034 ;
  assign n16571 = n8036 ^ n937 ^ 1'b0 ;
  assign n16572 = n16570 & ~n16571 ;
  assign n16573 = ~n3398 & n10968 ;
  assign n16574 = n15153 | n16573 ;
  assign n16575 = n16574 ^ n10216 ^ 1'b0 ;
  assign n16576 = n4006 & ~n6923 ;
  assign n16577 = ~n8960 & n16576 ;
  assign n16578 = ~n6708 & n16577 ;
  assign n16579 = n11859 ^ n1579 ^ 1'b0 ;
  assign n16580 = n7683 & ~n16579 ;
  assign n16581 = n14224 ^ n8027 ^ 1'b0 ;
  assign n16582 = n11474 & n16581 ;
  assign n16583 = n6800 ^ n4380 ^ 1'b0 ;
  assign n16589 = n15698 ^ n10700 ^ 1'b0 ;
  assign n16586 = n1219 | n4212 ;
  assign n16587 = n5533 | n16586 ;
  assign n16584 = n4098 ^ n351 ^ 1'b0 ;
  assign n16585 = n6061 & ~n16584 ;
  assign n16588 = n16587 ^ n16585 ^ n6841 ;
  assign n16590 = n16589 ^ n16588 ^ n16121 ;
  assign n16591 = n11051 & n15368 ;
  assign n16592 = n8864 & n16591 ;
  assign n16593 = n722 & ~n928 ;
  assign n16594 = n16593 ^ n9630 ^ 1'b0 ;
  assign n16595 = n3881 | n16594 ;
  assign n16596 = ~n1740 & n2271 ;
  assign n16597 = n8570 & ~n8760 ;
  assign n16598 = n16597 ^ n4875 ^ 1'b0 ;
  assign n16599 = n15202 ^ n6665 ^ 1'b0 ;
  assign n16600 = n2724 & n7300 ;
  assign n16601 = ~n16599 & n16600 ;
  assign n16602 = n12481 & n12966 ;
  assign n16603 = n3618 ^ n1070 ^ 1'b0 ;
  assign n16604 = n1811 | n12780 ;
  assign n16605 = n6153 & ~n16604 ;
  assign n16606 = ~n11353 & n16339 ;
  assign n16607 = ~n1230 & n16606 ;
  assign n16608 = n6696 ^ n3610 ^ 1'b0 ;
  assign n16609 = ~n5623 & n16608 ;
  assign n16610 = n16607 & n16609 ;
  assign n16611 = n3616 & n5492 ;
  assign n16612 = n9383 & n16611 ;
  assign n16613 = n2154 & ~n16612 ;
  assign n16614 = n15950 | n16613 ;
  assign n16615 = n13821 ^ n9865 ^ 1'b0 ;
  assign n16616 = n11908 & ~n12602 ;
  assign n16617 = ~n13099 & n16616 ;
  assign n16618 = n10803 ^ n10715 ^ n471 ;
  assign n16619 = n16618 ^ n593 ^ 1'b0 ;
  assign n16620 = n10237 & ~n16619 ;
  assign n16621 = n9322 ^ n3381 ^ 1'b0 ;
  assign n16622 = n7802 & ~n16621 ;
  assign n16623 = n7610 & ~n16622 ;
  assign n16624 = ( n7030 & n13393 ) | ( n7030 & ~n15020 ) | ( n13393 & ~n15020 ) ;
  assign n16625 = n11322 ^ n2924 ^ 1'b0 ;
  assign n16626 = n14298 | n16625 ;
  assign n16627 = n14028 & n16000 ;
  assign n16628 = n732 & ~n11544 ;
  assign n16629 = n16628 ^ n13683 ^ 1'b0 ;
  assign n16630 = n6869 & ~n7624 ;
  assign n16631 = ~x38 & n16630 ;
  assign n16632 = n3313 | n16631 ;
  assign n16633 = n16629 & ~n16632 ;
  assign n16634 = n499 | n15094 ;
  assign n16635 = n16634 ^ n2829 ^ 1'b0 ;
  assign n16636 = n11868 ^ n8841 ^ n2156 ;
  assign n16637 = n1295 & n13294 ;
  assign n16638 = n16637 ^ n15334 ^ 1'b0 ;
  assign n16639 = n5960 ^ n481 ^ 1'b0 ;
  assign n16640 = ~n7826 & n16639 ;
  assign n16641 = n15266 & n16640 ;
  assign n16642 = ~n9957 & n15550 ;
  assign n16643 = ~n10205 & n16642 ;
  assign n16644 = n4753 | n12940 ;
  assign n16645 = n7757 | n15995 ;
  assign n16646 = n16645 ^ n6188 ^ 1'b0 ;
  assign n16647 = n16646 ^ n6187 ^ 1'b0 ;
  assign n16648 = ~n5647 & n16647 ;
  assign n16649 = ~n4395 & n16648 ;
  assign n16650 = ~n2827 & n16649 ;
  assign n16651 = n1304 | n12807 ;
  assign n16652 = n16651 ^ n1596 ^ 1'b0 ;
  assign n16653 = n2849 & ~n6053 ;
  assign n16654 = n16653 ^ n4578 ^ 1'b0 ;
  assign n16655 = n16539 ^ n6574 ^ 1'b0 ;
  assign n16656 = n16654 | n16655 ;
  assign n16657 = n4113 | n11274 ;
  assign n16658 = n3167 & ~n16657 ;
  assign n16659 = n2388 & ~n3832 ;
  assign n16660 = n16658 & n16659 ;
  assign n16662 = n3364 | n4722 ;
  assign n16663 = ( ~n7842 & n10301 ) | ( ~n7842 & n16662 ) | ( n10301 & n16662 ) ;
  assign n16661 = x110 & ~n5590 ;
  assign n16664 = n16663 ^ n16661 ^ n14240 ;
  assign n16665 = n5859 & ~n12226 ;
  assign n16666 = n8371 ^ n6331 ^ 1'b0 ;
  assign n16667 = ~n6105 & n16666 ;
  assign n16668 = n16667 ^ n5966 ^ 1'b0 ;
  assign n16669 = ~n12308 & n16668 ;
  assign n16670 = n5586 & ~n6633 ;
  assign n16671 = n16670 ^ n9012 ^ 1'b0 ;
  assign n16678 = n13054 ^ n2407 ^ n293 ;
  assign n16679 = n7734 | n8335 ;
  assign n16680 = n16678 & ~n16679 ;
  assign n16681 = ~n9275 & n16680 ;
  assign n16672 = n7603 | n12153 ;
  assign n16673 = ~n3511 & n16672 ;
  assign n16674 = n16673 ^ n4257 ^ 1'b0 ;
  assign n16675 = n16674 ^ n6614 ^ 1'b0 ;
  assign n16676 = n8980 & n16675 ;
  assign n16677 = ~n903 & n16676 ;
  assign n16682 = n16681 ^ n16677 ^ 1'b0 ;
  assign n16683 = ( n2213 & n5859 ) | ( n2213 & ~n10573 ) | ( n5859 & ~n10573 ) ;
  assign n16684 = n9578 ^ n8045 ^ 1'b0 ;
  assign n16685 = n16683 & ~n16684 ;
  assign n16686 = n9528 & ~n9982 ;
  assign n16687 = n16686 ^ n10840 ^ 1'b0 ;
  assign n16691 = n3115 & ~n8003 ;
  assign n16688 = n4897 ^ n3225 ^ 1'b0 ;
  assign n16689 = n1021 | n16688 ;
  assign n16690 = n1163 & ~n16689 ;
  assign n16692 = n16691 ^ n16690 ^ 1'b0 ;
  assign n16693 = n16692 ^ n5064 ^ 1'b0 ;
  assign n16694 = n8695 ^ x4 ^ 1'b0 ;
  assign n16695 = n11635 | n16694 ;
  assign n16696 = n5970 & n16695 ;
  assign n16697 = n1503 & n12790 ;
  assign n16701 = n1652 & ~n12218 ;
  assign n16698 = n506 | n10265 ;
  assign n16699 = n16698 ^ n2990 ^ 1'b0 ;
  assign n16700 = ~n12141 & n16699 ;
  assign n16702 = n16701 ^ n16700 ^ 1'b0 ;
  assign n16703 = n16697 & ~n16702 ;
  assign n16704 = n10283 & n10310 ;
  assign n16705 = n632 & n16704 ;
  assign n16706 = n556 & ~n14372 ;
  assign n16707 = n5323 & n16706 ;
  assign n16708 = n11105 ^ n9950 ^ 1'b0 ;
  assign n16709 = n2308 | n6404 ;
  assign n16710 = n16157 ^ n423 ^ 1'b0 ;
  assign n16711 = n12009 ^ n4844 ^ 1'b0 ;
  assign n16714 = n6377 ^ n3398 ^ n2832 ;
  assign n16715 = n13494 & n16714 ;
  assign n16712 = n1588 | n10039 ;
  assign n16713 = n2370 | n16712 ;
  assign n16716 = n16715 ^ n16713 ^ 1'b0 ;
  assign n16718 = n636 ^ n605 ^ 1'b0 ;
  assign n16719 = n7973 & ~n16718 ;
  assign n16717 = n7964 | n8643 ;
  assign n16720 = n16719 ^ n16717 ^ 1'b0 ;
  assign n16721 = n9766 ^ n7806 ^ 1'b0 ;
  assign n16722 = n13268 | n16721 ;
  assign n16723 = n1615 | n16722 ;
  assign n16724 = n3641 ^ n2135 ^ 1'b0 ;
  assign n16725 = n8733 | n16724 ;
  assign n16726 = n16723 | n16725 ;
  assign n16727 = n16720 | n16726 ;
  assign n16730 = n4578 ^ n2280 ^ 1'b0 ;
  assign n16731 = ~n10960 & n16730 ;
  assign n16728 = n5526 | n6497 ;
  assign n16729 = n4252 & n16728 ;
  assign n16732 = n16731 ^ n16729 ^ 1'b0 ;
  assign n16733 = n12267 & ~n16732 ;
  assign n16734 = n4045 & n7951 ;
  assign n16735 = ~n8240 & n16734 ;
  assign n16736 = n16735 ^ n5511 ^ 1'b0 ;
  assign n16737 = n1497 | n16736 ;
  assign n16738 = n4126 & n11807 ;
  assign n16739 = n16738 ^ n9554 ^ 1'b0 ;
  assign n16740 = ( ~n882 & n2617 ) | ( ~n882 & n9195 ) | ( n2617 & n9195 ) ;
  assign n16741 = n4817 ^ n2776 ^ n549 ;
  assign n16742 = n3981 ^ n3304 ^ 1'b0 ;
  assign n16746 = n2517 & n4860 ;
  assign n16747 = ~n1396 & n16746 ;
  assign n16748 = n12370 ^ n11747 ^ 1'b0 ;
  assign n16749 = n16747 | n16748 ;
  assign n16743 = n10946 ^ n5102 ^ 1'b0 ;
  assign n16744 = n3405 | n16743 ;
  assign n16745 = n16744 ^ n15667 ^ 1'b0 ;
  assign n16750 = n16749 ^ n16745 ^ n7264 ;
  assign n16751 = ( n16741 & ~n16742 ) | ( n16741 & n16750 ) | ( ~n16742 & n16750 ) ;
  assign n16752 = ~n4609 & n10552 ;
  assign n16753 = n16752 ^ n7158 ^ 1'b0 ;
  assign n16755 = ~n3850 & n8534 ;
  assign n16754 = n5043 ^ n3051 ^ 1'b0 ;
  assign n16756 = n16755 ^ n16754 ^ n3257 ;
  assign n16757 = n16756 ^ n7230 ^ 1'b0 ;
  assign n16758 = n4923 ^ n1761 ^ 1'b0 ;
  assign n16759 = n5465 | n16758 ;
  assign n16760 = n13384 & ~n16759 ;
  assign n16761 = n7985 | n13046 ;
  assign n16762 = n8534 | n16761 ;
  assign n16763 = ~n209 & n6419 ;
  assign n16764 = n16763 ^ n14143 ^ 1'b0 ;
  assign n16765 = n10146 ^ n2109 ^ 1'b0 ;
  assign n16766 = n4224 & n4308 ;
  assign n16767 = n15415 ^ n6018 ^ n1541 ;
  assign n16768 = n1133 & n2670 ;
  assign n16769 = ( n1681 & n2138 ) | ( n1681 & ~n16768 ) | ( n2138 & ~n16768 ) ;
  assign n16770 = n954 & n16769 ;
  assign n16772 = n10368 ^ n8401 ^ 1'b0 ;
  assign n16773 = n1552 & n16772 ;
  assign n16774 = n16773 ^ n5834 ^ 1'b0 ;
  assign n16771 = n4767 | n8074 ;
  assign n16775 = n16774 ^ n16771 ^ 1'b0 ;
  assign n16776 = n1250 & ~n10208 ;
  assign n16777 = ~n16775 & n16776 ;
  assign n16778 = x34 | n992 ;
  assign n16779 = n3844 ^ n2717 ^ 1'b0 ;
  assign n16780 = n403 & ~n16779 ;
  assign n16781 = ~n16778 & n16780 ;
  assign n16782 = n10592 & n16781 ;
  assign n16783 = ~n747 & n4851 ;
  assign n16784 = n4906 & n16783 ;
  assign n16785 = n16784 ^ n3219 ^ 1'b0 ;
  assign n16786 = n1432 & n16674 ;
  assign n16788 = n2151 & ~n5997 ;
  assign n16789 = n16788 ^ n9796 ^ n2561 ;
  assign n16787 = n4647 & ~n7050 ;
  assign n16790 = n16789 ^ n16787 ^ 1'b0 ;
  assign n16791 = ( ~n747 & n3336 ) | ( ~n747 & n4757 ) | ( n3336 & n4757 ) ;
  assign n16792 = n2985 & n10189 ;
  assign n16793 = n1190 & n14586 ;
  assign n16794 = n16793 ^ n9323 ^ 1'b0 ;
  assign n16795 = n16792 & ~n16794 ;
  assign n16796 = n1531 | n6273 ;
  assign n16797 = ~n10861 & n16796 ;
  assign n16798 = n16797 ^ n7934 ^ 1'b0 ;
  assign n16799 = n8952 ^ n8841 ^ 1'b0 ;
  assign n16800 = ~n11181 & n16799 ;
  assign n16801 = ~n13680 & n16800 ;
  assign n16802 = n7102 & ~n14587 ;
  assign n16803 = ~n6206 & n10462 ;
  assign n16804 = n16803 ^ n6457 ^ 1'b0 ;
  assign n16805 = n15696 ^ n6122 ^ 1'b0 ;
  assign n16806 = n2170 & n16805 ;
  assign n16807 = n1259 ^ n453 ^ 1'b0 ;
  assign n16808 = n16806 & ~n16807 ;
  assign n16809 = n2676 & n7920 ;
  assign n16810 = ~n6189 & n15793 ;
  assign n16811 = n16810 ^ n10342 ^ 1'b0 ;
  assign n16812 = n13739 ^ n6321 ^ 1'b0 ;
  assign n16813 = n2987 & n3350 ;
  assign n16814 = n9775 & ~n16813 ;
  assign n16815 = n16814 ^ n9939 ^ 1'b0 ;
  assign n16816 = n8849 & n16691 ;
  assign n16817 = n10934 | n11117 ;
  assign n16818 = n16816 | n16817 ;
  assign n16819 = n461 | n9781 ;
  assign n16820 = n16819 ^ n11891 ^ 1'b0 ;
  assign n16821 = n833 & ~n16820 ;
  assign n16822 = n2289 | n3234 ;
  assign n16823 = n9362 & ~n9471 ;
  assign n16826 = n5968 ^ n1558 ^ 1'b0 ;
  assign n16824 = n8714 | n11410 ;
  assign n16825 = n874 | n16824 ;
  assign n16827 = n16826 ^ n16825 ^ 1'b0 ;
  assign n16828 = n4581 & ~n16827 ;
  assign n16829 = ~n14037 & n16828 ;
  assign n16833 = n4441 ^ x18 ^ 1'b0 ;
  assign n16830 = n2983 | n3403 ;
  assign n16831 = n16830 ^ n3674 ^ 1'b0 ;
  assign n16832 = ~n4883 & n16831 ;
  assign n16834 = n16833 ^ n16832 ^ 1'b0 ;
  assign n16837 = n538 & ~n10338 ;
  assign n16835 = n11650 ^ n7771 ^ 1'b0 ;
  assign n16836 = n1256 & n16835 ;
  assign n16838 = n16837 ^ n16836 ^ n8339 ;
  assign n16839 = n16838 ^ n13242 ^ 1'b0 ;
  assign n16840 = n16834 & n16839 ;
  assign n16841 = n4082 ^ n1380 ^ 1'b0 ;
  assign n16842 = n13992 ^ n13736 ^ n918 ;
  assign n16843 = n16842 ^ n5211 ^ n190 ;
  assign n16844 = n12790 ^ n10377 ^ n4813 ;
  assign n16845 = n6751 ^ n1215 ^ 1'b0 ;
  assign n16846 = ~n1553 & n16845 ;
  assign n16847 = n8688 & n16846 ;
  assign n16848 = n11474 & n13491 ;
  assign n16849 = n11971 & ~n13994 ;
  assign n16850 = n1271 & n2796 ;
  assign n16851 = n16850 ^ n6751 ^ 1'b0 ;
  assign n16852 = n16851 ^ n14832 ^ 1'b0 ;
  assign n16853 = n6364 | n13502 ;
  assign n16854 = n16853 ^ n16389 ^ n3573 ;
  assign n16855 = n11067 ^ n9845 ^ 1'b0 ;
  assign n16856 = n3978 & n8585 ;
  assign n16857 = ~n1770 & n12977 ;
  assign n16858 = ~n3965 & n5275 ;
  assign n16859 = n4649 ^ n3972 ^ 1'b0 ;
  assign n16860 = n3626 & ~n16859 ;
  assign n16861 = ( n5345 & n16858 ) | ( n5345 & n16860 ) | ( n16858 & n16860 ) ;
  assign n16862 = n15852 ^ n3011 ^ n595 ;
  assign n16863 = n10752 ^ n6307 ^ n2289 ;
  assign n16864 = n3965 & n16863 ;
  assign n16865 = n6929 & ~n14997 ;
  assign n16866 = n16865 ^ n8762 ^ 1'b0 ;
  assign n16867 = ~n1619 & n6356 ;
  assign n16868 = n16867 ^ n1973 ^ 1'b0 ;
  assign n16869 = n16868 ^ n11851 ^ 1'b0 ;
  assign n16870 = n7816 & n16869 ;
  assign n16872 = n13994 ^ n3365 ^ 1'b0 ;
  assign n16871 = n2481 & n14827 ;
  assign n16873 = n16872 ^ n16871 ^ 1'b0 ;
  assign n16874 = n2998 & ~n13427 ;
  assign n16875 = n11260 | n13466 ;
  assign n16876 = ~n2644 & n2912 ;
  assign n16877 = n12369 | n16876 ;
  assign n16878 = n8144 ^ n3880 ^ n425 ;
  assign n16879 = n14240 ^ n2814 ^ 1'b0 ;
  assign n16880 = n16879 ^ n1601 ^ 1'b0 ;
  assign n16881 = n16878 & n16880 ;
  assign n16882 = x27 & n16881 ;
  assign n16883 = n13804 & ~n15042 ;
  assign n16888 = n15802 ^ n13027 ^ 1'b0 ;
  assign n16889 = x71 & n16888 ;
  assign n16884 = x9 & ~n3447 ;
  assign n16885 = n16884 ^ n2769 ^ 1'b0 ;
  assign n16886 = n6676 & n16885 ;
  assign n16887 = ( ~n10615 & n12731 ) | ( ~n10615 & n16886 ) | ( n12731 & n16886 ) ;
  assign n16890 = n16889 ^ n16887 ^ 1'b0 ;
  assign n16891 = ~n15428 & n16890 ;
  assign n16892 = n15731 ^ n7514 ^ 1'b0 ;
  assign n16893 = n10730 & n16892 ;
  assign n16894 = n16893 ^ n2341 ^ 1'b0 ;
  assign n16895 = n1746 & ~n16894 ;
  assign n16896 = n16895 ^ n8776 ^ n5703 ;
  assign n16897 = ~n6084 & n15804 ;
  assign n16898 = n16897 ^ n12145 ^ 1'b0 ;
  assign n16899 = n960 & ~n3276 ;
  assign n16900 = n16899 ^ n4292 ^ n609 ;
  assign n16901 = ~n15030 & n16900 ;
  assign n16902 = x55 & ~n1488 ;
  assign n16903 = n1488 & n16902 ;
  assign n16904 = ~n7483 & n16903 ;
  assign n16905 = ~n2144 & n8634 ;
  assign n16906 = ~n8634 & n16905 ;
  assign n16907 = n911 & ~n16906 ;
  assign n16908 = ~n911 & n16907 ;
  assign n16909 = n16908 ^ n4217 ^ 1'b0 ;
  assign n16910 = ~n16904 & n16909 ;
  assign n16911 = n16904 & n16910 ;
  assign n16912 = n2960 | n4666 ;
  assign n16913 = n16912 ^ n7928 ^ 1'b0 ;
  assign n16914 = ( ~n1019 & n5552 ) | ( ~n1019 & n16913 ) | ( n5552 & n16913 ) ;
  assign n16915 = n16914 ^ n6753 ^ 1'b0 ;
  assign n16916 = n16915 ^ n1353 ^ 1'b0 ;
  assign n16917 = ~n12395 & n16916 ;
  assign n16918 = n4516 & ~n9949 ;
  assign n16919 = n16918 ^ n2566 ^ 1'b0 ;
  assign n16920 = n7267 | n16919 ;
  assign n16921 = ~n252 & n10043 ;
  assign n16922 = n16921 ^ n11737 ^ 1'b0 ;
  assign n16923 = n13330 ^ n7075 ^ 1'b0 ;
  assign n16924 = n16923 ^ n7329 ^ 1'b0 ;
  assign n16928 = n8502 & ~n13882 ;
  assign n16925 = x115 & ~n373 ;
  assign n16926 = n16925 ^ n15406 ^ 1'b0 ;
  assign n16927 = n9620 | n16926 ;
  assign n16929 = n16928 ^ n16927 ^ 1'b0 ;
  assign n16930 = n317 | n821 ;
  assign n16931 = ~n5052 & n5725 ;
  assign n16932 = n4055 | n9026 ;
  assign n16933 = n10836 & ~n16932 ;
  assign n16934 = n16931 & n16933 ;
  assign n16935 = ( ~n1661 & n1718 ) | ( ~n1661 & n16470 ) | ( n1718 & n16470 ) ;
  assign n16936 = n16935 ^ n14208 ^ 1'b0 ;
  assign n16937 = n4547 ^ n1738 ^ 1'b0 ;
  assign n16938 = n2228 | n14610 ;
  assign n16939 = n9103 ^ n5905 ^ 1'b0 ;
  assign n16940 = n13019 & ~n16939 ;
  assign n16941 = ~n1225 & n3647 ;
  assign n16942 = n16941 ^ n3635 ^ 1'b0 ;
  assign n16943 = ( n5355 & n14333 ) | ( n5355 & n16942 ) | ( n14333 & n16942 ) ;
  assign n16944 = n2293 & n16943 ;
  assign n16945 = n10801 ^ n9966 ^ 1'b0 ;
  assign n16946 = n16945 ^ n14260 ^ 1'b0 ;
  assign n16947 = n391 & ~n3973 ;
  assign n16948 = n13834 & n16947 ;
  assign n16949 = n1391 & n3815 ;
  assign n16950 = n16949 ^ n2103 ^ 1'b0 ;
  assign n16951 = x37 & n4069 ;
  assign n16952 = ~n14166 & n16951 ;
  assign n16953 = n6376 ^ n5168 ^ 1'b0 ;
  assign n16954 = n4764 ^ n2285 ^ 1'b0 ;
  assign n16955 = n3360 | n5244 ;
  assign n16956 = n16955 ^ n2824 ^ 1'b0 ;
  assign n16957 = n16956 ^ n1828 ^ 1'b0 ;
  assign n16958 = ~n15949 & n16957 ;
  assign n16959 = n6864 | n14687 ;
  assign n16960 = ~n6043 & n7102 ;
  assign n16961 = n7404 & n13972 ;
  assign n16962 = n10401 & ~n15966 ;
  assign n16963 = n16962 ^ n13760 ^ 1'b0 ;
  assign n16964 = n16963 ^ n5578 ^ 1'b0 ;
  assign n16965 = n13780 & ~n16964 ;
  assign n16966 = n7834 & n16965 ;
  assign n16967 = n5868 ^ n1536 ^ 1'b0 ;
  assign n16968 = n11872 | n16967 ;
  assign n16971 = n7525 & ~n9532 ;
  assign n16969 = n4510 | n5758 ;
  assign n16970 = n2156 & n16969 ;
  assign n16972 = n16971 ^ n16970 ^ 1'b0 ;
  assign n16973 = n2776 | n8020 ;
  assign n16974 = n6665 ^ n4776 ^ 1'b0 ;
  assign n16975 = ( n6120 & ~n12336 ) | ( n6120 & n16974 ) | ( ~n12336 & n16974 ) ;
  assign n16976 = n16975 ^ n3823 ^ 1'b0 ;
  assign n16977 = n1716 & n16976 ;
  assign n16978 = ~n14701 & n16977 ;
  assign n16979 = ~n16973 & n16978 ;
  assign n16980 = n16166 ^ n2970 ^ 1'b0 ;
  assign n16981 = n1442 & n16980 ;
  assign n16982 = n10885 & n16981 ;
  assign n16983 = n16982 ^ n7964 ^ 1'b0 ;
  assign n16984 = ~x6 & n16885 ;
  assign n16985 = n3203 ^ n1529 ^ 1'b0 ;
  assign n16986 = ~n8550 & n15255 ;
  assign n16987 = ~n16166 & n16986 ;
  assign n16988 = n10171 ^ n1772 ^ 1'b0 ;
  assign n16989 = ( n1121 & n13933 ) | ( n1121 & ~n15474 ) | ( n13933 & ~n15474 ) ;
  assign n16990 = ( ~n2118 & n6087 ) | ( ~n2118 & n6901 ) | ( n6087 & n6901 ) ;
  assign n16991 = n15388 | n16990 ;
  assign n16992 = n6523 & n9988 ;
  assign n16993 = n16992 ^ n10820 ^ 1'b0 ;
  assign n16994 = n4065 & ~n16993 ;
  assign n16995 = ~n1538 & n15312 ;
  assign n16996 = n2575 & n14846 ;
  assign n16997 = n16996 ^ n1865 ^ 1'b0 ;
  assign n16998 = n14201 | n16997 ;
  assign n16999 = n2470 & ~n3089 ;
  assign n17000 = n16999 ^ x69 ^ 1'b0 ;
  assign n17001 = n1761 & n6145 ;
  assign n17002 = n2020 & n8240 ;
  assign n17003 = ~n7538 & n17002 ;
  assign n17004 = n17003 ^ n1433 ^ 1'b0 ;
  assign n17005 = n7250 ^ n6044 ^ 1'b0 ;
  assign n17006 = n4130 | n17005 ;
  assign n17007 = n5135 | n17006 ;
  assign n17008 = n2029 & ~n17007 ;
  assign n17009 = n9638 & ~n15049 ;
  assign n17010 = ~n11737 & n17009 ;
  assign n17014 = n676 | n2670 ;
  assign n17015 = n17014 ^ n5044 ^ 1'b0 ;
  assign n17016 = x82 & n3815 ;
  assign n17017 = ~n17015 & n17016 ;
  assign n17018 = n12717 | n17017 ;
  assign n17019 = n17018 ^ n16095 ^ 1'b0 ;
  assign n17020 = n8198 & ~n17019 ;
  assign n17011 = n9291 ^ n6932 ^ 1'b0 ;
  assign n17012 = n4588 | n17011 ;
  assign n17013 = n5481 | n17012 ;
  assign n17021 = n17020 ^ n17013 ^ 1'b0 ;
  assign n17024 = n8129 & ~n12686 ;
  assign n17022 = n2694 | n9303 ;
  assign n17023 = n3569 | n17022 ;
  assign n17025 = n17024 ^ n17023 ^ 1'b0 ;
  assign n17026 = n7160 | n17025 ;
  assign n17027 = n2308 & ~n3124 ;
  assign n17028 = n4044 ^ n2447 ^ 1'b0 ;
  assign n17029 = n15391 & ~n17028 ;
  assign n17030 = n5238 & n17029 ;
  assign n17031 = ~n4018 & n17030 ;
  assign n17032 = n6188 | n17031 ;
  assign n17033 = ~n6114 & n6472 ;
  assign n17034 = n9801 & n17033 ;
  assign n17035 = n17034 ^ n1346 ^ 1'b0 ;
  assign n17036 = ~n2810 & n3795 ;
  assign n17037 = n17036 ^ n444 ^ 1'b0 ;
  assign n17038 = n8686 & ~n11578 ;
  assign n17039 = ~n5040 & n17038 ;
  assign n17040 = n9706 & n17039 ;
  assign n17041 = n4879 | n17040 ;
  assign n17042 = n8299 ^ n777 ^ 1'b0 ;
  assign n17043 = ~n4777 & n17042 ;
  assign n17044 = n488 | n5183 ;
  assign n17045 = n488 & ~n17044 ;
  assign n17046 = n981 & ~n17045 ;
  assign n17047 = n17046 ^ n844 ^ 1'b0 ;
  assign n17048 = ~n15431 & n17047 ;
  assign n17049 = ~n2203 & n4574 ;
  assign n17050 = n17049 ^ n4408 ^ 1'b0 ;
  assign n17051 = n10041 ^ n4309 ^ 1'b0 ;
  assign n17052 = n17050 & ~n17051 ;
  assign n17053 = n17052 ^ n8081 ^ 1'b0 ;
  assign n17054 = n3925 | n17053 ;
  assign n17055 = n15058 ^ n3229 ^ 1'b0 ;
  assign n17056 = n10392 & ~n11822 ;
  assign n17058 = n10397 & ~n13469 ;
  assign n17059 = n17058 ^ n1155 ^ 1'b0 ;
  assign n17060 = n4004 & n17059 ;
  assign n17057 = n4700 & ~n6724 ;
  assign n17061 = n17060 ^ n17057 ^ 1'b0 ;
  assign n17062 = n17056 & n17061 ;
  assign n17063 = n17062 ^ n9452 ^ 1'b0 ;
  assign n17064 = n8619 ^ n7568 ^ 1'b0 ;
  assign n17065 = n8677 ^ n2853 ^ 1'b0 ;
  assign n17066 = n17064 & ~n17065 ;
  assign n17067 = n17066 ^ n13803 ^ 1'b0 ;
  assign n17068 = ~n2856 & n17067 ;
  assign n17069 = n8795 ^ n1970 ^ 1'b0 ;
  assign n17070 = n13162 & n17069 ;
  assign n17071 = n2067 | n2178 ;
  assign n17072 = n3212 | n17071 ;
  assign n17073 = n17072 ^ n4579 ^ 1'b0 ;
  assign n17074 = n11333 ^ n5370 ^ 1'b0 ;
  assign n17075 = n17073 & ~n17074 ;
  assign n17076 = n1019 | n1166 ;
  assign n17077 = n12926 & ~n17076 ;
  assign n17078 = ( n1654 & ~n17075 ) | ( n1654 & n17077 ) | ( ~n17075 & n17077 ) ;
  assign n17079 = n13516 | n15985 ;
  assign n17080 = n4554 | n17079 ;
  assign n17081 = n2156 | n17080 ;
  assign n17082 = ~n1235 & n15544 ;
  assign n17083 = n11208 ^ n5513 ^ 1'b0 ;
  assign n17084 = n17082 & n17083 ;
  assign n17085 = ~x103 & n878 ;
  assign n17086 = n11399 & ~n17085 ;
  assign n17087 = n15294 & n17086 ;
  assign n17088 = n3118 & ~n9570 ;
  assign n17089 = n3494 & n14941 ;
  assign n17090 = n17088 & n17089 ;
  assign n17091 = n11121 ^ n9600 ^ 1'b0 ;
  assign n17093 = n6861 ^ n3863 ^ 1'b0 ;
  assign n17094 = ~n560 & n17093 ;
  assign n17095 = n17094 ^ n5533 ^ 1'b0 ;
  assign n17092 = n3804 | n11921 ;
  assign n17096 = n17095 ^ n17092 ^ 1'b0 ;
  assign n17097 = n14159 | n17096 ;
  assign n17098 = n7279 | n17097 ;
  assign n17099 = n9587 | n10039 ;
  assign n17100 = n17099 ^ n7705 ^ 1'b0 ;
  assign n17101 = n17100 ^ n9225 ^ 1'b0 ;
  assign n17102 = n3072 | n17101 ;
  assign n17103 = ~n15134 & n15352 ;
  assign n17104 = n17103 ^ n2527 ^ 1'b0 ;
  assign n17105 = n4851 & n6101 ;
  assign n17106 = n9273 & n17105 ;
  assign n17107 = n9084 ^ n1081 ^ 1'b0 ;
  assign n17108 = n17107 ^ n12213 ^ n6644 ;
  assign n17109 = n17108 ^ n709 ^ 1'b0 ;
  assign n17110 = n15359 | n17109 ;
  assign n17111 = n16242 ^ n2445 ^ 1'b0 ;
  assign n17112 = n14296 ^ n1105 ^ 1'b0 ;
  assign n17113 = n311 & n17112 ;
  assign n17114 = n15106 & n17113 ;
  assign n17115 = n17114 ^ n1920 ^ 1'b0 ;
  assign n17116 = n7925 | n11324 ;
  assign n17117 = n17115 | n17116 ;
  assign n17118 = x24 & ~n12678 ;
  assign n17119 = n6212 ^ n2340 ^ 1'b0 ;
  assign n17120 = n9955 ^ n5034 ^ 1'b0 ;
  assign n17121 = ~n14089 & n17120 ;
  assign n17122 = ~n8413 & n17121 ;
  assign n17123 = n369 | n17122 ;
  assign n17124 = n8386 & n13346 ;
  assign n17125 = x83 & n6159 ;
  assign n17126 = n179 & ~n10573 ;
  assign n17127 = n9452 & n17126 ;
  assign n17128 = ( n5829 & ~n8597 ) | ( n5829 & n17127 ) | ( ~n8597 & n17127 ) ;
  assign n17129 = n7531 ^ n2694 ^ 1'b0 ;
  assign n17130 = n3174 & ~n12487 ;
  assign n17131 = ~n9810 & n17130 ;
  assign n17133 = n6781 ^ n5459 ^ n3646 ;
  assign n17134 = n7075 ^ n5150 ^ 1'b0 ;
  assign n17135 = ~n17133 & n17134 ;
  assign n17132 = n11703 | n11985 ;
  assign n17136 = n17135 ^ n17132 ^ 1'b0 ;
  assign n17137 = n17136 ^ n5715 ^ 1'b0 ;
  assign n17138 = n11000 & n17137 ;
  assign n17139 = n12409 & ~n14732 ;
  assign n17140 = n17139 ^ n12491 ^ 1'b0 ;
  assign n17141 = n16414 | n17140 ;
  assign n17142 = n14016 ^ n4924 ^ 1'b0 ;
  assign n17143 = ( n3587 & ~n6111 ) | ( n3587 & n6386 ) | ( ~n6111 & n6386 ) ;
  assign n17144 = n17143 ^ n12458 ^ n6440 ;
  assign n17145 = n10797 & n13425 ;
  assign n17146 = n3839 | n7527 ;
  assign n17147 = ~n6535 & n17146 ;
  assign n17148 = n14923 & n17147 ;
  assign n17149 = n905 & n12974 ;
  assign n17150 = n3367 & n6753 ;
  assign n17151 = ~n17149 & n17150 ;
  assign n17152 = n6110 & ~n11575 ;
  assign n17153 = n3364 | n6281 ;
  assign n17154 = n17153 ^ n2213 ^ 1'b0 ;
  assign n17155 = n17154 ^ n1289 ^ 1'b0 ;
  assign n17156 = n157 & ~n17155 ;
  assign n17157 = n17156 ^ n11996 ^ 1'b0 ;
  assign n17158 = ( n2053 & n2489 ) | ( n2053 & n3662 ) | ( n2489 & n3662 ) ;
  assign n17159 = n4523 & ~n8915 ;
  assign n17160 = n17159 ^ n2014 ^ 1'b0 ;
  assign n17161 = n2542 & ~n5142 ;
  assign n17162 = n11650 ^ n7797 ^ 1'b0 ;
  assign n17163 = n7300 & ~n17162 ;
  assign n17164 = ~n786 & n2027 ;
  assign n17165 = n883 & ~n17164 ;
  assign n17166 = n17165 ^ n14079 ^ 1'b0 ;
  assign n17167 = n17163 & n17166 ;
  assign n17168 = ~n3300 & n3717 ;
  assign n17169 = n9295 & n17168 ;
  assign n17170 = n3931 & n4377 ;
  assign n17171 = n17170 ^ n15078 ^ n7711 ;
  assign n17173 = n4077 | n8191 ;
  assign n17172 = ~n6002 & n8996 ;
  assign n17174 = n17173 ^ n17172 ^ 1'b0 ;
  assign n17175 = n888 & ~n4441 ;
  assign n17176 = ( n4648 & n5129 ) | ( n4648 & n13771 ) | ( n5129 & n13771 ) ;
  assign n17177 = n17176 ^ n14085 ^ n12974 ;
  assign n17178 = n17175 & ~n17177 ;
  assign n17179 = ~n2374 & n3808 ;
  assign n17180 = n11389 & n17179 ;
  assign n17181 = n13112 & n14803 ;
  assign n17182 = n17181 ^ n9517 ^ n2042 ;
  assign n17184 = n4273 ^ n3148 ^ 1'b0 ;
  assign n17185 = ~n13083 & n17184 ;
  assign n17183 = n1054 & n10992 ;
  assign n17186 = n17185 ^ n17183 ^ 1'b0 ;
  assign n17187 = n5374 | n17186 ;
  assign n17188 = n17187 ^ n5127 ^ 1'b0 ;
  assign n17189 = n7114 ^ n5385 ^ 1'b0 ;
  assign n17190 = ( n2470 & n2901 ) | ( n2470 & n5874 ) | ( n2901 & n5874 ) ;
  assign n17191 = n17190 ^ n5487 ^ 1'b0 ;
  assign n17192 = n3460 & ~n17191 ;
  assign n17193 = x97 & n3478 ;
  assign n17194 = n17193 ^ n1116 ^ 1'b0 ;
  assign n17195 = n15955 ^ n8776 ^ 1'b0 ;
  assign n17196 = n3019 & n17195 ;
  assign n17197 = n1570 & n2961 ;
  assign n17198 = n12813 & n17197 ;
  assign n17199 = n2259 | n3884 ;
  assign n17200 = n5665 ^ n525 ^ 1'b0 ;
  assign n17201 = n17200 ^ n10399 ^ n338 ;
  assign n17202 = ( ~n5846 & n17199 ) | ( ~n5846 & n17201 ) | ( n17199 & n17201 ) ;
  assign n17203 = n5910 & ~n15002 ;
  assign n17204 = n9603 ^ n5643 ^ 1'b0 ;
  assign n17206 = n9132 ^ n4085 ^ 1'b0 ;
  assign n17207 = n17206 ^ n8189 ^ 1'b0 ;
  assign n17208 = ~n3635 & n17207 ;
  assign n17205 = n1722 | n2899 ;
  assign n17209 = n17208 ^ n17205 ^ 1'b0 ;
  assign n17210 = n8971 ^ n6148 ^ 1'b0 ;
  assign n17211 = ( ~n261 & n6321 ) | ( ~n261 & n16768 ) | ( n6321 & n16768 ) ;
  assign n17212 = n17211 ^ n2622 ^ 1'b0 ;
  assign n17213 = n1847 ^ n477 ^ 1'b0 ;
  assign n17214 = n4008 | n17213 ;
  assign n17215 = n17214 ^ n16234 ^ 1'b0 ;
  assign n17216 = n13360 | n17215 ;
  assign n17217 = n14316 ^ n551 ^ 1'b0 ;
  assign n17218 = n13050 & ~n13323 ;
  assign n17219 = n5954 & n16691 ;
  assign n17220 = ~n13279 & n17219 ;
  assign n17221 = ( ~n17217 & n17218 ) | ( ~n17217 & n17220 ) | ( n17218 & n17220 ) ;
  assign n17222 = n3993 ^ n1776 ^ 1'b0 ;
  assign n17223 = n3685 | n17222 ;
  assign n17224 = n8509 & ~n16031 ;
  assign n17225 = n15383 & ~n17224 ;
  assign n17226 = n17225 ^ n7674 ^ 1'b0 ;
  assign n17227 = n3217 & n14839 ;
  assign n17228 = ~n6981 & n17227 ;
  assign n17229 = n5297 & ~n17228 ;
  assign n17230 = n17229 ^ n1066 ^ 1'b0 ;
  assign n17231 = n14543 & ~n17230 ;
  assign n17232 = ~n17226 & n17231 ;
  assign n17233 = n17126 ^ n5238 ^ n3505 ;
  assign n17234 = n6762 & n17233 ;
  assign n17235 = n986 & n2693 ;
  assign n17236 = n17235 ^ n16636 ^ 1'b0 ;
  assign n17237 = n4006 & ~n6984 ;
  assign n17238 = n9837 | n17237 ;
  assign n17239 = n14298 | n15378 ;
  assign n17240 = n1133 | n17239 ;
  assign n17243 = n5960 | n13854 ;
  assign n17244 = n12734 | n17243 ;
  assign n17245 = ( ~n1910 & n10891 ) | ( ~n1910 & n17244 ) | ( n10891 & n17244 ) ;
  assign n17241 = n3476 & ~n6680 ;
  assign n17242 = n8237 | n17241 ;
  assign n17246 = n17245 ^ n17242 ^ 1'b0 ;
  assign n17250 = n8583 ^ n1865 ^ x98 ;
  assign n17251 = ~n5315 & n17250 ;
  assign n17252 = n17251 ^ n9794 ^ 1'b0 ;
  assign n17249 = ~n2228 & n6608 ;
  assign n17253 = n17252 ^ n17249 ^ 1'b0 ;
  assign n17247 = n10999 & n16816 ;
  assign n17248 = n2645 & n17247 ;
  assign n17254 = n17253 ^ n17248 ^ 1'b0 ;
  assign n17255 = n2689 | n3651 ;
  assign n17256 = ~n8490 & n12912 ;
  assign n17257 = n14138 ^ n6796 ^ 1'b0 ;
  assign n17258 = n3058 & n9413 ;
  assign n17259 = n2936 & n17258 ;
  assign n17260 = n1484 | n17259 ;
  assign n17261 = n17260 ^ n1742 ^ 1'b0 ;
  assign n17262 = n3704 & ~n17261 ;
  assign n17263 = n5451 ^ n2261 ^ 1'b0 ;
  assign n17264 = n12083 & n17263 ;
  assign n17265 = n17264 ^ n6667 ^ 1'b0 ;
  assign n17266 = ( ~n706 & n8880 ) | ( ~n706 & n9396 ) | ( n8880 & n9396 ) ;
  assign n17267 = n4266 & n17266 ;
  assign n17268 = n8146 & n17267 ;
  assign n17269 = n11004 | n17268 ;
  assign n17270 = n8867 ^ n759 ^ 1'b0 ;
  assign n17271 = n5206 | n17270 ;
  assign n17272 = n13817 | n17271 ;
  assign n17273 = ~n9132 & n15941 ;
  assign n17274 = n9383 ^ n2054 ^ 1'b0 ;
  assign n17275 = n239 & ~n8803 ;
  assign n17276 = n17275 ^ n3145 ^ 1'b0 ;
  assign n17277 = ( n7024 & ~n10305 ) | ( n7024 & n17276 ) | ( ~n10305 & n17276 ) ;
  assign n17278 = n7315 & n7345 ;
  assign n17279 = n17278 ^ n14592 ^ 1'b0 ;
  assign n17280 = n17279 ^ x46 ^ 1'b0 ;
  assign n17281 = n9690 & n17280 ;
  assign n17282 = n4388 ^ n1479 ^ 1'b0 ;
  assign n17283 = n530 & ~n17282 ;
  assign n17284 = n7049 ^ n448 ^ 1'b0 ;
  assign n17285 = n17283 & ~n17284 ;
  assign n17286 = n9610 ^ n6991 ^ 1'b0 ;
  assign n17287 = n10571 & n17286 ;
  assign n17288 = n3795 ^ n1746 ^ n143 ;
  assign n17289 = n17288 ^ n1787 ^ 1'b0 ;
  assign n17290 = n2607 | n9089 ;
  assign n17291 = n8966 & ~n17290 ;
  assign n17292 = n17291 ^ n2312 ^ 1'b0 ;
  assign n17293 = n14662 & n15736 ;
  assign n17294 = n17293 ^ n14990 ^ 1'b0 ;
  assign n17295 = n16206 ^ n5344 ^ 1'b0 ;
  assign n17296 = n14875 ^ n2261 ^ 1'b0 ;
  assign n17297 = n12023 & ~n17296 ;
  assign n17298 = n16532 ^ n4018 ^ x98 ;
  assign n17299 = n4126 & ~n17298 ;
  assign n17300 = n17299 ^ n8660 ^ 1'b0 ;
  assign n17301 = n2798 & n17300 ;
  assign n17302 = n8810 & n17301 ;
  assign n17303 = n8415 ^ n260 ^ 1'b0 ;
  assign n17304 = n6786 & n17303 ;
  assign n17305 = n3778 & ~n4107 ;
  assign n17306 = n17305 ^ n12471 ^ n11902 ;
  assign n17307 = n3215 | n16434 ;
  assign n17308 = n7022 ^ n2382 ^ 1'b0 ;
  assign n17309 = ~n157 & n7930 ;
  assign n17310 = n2636 & n17309 ;
  assign n17311 = n17310 ^ n12980 ^ 1'b0 ;
  assign n17312 = n17311 ^ n15605 ^ n13505 ;
  assign n17313 = n9892 & ~n12634 ;
  assign n17314 = n2652 & n17313 ;
  assign n17315 = n1612 | n5187 ;
  assign n17316 = n17314 & ~n17315 ;
  assign n17320 = ( x41 & ~n2140 ) | ( x41 & n4335 ) | ( ~n2140 & n4335 ) ;
  assign n17321 = n5904 | n7559 ;
  assign n17322 = n17320 | n17321 ;
  assign n17323 = ( n7793 & n15567 ) | ( n7793 & ~n17322 ) | ( n15567 & ~n17322 ) ;
  assign n17317 = n15576 ^ n12735 ^ 1'b0 ;
  assign n17318 = n6147 & n17317 ;
  assign n17319 = n10859 & n17318 ;
  assign n17324 = n17323 ^ n17319 ^ 1'b0 ;
  assign n17326 = n11244 ^ n9676 ^ 1'b0 ;
  assign n17327 = ~n756 & n17326 ;
  assign n17325 = x11 | n7575 ;
  assign n17328 = n17327 ^ n17325 ^ n7942 ;
  assign n17329 = n8306 & ~n17328 ;
  assign n17331 = ~n2893 & n3996 ;
  assign n17332 = n17331 ^ n7160 ^ 1'b0 ;
  assign n17330 = n11749 ^ n9768 ^ n1576 ;
  assign n17333 = n17332 ^ n17330 ^ n243 ;
  assign n17334 = n15171 ^ n8237 ^ 1'b0 ;
  assign n17335 = n10357 | n17334 ;
  assign n17336 = n799 & ~n6459 ;
  assign n17337 = n17336 ^ n8699 ^ 1'b0 ;
  assign n17338 = n17337 ^ n7534 ^ 1'b0 ;
  assign n17339 = n11477 & n17338 ;
  assign n17340 = ~n6258 & n11706 ;
  assign n17341 = n17340 ^ n13173 ^ 1'b0 ;
  assign n17342 = n13425 ^ n6558 ^ 1'b0 ;
  assign n17343 = n14357 & ~n16460 ;
  assign n17344 = n17343 ^ n13882 ^ 1'b0 ;
  assign n17345 = n10803 ^ n1150 ^ 1'b0 ;
  assign n17346 = n4639 | n9573 ;
  assign n17347 = ~n3030 & n3649 ;
  assign n17348 = ~n4581 & n17347 ;
  assign n17352 = n3947 & n11519 ;
  assign n17353 = n3086 & n17352 ;
  assign n17349 = n9964 & n16483 ;
  assign n17350 = ( ~n468 & n9884 ) | ( ~n468 & n11732 ) | ( n9884 & n11732 ) ;
  assign n17351 = n17349 & ~n17350 ;
  assign n17354 = n17353 ^ n17351 ^ 1'b0 ;
  assign n17357 = ( n2111 & n3674 ) | ( n2111 & n8000 ) | ( n3674 & n8000 ) ;
  assign n17355 = ~n2958 & n13459 ;
  assign n17356 = n17355 ^ n4944 ^ 1'b0 ;
  assign n17358 = n17357 ^ n17356 ^ 1'b0 ;
  assign n17359 = ~n10431 & n17358 ;
  assign n17360 = n16926 & n17359 ;
  assign n17361 = ~n763 & n5492 ;
  assign n17362 = n16217 ^ n2222 ^ 1'b0 ;
  assign n17363 = n8269 & n17362 ;
  assign n17364 = n6895 & ~n12380 ;
  assign n17365 = n1693 & ~n4866 ;
  assign n17366 = n17365 ^ n947 ^ 1'b0 ;
  assign n17367 = ~n504 & n17366 ;
  assign n17368 = n2992 & n8391 ;
  assign n17369 = n17368 ^ n2425 ^ 1'b0 ;
  assign n17370 = n17367 & ~n17369 ;
  assign n17371 = n14066 | n14372 ;
  assign n17372 = n13187 ^ n8939 ^ n1587 ;
  assign n17373 = n6114 | n13586 ;
  assign n17374 = n17373 ^ n11727 ^ 1'b0 ;
  assign n17375 = n487 | n4603 ;
  assign n17376 = n10732 ^ n5899 ^ 1'b0 ;
  assign n17377 = ~n15001 & n17376 ;
  assign n17378 = n11845 & ~n17377 ;
  assign n17379 = n9164 & ~n11099 ;
  assign n17380 = n16024 ^ n6009 ^ 1'b0 ;
  assign n17381 = ( n1865 & n3990 ) | ( n1865 & n7612 ) | ( n3990 & n7612 ) ;
  assign n17382 = n17381 ^ n12368 ^ 1'b0 ;
  assign n17383 = n4379 | n6919 ;
  assign n17384 = n17383 ^ n1627 ^ 1'b0 ;
  assign n17385 = ( n4468 & n14409 ) | ( n4468 & ~n17384 ) | ( n14409 & ~n17384 ) ;
  assign n17386 = n16858 | n17385 ;
  assign n17387 = n165 | n15144 ;
  assign n17388 = n16104 & ~n17387 ;
  assign n17389 = n1853 & ~n4753 ;
  assign n17390 = n2984 & n17389 ;
  assign n17391 = n17390 ^ n2070 ^ 1'b0 ;
  assign n17392 = n16612 ^ n11437 ^ n3280 ;
  assign n17393 = n3460 ^ n2222 ^ 1'b0 ;
  assign n17394 = n8800 | n17393 ;
  assign n17395 = n10979 | n15667 ;
  assign n17396 = n11985 & ~n17395 ;
  assign n17397 = n5669 & ~n12774 ;
  assign n17398 = n10105 & n17397 ;
  assign n17399 = n10577 ^ n1847 ^ 1'b0 ;
  assign n17400 = ~n13008 & n17399 ;
  assign n17401 = n16102 & n17400 ;
  assign n17402 = n11995 & n17401 ;
  assign n17407 = n2116 ^ n1619 ^ 1'b0 ;
  assign n17408 = n2848 & ~n17407 ;
  assign n17403 = n5857 & n7851 ;
  assign n17404 = n8682 ^ n4834 ^ 1'b0 ;
  assign n17405 = n17403 & n17404 ;
  assign n17406 = ~n10627 & n17405 ;
  assign n17409 = n17408 ^ n17406 ^ 1'b0 ;
  assign n17410 = n2882 & ~n5632 ;
  assign n17411 = n6715 & n17410 ;
  assign n17412 = n15935 ^ n7788 ^ n4287 ;
  assign n17413 = n4352 & ~n17412 ;
  assign n17414 = ~n11797 & n17413 ;
  assign n17415 = n8504 ^ n3690 ^ 1'b0 ;
  assign n17416 = n738 & n8719 ;
  assign n17417 = ~n17415 & n17416 ;
  assign n17418 = n9053 & ~n17417 ;
  assign n17419 = n1229 & n7192 ;
  assign n17420 = n3365 ^ n1899 ^ 1'b0 ;
  assign n17421 = n3662 & ~n17420 ;
  assign n17422 = ~n5992 & n9520 ;
  assign n17423 = n17421 & ~n17422 ;
  assign n17424 = n17423 ^ n894 ^ 1'b0 ;
  assign n17425 = n17228 ^ n6478 ^ n4021 ;
  assign n17426 = n521 & ~n2026 ;
  assign n17427 = n11870 & ~n17426 ;
  assign n17428 = n17421 ^ n12565 ^ 1'b0 ;
  assign n17429 = n4506 | n17428 ;
  assign n17430 = n17429 ^ n5404 ^ 1'b0 ;
  assign n17431 = ~n3572 & n17430 ;
  assign n17432 = ~n732 & n6871 ;
  assign n17433 = n1957 & n17432 ;
  assign n17434 = n13253 & ~n17433 ;
  assign n17435 = ~n2024 & n3859 ;
  assign n17436 = n10040 ^ n792 ^ 1'b0 ;
  assign n17438 = n7036 ^ n4145 ^ 1'b0 ;
  assign n17437 = ~n10368 & n12728 ;
  assign n17439 = n17438 ^ n17437 ^ n3474 ;
  assign n17440 = n3300 ^ n1880 ^ 1'b0 ;
  assign n17441 = n7217 & n17440 ;
  assign n17442 = n4520 & ~n13692 ;
  assign n17443 = n1250 & n17442 ;
  assign n17444 = ~n1537 & n17443 ;
  assign n17445 = n17444 ^ n7043 ^ 1'b0 ;
  assign n17446 = n17445 ^ n4334 ^ 1'b0 ;
  assign n17447 = n11916 ^ n4370 ^ 1'b0 ;
  assign n17448 = n11131 ^ n4323 ^ 1'b0 ;
  assign n17449 = n6277 ^ n5349 ^ 1'b0 ;
  assign n17450 = n5791 & n17449 ;
  assign n17451 = n10758 ^ n1040 ^ 1'b0 ;
  assign n17452 = n17451 ^ n7298 ^ 1'b0 ;
  assign n17453 = n6414 | n17452 ;
  assign n17455 = n1308 & ~n8946 ;
  assign n17456 = n17455 ^ n5061 ^ 1'b0 ;
  assign n17454 = n5666 & n6785 ;
  assign n17457 = n17456 ^ n17454 ^ 1'b0 ;
  assign n17458 = n14147 ^ n7816 ^ 1'b0 ;
  assign n17459 = n17457 & ~n17458 ;
  assign n17460 = n1235 | n17459 ;
  assign n17461 = n1277 & ~n8310 ;
  assign n17462 = ( n662 & n5358 ) | ( n662 & n15310 ) | ( n5358 & n15310 ) ;
  assign n17463 = n208 | n6863 ;
  assign n17464 = n2890 & n10338 ;
  assign n17465 = n17464 ^ n3391 ^ 1'b0 ;
  assign n17466 = n12425 | n17465 ;
  assign n17467 = n6133 & ~n17466 ;
  assign n17468 = n14596 ^ n7688 ^ 1'b0 ;
  assign n17469 = ~n1329 & n3697 ;
  assign n17470 = ~n8691 & n17469 ;
  assign n17471 = n138 & ~n6474 ;
  assign n17472 = n17471 ^ n16667 ^ 1'b0 ;
  assign n17473 = ~n17470 & n17472 ;
  assign n17474 = n2340 & n7987 ;
  assign n17475 = n17474 ^ n15827 ^ 1'b0 ;
  assign n17476 = ( n1995 & ~n3888 ) | ( n1995 & n17475 ) | ( ~n3888 & n17475 ) ;
  assign n17477 = n7644 | n17476 ;
  assign n17478 = n17477 ^ n10173 ^ n2365 ;
  assign n17479 = n5813 & ~n10401 ;
  assign n17480 = ~n9850 & n16269 ;
  assign n17481 = n13754 ^ n5374 ^ 1'b0 ;
  assign n17482 = n342 & n12491 ;
  assign n17483 = n17482 ^ n11406 ^ 1'b0 ;
  assign n17484 = n1920 | n3229 ;
  assign n17485 = n17484 ^ n9265 ^ 1'b0 ;
  assign n17486 = n3289 | n4153 ;
  assign n17487 = n17486 ^ n565 ^ 1'b0 ;
  assign n17488 = n17487 ^ n2953 ^ n1537 ;
  assign n17489 = n9066 & n10469 ;
  assign n17490 = n7788 | n15260 ;
  assign n17491 = n17489 | n17490 ;
  assign n17492 = ~n2633 & n10433 ;
  assign n17493 = n17492 ^ n6787 ^ 1'b0 ;
  assign n17494 = n11961 ^ n9555 ^ 1'b0 ;
  assign n17495 = ~n7288 & n17494 ;
  assign n17496 = n15415 ^ n11181 ^ 1'b0 ;
  assign n17497 = n13713 ^ n3731 ^ n2924 ;
  assign n17498 = n1325 & ~n13933 ;
  assign n17499 = n10453 & ~n17498 ;
  assign n17500 = n15701 ^ n7693 ^ 1'b0 ;
  assign n17501 = n347 & n6790 ;
  assign n17502 = n17501 ^ n395 ^ 1'b0 ;
  assign n17503 = n10408 | n14688 ;
  assign n17504 = n17503 ^ n5592 ^ 1'b0 ;
  assign n17505 = n12391 & n17504 ;
  assign n17506 = n17502 & n17505 ;
  assign n17507 = n5000 & n15884 ;
  assign n17508 = n2082 & n17507 ;
  assign n17510 = n8309 ^ n5311 ^ 1'b0 ;
  assign n17509 = ~n4730 & n6437 ;
  assign n17511 = n17510 ^ n17509 ^ 1'b0 ;
  assign n17512 = ( n773 & ~n3367 ) | ( n773 & n5564 ) | ( ~n3367 & n5564 ) ;
  assign n17513 = n3219 ^ n1115 ^ 1'b0 ;
  assign n17514 = n1159 | n3489 ;
  assign n17515 = n9365 ^ n2348 ^ 1'b0 ;
  assign n17516 = n17514 | n17515 ;
  assign n17517 = n1467 | n9246 ;
  assign n17518 = n13358 ^ n1359 ^ 1'b0 ;
  assign n17519 = n17517 | n17518 ;
  assign n17520 = n16789 ^ n6109 ^ 1'b0 ;
  assign n17521 = n11645 | n13798 ;
  assign n17522 = n17521 ^ n4287 ^ 1'b0 ;
  assign n17523 = n8490 & n14732 ;
  assign n17524 = ~n2371 & n8608 ;
  assign n17525 = ~n950 & n6355 ;
  assign n17526 = ~n14189 & n15474 ;
  assign n17527 = ( ~n9025 & n12057 ) | ( ~n9025 & n17526 ) | ( n12057 & n17526 ) ;
  assign n17528 = n8588 ^ n3434 ^ 1'b0 ;
  assign n17529 = n6249 & ~n12865 ;
  assign n17530 = n7380 ^ n2020 ^ 1'b0 ;
  assign n17531 = n2084 ^ n651 ^ 1'b0 ;
  assign n17532 = n7249 | n17531 ;
  assign n17533 = n17532 ^ n7432 ^ 1'b0 ;
  assign n17534 = n3945 & ~n11275 ;
  assign n17535 = n17534 ^ x58 ^ 1'b0 ;
  assign n17536 = ~n17533 & n17535 ;
  assign n17537 = ~n6827 & n14969 ;
  assign n17538 = n17537 ^ n5952 ^ 1'b0 ;
  assign n17539 = n13027 ^ n1040 ^ 1'b0 ;
  assign n17540 = n614 & n16595 ;
  assign n17541 = n17540 ^ n6504 ^ 1'b0 ;
  assign n17542 = n17541 ^ n4876 ^ 1'b0 ;
  assign n17543 = n14708 & ~n17542 ;
  assign n17544 = n12964 ^ n9632 ^ 1'b0 ;
  assign n17545 = n10429 ^ n4215 ^ 1'b0 ;
  assign n17546 = ~n6331 & n17545 ;
  assign n17547 = ( ~n646 & n740 ) | ( ~n646 & n1289 ) | ( n740 & n1289 ) ;
  assign n17548 = n3310 & n17547 ;
  assign n17549 = ~n17546 & n17548 ;
  assign n17550 = n17549 ^ n10970 ^ n7649 ;
  assign n17553 = n5086 & ~n6037 ;
  assign n17554 = n17553 ^ n9596 ^ 1'b0 ;
  assign n17551 = n16485 ^ n231 ^ 1'b0 ;
  assign n17552 = ~n9097 & n17551 ;
  assign n17555 = n17554 ^ n17552 ^ x98 ;
  assign n17556 = n5368 | n6575 ;
  assign n17557 = n12240 ^ n3936 ^ 1'b0 ;
  assign n17558 = n9949 & ~n17557 ;
  assign n17559 = n13817 ^ n7805 ^ 1'b0 ;
  assign n17560 = n17559 ^ n5644 ^ n4640 ;
  assign n17561 = n7720 ^ n5243 ^ 1'b0 ;
  assign n17562 = n4419 & ~n17561 ;
  assign n17564 = ~n3053 & n8887 ;
  assign n17565 = n6608 & n17564 ;
  assign n17566 = n17565 ^ n7259 ^ 1'b0 ;
  assign n17563 = n1159 & ~n2685 ;
  assign n17567 = n17566 ^ n17563 ^ 1'b0 ;
  assign n17568 = ~n1637 & n7527 ;
  assign n17569 = n6415 | n17411 ;
  assign n17570 = n17569 ^ n15201 ^ 1'b0 ;
  assign n17571 = n7485 | n13153 ;
  assign n17572 = n17571 ^ n7587 ^ 1'b0 ;
  assign n17573 = n6695 & n13465 ;
  assign n17574 = n17573 ^ n7612 ^ 1'b0 ;
  assign n17575 = n3248 ^ n2824 ^ 1'b0 ;
  assign n17576 = n5232 | n17575 ;
  assign n17577 = ~n7042 & n13941 ;
  assign n17578 = n17577 ^ x37 ^ 1'b0 ;
  assign n17579 = n16354 ^ n12300 ^ 1'b0 ;
  assign n17580 = n12541 ^ n1217 ^ 1'b0 ;
  assign n17581 = n17579 & ~n17580 ;
  assign n17582 = n8541 ^ n3672 ^ n3215 ;
  assign n17583 = n12816 ^ n2638 ^ 1'b0 ;
  assign n17584 = n11246 ^ n5297 ^ 1'b0 ;
  assign n17585 = n7578 ^ n4949 ^ 1'b0 ;
  assign n17586 = n17585 ^ n4979 ^ 1'b0 ;
  assign n17587 = n17584 | n17586 ;
  assign n17588 = ~n5294 & n12734 ;
  assign n17589 = n11125 & n17588 ;
  assign n17590 = n16181 ^ n7419 ^ 1'b0 ;
  assign n17591 = n17590 ^ n1676 ^ 1'b0 ;
  assign n17592 = ( n1718 & n17385 ) | ( n1718 & n17591 ) | ( n17385 & n17591 ) ;
  assign n17593 = ( ~n3842 & n5018 ) | ( ~n3842 & n17592 ) | ( n5018 & n17592 ) ;
  assign n17594 = n11766 ^ n1355 ^ 1'b0 ;
  assign n17595 = n16981 ^ n2489 ^ 1'b0 ;
  assign n17596 = n10226 | n17595 ;
  assign n17597 = n2984 & n12481 ;
  assign n17598 = n17597 ^ n16378 ^ 1'b0 ;
  assign n17599 = n14960 ^ n10131 ^ 1'b0 ;
  assign n17600 = n10665 & ~n12564 ;
  assign n17601 = ~n11327 & n17600 ;
  assign n17602 = n1878 & ~n10106 ;
  assign n17603 = n4696 & n11034 ;
  assign n17604 = n17477 ^ n16267 ^ n634 ;
  assign n17605 = n4555 & ~n5048 ;
  assign n17606 = n17605 ^ n1824 ^ 1'b0 ;
  assign n17607 = n4759 & ~n17606 ;
  assign n17608 = n5983 ^ n3404 ^ 1'b0 ;
  assign n17609 = n7893 & n17608 ;
  assign n17610 = n4097 & ~n5747 ;
  assign n17611 = ~n3674 & n17610 ;
  assign n17612 = ~n17609 & n17611 ;
  assign n17613 = ~n1438 & n9151 ;
  assign n17614 = n5732 & ~n12453 ;
  assign n17615 = n4253 ^ n2543 ^ 1'b0 ;
  assign n17616 = n9522 ^ n3722 ^ 1'b0 ;
  assign n17617 = n16015 & n17616 ;
  assign n17618 = n11677 ^ n3054 ^ n324 ;
  assign n17619 = x42 | n2185 ;
  assign n17620 = n8911 ^ n8331 ^ 1'b0 ;
  assign n17621 = n14673 & n17620 ;
  assign n17622 = ~n3762 & n17621 ;
  assign n17623 = n15696 & n17622 ;
  assign n17624 = n540 & n2042 ;
  assign n17625 = n5037 & n17624 ;
  assign n17626 = ~n10526 & n13377 ;
  assign n17627 = ~n4979 & n17626 ;
  assign n17628 = ( ~n2196 & n12970 ) | ( ~n2196 & n17627 ) | ( n12970 & n17627 ) ;
  assign n17629 = n676 | n2278 ;
  assign n17630 = n676 & ~n17629 ;
  assign n17631 = n7303 ^ n2228 ^ 1'b0 ;
  assign n17632 = n2828 & ~n16437 ;
  assign n17633 = n4662 & ~n15320 ;
  assign n17634 = ~n4831 & n17633 ;
  assign n17635 = n4447 ^ n4045 ^ 1'b0 ;
  assign n17636 = n6649 | n17635 ;
  assign n17637 = n2405 & ~n17636 ;
  assign n17638 = ~n7755 & n17637 ;
  assign n17639 = n17638 ^ n6108 ^ n1992 ;
  assign n17640 = n17639 ^ n12625 ^ n3653 ;
  assign n17641 = n851 & ~n15789 ;
  assign n17642 = ~n6639 & n17641 ;
  assign n17643 = ( n8458 & ~n17640 ) | ( n8458 & n17642 ) | ( ~n17640 & n17642 ) ;
  assign n17644 = n2491 & n3321 ;
  assign n17645 = n1079 | n5739 ;
  assign n17646 = n17645 ^ n2434 ^ 1'b0 ;
  assign n17647 = n9101 | n9694 ;
  assign n17648 = n8820 ^ n2042 ^ n464 ;
  assign n17649 = n15708 ^ n11121 ^ 1'b0 ;
  assign n17650 = n10246 | n17649 ;
  assign n17651 = n7100 & ~n13754 ;
  assign n17652 = n17650 & ~n17651 ;
  assign n17653 = ~n5214 & n17652 ;
  assign n17654 = n17653 ^ n10552 ^ 1'b0 ;
  assign n17655 = n719 & n8946 ;
  assign n17656 = n3962 & n17655 ;
  assign n17657 = ~n8801 & n11577 ;
  assign n17658 = n9823 & n17657 ;
  assign n17659 = n13285 | n17658 ;
  assign n17660 = n3601 & ~n17659 ;
  assign n17661 = n14381 ^ n1943 ^ 1'b0 ;
  assign n17662 = ( x99 & x107 ) | ( x99 & n10276 ) | ( x107 & n10276 ) ;
  assign n17663 = n11828 ^ n8123 ^ n2958 ;
  assign n17664 = ~n3138 & n17663 ;
  assign n17665 = n12736 ^ n7529 ^ n5840 ;
  assign n17666 = n5963 ^ n3798 ^ 1'b0 ;
  assign n17667 = n17665 & n17666 ;
  assign n17668 = n5288 | n6206 ;
  assign n17669 = n6791 & ~n17668 ;
  assign n17670 = n17669 ^ n7447 ^ 1'b0 ;
  assign n17671 = n8637 ^ n5974 ^ 1'b0 ;
  assign n17672 = n525 & n17671 ;
  assign n17673 = n3542 | n17672 ;
  assign n17681 = x59 & ~n5362 ;
  assign n17674 = ( n1229 & n8181 ) | ( n1229 & ~n10399 ) | ( n8181 & ~n10399 ) ;
  assign n17675 = ( n525 & n9800 ) | ( n525 & ~n17674 ) | ( n9800 & ~n17674 ) ;
  assign n17676 = ~n1398 & n17675 ;
  assign n17677 = n9960 & n17676 ;
  assign n17678 = ( n5248 & ~n14123 ) | ( n5248 & n17677 ) | ( ~n14123 & n17677 ) ;
  assign n17679 = ~n9985 & n17678 ;
  assign n17680 = n1840 & n17679 ;
  assign n17682 = n17681 ^ n17680 ^ 1'b0 ;
  assign n17683 = n1211 & ~n17682 ;
  assign n17684 = n14348 ^ n8119 ^ 1'b0 ;
  assign n17685 = ~n15500 & n17684 ;
  assign n17686 = n8435 & n10109 ;
  assign n17687 = ~n4979 & n17686 ;
  assign n17688 = ( n1308 & n6490 ) | ( n1308 & n9915 ) | ( n6490 & n9915 ) ;
  assign n17689 = x112 & ~n14713 ;
  assign n17690 = n17689 ^ n1495 ^ 1'b0 ;
  assign n17691 = n13002 ^ n3714 ^ 1'b0 ;
  assign n17692 = n7863 | n17691 ;
  assign n17700 = n4652 | n5883 ;
  assign n17701 = n10952 | n17700 ;
  assign n17693 = n1027 & ~n6936 ;
  assign n17694 = ~n1027 & n17693 ;
  assign n17695 = n6340 & ~n17694 ;
  assign n17696 = n3651 & n17695 ;
  assign n17697 = n3583 & ~n17696 ;
  assign n17698 = n13569 & n17697 ;
  assign n17699 = n5419 & ~n17698 ;
  assign n17702 = n17701 ^ n17699 ^ 1'b0 ;
  assign n17703 = n9141 | n11114 ;
  assign n17704 = n17703 ^ n2235 ^ 1'b0 ;
  assign n17705 = n17704 ^ n7449 ^ 1'b0 ;
  assign n17706 = n13144 & ~n17705 ;
  assign n17708 = n5211 | n5522 ;
  assign n17707 = n323 & ~n15867 ;
  assign n17709 = n17708 ^ n17707 ^ 1'b0 ;
  assign n17710 = n13957 ^ n9021 ^ 1'b0 ;
  assign n17711 = n17709 & ~n17710 ;
  assign n17712 = n9301 ^ n8496 ^ 1'b0 ;
  assign n17713 = ( n2636 & ~n12737 ) | ( n2636 & n17712 ) | ( ~n12737 & n17712 ) ;
  assign n17714 = ~n2240 & n17713 ;
  assign n17715 = n1408 & n17714 ;
  assign n17716 = ~n4205 & n5652 ;
  assign n17717 = n17716 ^ n177 ^ 1'b0 ;
  assign n17718 = n5370 & n5906 ;
  assign n17719 = n6807 ^ n6124 ^ 1'b0 ;
  assign n17720 = n9624 | n12796 ;
  assign n17721 = n5205 & ~n6862 ;
  assign n17722 = ~n2466 & n17721 ;
  assign n17723 = n2235 & n2619 ;
  assign n17724 = ~n10683 & n13794 ;
  assign n17725 = ~n5410 & n17724 ;
  assign n17726 = ( n10860 & n17723 ) | ( n10860 & ~n17725 ) | ( n17723 & ~n17725 ) ;
  assign n17727 = n10752 ^ n1686 ^ 1'b0 ;
  assign n17728 = n16720 ^ n8513 ^ 1'b0 ;
  assign n17729 = x117 & ~n1089 ;
  assign n17730 = ~n7488 & n17729 ;
  assign n17731 = n3528 & n17730 ;
  assign n17732 = n2389 ^ n1392 ^ 1'b0 ;
  assign n17733 = ~n17731 & n17732 ;
  assign n17735 = ( n3597 & n7032 ) | ( n3597 & ~n7386 ) | ( n7032 & ~n7386 ) ;
  assign n17734 = ~n2134 & n2996 ;
  assign n17736 = n17735 ^ n17734 ^ 1'b0 ;
  assign n17737 = n630 ^ x65 ^ 1'b0 ;
  assign n17739 = ~n6120 & n9892 ;
  assign n17738 = ~n5310 & n11577 ;
  assign n17740 = n17739 ^ n17738 ^ 1'b0 ;
  assign n17741 = ~n17737 & n17740 ;
  assign n17744 = n5576 ^ n1642 ^ 1'b0 ;
  assign n17745 = x13 & ~n17744 ;
  assign n17746 = n17745 ^ n5463 ^ 1'b0 ;
  assign n17742 = n7705 ^ n7187 ^ 1'b0 ;
  assign n17743 = n13249 & n17742 ;
  assign n17747 = n17746 ^ n17743 ^ n10554 ;
  assign n17748 = n6741 & ~n16184 ;
  assign n17749 = n3203 | n11560 ;
  assign n17750 = ( n3881 & n7343 ) | ( n3881 & ~n11036 ) | ( n7343 & ~n11036 ) ;
  assign n17751 = ~n4923 & n12422 ;
  assign n17752 = n3112 & n17751 ;
  assign n17753 = ~n17750 & n17752 ;
  assign n17755 = n12935 ^ n2103 ^ 1'b0 ;
  assign n17756 = n4048 | n17755 ;
  assign n17754 = ( n11071 & n11574 ) | ( n11071 & ~n17120 ) | ( n11574 & ~n17120 ) ;
  assign n17757 = n17756 ^ n17754 ^ n7606 ;
  assign n17758 = n1747 | n6451 ;
  assign n17759 = n17758 ^ n2998 ^ 1'b0 ;
  assign n17760 = n2210 & n8722 ;
  assign n17761 = n17760 ^ n8613 ^ 1'b0 ;
  assign n17762 = n15152 | n17316 ;
  assign n17763 = n2523 & ~n17762 ;
  assign n17764 = n8377 ^ n6207 ^ 1'b0 ;
  assign n17765 = n17764 ^ n12349 ^ 1'b0 ;
  assign n17766 = n882 & n5752 ;
  assign n17771 = n4233 | n16974 ;
  assign n17772 = n17771 ^ n4917 ^ 1'b0 ;
  assign n17767 = n2872 | n12034 ;
  assign n17768 = n17767 ^ n5161 ^ 1'b0 ;
  assign n17769 = n6333 & n17768 ;
  assign n17770 = n2742 & n17769 ;
  assign n17773 = n17772 ^ n17770 ^ 1'b0 ;
  assign n17774 = ( n2628 & n4798 ) | ( n2628 & ~n5357 ) | ( n4798 & ~n5357 ) ;
  assign n17775 = n14204 & n17774 ;
  assign n17776 = n17775 ^ n16893 ^ 1'b0 ;
  assign n17777 = n2595 ^ n1716 ^ 1'b0 ;
  assign n17778 = n7475 ^ n3207 ^ n1077 ;
  assign n17779 = n5623 ^ n1338 ^ 1'b0 ;
  assign n17780 = n17778 & ~n17779 ;
  assign n17781 = n2693 ^ n1566 ^ 1'b0 ;
  assign n17782 = n3841 | n17781 ;
  assign n17783 = n17782 ^ n6403 ^ 1'b0 ;
  assign n17784 = n16413 ^ n7042 ^ n5079 ;
  assign n17785 = n15706 ^ n11107 ^ 1'b0 ;
  assign n17786 = n2611 | n9666 ;
  assign n17787 = n560 | n17786 ;
  assign n17788 = n16382 ^ n16113 ^ 1'b0 ;
  assign n17789 = n17787 & n17788 ;
  assign n17790 = n7643 ^ n3603 ^ 1'b0 ;
  assign n17791 = ( n9781 & n12782 ) | ( n9781 & n17790 ) | ( n12782 & n17790 ) ;
  assign n17792 = ~n6053 & n11537 ;
  assign n17793 = n17792 ^ n4575 ^ 1'b0 ;
  assign n17794 = n5944 & n17793 ;
  assign n17795 = n8062 ^ n2222 ^ 1'b0 ;
  assign n17796 = ~n7258 & n17795 ;
  assign n17797 = n17796 ^ n11928 ^ 1'b0 ;
  assign n17798 = n4105 ^ n3974 ^ 1'b0 ;
  assign n17799 = n7360 | n17798 ;
  assign n17800 = ~n5634 & n9724 ;
  assign n17801 = n2353 ^ n1529 ^ 1'b0 ;
  assign n17802 = n17801 ^ n1740 ^ 1'b0 ;
  assign n17803 = n14163 ^ n8906 ^ n2702 ;
  assign n17804 = n15406 ^ n1562 ^ 1'b0 ;
  assign n17805 = n4037 & ~n13274 ;
  assign n17806 = n8569 & n17805 ;
  assign n17807 = n240 & ~n799 ;
  assign n17808 = n11308 & ~n17807 ;
  assign n17809 = ~n17504 & n17808 ;
  assign n17810 = n17809 ^ n1700 ^ 1'b0 ;
  assign n17811 = n17806 & n17810 ;
  assign n17812 = n7465 & n17029 ;
  assign n17813 = n10885 & n17812 ;
  assign n17814 = n5840 & n8454 ;
  assign n17815 = n11512 & n17814 ;
  assign n17816 = n3407 & ~n14161 ;
  assign n17817 = ( n16165 & n17815 ) | ( n16165 & n17816 ) | ( n17815 & n17816 ) ;
  assign n17818 = n718 & n7457 ;
  assign n17819 = n13904 & n17818 ;
  assign n17820 = n14480 ^ n131 ^ 1'b0 ;
  assign n17821 = n5791 & n17820 ;
  assign n17823 = n10997 ^ n5762 ^ 1'b0 ;
  assign n17822 = n4063 & n8936 ;
  assign n17824 = n17823 ^ n17822 ^ 1'b0 ;
  assign n17825 = n10457 & ~n17824 ;
  assign n17826 = n8468 & n13853 ;
  assign n17827 = n17826 ^ n5551 ^ 1'b0 ;
  assign n17828 = n623 & ~n11208 ;
  assign n17829 = ( ~n632 & n9146 ) | ( ~n632 & n17828 ) | ( n9146 & n17828 ) ;
  assign n17830 = ( x71 & n254 ) | ( x71 & n16351 ) | ( n254 & n16351 ) ;
  assign n17831 = n9847 ^ n468 ^ 1'b0 ;
  assign n17832 = n15164 & n17831 ;
  assign n17833 = n3458 & ~n9942 ;
  assign n17834 = ~n13971 & n17833 ;
  assign n17835 = n3772 & n17834 ;
  assign n17836 = n16360 | n17835 ;
  assign n17837 = n11032 & ~n17836 ;
  assign n17838 = n6399 & ~n7436 ;
  assign n17839 = n17838 ^ n3226 ^ 1'b0 ;
  assign n17840 = ( n11096 & ~n12409 ) | ( n11096 & n17839 ) | ( ~n12409 & n17839 ) ;
  assign n17841 = n7641 & n12391 ;
  assign n17842 = n7727 ^ n5733 ^ 1'b0 ;
  assign n17843 = ~n16053 & n17842 ;
  assign n17844 = n1691 & n4564 ;
  assign n17845 = n17844 ^ n9066 ^ 1'b0 ;
  assign n17846 = n13565 & ~n17845 ;
  assign n17847 = n17846 ^ n6844 ^ 1'b0 ;
  assign n17848 = n6013 ^ n1015 ^ 1'b0 ;
  assign n17849 = n4200 ^ n3016 ^ 1'b0 ;
  assign n17850 = n5253 & n17849 ;
  assign n17851 = n5494 | n17850 ;
  assign n17853 = n888 & n9511 ;
  assign n17854 = n17853 ^ n9529 ^ 1'b0 ;
  assign n17852 = ~n1263 & n15860 ;
  assign n17855 = n17854 ^ n17852 ^ 1'b0 ;
  assign n17856 = n17855 ^ n8565 ^ 1'b0 ;
  assign n17857 = n17851 & ~n17856 ;
  assign n17858 = n12025 & n17857 ;
  assign n17859 = ~n6227 & n7401 ;
  assign n17860 = n17859 ^ n4606 ^ n973 ;
  assign n17861 = n2327 & ~n3590 ;
  assign n17862 = n8396 & n17861 ;
  assign n17863 = ~n15178 & n17862 ;
  assign n17864 = n8282 & n15338 ;
  assign n17865 = n17864 ^ n15392 ^ 1'b0 ;
  assign n17866 = n9651 ^ n767 ^ 1'b0 ;
  assign n17867 = n13005 & ~n13417 ;
  assign n17871 = x69 & ~n11056 ;
  assign n17868 = ~n3240 & n6688 ;
  assign n17869 = n17868 ^ n3518 ^ 1'b0 ;
  assign n17870 = n7840 & n17869 ;
  assign n17872 = n17871 ^ n17870 ^ 1'b0 ;
  assign n17873 = n11948 ^ n4307 ^ 1'b0 ;
  assign n17874 = n11750 ^ n1982 ^ n334 ;
  assign n17875 = n883 & ~n2972 ;
  assign n17876 = n1767 & n17875 ;
  assign n17877 = n1401 | n5678 ;
  assign n17878 = n17876 & ~n17877 ;
  assign n17879 = ~n4324 & n8086 ;
  assign n17880 = n9616 ^ n362 ^ 1'b0 ;
  assign n17881 = n17879 & n17880 ;
  assign n17882 = n3033 | n11339 ;
  assign n17883 = n13608 ^ n11081 ^ n5302 ;
  assign n17884 = n4938 | n17883 ;
  assign n17885 = n801 | n17884 ;
  assign n17886 = n6454 ^ n4553 ^ n423 ;
  assign n17887 = ( n2222 & ~n3582 ) | ( n2222 & n17886 ) | ( ~n3582 & n17886 ) ;
  assign n17888 = ~n1306 & n1853 ;
  assign n17889 = n17888 ^ n5034 ^ n641 ;
  assign n17890 = ( n297 & n4798 ) | ( n297 & ~n17154 ) | ( n4798 & ~n17154 ) ;
  assign n17891 = ( ~n2961 & n17889 ) | ( ~n2961 & n17890 ) | ( n17889 & n17890 ) ;
  assign n17892 = n10888 ^ n1378 ^ 1'b0 ;
  assign n17893 = n15339 & n17892 ;
  assign n17894 = ~n6557 & n14369 ;
  assign n17895 = n3973 & n17894 ;
  assign n17896 = n17895 ^ n6754 ^ 1'b0 ;
  assign n17897 = n7739 | n17896 ;
  assign n17898 = n12799 ^ n5687 ^ 1'b0 ;
  assign n17899 = ~n7030 & n12287 ;
  assign n17900 = n17899 ^ n4957 ^ 1'b0 ;
  assign n17901 = n17900 ^ n10689 ^ 1'b0 ;
  assign n17902 = n13289 ^ n5064 ^ 1'b0 ;
  assign n17903 = n12724 ^ n5261 ^ 1'b0 ;
  assign n17904 = n2742 & ~n17903 ;
  assign n17905 = n17902 & n17904 ;
  assign n17906 = n17905 ^ n3405 ^ 1'b0 ;
  assign n17907 = x107 | n13370 ;
  assign n17908 = n4142 ^ n2673 ^ 1'b0 ;
  assign n17909 = n8215 & n13215 ;
  assign n17910 = n17909 ^ n6814 ^ 1'b0 ;
  assign n17911 = n10008 & ~n16824 ;
  assign n17912 = n17911 ^ n8396 ^ 1'b0 ;
  assign n17913 = n15750 ^ n13249 ^ 1'b0 ;
  assign n17914 = n14085 ^ n6321 ^ n357 ;
  assign n17915 = n9389 | n17914 ;
  assign n17916 = n3965 | n4039 ;
  assign n17917 = n17915 & n17916 ;
  assign n17918 = n2280 & ~n8719 ;
  assign n17919 = n17855 ^ n8476 ^ 1'b0 ;
  assign n17920 = ~n8864 & n17919 ;
  assign n17921 = ( ~n4327 & n7876 ) | ( ~n4327 & n9503 ) | ( n7876 & n9503 ) ;
  assign n17922 = n17921 ^ n12291 ^ 1'b0 ;
  assign n17923 = n16104 & n17922 ;
  assign n17927 = n4121 ^ n2356 ^ n1204 ;
  assign n17928 = n3183 | n17927 ;
  assign n17929 = n5020 ^ x70 ^ 1'b0 ;
  assign n17930 = n17928 & ~n17929 ;
  assign n17925 = n3950 & ~n15500 ;
  assign n17926 = ~n2790 & n17925 ;
  assign n17931 = n17930 ^ n17926 ^ n2832 ;
  assign n17932 = ( n9033 & n10111 ) | ( n9033 & ~n17931 ) | ( n10111 & ~n17931 ) ;
  assign n17933 = n5855 & n17932 ;
  assign n17934 = ~n10472 & n17933 ;
  assign n17924 = n4832 | n11224 ;
  assign n17935 = n17934 ^ n17924 ^ 1'b0 ;
  assign n17936 = n4507 & ~n8073 ;
  assign n17937 = n2963 | n6156 ;
  assign n17938 = n17937 ^ n406 ^ 1'b0 ;
  assign n17939 = ~n8167 & n13788 ;
  assign n17940 = n15473 & n17939 ;
  assign n17941 = n7512 ^ n5654 ^ 1'b0 ;
  assign n17942 = ~n709 & n10029 ;
  assign n17943 = ~n17941 & n17942 ;
  assign n17944 = n5914 ^ n3278 ^ 1'b0 ;
  assign n17945 = n3477 & n17944 ;
  assign n17946 = n11339 | n17945 ;
  assign n17947 = n1489 & ~n6597 ;
  assign n17948 = ~n17946 & n17947 ;
  assign n17949 = n12887 ^ x30 ^ 1'b0 ;
  assign n17950 = n2401 | n17949 ;
  assign n17951 = n17859 | n17950 ;
  assign n17952 = n11488 | n17951 ;
  assign n17953 = n5725 ^ n453 ^ 1'b0 ;
  assign n17954 = n7998 & n17953 ;
  assign n17955 = n6354 & n17954 ;
  assign n17956 = n17955 ^ n9048 ^ 1'b0 ;
  assign n17957 = n9865 & n17956 ;
  assign n17958 = n8292 ^ n4592 ^ 1'b0 ;
  assign n17959 = n1197 | n7991 ;
  assign n17960 = n17959 ^ n4645 ^ 1'b0 ;
  assign n17961 = n17960 ^ n303 ^ 1'b0 ;
  assign n17962 = n17961 ^ n1812 ^ 1'b0 ;
  assign n17963 = n17962 ^ n12309 ^ 1'b0 ;
  assign n17964 = n15056 | n15454 ;
  assign n17965 = n17963 & ~n17964 ;
  assign n17966 = ~n4032 & n10657 ;
  assign n17970 = ( ~n556 & n3908 ) | ( ~n556 & n4768 ) | ( n3908 & n4768 ) ;
  assign n17971 = n6805 & n17970 ;
  assign n17972 = ~n7025 & n17971 ;
  assign n17967 = n16680 ^ n4468 ^ 1'b0 ;
  assign n17968 = n10779 & n17967 ;
  assign n17969 = n12763 & n17968 ;
  assign n17973 = n17972 ^ n17969 ^ 1'b0 ;
  assign n17974 = n1790 | n8126 ;
  assign n17975 = ~n10967 & n17974 ;
  assign n17976 = n15755 & n17975 ;
  assign n17977 = n3130 ^ n874 ^ 1'b0 ;
  assign n17978 = n5971 & ~n17977 ;
  assign n17979 = n17978 ^ n8476 ^ 1'b0 ;
  assign n17980 = n13458 ^ n11562 ^ n10656 ;
  assign n17981 = ( ~n281 & n3495 ) | ( ~n281 & n8244 ) | ( n3495 & n8244 ) ;
  assign n17983 = n1941 | n16588 ;
  assign n17984 = n3472 | n17983 ;
  assign n17982 = n3021 & n9696 ;
  assign n17985 = n17984 ^ n17982 ^ 1'b0 ;
  assign n17989 = n6121 ^ n377 ^ 1'b0 ;
  assign n17990 = n13937 ^ n13087 ^ 1'b0 ;
  assign n17991 = n17989 & ~n17990 ;
  assign n17986 = n3087 ^ x0 ^ 1'b0 ;
  assign n17987 = n384 & n17986 ;
  assign n17988 = n17987 ^ n9460 ^ 1'b0 ;
  assign n17992 = n17991 ^ n17988 ^ 1'b0 ;
  assign n17993 = n8880 & n17992 ;
  assign n17994 = n11829 & n15506 ;
  assign n17996 = n8799 ^ n692 ^ 1'b0 ;
  assign n17997 = n400 | n17996 ;
  assign n17995 = ~n8764 & n9215 ;
  assign n17998 = n17997 ^ n17995 ^ 1'b0 ;
  assign n17999 = x45 & ~n5948 ;
  assign n18000 = n16486 ^ n2170 ^ n1159 ;
  assign n18001 = ( n5429 & n17999 ) | ( n5429 & ~n18000 ) | ( n17999 & ~n18000 ) ;
  assign n18002 = n14863 ^ n4647 ^ 1'b0 ;
  assign n18003 = n398 | n18002 ;
  assign n18004 = n18003 ^ n560 ^ 1'b0 ;
  assign n18005 = n4043 | n4117 ;
  assign n18006 = n1971 | n18005 ;
  assign n18007 = n6347 ^ n3491 ^ 1'b0 ;
  assign n18008 = ~n12236 & n18007 ;
  assign n18009 = n18008 ^ n7689 ^ 1'b0 ;
  assign n18010 = n18006 & ~n18009 ;
  assign n18011 = n2788 | n2976 ;
  assign n18012 = n12011 & n15370 ;
  assign n18013 = n7932 ^ n3021 ^ n2436 ;
  assign n18014 = n18013 ^ n400 ^ 1'b0 ;
  assign n18015 = n18014 ^ n12552 ^ n3685 ;
  assign n18016 = n165 & n14969 ;
  assign n18017 = n2339 & n12923 ;
  assign n18018 = n5781 ^ n1129 ^ 1'b0 ;
  assign n18019 = ~n16830 & n18018 ;
  assign n18020 = n3560 & ~n7041 ;
  assign n18021 = ~n15404 & n18020 ;
  assign n18022 = n18021 ^ n4785 ^ 1'b0 ;
  assign n18023 = n6932 & n18022 ;
  assign n18024 = n384 & n7967 ;
  assign n18025 = n13592 ^ n3572 ^ 1'b0 ;
  assign n18026 = ( n3594 & n4251 ) | ( n3594 & ~n6132 ) | ( n4251 & ~n6132 ) ;
  assign n18027 = ( n15197 & n18025 ) | ( n15197 & ~n18026 ) | ( n18025 & ~n18026 ) ;
  assign n18028 = ~n9041 & n15546 ;
  assign n18029 = n18028 ^ n12848 ^ 1'b0 ;
  assign n18030 = n18029 ^ n1722 ^ 1'b0 ;
  assign n18031 = ~n9290 & n18030 ;
  assign n18032 = n6974 ^ n393 ^ 1'b0 ;
  assign n18033 = n4985 & n18032 ;
  assign n18034 = ~n5486 & n18033 ;
  assign n18035 = n3224 ^ n1683 ^ 1'b0 ;
  assign n18036 = n8268 & n18035 ;
  assign n18037 = n10571 ^ n1155 ^ 1'b0 ;
  assign n18038 = n175 | n18037 ;
  assign n18039 = n18036 | n18038 ;
  assign n18040 = ~n2960 & n5093 ;
  assign n18041 = n18040 ^ n17250 ^ 1'b0 ;
  assign n18042 = n6596 ^ n2267 ^ 1'b0 ;
  assign n18043 = n6273 & n18042 ;
  assign n18044 = n18043 ^ n13157 ^ n182 ;
  assign n18045 = n5093 & n13806 ;
  assign n18046 = n18044 & n18045 ;
  assign n18051 = ~n3017 & n9106 ;
  assign n18047 = n192 & n1688 ;
  assign n18048 = n18047 ^ n794 ^ 1'b0 ;
  assign n18049 = n6991 | n14621 ;
  assign n18050 = n18048 & n18049 ;
  assign n18052 = n18051 ^ n18050 ^ 1'b0 ;
  assign n18053 = n6888 & ~n13083 ;
  assign n18054 = n18053 ^ n1526 ^ 1'b0 ;
  assign n18055 = n18052 & n18054 ;
  assign n18059 = ~n3762 & n11258 ;
  assign n18056 = n4997 & n6871 ;
  assign n18057 = ~n5198 & n18056 ;
  assign n18058 = n6403 & ~n18057 ;
  assign n18060 = n18059 ^ n18058 ^ 1'b0 ;
  assign n18061 = n2676 & n5447 ;
  assign n18062 = ~n669 & n18061 ;
  assign n18063 = n411 | n7548 ;
  assign n18064 = n18062 & ~n18063 ;
  assign n18065 = n3873 ^ n476 ^ 1'b0 ;
  assign n18066 = n15966 & ~n18065 ;
  assign n18067 = n4828 ^ n1555 ^ 1'b0 ;
  assign n18068 = n8920 ^ n1588 ^ 1'b0 ;
  assign n18069 = n5516 & ~n10360 ;
  assign n18070 = n18069 ^ n6504 ^ 1'b0 ;
  assign n18071 = n6757 & ~n10043 ;
  assign n18072 = n2632 & n18071 ;
  assign n18073 = n6753 & n10900 ;
  assign n18074 = n1493 & ~n3408 ;
  assign n18075 = n18074 ^ n1027 ^ 1'b0 ;
  assign n18076 = n3804 | n5125 ;
  assign n18077 = n5243 | n18076 ;
  assign n18078 = ( ~n2323 & n18075 ) | ( ~n2323 & n18077 ) | ( n18075 & n18077 ) ;
  assign n18079 = n18078 ^ n8838 ^ 1'b0 ;
  assign n18080 = n16151 ^ n10891 ^ 1'b0 ;
  assign n18081 = n15116 | n18080 ;
  assign n18084 = n3468 ^ n1028 ^ 1'b0 ;
  assign n18082 = n1475 | n2477 ;
  assign n18083 = ~n5941 & n18082 ;
  assign n18085 = n18084 ^ n18083 ^ 1'b0 ;
  assign n18086 = n8695 & n9162 ;
  assign n18087 = n2401 | n4024 ;
  assign n18088 = n18086 | n18087 ;
  assign n18089 = n2905 | n12087 ;
  assign n18090 = n18089 ^ n6233 ^ 1'b0 ;
  assign n18091 = n6889 ^ n5605 ^ 1'b0 ;
  assign n18092 = n2613 & ~n5513 ;
  assign n18093 = n7575 & n18092 ;
  assign n18094 = n4664 | n18093 ;
  assign n18095 = n18094 ^ n10343 ^ 1'b0 ;
  assign n18096 = n3916 & ~n18095 ;
  assign n18097 = n3124 & ~n18096 ;
  assign n18098 = n7130 & n18097 ;
  assign n18099 = n1713 ^ n1476 ^ 1'b0 ;
  assign n18100 = n17270 | n18099 ;
  assign n18101 = ~n3167 & n9000 ;
  assign n18102 = ~n5806 & n18101 ;
  assign n18103 = n730 | n3557 ;
  assign n18104 = n18103 ^ n702 ^ 1'b0 ;
  assign n18105 = n11650 ^ n5776 ^ 1'b0 ;
  assign n18106 = n16397 ^ n15426 ^ 1'b0 ;
  assign n18107 = ~n18105 & n18106 ;
  assign n18108 = n13804 ^ n10045 ^ 1'b0 ;
  assign n18109 = n18107 & n18108 ;
  assign n18110 = n5414 ^ n4638 ^ n2893 ;
  assign n18111 = n3614 & ~n3648 ;
  assign n18112 = x6 | n18111 ;
  assign n18113 = n18110 & ~n18112 ;
  assign n18114 = n15474 ^ n1070 ^ 1'b0 ;
  assign n18115 = n11308 & n18114 ;
  assign n18116 = ~n1624 & n10416 ;
  assign n18117 = n18116 ^ n8657 ^ n1876 ;
  assign n18118 = n12182 & n18117 ;
  assign n18119 = ~n8552 & n16272 ;
  assign n18120 = n18119 ^ n7432 ^ 1'b0 ;
  assign n18121 = n305 & n18120 ;
  assign n18122 = n7865 & ~n15433 ;
  assign n18123 = n2134 & n18122 ;
  assign n18124 = n437 | n18123 ;
  assign n18125 = n1024 & ~n18124 ;
  assign n18126 = n18125 ^ n6156 ^ n6036 ;
  assign n18127 = ~n8442 & n11740 ;
  assign n18128 = ~n7478 & n18127 ;
  assign n18129 = n1483 & ~n11280 ;
  assign n18130 = n505 & n18129 ;
  assign n18131 = ~n3729 & n18130 ;
  assign n18132 = n7048 & ~n9692 ;
  assign n18133 = ~n9868 & n18132 ;
  assign n18134 = n3533 | n3757 ;
  assign n18135 = n5972 & n9200 ;
  assign n18136 = n18135 ^ n3962 ^ 1'b0 ;
  assign n18137 = n12651 ^ n8271 ^ 1'b0 ;
  assign n18138 = n3205 & ~n4448 ;
  assign n18139 = ~n6914 & n18138 ;
  assign n18140 = n3055 & ~n15500 ;
  assign n18141 = n18140 ^ n14022 ^ 1'b0 ;
  assign n18142 = n16640 & ~n18141 ;
  assign n18143 = n1393 & n18142 ;
  assign n18144 = ~n3336 & n14587 ;
  assign n18145 = n18144 ^ n7145 ^ 1'b0 ;
  assign n18146 = n13352 ^ n12913 ^ 1'b0 ;
  assign n18147 = n1241 & n18146 ;
  assign n18148 = n1769 | n14093 ;
  assign n18149 = n6450 | n11277 ;
  assign n18151 = n2195 & ~n13487 ;
  assign n18150 = n2567 & n8601 ;
  assign n18152 = n18151 ^ n18150 ^ n3690 ;
  assign n18153 = n5043 & ~n18152 ;
  assign n18154 = n1529 | n2167 ;
  assign n18155 = ( n9092 & n14299 ) | ( n9092 & n18154 ) | ( n14299 & n18154 ) ;
  assign n18156 = n11990 & ~n18155 ;
  assign n18157 = ~n3877 & n9233 ;
  assign n18158 = n6297 ^ n6124 ^ 1'b0 ;
  assign n18159 = n18157 & n18158 ;
  assign n18160 = n3750 | n4602 ;
  assign n18161 = n18159 | n18160 ;
  assign n18162 = n9402 & n16062 ;
  assign n18163 = n18162 ^ n3289 ^ 1'b0 ;
  assign n18164 = n13431 & n18163 ;
  assign n18165 = n11092 ^ n3350 ^ 1'b0 ;
  assign n18166 = n496 & ~n18165 ;
  assign n18167 = n1217 & ~n14142 ;
  assign n18168 = ~n13485 & n18167 ;
  assign n18169 = ~n10535 & n18168 ;
  assign n18170 = ~n18166 & n18169 ;
  assign n18171 = n10806 ^ n7577 ^ 1'b0 ;
  assign n18172 = ~n345 & n589 ;
  assign n18173 = n529 & n18172 ;
  assign n18174 = n5177 & n18173 ;
  assign n18175 = n7692 & n9847 ;
  assign n18176 = n18175 ^ n4808 ^ 1'b0 ;
  assign n18177 = n9367 ^ n4143 ^ 1'b0 ;
  assign n18178 = n1937 & n7321 ;
  assign n18179 = n18178 ^ n11868 ^ n9799 ;
  assign n18180 = n8985 ^ n7906 ^ n355 ;
  assign n18181 = n7612 & ~n14212 ;
  assign n18182 = n3968 & ~n18075 ;
  assign n18183 = n17264 | n17435 ;
  assign n18184 = n18183 ^ n6377 ^ 1'b0 ;
  assign n18185 = ~n14286 & n18136 ;
  assign n18186 = n6477 ^ n2745 ^ n198 ;
  assign n18187 = n3944 ^ n2632 ^ 1'b0 ;
  assign n18188 = ~n18186 & n18187 ;
  assign n18189 = n4336 ^ n699 ^ 1'b0 ;
  assign n18190 = n18189 ^ n10951 ^ n614 ;
  assign n18191 = n18190 ^ n2384 ^ 1'b0 ;
  assign n18192 = n6403 & n12879 ;
  assign n18193 = n4527 & n18192 ;
  assign n18194 = n3870 | n5088 ;
  assign n18195 = n3313 & n15276 ;
  assign n18196 = n8304 ^ n3408 ^ 1'b0 ;
  assign n18197 = n3567 & ~n9203 ;
  assign n18198 = ~n7643 & n18197 ;
  assign n18199 = ~n1529 & n2449 ;
  assign n18200 = ~n1079 & n9899 ;
  assign n18201 = n18199 & n18200 ;
  assign n18202 = n15788 & ~n18201 ;
  assign n18203 = n9481 & n18202 ;
  assign n18204 = n12471 ^ n4989 ^ 1'b0 ;
  assign n18205 = n6810 & n18204 ;
  assign n18206 = n652 & n14190 ;
  assign n18207 = n17845 ^ n10909 ^ 1'b0 ;
  assign n18210 = ~n3083 & n7676 ;
  assign n18208 = n3468 & n4581 ;
  assign n18209 = n4710 | n18208 ;
  assign n18211 = n18210 ^ n18209 ^ 1'b0 ;
  assign n18212 = n3182 ^ n1661 ^ n324 ;
  assign n18213 = n14565 | n17915 ;
  assign n18214 = n18213 ^ n14895 ^ 1'b0 ;
  assign n18215 = n1070 & n18214 ;
  assign n18216 = ~n2213 & n18215 ;
  assign n18217 = n1805 & n9186 ;
  assign n18218 = n666 | n5941 ;
  assign n18219 = n18218 ^ n10782 ^ 1'b0 ;
  assign n18220 = n1256 & n2754 ;
  assign n18221 = n16885 ^ n14293 ^ 1'b0 ;
  assign n18222 = x47 & ~n8895 ;
  assign n18223 = n1535 & ~n18222 ;
  assign n18224 = n18221 & n18223 ;
  assign n18225 = n6896 ^ n3370 ^ 1'b0 ;
  assign n18226 = n2198 ^ n656 ^ 1'b0 ;
  assign n18227 = ~n18093 & n18226 ;
  assign n18228 = n5145 ^ n3262 ^ 1'b0 ;
  assign n18229 = ~n5434 & n18228 ;
  assign n18230 = n7731 | n16990 ;
  assign n18231 = n11468 | n18230 ;
  assign n18232 = n18231 ^ n11255 ^ n832 ;
  assign n18233 = ~n1114 & n7801 ;
  assign n18234 = n18233 ^ n630 ^ 1'b0 ;
  assign n18235 = n7794 | n7968 ;
  assign n18236 = n18235 ^ n1642 ^ 1'b0 ;
  assign n18237 = n3991 & n18236 ;
  assign n18238 = ~n8454 & n18237 ;
  assign n18239 = ~n10487 & n12313 ;
  assign n18240 = n4318 | n14001 ;
  assign n18241 = n18240 ^ n13298 ^ 1'b0 ;
  assign n18242 = ~n6052 & n18241 ;
  assign n18243 = ~n6531 & n18242 ;
  assign n18244 = n18243 ^ n15049 ^ 1'b0 ;
  assign n18245 = n1828 | n13281 ;
  assign n18246 = n2776 & n13246 ;
  assign n18247 = ~n18245 & n18246 ;
  assign n18248 = n10157 ^ n4432 ^ n521 ;
  assign n18250 = n4335 & ~n5111 ;
  assign n18251 = n18250 ^ n17745 ^ 1'b0 ;
  assign n18249 = n12410 ^ n10379 ^ 1'b0 ;
  assign n18252 = n18251 ^ n18249 ^ n6188 ;
  assign n18253 = n9433 | n13092 ;
  assign n18254 = n18253 ^ n3630 ^ 1'b0 ;
  assign n18255 = ~n12235 & n18254 ;
  assign n18256 = n14201 ^ n7984 ^ 1'b0 ;
  assign n18257 = n18256 ^ n2750 ^ 1'b0 ;
  assign n18258 = n2435 & n18257 ;
  assign n18259 = ( n3714 & n3952 ) | ( n3714 & n14187 ) | ( n3952 & n14187 ) ;
  assign n18260 = n5381 ^ n1534 ^ 1'b0 ;
  assign n18261 = ( n1796 & n12014 ) | ( n1796 & ~n18260 ) | ( n12014 & ~n18260 ) ;
  assign n18262 = n17353 ^ n8168 ^ 1'b0 ;
  assign n18263 = n6024 & ~n7798 ;
  assign n18264 = n18263 ^ n5156 ^ 1'b0 ;
  assign n18265 = ~n4571 & n7589 ;
  assign n18266 = n4045 & n8435 ;
  assign n18267 = n4567 ^ n3122 ^ 1'b0 ;
  assign n18268 = n6352 | n18267 ;
  assign n18269 = n2228 & ~n3362 ;
  assign n18270 = n18269 ^ x15 ^ 1'b0 ;
  assign n18271 = n5170 & n6940 ;
  assign n18272 = n4773 & ~n18271 ;
  assign n18273 = ~n1939 & n2105 ;
  assign n18274 = n12402 & ~n13699 ;
  assign n18275 = n11555 ^ n3356 ^ 1'b0 ;
  assign n18276 = n6713 | n8278 ;
  assign n18277 = n10304 & ~n18276 ;
  assign n18278 = n7016 ^ n4987 ^ 1'b0 ;
  assign n18279 = n18277 | n18278 ;
  assign n18280 = n18279 ^ n13674 ^ 1'b0 ;
  assign n18281 = n17457 ^ x2 ^ 1'b0 ;
  assign n18282 = n17517 ^ n7216 ^ 1'b0 ;
  assign n18283 = ~n9474 & n18282 ;
  assign n18284 = n18283 ^ n3937 ^ 1'b0 ;
  assign n18285 = ~n14286 & n18284 ;
  assign n18286 = ~n3029 & n10577 ;
  assign n18287 = n18286 ^ n13710 ^ 1'b0 ;
  assign n18288 = ~n2840 & n18287 ;
  assign n18289 = ~n11088 & n18288 ;
  assign n18290 = ( n7645 & ~n15731 ) | ( n7645 & n18289 ) | ( ~n15731 & n18289 ) ;
  assign n18291 = ~n4251 & n10616 ;
  assign n18292 = x62 & ~n16428 ;
  assign n18293 = n7559 | n14889 ;
  assign n18294 = n9650 ^ n9189 ^ 1'b0 ;
  assign n18295 = n2670 ^ n690 ^ 1'b0 ;
  assign n18296 = n3438 & n3722 ;
  assign n18297 = n18295 & n18296 ;
  assign n18298 = n15063 | n18297 ;
  assign n18299 = n6942 & ~n18298 ;
  assign n18300 = n16463 ^ n2111 ^ 1'b0 ;
  assign n18301 = ~n8850 & n18300 ;
  assign n18302 = n5552 | n16693 ;
  assign n18303 = n18302 ^ n5854 ^ 1'b0 ;
  assign n18304 = n998 | n9884 ;
  assign n18305 = n12887 & ~n18304 ;
  assign n18306 = n18305 ^ n8558 ^ n1575 ;
  assign n18307 = n18306 ^ n10858 ^ 1'b0 ;
  assign n18308 = n11455 ^ n5093 ^ 1'b0 ;
  assign n18309 = n8257 & n18308 ;
  assign n18310 = n5948 ^ n5135 ^ 1'b0 ;
  assign n18311 = ~n15433 & n18310 ;
  assign n18312 = n18311 ^ n3295 ^ 1'b0 ;
  assign n18313 = n5671 | n12031 ;
  assign n18314 = x48 | n18313 ;
  assign n18315 = n8890 & n18314 ;
  assign n18316 = ~n18312 & n18315 ;
  assign n18317 = n11255 ^ n8747 ^ 1'b0 ;
  assign n18318 = n3521 & ~n18317 ;
  assign n18319 = ~n10669 & n18318 ;
  assign n18320 = n9476 ^ n3116 ^ 1'b0 ;
  assign n18321 = ~n2357 & n18320 ;
  assign n18322 = n11244 ^ n4793 ^ 1'b0 ;
  assign n18323 = n18321 & ~n18322 ;
  assign n18324 = n4903 ^ n4068 ^ n1534 ;
  assign n18325 = n18324 ^ n2989 ^ 1'b0 ;
  assign n18326 = n18323 & n18325 ;
  assign n18327 = n6829 ^ n3182 ^ 1'b0 ;
  assign n18328 = n3565 & ~n18327 ;
  assign n18329 = n5934 ^ n2988 ^ 1'b0 ;
  assign n18330 = n3056 | n18329 ;
  assign n18331 = ( n13658 & n14250 ) | ( n13658 & n18330 ) | ( n14250 & n18330 ) ;
  assign n18332 = n10069 ^ n5949 ^ 1'b0 ;
  assign n18333 = n10897 & n18332 ;
  assign n18334 = n18333 ^ n5178 ^ n2748 ;
  assign n18336 = n3976 & ~n15457 ;
  assign n18337 = n5336 & n18336 ;
  assign n18335 = n16676 & ~n17566 ;
  assign n18338 = n18337 ^ n18335 ^ 1'b0 ;
  assign n18339 = n334 & n377 ;
  assign n18340 = ~n2198 & n18339 ;
  assign n18341 = n1204 & ~n4934 ;
  assign n18342 = n17941 ^ n13202 ^ n2810 ;
  assign n18348 = n3148 ^ n2388 ^ 1'b0 ;
  assign n18349 = n7014 & ~n18348 ;
  assign n18350 = ~n7045 & n18349 ;
  assign n18351 = n7213 & n18350 ;
  assign n18343 = ( n3734 & ~n3935 ) | ( n3734 & n5549 ) | ( ~n3935 & n5549 ) ;
  assign n18344 = ~n1937 & n18343 ;
  assign n18345 = n18344 ^ n15400 ^ 1'b0 ;
  assign n18346 = n10541 & ~n18345 ;
  assign n18347 = ~n17138 & n18346 ;
  assign n18352 = n18351 ^ n18347 ^ 1'b0 ;
  assign n18353 = n7588 & n18352 ;
  assign n18354 = ~n1073 & n1873 ;
  assign n18355 = n14223 ^ n7377 ^ n4290 ;
  assign n18356 = ~n1797 & n3190 ;
  assign n18357 = n6311 ^ n5948 ^ 1'b0 ;
  assign n18358 = n6989 & ~n7719 ;
  assign n18359 = n18358 ^ n11849 ^ 1'b0 ;
  assign n18360 = n14527 ^ n1079 ^ 1'b0 ;
  assign n18361 = ~n5451 & n18360 ;
  assign n18362 = n11316 ^ n6050 ^ 1'b0 ;
  assign n18363 = ( n14615 & ~n14966 ) | ( n14615 & n17934 ) | ( ~n14966 & n17934 ) ;
  assign n18364 = n3517 | n11284 ;
  assign n18365 = n14540 ^ n7037 ^ 1'b0 ;
  assign n18366 = ~n3956 & n5167 ;
  assign n18367 = n1743 | n1933 ;
  assign n18368 = ~n18366 & n18367 ;
  assign n18369 = n1835 ^ n653 ^ 1'b0 ;
  assign n18370 = n7019 ^ n1790 ^ 1'b0 ;
  assign n18371 = n5220 & n18370 ;
  assign n18374 = n4558 ^ n4320 ^ 1'b0 ;
  assign n18372 = n8341 ^ n3316 ^ 1'b0 ;
  assign n18373 = n15034 | n18372 ;
  assign n18375 = n18374 ^ n18373 ^ 1'b0 ;
  assign n18376 = n4659 | n5148 ;
  assign n18377 = n18376 ^ n3924 ^ 1'b0 ;
  assign n18378 = n15557 & ~n18377 ;
  assign n18379 = ~n8158 & n18378 ;
  assign n18380 = n18379 ^ n11178 ^ 1'b0 ;
  assign n18381 = n666 | n5049 ;
  assign n18382 = n13757 & ~n18381 ;
  assign n18383 = ~n1572 & n18382 ;
  assign n18384 = n4046 & ~n18383 ;
  assign n18385 = n10794 & n18384 ;
  assign n18387 = n4929 ^ n258 ^ 1'b0 ;
  assign n18388 = ~n7261 & n18387 ;
  assign n18386 = n6696 ^ n4987 ^ 1'b0 ;
  assign n18389 = n18388 ^ n18386 ^ 1'b0 ;
  assign n18390 = n3037 & ~n18389 ;
  assign n18391 = n5492 ^ n1361 ^ 1'b0 ;
  assign n18392 = n708 | n18391 ;
  assign n18393 = n18392 ^ n3850 ^ 1'b0 ;
  assign n18394 = n18251 ^ n2414 ^ 1'b0 ;
  assign n18395 = n5711 & n7288 ;
  assign n18396 = n5398 ^ n3746 ^ 1'b0 ;
  assign n18397 = ~n1089 & n18396 ;
  assign n18398 = ~x6 & n1092 ;
  assign n18399 = n18398 ^ n10808 ^ 1'b0 ;
  assign n18400 = ~n18397 & n18399 ;
  assign n18401 = n18395 | n18400 ;
  assign n18402 = n2491 ^ n844 ^ 1'b0 ;
  assign n18403 = n18402 ^ n3622 ^ 1'b0 ;
  assign n18404 = n18403 ^ n7118 ^ 1'b0 ;
  assign n18405 = n3532 & n13483 ;
  assign n18406 = ~n2487 & n7137 ;
  assign n18407 = n18406 ^ n9025 ^ 1'b0 ;
  assign n18408 = n250 | n7380 ;
  assign n18409 = n3809 | n18408 ;
  assign n18410 = ~n5408 & n18409 ;
  assign n18411 = n9587 & n10053 ;
  assign n18412 = n14635 ^ n2328 ^ 1'b0 ;
  assign n18413 = ( n3210 & n4175 ) | ( n3210 & n5044 ) | ( n4175 & n5044 ) ;
  assign n18414 = x110 & ~n18413 ;
  assign n18415 = n11417 | n18414 ;
  assign n18416 = ~n4001 & n8315 ;
  assign n18417 = n18416 ^ n7261 ^ 1'b0 ;
  assign n18418 = n652 & n13032 ;
  assign n18419 = ~n3787 & n18418 ;
  assign n18420 = n2723 | n8940 ;
  assign n18421 = n18419 & ~n18420 ;
  assign n18422 = n6992 ^ n5129 ^ 1'b0 ;
  assign n18423 = x70 | n18422 ;
  assign n18424 = n10843 ^ n6066 ^ 1'b0 ;
  assign n18425 = ~n3678 & n13937 ;
  assign n18426 = n18424 | n18425 ;
  assign n18427 = n18426 ^ n8236 ^ 1'b0 ;
  assign n18428 = n4467 ^ n1884 ^ 1'b0 ;
  assign n18429 = ( n4250 & ~n4879 ) | ( n4250 & n18428 ) | ( ~n4879 & n18428 ) ;
  assign n18430 = n18429 ^ n3924 ^ 1'b0 ;
  assign n18431 = n5075 & ~n5578 ;
  assign n18432 = n2602 & n18431 ;
  assign n18433 = n18432 ^ n12696 ^ n7695 ;
  assign n18434 = n5246 & ~n8237 ;
  assign n18435 = ~n3073 & n18434 ;
  assign n18436 = ( ~n10775 & n18433 ) | ( ~n10775 & n18435 ) | ( n18433 & n18435 ) ;
  assign n18437 = n3338 | n18404 ;
  assign n18438 = n18437 ^ n7116 ^ 1'b0 ;
  assign n18439 = n12727 ^ n593 ^ 1'b0 ;
  assign n18440 = n8863 ^ n672 ^ 1'b0 ;
  assign n18441 = n9389 ^ n369 ^ 1'b0 ;
  assign n18442 = ~n4759 & n18441 ;
  assign n18443 = n4380 | n16879 ;
  assign n18444 = ~n4081 & n10546 ;
  assign n18445 = n9843 | n16050 ;
  assign n18446 = n15002 ^ n10528 ^ 1'b0 ;
  assign n18447 = ( n9724 & ~n18445 ) | ( n9724 & n18446 ) | ( ~n18445 & n18446 ) ;
  assign n18448 = n13786 ^ n8747 ^ 1'b0 ;
  assign n18449 = n17497 ^ n15486 ^ 1'b0 ;
  assign n18450 = ~n15704 & n18449 ;
  assign n18451 = n5949 ^ n1295 ^ 1'b0 ;
  assign n18452 = n9438 & n18451 ;
  assign n18453 = n16364 & n18452 ;
  assign n18454 = ~n18450 & n18453 ;
  assign n18455 = n9058 ^ n5108 ^ 1'b0 ;
  assign n18456 = n9753 ^ n7636 ^ 1'b0 ;
  assign n18457 = n4549 & ~n18456 ;
  assign n18458 = ( n3749 & n7155 ) | ( n3749 & n18457 ) | ( n7155 & n18457 ) ;
  assign n18459 = n14800 & ~n15147 ;
  assign n18460 = ~n18458 & n18459 ;
  assign n18461 = n3167 | n6693 ;
  assign n18462 = n18461 ^ n4095 ^ 1'b0 ;
  assign n18463 = ~n920 & n4576 ;
  assign n18464 = n18463 ^ n5228 ^ 1'b0 ;
  assign n18466 = n1244 & ~n7518 ;
  assign n18467 = n18466 ^ n6990 ^ 1'b0 ;
  assign n18468 = ( n7865 & n11782 ) | ( n7865 & n18467 ) | ( n11782 & n18467 ) ;
  assign n18465 = n1164 | n5495 ;
  assign n18469 = n18468 ^ n18465 ^ 1'b0 ;
  assign n18470 = n1128 & n9482 ;
  assign n18471 = ( n5495 & n10170 ) | ( n5495 & n11308 ) | ( n10170 & n11308 ) ;
  assign n18472 = n6933 & ~n18471 ;
  assign n18473 = n2911 & n18472 ;
  assign n18474 = n7360 ^ n6356 ^ n2861 ;
  assign n18476 = ~n1937 & n16445 ;
  assign n18475 = n5443 | n11995 ;
  assign n18477 = n18476 ^ n18475 ^ 1'b0 ;
  assign n18478 = ~n1865 & n6343 ;
  assign n18479 = n18478 ^ n2951 ^ 1'b0 ;
  assign n18480 = n10026 ^ n7863 ^ 1'b0 ;
  assign n18481 = ~n4666 & n18480 ;
  assign n18482 = n9928 & n14785 ;
  assign n18483 = n18482 ^ n412 ^ 1'b0 ;
  assign n18484 = ~n12345 & n18483 ;
  assign n18485 = n4362 & n8425 ;
  assign n18486 = n18485 ^ x94 ^ 1'b0 ;
  assign n18487 = n18486 ^ n12124 ^ n6103 ;
  assign n18488 = ~n1224 & n7760 ;
  assign n18489 = ~n198 & n18488 ;
  assign n18490 = n8493 ^ n5727 ^ 1'b0 ;
  assign n18491 = ~n18489 & n18490 ;
  assign n18492 = n12293 | n17096 ;
  assign n18493 = n460 | n18492 ;
  assign n18494 = n1512 ^ n313 ^ 1'b0 ;
  assign n18495 = n1714 & ~n2558 ;
  assign n18496 = n18495 ^ n7689 ^ 1'b0 ;
  assign n18497 = x92 & n18496 ;
  assign n18498 = n18497 ^ n7991 ^ 1'b0 ;
  assign n18499 = ~n14892 & n18498 ;
  assign n18500 = x105 & n2551 ;
  assign n18501 = n18500 ^ n15782 ^ 1'b0 ;
  assign n18502 = n5251 & n15588 ;
  assign n18503 = n2634 & n18502 ;
  assign n18504 = ( n3744 & n11333 ) | ( n3744 & n18503 ) | ( n11333 & n18503 ) ;
  assign n18505 = n3671 ^ n1705 ^ x47 ;
  assign n18506 = ~n2756 & n4505 ;
  assign n18507 = ~n3205 & n18506 ;
  assign n18508 = n18507 ^ n14469 ^ n4064 ;
  assign n18509 = n9869 & ~n18508 ;
  assign n18510 = n18509 ^ n653 ^ 1'b0 ;
  assign n18511 = n12400 ^ n769 ^ 1'b0 ;
  assign n18512 = n3190 & ~n18511 ;
  assign n18513 = n18512 ^ n13961 ^ 1'b0 ;
  assign n18514 = n7549 ^ n5533 ^ 1'b0 ;
  assign n18515 = n4609 | n18514 ;
  assign n18516 = n2261 & n7110 ;
  assign n18517 = n18516 ^ n4020 ^ 1'b0 ;
  assign n18518 = n18517 ^ n5144 ^ 1'b0 ;
  assign n18519 = ~n3472 & n18518 ;
  assign n18520 = n13124 | n18519 ;
  assign n18521 = n18520 ^ n17224 ^ 1'b0 ;
  assign n18523 = n2109 | n2123 ;
  assign n18524 = n2123 & ~n18523 ;
  assign n18525 = n18524 ^ n805 ^ 1'b0 ;
  assign n18526 = n217 & n4149 ;
  assign n18527 = ~n4149 & n18526 ;
  assign n18528 = n18527 ^ n2246 ^ 1'b0 ;
  assign n18529 = x84 & ~n10745 ;
  assign n18530 = ~x84 & n18529 ;
  assign n18531 = ( n18525 & ~n18528 ) | ( n18525 & n18530 ) | ( ~n18528 & n18530 ) ;
  assign n18522 = n3604 & ~n6366 ;
  assign n18532 = n18531 ^ n18522 ^ 1'b0 ;
  assign n18534 = n6916 ^ n521 ^ 1'b0 ;
  assign n18535 = n5202 & n18534 ;
  assign n18536 = ~n2128 & n18535 ;
  assign n18533 = n362 & n2662 ;
  assign n18537 = n18536 ^ n18533 ^ 1'b0 ;
  assign n18538 = n9269 | n18537 ;
  assign n18539 = n18532 | n18538 ;
  assign n18540 = n836 & n18539 ;
  assign n18541 = n18078 ^ n12378 ^ 1'b0 ;
  assign n18542 = n4633 ^ n3579 ^ 1'b0 ;
  assign n18543 = n11845 & n18542 ;
  assign n18544 = n18543 ^ n7629 ^ 1'b0 ;
  assign n18545 = n2909 ^ n755 ^ 1'b0 ;
  assign n18548 = ~n4324 & n6504 ;
  assign n18549 = n18548 ^ n8440 ^ 1'b0 ;
  assign n18546 = ~n655 & n1058 ;
  assign n18547 = n14777 & ~n18546 ;
  assign n18550 = n18549 ^ n18547 ^ n3429 ;
  assign n18551 = n2746 & ~n18550 ;
  assign n18552 = n18551 ^ n2633 ^ 1'b0 ;
  assign n18553 = n3381 ^ n1710 ^ 1'b0 ;
  assign n18554 = n18553 ^ n16050 ^ n7279 ;
  assign n18555 = n7170 | n18554 ;
  assign n18556 = ~n3958 & n9554 ;
  assign n18557 = n7353 ^ n4602 ^ 1'b0 ;
  assign n18558 = ~n3391 & n18557 ;
  assign n18559 = ( ~n15045 & n18358 ) | ( ~n15045 & n18558 ) | ( n18358 & n18558 ) ;
  assign n18560 = n6133 ^ n218 ^ 1'b0 ;
  assign n18561 = n7486 | n14505 ;
  assign n18562 = n3017 & n12748 ;
  assign n18563 = ~n5011 & n8464 ;
  assign n18564 = n3160 | n8998 ;
  assign n18565 = n4635 & ~n4777 ;
  assign n18566 = n1469 & n18565 ;
  assign n18567 = n6919 & ~n11522 ;
  assign n18568 = ( n453 & ~n2928 ) | ( n453 & n7026 ) | ( ~n2928 & n7026 ) ;
  assign n18569 = n14147 & n18568 ;
  assign n18570 = ~n1512 & n17493 ;
  assign n18572 = n10357 ^ n7177 ^ n7157 ;
  assign n18571 = n4925 ^ n3474 ^ n1520 ;
  assign n18573 = n18572 ^ n18571 ^ n1475 ;
  assign n18575 = n6172 & ~n8114 ;
  assign n18576 = n18575 ^ n9503 ^ 1'b0 ;
  assign n18574 = n6403 & ~n13195 ;
  assign n18577 = n18576 ^ n18574 ^ 1'b0 ;
  assign n18578 = n13119 ^ n5381 ^ 1'b0 ;
  assign n18579 = n18578 ^ n12000 ^ 1'b0 ;
  assign n18580 = n6815 & n18579 ;
  assign n18581 = n18580 ^ n4710 ^ 1'b0 ;
  assign n18582 = n1661 | n4292 ;
  assign n18583 = n18582 ^ n875 ^ 1'b0 ;
  assign n18584 = n11234 ^ n3433 ^ 1'b0 ;
  assign n18585 = n18584 ^ n15717 ^ 1'b0 ;
  assign n18586 = ~n11369 & n11775 ;
  assign n18587 = n3921 | n8656 ;
  assign n18588 = n18587 ^ n9055 ^ 1'b0 ;
  assign n18589 = n14543 ^ n4728 ^ 1'b0 ;
  assign n18590 = n3138 | n6791 ;
  assign n18591 = n18590 ^ n840 ^ 1'b0 ;
  assign n18592 = n3338 ^ n1772 ^ 1'b0 ;
  assign n18593 = n6293 ^ n4626 ^ 1'b0 ;
  assign n18594 = n2297 ^ n852 ^ 1'b0 ;
  assign n18595 = ~n5890 & n18594 ;
  assign n18596 = n12023 ^ n1070 ^ 1'b0 ;
  assign n18597 = ~n18595 & n18596 ;
  assign n18598 = n8052 ^ n726 ^ 1'b0 ;
  assign n18599 = n11793 ^ n1303 ^ 1'b0 ;
  assign n18600 = ~n18598 & n18599 ;
  assign n18601 = n4973 & ~n12374 ;
  assign n18602 = n18601 ^ n3677 ^ 1'b0 ;
  assign n18603 = n15760 ^ n2489 ^ 1'b0 ;
  assign n18604 = ~n3442 & n13529 ;
  assign n18605 = n18604 ^ n11055 ^ 1'b0 ;
  assign n18606 = n3515 & ~n14713 ;
  assign n18607 = ~n8836 & n18606 ;
  assign n18608 = ~n18605 & n18607 ;
  assign n18609 = n5430 ^ n2908 ^ 1'b0 ;
  assign n18610 = n987 | n17066 ;
  assign n18611 = ( n3785 & ~n9380 ) | ( n3785 & n12460 ) | ( ~n9380 & n12460 ) ;
  assign n18612 = n799 ^ n224 ^ 1'b0 ;
  assign n18613 = n18612 ^ n12587 ^ n2704 ;
  assign n18614 = n12879 ^ n12696 ^ 1'b0 ;
  assign n18615 = n163 | n690 ;
  assign n18616 = n15603 ^ n13271 ^ 1'b0 ;
  assign n18617 = ~n4344 & n11701 ;
  assign n18618 = n1392 ^ n1015 ^ 1'b0 ;
  assign n18619 = x62 & n18618 ;
  assign n18620 = n18619 ^ n4777 ^ 1'b0 ;
  assign n18621 = n17015 ^ n6158 ^ 1'b0 ;
  assign n18622 = n12009 | n18621 ;
  assign n18623 = n16515 & n16691 ;
  assign n18624 = n3273 | n12218 ;
  assign n18625 = n18623 | n18624 ;
  assign n18626 = ~n533 & n14951 ;
  assign n18627 = n18626 ^ n11905 ^ n4318 ;
  assign n18628 = n7187 | n8236 ;
  assign n18629 = n14298 & ~n18628 ;
  assign n18630 = n13469 ^ n5969 ^ 1'b0 ;
  assign n18631 = n2243 | n18630 ;
  assign n18632 = n209 & n6430 ;
  assign n18633 = n5074 ^ n3869 ^ 1'b0 ;
  assign n18634 = n3376 | n18633 ;
  assign n18635 = ~n856 & n18634 ;
  assign n18636 = n18632 & n18635 ;
  assign n18637 = n3485 ^ n560 ^ 1'b0 ;
  assign n18638 = n7191 & ~n18637 ;
  assign n18639 = n13960 | n18638 ;
  assign n18640 = n883 & ~n9725 ;
  assign n18641 = n17475 & n18640 ;
  assign n18642 = n4408 | n18641 ;
  assign n18643 = n14100 & ~n18642 ;
  assign n18644 = n6174 | n12408 ;
  assign n18645 = n18643 & ~n18644 ;
  assign n18646 = n3778 & ~n18645 ;
  assign n18647 = n3899 & ~n11307 ;
  assign n18648 = ~n6187 & n18647 ;
  assign n18649 = n898 & n6714 ;
  assign n18650 = ( n9805 & ~n13271 ) | ( n9805 & n18649 ) | ( ~n13271 & n18649 ) ;
  assign n18651 = n6707 | n9852 ;
  assign n18652 = n10606 | n11611 ;
  assign n18653 = n4216 & ~n12707 ;
  assign n18654 = ~x73 & n18653 ;
  assign n18655 = n18654 ^ n1773 ^ 1'b0 ;
  assign n18656 = n11730 ^ n3629 ^ 1'b0 ;
  assign n18657 = ~n2676 & n9032 ;
  assign n18658 = n14433 ^ n3086 ^ 1'b0 ;
  assign n18659 = ~n9045 & n18658 ;
  assign n18660 = n8918 | n11818 ;
  assign n18661 = n9176 & ~n18660 ;
  assign n18662 = n1015 | n6779 ;
  assign n18663 = n18662 ^ n4767 ^ 1'b0 ;
  assign n18664 = n11051 & n18663 ;
  assign n18665 = n3417 & n11567 ;
  assign n18666 = n18664 & n18665 ;
  assign n18667 = x110 & ~n3120 ;
  assign n18668 = n18667 ^ n902 ^ 1'b0 ;
  assign n18669 = n1184 | n1420 ;
  assign n18670 = n14808 & ~n18669 ;
  assign n18671 = n14985 | n18670 ;
  assign n18672 = n5971 & n18671 ;
  assign n18673 = n14280 & n18672 ;
  assign n18674 = n4543 & ~n4899 ;
  assign n18675 = n7126 & n18674 ;
  assign n18676 = n12475 & n18675 ;
  assign n18677 = x30 | n7794 ;
  assign n18678 = n9147 ^ n7382 ^ 1'b0 ;
  assign n18679 = ~n8891 & n18678 ;
  assign n18680 = n1774 & n2463 ;
  assign n18681 = n8437 ^ n1937 ^ 1'b0 ;
  assign n18682 = n18671 & ~n18681 ;
  assign n18683 = ( n1145 & n8106 ) | ( n1145 & n14808 ) | ( n8106 & n14808 ) ;
  assign n18684 = n9132 ^ n8820 ^ 1'b0 ;
  assign n18685 = n5413 & ~n18684 ;
  assign n18688 = ~n6439 & n7987 ;
  assign n18689 = n18688 ^ n4876 ^ 1'b0 ;
  assign n18686 = n184 | n521 ;
  assign n18687 = n18686 ^ n7256 ^ 1'b0 ;
  assign n18690 = n18689 ^ n18687 ^ 1'b0 ;
  assign n18691 = n2131 & n9942 ;
  assign n18693 = n973 & ~n3887 ;
  assign n18692 = n12640 ^ n8916 ^ 1'b0 ;
  assign n18694 = n18693 ^ n18692 ^ 1'b0 ;
  assign n18695 = ~n18691 & n18694 ;
  assign n18696 = n6242 ^ n5321 ^ 1'b0 ;
  assign n18697 = n18696 ^ n15613 ^ n10527 ;
  assign n18698 = n8368 ^ n1195 ^ 1'b0 ;
  assign n18699 = n13054 & ~n18698 ;
  assign n18700 = n7382 & ~n10699 ;
  assign n18701 = ~n1225 & n3065 ;
  assign n18702 = n18701 ^ n16631 ^ 1'b0 ;
  assign n18703 = ( n1208 & n12135 ) | ( n1208 & n17915 ) | ( n12135 & n17915 ) ;
  assign n18704 = n14254 ^ n10603 ^ 1'b0 ;
  assign n18705 = ~n4018 & n6201 ;
  assign n18706 = n18705 ^ n8403 ^ 1'b0 ;
  assign n18707 = n18292 ^ n12994 ^ 1'b0 ;
  assign n18708 = ~n5499 & n9066 ;
  assign n18709 = ~n10947 & n18201 ;
  assign n18710 = n3153 & ~n15623 ;
  assign n18711 = n18710 ^ n836 ^ 1'b0 ;
  assign n18712 = ~n3357 & n10903 ;
  assign n18713 = n18712 ^ n1426 ^ 1'b0 ;
  assign n18714 = n8383 ^ n5152 ^ 1'b0 ;
  assign n18715 = n11259 & n18714 ;
  assign n18716 = n9935 & n10885 ;
  assign n18717 = n13593 ^ n2397 ^ 1'b0 ;
  assign n18718 = n18717 ^ n15642 ^ 1'b0 ;
  assign n18719 = n13094 ^ n11380 ^ n2832 ;
  assign n18720 = ( n863 & n4983 ) | ( n863 & ~n18719 ) | ( n4983 & ~n18719 ) ;
  assign n18721 = n9377 ^ n8990 ^ 1'b0 ;
  assign n18722 = n9668 | n18721 ;
  assign n18723 = n2456 | n18722 ;
  assign n18724 = n18723 ^ n1184 ^ 1'b0 ;
  assign n18725 = n9256 & n11013 ;
  assign n18726 = ~n7210 & n15727 ;
  assign n18731 = n3790 & ~n6681 ;
  assign n18732 = n11011 ^ n6966 ^ 1'b0 ;
  assign n18733 = n18731 & ~n18732 ;
  assign n18727 = n12336 & ~n16990 ;
  assign n18728 = ~n3792 & n9879 ;
  assign n18729 = n18727 & n18728 ;
  assign n18730 = n8888 & ~n18729 ;
  assign n18734 = n18733 ^ n18730 ^ 1'b0 ;
  assign n18735 = n18734 ^ n6308 ^ n3237 ;
  assign n18736 = n521 | n11649 ;
  assign n18737 = n18736 ^ n8925 ^ 1'b0 ;
  assign n18738 = n7219 | n18737 ;
  assign n18739 = ~n2380 & n11910 ;
  assign n18740 = n12778 | n18546 ;
  assign n18741 = n15369 | n18740 ;
  assign n18742 = n10818 ^ n9671 ^ 1'b0 ;
  assign n18743 = x23 & n18742 ;
  assign n18744 = n7716 | n10950 ;
  assign n18745 = n1897 | n18744 ;
  assign n18746 = ( ~n788 & n875 ) | ( ~n788 & n18388 ) | ( n875 & n18388 ) ;
  assign n18747 = n3606 ^ n756 ^ 1'b0 ;
  assign n18748 = n2663 | n18747 ;
  assign n18749 = n18748 ^ n9005 ^ n1689 ;
  assign n18750 = ( ~n4384 & n6756 ) | ( ~n4384 & n18749 ) | ( n6756 & n18749 ) ;
  assign n18751 = n900 & ~n9411 ;
  assign n18752 = ~n17989 & n18751 ;
  assign n18753 = n2558 & ~n8232 ;
  assign n18754 = n1680 & ~n18753 ;
  assign n18755 = n3403 | n12917 ;
  assign n18756 = n18755 ^ n13285 ^ 1'b0 ;
  assign n18757 = n12101 & n18756 ;
  assign n18758 = n10271 ^ n6569 ^ 1'b0 ;
  assign n18759 = n13824 ^ n3961 ^ 1'b0 ;
  assign n18760 = ~n9568 & n13663 ;
  assign n18761 = n18759 & n18760 ;
  assign n18762 = ~n1774 & n11875 ;
  assign n18763 = n10457 & ~n18762 ;
  assign n18764 = n2622 & ~n5357 ;
  assign n18765 = n18764 ^ n4024 ^ 1'b0 ;
  assign n18766 = n18279 | n18765 ;
  assign n18767 = n1017 | n8006 ;
  assign n18768 = n5530 & ~n12591 ;
  assign n18769 = n18767 & n18768 ;
  assign n18770 = n12715 & n18769 ;
  assign n18771 = n8601 & ~n11921 ;
  assign n18772 = n5443 & n18771 ;
  assign n18773 = n18772 ^ n5671 ^ 1'b0 ;
  assign n18774 = n7971 ^ n4767 ^ 1'b0 ;
  assign n18775 = ~n3111 & n11996 ;
  assign n18776 = n17421 ^ n1189 ^ 1'b0 ;
  assign n18777 = n12387 ^ n169 ^ 1'b0 ;
  assign n18778 = n18021 | n18777 ;
  assign n18779 = ~n569 & n14574 ;
  assign n18780 = n3322 & n18779 ;
  assign n18781 = n7787 ^ n1683 ^ 1'b0 ;
  assign n18782 = n18780 | n18781 ;
  assign n18783 = n8187 | n18782 ;
  assign n18784 = n8925 ^ n1268 ^ 1'b0 ;
  assign n18785 = n13301 & ~n18784 ;
  assign n18786 = n7652 ^ n2901 ^ 1'b0 ;
  assign n18787 = ~n6293 & n18786 ;
  assign n18788 = n1526 & n4678 ;
  assign n18789 = n3226 | n18788 ;
  assign n18790 = n6107 ^ n861 ^ 1'b0 ;
  assign n18791 = n18789 & ~n18790 ;
  assign n18792 = n7483 ^ n180 ^ 1'b0 ;
  assign n18793 = n15046 ^ n2670 ^ 1'b0 ;
  assign n18794 = n8122 & ~n9184 ;
  assign n18795 = ( n6885 & n8006 ) | ( n6885 & ~n8962 ) | ( n8006 & ~n8962 ) ;
  assign n18796 = n5238 & n14685 ;
  assign n18797 = n18795 & n18796 ;
  assign n18798 = ~n9808 & n14969 ;
  assign n18799 = ~n15148 & n18798 ;
  assign n18800 = n18799 ^ n8958 ^ 1'b0 ;
  assign n18801 = ~n18797 & n18800 ;
  assign n18802 = ~n4793 & n10923 ;
  assign n18803 = n7813 | n12422 ;
  assign n18804 = n4071 ^ n1578 ^ n874 ;
  assign n18805 = ~n758 & n1266 ;
  assign n18806 = n15467 & n18805 ;
  assign n18807 = n16118 ^ n8840 ^ 1'b0 ;
  assign n18808 = ~n5755 & n18807 ;
  assign n18809 = ~n5523 & n8752 ;
  assign n18810 = n17465 & n18809 ;
  assign n18811 = n2826 & ~n8823 ;
  assign n18813 = n6538 ^ n1615 ^ n392 ;
  assign n18812 = n12261 | n13266 ;
  assign n18814 = n18813 ^ n18812 ^ 1'b0 ;
  assign n18817 = ( n637 & n1204 ) | ( n637 & n6090 ) | ( n1204 & n6090 ) ;
  assign n18815 = n3164 & n9167 ;
  assign n18816 = n18815 ^ n1791 ^ 1'b0 ;
  assign n18818 = n18817 ^ n18816 ^ 1'b0 ;
  assign n18819 = n18818 ^ n11855 ^ 1'b0 ;
  assign n18820 = n4956 & ~n18819 ;
  assign n18821 = ~n1725 & n3398 ;
  assign n18822 = n11296 & ~n18821 ;
  assign n18823 = n14908 ^ n6630 ^ 1'b0 ;
  assign n18824 = n17322 ^ n10551 ^ 1'b0 ;
  assign n18825 = n11160 | n12601 ;
  assign n18826 = n18825 ^ x54 ^ 1'b0 ;
  assign n18827 = ~n18824 & n18826 ;
  assign n18828 = n18827 ^ n17792 ^ 1'b0 ;
  assign n18829 = n4323 | n10261 ;
  assign n18830 = n18829 ^ n8805 ^ 1'b0 ;
  assign n18831 = ~n11593 & n18830 ;
  assign n18832 = n18831 ^ n2844 ^ 1'b0 ;
  assign n18833 = n4664 & ~n18832 ;
  assign n18834 = n709 | n13119 ;
  assign n18835 = n9367 | n9942 ;
  assign n18836 = n11963 ^ n3649 ^ 1'b0 ;
  assign n18837 = n7426 & n18836 ;
  assign n18838 = n8623 ^ n468 ^ 1'b0 ;
  assign n18839 = n16663 ^ n5537 ^ 1'b0 ;
  assign n18840 = ~n3653 & n14145 ;
  assign n18841 = n12840 & n13686 ;
  assign n18842 = n5064 & ~n6151 ;
  assign n18843 = n18842 ^ n2931 ^ 1'b0 ;
  assign n18844 = n18843 ^ n639 ^ 1'b0 ;
  assign n18845 = ~n13779 & n18844 ;
  assign n18846 = ~n3511 & n9077 ;
  assign n18847 = ~n13293 & n18846 ;
  assign n18848 = n10399 & ~n18207 ;
  assign n18849 = n5634 ^ n4604 ^ 1'b0 ;
  assign n18850 = n14847 & n18849 ;
  assign n18851 = n3290 | n18850 ;
  assign n18852 = n5104 & n11267 ;
  assign n18853 = ~n2111 & n18852 ;
  assign n18854 = n18853 ^ n4875 ^ 1'b0 ;
  assign n18855 = n3859 ^ n3690 ^ 1'b0 ;
  assign n18856 = n10496 ^ n8348 ^ n2884 ;
  assign n18857 = n18856 ^ n11131 ^ 1'b0 ;
  assign n18858 = n18855 & ~n18857 ;
  assign n18859 = n2168 & n11130 ;
  assign n18860 = ( n9295 & n14625 ) | ( n9295 & n18859 ) | ( n14625 & n18859 ) ;
  assign n18861 = x49 & ~n9890 ;
  assign n18862 = n8092 ^ n5946 ^ n5859 ;
  assign n18863 = n1962 | n7226 ;
  assign n18864 = ( ~n4701 & n8500 ) | ( ~n4701 & n18863 ) | ( n8500 & n18863 ) ;
  assign n18865 = n18864 ^ n6634 ^ 1'b0 ;
  assign n18866 = n4482 & n18865 ;
  assign n18867 = n6763 & ~n17007 ;
  assign n18868 = n692 & n1738 ;
  assign n18869 = ~n2510 & n18868 ;
  assign n18870 = n11778 & ~n18869 ;
  assign n18871 = ~n733 & n18870 ;
  assign n18872 = ~n1383 & n13797 ;
  assign n18873 = n10759 ^ n2945 ^ 1'b0 ;
  assign n18874 = n18872 & ~n18873 ;
  assign n18875 = n8005 ^ n6577 ^ 1'b0 ;
  assign n18876 = n3641 & n18875 ;
  assign n18877 = ( n5402 & ~n16697 ) | ( n5402 & n18876 ) | ( ~n16697 & n18876 ) ;
  assign n18879 = n12706 ^ n12541 ^ 1'b0 ;
  assign n18878 = ~n285 & n16221 ;
  assign n18880 = n18879 ^ n18878 ^ 1'b0 ;
  assign n18881 = n16396 ^ n10104 ^ 1'b0 ;
  assign n18882 = ~n11680 & n18881 ;
  assign n18883 = n12976 & n18882 ;
  assign n18884 = ~n15259 & n18883 ;
  assign n18885 = n2634 | n7967 ;
  assign n18886 = n1300 | n18885 ;
  assign n18887 = n18188 ^ n5647 ^ 1'b0 ;
  assign n18888 = n5390 ^ n1689 ^ 1'b0 ;
  assign n18889 = n1487 & ~n3015 ;
  assign n18890 = n1718 & n18889 ;
  assign n18891 = n18890 ^ x79 ^ 1'b0 ;
  assign n18892 = n7603 & n18891 ;
  assign n18893 = n9958 ^ n2809 ^ 1'b0 ;
  assign n18894 = ~n2159 & n3339 ;
  assign n18895 = n18894 ^ n208 ^ 1'b0 ;
  assign n18896 = n18893 & n18895 ;
  assign n18897 = n9478 | n13659 ;
  assign n18898 = ( n5766 & n7678 ) | ( n5766 & ~n10818 ) | ( n7678 & ~n10818 ) ;
  assign n18899 = n15456 & ~n18898 ;
  assign n18900 = ~n18897 & n18899 ;
  assign n18901 = ~n9990 & n10564 ;
  assign n18902 = ~x63 & n18901 ;
  assign n18903 = n18902 ^ n7267 ^ 1'b0 ;
  assign n18904 = n14333 ^ n7094 ^ 1'b0 ;
  assign n18905 = n556 & n10450 ;
  assign n18906 = n2442 & n18905 ;
  assign n18907 = n1276 | n18906 ;
  assign n18908 = n18907 ^ n12609 ^ 1'b0 ;
  assign n18909 = n7453 | n14923 ;
  assign n18910 = n5457 | n13625 ;
  assign n18911 = n13625 & ~n18910 ;
  assign n18912 = x14 & n518 ;
  assign n18913 = ~n518 & n18912 ;
  assign n18914 = n3792 & ~n18913 ;
  assign n18915 = n18913 & n18914 ;
  assign n18916 = x123 & ~n18915 ;
  assign n18917 = ~x123 & n18916 ;
  assign n18918 = n8429 & ~n18917 ;
  assign n18919 = ~n8429 & n18918 ;
  assign n18920 = ~n2579 & n11538 ;
  assign n18921 = n18919 & n18920 ;
  assign n18922 = n18911 | n18921 ;
  assign n18923 = n18911 & ~n18922 ;
  assign n18924 = n9632 | n15113 ;
  assign n18925 = n18924 ^ n6719 ^ 1'b0 ;
  assign n18926 = ( ~n6284 & n18923 ) | ( ~n6284 & n18925 ) | ( n18923 & n18925 ) ;
  assign n18927 = n6382 ^ n5574 ^ 1'b0 ;
  assign n18928 = ~n9307 & n18927 ;
  assign n18929 = n3323 & ~n18928 ;
  assign n18930 = n4147 & n18929 ;
  assign n18931 = n10075 ^ n7371 ^ 1'b0 ;
  assign n18932 = n7330 & ~n15921 ;
  assign n18933 = n18931 & n18932 ;
  assign n18934 = ~n18931 & n18933 ;
  assign n18935 = n12391 ^ n742 ^ 1'b0 ;
  assign n18936 = n5256 & ~n18935 ;
  assign n18937 = ~n13622 & n18936 ;
  assign n18938 = n11717 ^ n11709 ^ 1'b0 ;
  assign n18939 = n14683 ^ n10402 ^ 1'b0 ;
  assign n18940 = ~n8987 & n18939 ;
  assign n18942 = n8431 ^ n3214 ^ 1'b0 ;
  assign n18941 = ~n756 & n3476 ;
  assign n18943 = n18942 ^ n18941 ^ n7029 ;
  assign n18944 = n16521 & ~n17415 ;
  assign n18945 = ( n5422 & n10931 ) | ( n5422 & ~n11334 ) | ( n10931 & ~n11334 ) ;
  assign n18946 = n262 & ~n1642 ;
  assign n18947 = ~n4769 & n8803 ;
  assign n18948 = ~n7111 & n18947 ;
  assign n18949 = n11607 & n12041 ;
  assign n18950 = n18949 ^ n5931 ^ 1'b0 ;
  assign n18951 = n2743 | n18950 ;
  assign n18952 = n1211 | n4252 ;
  assign n18953 = n18952 ^ n10718 ^ 1'b0 ;
  assign n18954 = ~n1725 & n18953 ;
  assign n18955 = n14489 ^ n10952 ^ 1'b0 ;
  assign n18956 = n3974 ^ n1457 ^ 1'b0 ;
  assign n18957 = n2998 & ~n6885 ;
  assign n18958 = n18957 ^ n597 ^ 1'b0 ;
  assign n18959 = n4433 & n9586 ;
  assign n18960 = n12899 ^ n5547 ^ n5049 ;
  assign n18961 = ~n2504 & n4461 ;
  assign n18962 = n18961 ^ n9465 ^ 1'b0 ;
  assign n18963 = n6917 & n9931 ;
  assign n18964 = n10417 ^ n8113 ^ n6114 ;
  assign n18967 = n8885 ^ n1606 ^ 1'b0 ;
  assign n18965 = n13120 ^ n9006 ^ 1'b0 ;
  assign n18966 = x17 & ~n18965 ;
  assign n18968 = n18967 ^ n18966 ^ 1'b0 ;
  assign n18969 = n5324 | n17259 ;
  assign n18970 = n18969 ^ n17555 ^ 1'b0 ;
  assign n18971 = n7932 ^ n7581 ^ 1'b0 ;
  assign n18972 = ~n7705 & n18971 ;
  assign n18973 = ~n1590 & n18972 ;
  assign n18974 = n15048 ^ n14561 ^ 1'b0 ;
  assign n18975 = n6362 | n18974 ;
  assign n18976 = n15401 ^ n5378 ^ n876 ;
  assign n18977 = n4898 ^ x79 ^ 1'b0 ;
  assign n18978 = ~n4893 & n18977 ;
  assign n18979 = n11506 | n18630 ;
  assign n18980 = n1088 & ~n9148 ;
  assign n18981 = ( n6605 & n6641 ) | ( n6605 & ~n18402 ) | ( n6641 & ~n18402 ) ;
  assign n18982 = ~n2054 & n6606 ;
  assign n18983 = ~n10905 & n18982 ;
  assign n18984 = n18983 ^ n2341 ^ 1'b0 ;
  assign n18985 = n18984 ^ n9472 ^ n232 ;
  assign n18986 = n18985 ^ n10426 ^ 1'b0 ;
  assign n18987 = n1128 & ~n11032 ;
  assign n18988 = n18987 ^ n8873 ^ 1'b0 ;
  assign n18989 = n18988 ^ n18045 ^ 1'b0 ;
  assign n18990 = n3035 | n15981 ;
  assign n18991 = n7880 & ~n18990 ;
  assign n18992 = n4200 & ~n8332 ;
  assign n18993 = n18992 ^ n11489 ^ 1'b0 ;
  assign n18995 = n8847 ^ n2299 ^ 1'b0 ;
  assign n18996 = ~n2078 & n18995 ;
  assign n18994 = ~n2221 & n2726 ;
  assign n18997 = n18996 ^ n18994 ^ 1'b0 ;
  assign n18998 = n2484 & ~n7673 ;
  assign n18999 = ~n6900 & n18998 ;
  assign n19000 = n2730 & n14387 ;
  assign n19001 = ~n10558 & n19000 ;
  assign n19002 = ~n4319 & n19001 ;
  assign n19003 = n18584 ^ n7106 ^ n4947 ;
  assign n19004 = n9261 ^ n3920 ^ 1'b0 ;
  assign n19005 = n5897 | n19004 ;
  assign n19006 = ( n11477 & ~n12026 ) | ( n11477 & n16287 ) | ( ~n12026 & n16287 ) ;
  assign n19007 = n19005 & n19006 ;
  assign n19008 = n17708 ^ n10026 ^ 1'b0 ;
  assign n19009 = n6437 ^ n623 ^ 1'b0 ;
  assign n19010 = n6012 ^ n5062 ^ n2118 ;
  assign n19011 = n10149 & ~n10818 ;
  assign n19012 = n658 & ~n4125 ;
  assign n19013 = n6877 ^ n1575 ^ n1257 ;
  assign n19014 = n6963 ^ n3644 ^ 1'b0 ;
  assign n19015 = n19013 | n19014 ;
  assign n19016 = n5315 | n19015 ;
  assign n19017 = n19016 ^ n13397 ^ 1'b0 ;
  assign n19018 = n10109 & n14344 ;
  assign n19019 = n19017 & n19018 ;
  assign n19020 = n13741 ^ n5062 ^ 1'b0 ;
  assign n19021 = n8714 ^ n2312 ^ 1'b0 ;
  assign n19022 = n14742 & n19021 ;
  assign n19025 = ( n2235 & n5885 ) | ( n2235 & ~n7698 ) | ( n5885 & ~n7698 ) ;
  assign n19023 = ~n3526 & n15599 ;
  assign n19024 = n6233 & ~n19023 ;
  assign n19026 = n19025 ^ n19024 ^ 1'b0 ;
  assign n19027 = n11156 ^ n9184 ^ 1'b0 ;
  assign n19028 = n16280 ^ n11449 ^ 1'b0 ;
  assign n19029 = n2970 & ~n19028 ;
  assign n19030 = n3294 & n13794 ;
  assign n19031 = n1300 & n19030 ;
  assign n19032 = n2249 & n3008 ;
  assign n19033 = n19032 ^ n2705 ^ 1'b0 ;
  assign n19034 = ( n6075 & n11320 ) | ( n6075 & ~n19033 ) | ( n11320 & ~n19033 ) ;
  assign n19035 = ~n15305 & n17902 ;
  assign n19036 = n15143 & n19035 ;
  assign n19037 = n1219 | n6207 ;
  assign n19038 = n19037 ^ n8613 ^ 1'b0 ;
  assign n19039 = n612 & n5200 ;
  assign n19040 = n19038 & n19039 ;
  assign n19041 = n14484 ^ n900 ^ 1'b0 ;
  assign n19042 = n5688 & n19041 ;
  assign n19043 = ~n10747 & n12369 ;
  assign n19044 = n2452 & ~n18062 ;
  assign n19045 = ~n9890 & n19044 ;
  assign n19046 = n7291 | n19045 ;
  assign n19047 = n6981 & n17149 ;
  assign n19048 = n19047 ^ n10189 ^ 1'b0 ;
  assign n19049 = n1541 & n3354 ;
  assign n19050 = n3056 & n19049 ;
  assign n19051 = ( n1266 & ~n8059 ) | ( n1266 & n9207 ) | ( ~n8059 & n9207 ) ;
  assign n19052 = n19051 ^ n7968 ^ 1'b0 ;
  assign n19053 = ~n19050 & n19052 ;
  assign n19054 = n13087 & ~n16434 ;
  assign n19055 = n11018 ^ n7425 ^ 1'b0 ;
  assign n19056 = ( ~n753 & n1143 ) | ( ~n753 & n19055 ) | ( n1143 & n19055 ) ;
  assign n19057 = n6606 ^ n4319 ^ 1'b0 ;
  assign n19058 = ~n6348 & n19057 ;
  assign n19059 = n19058 ^ n7413 ^ 1'b0 ;
  assign n19060 = n19056 & ~n19059 ;
  assign n19061 = n4922 & n8947 ;
  assign n19062 = n8845 ^ n900 ^ 1'b0 ;
  assign n19063 = n19061 & n19062 ;
  assign n19068 = n6153 | n13360 ;
  assign n19066 = n10668 | n15842 ;
  assign n19067 = n19066 ^ n2312 ^ 1'b0 ;
  assign n19064 = n12978 & ~n13502 ;
  assign n19065 = n4281 & n19064 ;
  assign n19069 = n19068 ^ n19067 ^ n19065 ;
  assign n19070 = n12147 | n18366 ;
  assign n19071 = n5789 ^ n5317 ^ n2953 ;
  assign n19072 = n11224 & ~n19071 ;
  assign n19073 = n19072 ^ n3259 ^ 1'b0 ;
  assign n19074 = n5860 & n19073 ;
  assign n19075 = n9904 ^ n7163 ^ 1'b0 ;
  assign n19076 = ~n14585 & n19075 ;
  assign n19077 = n9882 & ~n12224 ;
  assign n19078 = n15600 ^ n6590 ^ 1'b0 ;
  assign n19081 = n5264 ^ n2557 ^ 1'b0 ;
  assign n19082 = ~n2758 & n19081 ;
  assign n19079 = ~n2945 & n16495 ;
  assign n19080 = n11913 & ~n19079 ;
  assign n19083 = n19082 ^ n19080 ^ n10284 ;
  assign n19084 = n19083 ^ n14187 ^ n12191 ;
  assign n19085 = ~n5594 & n19084 ;
  assign n19086 = ~n12091 & n19085 ;
  assign n19087 = n8738 | n13802 ;
  assign n19088 = n15531 & ~n19087 ;
  assign n19089 = n4781 & ~n19088 ;
  assign n19090 = ~n1632 & n13356 ;
  assign n19091 = n17122 & n19090 ;
  assign n19092 = n17073 ^ n3426 ^ 1'b0 ;
  assign n19093 = n3897 & ~n19092 ;
  assign n19094 = n928 & n19093 ;
  assign n19095 = n9960 ^ n560 ^ 1'b0 ;
  assign n19096 = n9920 ^ n5501 ^ 1'b0 ;
  assign n19097 = n3148 & ~n8801 ;
  assign n19098 = n8850 & ~n12707 ;
  assign n19099 = n14505 ^ n3687 ^ 1'b0 ;
  assign n19100 = n7208 | n19099 ;
  assign n19101 = n11369 ^ n456 ^ 1'b0 ;
  assign n19102 = n19100 | n19101 ;
  assign n19103 = n7872 | n9263 ;
  assign n19104 = n19103 ^ n1212 ^ 1'b0 ;
  assign n19105 = ~n2330 & n8868 ;
  assign n19106 = n19105 ^ n18749 ^ n4981 ;
  assign n19108 = n4814 ^ n3086 ^ 1'b0 ;
  assign n19107 = n3058 & n3908 ;
  assign n19109 = n19108 ^ n19107 ^ 1'b0 ;
  assign n19110 = n11453 ^ n10549 ^ 1'b0 ;
  assign n19111 = ~n11964 & n19110 ;
  assign n19112 = n19111 ^ n11596 ^ 1'b0 ;
  assign n19113 = n15328 ^ n14781 ^ 1'b0 ;
  assign n19114 = n6013 & ~n15249 ;
  assign n19115 = n19114 ^ n13474 ^ 1'b0 ;
  assign n19116 = n788 & ~n6407 ;
  assign n19117 = ~n2948 & n19116 ;
  assign n19118 = n19117 ^ n8268 ^ 1'b0 ;
  assign n19119 = n19118 ^ n7709 ^ 1'b0 ;
  assign n19120 = n16508 & n19119 ;
  assign n19121 = n19120 ^ n13643 ^ n7578 ;
  assign n19122 = ~n1225 & n5435 ;
  assign n19123 = n19122 ^ n2872 ^ 1'b0 ;
  assign n19124 = n4020 & ~n19123 ;
  assign n19125 = n3082 | n5755 ;
  assign n19126 = n19124 | n19125 ;
  assign n19127 = n8817 ^ n1396 ^ 1'b0 ;
  assign n19128 = n19126 & n19127 ;
  assign n19129 = ~n4204 & n5055 ;
  assign n19130 = n19129 ^ n8027 ^ 1'b0 ;
  assign n19131 = n16816 & ~n19130 ;
  assign n19132 = n16282 ^ n3887 ^ n2787 ;
  assign n19134 = n2927 ^ n559 ^ n391 ;
  assign n19135 = n3601 & n19134 ;
  assign n19133 = n7247 | n18037 ;
  assign n19136 = n19135 ^ n19133 ^ 1'b0 ;
  assign n19137 = n3974 ^ n3528 ^ 1'b0 ;
  assign n19138 = n5475 & ~n19137 ;
  assign n19139 = n6472 | n19138 ;
  assign n19140 = n1211 ^ n821 ^ 1'b0 ;
  assign n19141 = n2228 & n10258 ;
  assign n19142 = ( n6749 & ~n14641 ) | ( n6749 & n19141 ) | ( ~n14641 & n19141 ) ;
  assign n19143 = n1888 ^ n1204 ^ 1'b0 ;
  assign n19144 = n9012 & ~n13599 ;
  assign n19145 = n6461 & n19144 ;
  assign n19147 = n5623 | n5850 ;
  assign n19148 = n19147 ^ n600 ^ 1'b0 ;
  assign n19146 = n2412 & n10343 ;
  assign n19149 = n19148 ^ n19146 ^ 1'b0 ;
  assign n19150 = n1911 & ~n3143 ;
  assign n19151 = n19150 ^ n11863 ^ 1'b0 ;
  assign n19152 = n10026 & ~n14994 ;
  assign n19153 = n505 & n9987 ;
  assign n19154 = ~n3526 & n11527 ;
  assign n19155 = n16566 & n19154 ;
  assign n19156 = n9146 | n11655 ;
  assign n19157 = ~n662 & n18252 ;
  assign n19158 = n14038 & ~n15978 ;
  assign n19159 = n9438 ^ n1601 ^ 1'b0 ;
  assign n19160 = n3895 & n6966 ;
  assign n19161 = n19160 ^ n11036 ^ n2967 ;
  assign n19162 = n18537 ^ n3702 ^ n2983 ;
  assign n19163 = n8706 ^ n3824 ^ 1'b0 ;
  assign n19164 = n13368 | n14225 ;
  assign n19165 = n15294 & ~n19164 ;
  assign n19166 = n14132 & ~n17349 ;
  assign n19167 = n15387 ^ n5187 ^ 1'b0 ;
  assign n19168 = n10878 | n19167 ;
  assign n19169 = n12031 & ~n19168 ;
  assign n19170 = n4800 & n12728 ;
  assign n19171 = n16098 ^ n2903 ^ 1'b0 ;
  assign n19172 = n8741 ^ n5306 ^ 1'b0 ;
  assign n19173 = n2818 | n19172 ;
  assign n19174 = n19173 ^ n17176 ^ 1'b0 ;
  assign n19176 = n5427 & ~n12682 ;
  assign n19177 = ~n7449 & n19176 ;
  assign n19175 = n3212 & ~n9768 ;
  assign n19178 = n19177 ^ n19175 ^ 1'b0 ;
  assign n19179 = n18692 ^ n923 ^ 1'b0 ;
  assign n19180 = n6054 & ~n19179 ;
  assign n19181 = ~n12043 & n17483 ;
  assign n19182 = n12535 ^ n8858 ^ 1'b0 ;
  assign n19183 = n13446 | n19182 ;
  assign n19184 = n5981 ^ n2151 ^ 1'b0 ;
  assign n19185 = n1599 & n3328 ;
  assign n19186 = n19184 & n19185 ;
  assign n19187 = n15080 & ~n19019 ;
  assign n19188 = n19187 ^ x46 ^ 1'b0 ;
  assign n19189 = n4308 & ~n9642 ;
  assign n19190 = n8711 & n19189 ;
  assign n19191 = n4694 | n18050 ;
  assign n19192 = n1812 & n8236 ;
  assign n19193 = n10794 & n19192 ;
  assign n19194 = n10554 & ~n15995 ;
  assign n19195 = n19194 ^ n11410 ^ 1'b0 ;
  assign n19196 = n6465 & n9236 ;
  assign n19197 = ( n2942 & ~n5667 ) | ( n2942 & n14036 ) | ( ~n5667 & n14036 ) ;
  assign n19198 = n19197 ^ n11381 ^ n3757 ;
  assign n19199 = n19198 ^ n4909 ^ 1'b0 ;
  assign n19200 = n531 | n2714 ;
  assign n19201 = n5885 | n19200 ;
  assign n19202 = ~x81 & n10747 ;
  assign n19203 = ( ~n2917 & n7595 ) | ( ~n2917 & n7953 ) | ( n7595 & n7953 ) ;
  assign n19204 = n17079 ^ n8856 ^ 1'b0 ;
  assign n19205 = n3543 & ~n5152 ;
  assign n19206 = n5951 & ~n19205 ;
  assign n19207 = ~n16244 & n19206 ;
  assign n19208 = n17876 | n18193 ;
  assign n19209 = n10198 | n14825 ;
  assign n19210 = n5985 | n19209 ;
  assign n19211 = ~n4022 & n8187 ;
  assign n19212 = ~n4678 & n19211 ;
  assign n19213 = n898 | n1425 ;
  assign n19214 = n3987 & ~n19213 ;
  assign n19215 = n10825 | n19214 ;
  assign n19216 = n19215 ^ n19143 ^ 1'b0 ;
  assign n19217 = n18289 & ~n19216 ;
  assign n19218 = n7988 ^ n6191 ^ 1'b0 ;
  assign n19219 = ~n7763 & n19218 ;
  assign n19220 = n19219 ^ n8119 ^ 1'b0 ;
  assign n19221 = n2952 & ~n19220 ;
  assign n19222 = n8284 ^ n6653 ^ 1'b0 ;
  assign n19223 = n4784 & n5485 ;
  assign n19224 = n17361 | n17571 ;
  assign n19225 = n19223 & ~n19224 ;
  assign n19226 = n1939 & ~n5453 ;
  assign n19227 = n9150 & n19226 ;
  assign n19228 = n7852 | n9240 ;
  assign n19229 = n19227 & ~n19228 ;
  assign n19230 = n209 | n1787 ;
  assign n19231 = n19230 ^ n17206 ^ 1'b0 ;
  assign n19232 = n2986 & n19231 ;
  assign n19233 = n19229 | n19232 ;
  assign n19234 = n12171 & ~n13012 ;
  assign n19235 = n5836 & ~n9488 ;
  assign n19236 = n4624 & ~n19235 ;
  assign n19237 = ~n15223 & n19236 ;
  assign n19238 = n4588 | n9012 ;
  assign n19239 = n1325 | n19238 ;
  assign n19240 = n4743 ^ n4448 ^ 1'b0 ;
  assign n19241 = n4430 & ~n19240 ;
  assign n19242 = n19241 ^ n2596 ^ 1'b0 ;
  assign n19245 = ~n5865 & n6497 ;
  assign n19246 = ~n706 & n2877 ;
  assign n19247 = n19246 ^ n184 ^ 1'b0 ;
  assign n19248 = n19245 | n19247 ;
  assign n19249 = n19248 ^ n13224 ^ 1'b0 ;
  assign n19243 = ~n5203 & n16840 ;
  assign n19244 = ~n12880 & n19243 ;
  assign n19250 = n19249 ^ n19244 ^ 1'b0 ;
  assign n19251 = n4868 ^ n1689 ^ 1'b0 ;
  assign n19252 = n4153 ^ n849 ^ 1'b0 ;
  assign n19253 = ~n2135 & n19252 ;
  assign n19254 = n19253 ^ n16034 ^ 1'b0 ;
  assign n19255 = n19254 ^ n3950 ^ 1'b0 ;
  assign n19256 = n9812 | n19255 ;
  assign n19262 = n435 & ~n2810 ;
  assign n19263 = ~n7038 & n19262 ;
  assign n19259 = n4953 ^ n1933 ^ 1'b0 ;
  assign n19260 = n7578 | n19259 ;
  assign n19261 = n19260 ^ n10301 ^ 1'b0 ;
  assign n19257 = n10024 ^ n7723 ^ n6545 ;
  assign n19258 = n19257 ^ n2313 ^ 1'b0 ;
  assign n19264 = n19263 ^ n19261 ^ n19258 ;
  assign n19265 = ( n1623 & ~n5808 ) | ( n1623 & n19264 ) | ( ~n5808 & n19264 ) ;
  assign n19266 = n6334 ^ n1028 ^ 1'b0 ;
  assign n19267 = n7221 & ~n19266 ;
  assign n19268 = n13495 ^ n2880 ^ 1'b0 ;
  assign n19269 = ( n639 & ~n2302 ) | ( n639 & n5632 ) | ( ~n2302 & n5632 ) ;
  assign n19270 = n10838 & ~n19015 ;
  assign n19271 = n8838 & ~n18341 ;
  assign n19272 = n13612 ^ n1579 ^ 1'b0 ;
  assign n19273 = n8749 ^ n5593 ^ 1'b0 ;
  assign n19274 = ~n19272 & n19273 ;
  assign n19275 = n5165 & n11195 ;
  assign n19276 = ~n6800 & n7646 ;
  assign n19277 = ~n4793 & n19276 ;
  assign n19278 = ~n6854 & n13808 ;
  assign n19279 = n4831 ^ n867 ^ 1'b0 ;
  assign n19280 = ~n2254 & n19279 ;
  assign n19281 = n808 & n19280 ;
  assign n19282 = n19281 ^ n7183 ^ 1'b0 ;
  assign n19283 = ~n5404 & n5972 ;
  assign n19284 = n19283 ^ n5151 ^ x74 ;
  assign n19285 = n8082 ^ n5429 ^ 1'b0 ;
  assign n19286 = n5625 & n19285 ;
  assign n19287 = n19286 ^ n2543 ^ 1'b0 ;
  assign n19288 = n10594 | n19287 ;
  assign n19289 = ~n1868 & n5442 ;
  assign n19290 = n2992 & ~n15721 ;
  assign n19291 = n9696 & ~n13017 ;
  assign n19292 = n16678 ^ n15778 ^ 1'b0 ;
  assign n19293 = n9532 & ~n12797 ;
  assign n19294 = ( n8132 & ~n13425 ) | ( n8132 & n19293 ) | ( ~n13425 & n19293 ) ;
  assign n19295 = n8176 & n19294 ;
  assign n19296 = n17754 ^ n9865 ^ 1'b0 ;
  assign n19299 = ~n7164 & n9141 ;
  assign n19297 = ~n1111 & n9833 ;
  assign n19298 = ~n10587 & n19297 ;
  assign n19300 = n19299 ^ n19298 ^ 1'b0 ;
  assign n19301 = ~n2752 & n18830 ;
  assign n19302 = ~n18830 & n19301 ;
  assign n19303 = ~n272 & n11527 ;
  assign n19304 = n19303 ^ n9703 ^ 1'b0 ;
  assign n19306 = n8797 ^ n4843 ^ 1'b0 ;
  assign n19305 = n2180 & n18129 ;
  assign n19307 = n19306 ^ n19305 ^ 1'b0 ;
  assign n19308 = n5967 & ~n19307 ;
  assign n19309 = n19308 ^ n2289 ^ 1'b0 ;
  assign n19310 = n5685 & n19309 ;
  assign n19311 = n3987 ^ x55 ^ 1'b0 ;
  assign n19312 = n4618 & ~n19311 ;
  assign n19313 = n17978 ^ n11011 ^ n2463 ;
  assign n19314 = ( ~n6477 & n9005 ) | ( ~n6477 & n14240 ) | ( n9005 & n14240 ) ;
  assign n19315 = n9731 ^ n2972 ^ 1'b0 ;
  assign n19316 = ~n1886 & n4558 ;
  assign n19317 = n11320 ^ n7371 ^ 1'b0 ;
  assign n19318 = n16789 & ~n19317 ;
  assign n19319 = n19318 ^ n10838 ^ 1'b0 ;
  assign n19320 = n3343 | n4987 ;
  assign n19321 = n19320 ^ n1689 ^ 1'b0 ;
  assign n19322 = n3654 | n11962 ;
  assign n19323 = ( n5183 & ~n9610 ) | ( n5183 & n18551 ) | ( ~n9610 & n18551 ) ;
  assign n19324 = ( n1470 & n19322 ) | ( n1470 & ~n19323 ) | ( n19322 & ~n19323 ) ;
  assign n19325 = n12686 & n19324 ;
  assign n19326 = ( n7023 & n19321 ) | ( n7023 & ~n19325 ) | ( n19321 & ~n19325 ) ;
  assign n19327 = n5079 & n19326 ;
  assign n19328 = n19327 ^ n4676 ^ 1'b0 ;
  assign n19329 = ~n1199 & n16157 ;
  assign n19330 = n19329 ^ n1244 ^ 1'b0 ;
  assign n19331 = n19254 ^ n8273 ^ 1'b0 ;
  assign n19332 = n14887 ^ n9066 ^ 1'b0 ;
  assign n19333 = n9949 ^ n844 ^ 1'b0 ;
  assign n19334 = n4800 & ~n19333 ;
  assign n19335 = n5756 & ~n15546 ;
  assign n19336 = n13794 ^ n11789 ^ 1'b0 ;
  assign n19337 = ~n180 & n8500 ;
  assign n19338 = ~n2621 & n19337 ;
  assign n19339 = n19338 ^ n14934 ^ 1'b0 ;
  assign n19340 = n7336 ^ n1792 ^ 1'b0 ;
  assign n19341 = n17989 & n19340 ;
  assign n19342 = n1200 & n10938 ;
  assign n19343 = ~n5674 & n19342 ;
  assign n19344 = n19343 ^ n9372 ^ 1'b0 ;
  assign n19345 = n19341 & n19344 ;
  assign n19346 = n19345 ^ n10993 ^ 1'b0 ;
  assign n19347 = n2556 | n3319 ;
  assign n19348 = n19347 ^ n853 ^ 1'b0 ;
  assign n19349 = n484 & ~n4753 ;
  assign n19350 = ~n4870 & n9392 ;
  assign n19351 = n9724 & n19350 ;
  assign n19352 = n2179 & ~n8687 ;
  assign n19353 = n18093 ^ n6152 ^ 1'b0 ;
  assign n19354 = n808 | n19353 ;
  assign n19355 = n19354 ^ n1645 ^ 1'b0 ;
  assign n19356 = ~n13516 & n19355 ;
  assign n19357 = n1212 & ~n1761 ;
  assign n19358 = ~n17904 & n19357 ;
  assign n19359 = ~n9865 & n17879 ;
  assign n19360 = n1079 & n19359 ;
  assign n19361 = n4051 & ~n7968 ;
  assign n19362 = n6069 ^ n3790 ^ n679 ;
  assign n19363 = n4433 ^ n2093 ^ 1'b0 ;
  assign n19364 = n3007 & ~n19363 ;
  assign n19365 = n2604 | n19364 ;
  assign n19366 = n3689 | n4455 ;
  assign n19367 = n19366 ^ n3580 ^ 1'b0 ;
  assign n19368 = ( n5727 & ~n6378 ) | ( n5727 & n18343 ) | ( ~n6378 & n18343 ) ;
  assign n19369 = n3543 | n3623 ;
  assign n19370 = n19369 ^ n5461 ^ 1'b0 ;
  assign n19371 = n11297 & ~n19370 ;
  assign n19372 = ~n9835 & n12967 ;
  assign n19373 = ~x52 & n19372 ;
  assign n19374 = n13397 ^ n3869 ^ 1'b0 ;
  assign n19375 = n10568 & n14187 ;
  assign n19376 = n983 | n16599 ;
  assign n19377 = n4820 ^ n2365 ^ 1'b0 ;
  assign n19378 = n3784 | n19377 ;
  assign n19379 = n3998 & ~n15776 ;
  assign n19380 = ~n3069 & n12920 ;
  assign n19381 = ~n1089 & n1378 ;
  assign n19382 = n19381 ^ n1103 ^ 1'b0 ;
  assign n19383 = n19382 ^ n4427 ^ 1'b0 ;
  assign n19384 = ~n13292 & n19383 ;
  assign n19385 = n6531 & n18843 ;
  assign n19386 = n5594 & ~n5672 ;
  assign n19387 = n7375 & n12583 ;
  assign n19388 = n1951 | n7866 ;
  assign n19389 = n11737 ^ n2494 ^ 1'b0 ;
  assign n19390 = n14920 ^ n11305 ^ n8146 ;
  assign n19391 = n2454 | n19390 ;
  assign n19392 = n1222 & n6886 ;
  assign n19393 = ~n9071 & n19392 ;
  assign n19394 = n7662 ^ n3334 ^ 1'b0 ;
  assign n19395 = ~n3095 & n3233 ;
  assign n19396 = ~n509 & n19395 ;
  assign n19397 = ~n358 & n2674 ;
  assign n19398 = n9820 | n15942 ;
  assign n19399 = n19397 | n19398 ;
  assign n19400 = n19399 ^ n2635 ^ 1'b0 ;
  assign n19401 = ~n3118 & n19400 ;
  assign n19402 = n2060 ^ n1244 ^ 1'b0 ;
  assign n19403 = ~n6364 & n11200 ;
  assign n19404 = n13992 & n19403 ;
  assign n19405 = n13549 & ~n19404 ;
  assign n19406 = n19405 ^ n16252 ^ 1'b0 ;
  assign n19407 = n19406 ^ n12243 ^ 1'b0 ;
  assign n19408 = n444 | n2621 ;
  assign n19409 = n7621 | n19408 ;
  assign n19410 = ~n2006 & n16515 ;
  assign n19411 = ( ~n3992 & n4659 ) | ( ~n3992 & n7558 ) | ( n4659 & n7558 ) ;
  assign n19412 = n17120 ^ n14587 ^ 1'b0 ;
  assign n19413 = ~n15802 & n19412 ;
  assign n19414 = n3326 & ~n19413 ;
  assign n19415 = n4578 ^ n190 ^ 1'b0 ;
  assign n19416 = ~n2018 & n19415 ;
  assign n19417 = n2545 ^ n2372 ^ 1'b0 ;
  assign n19418 = n4292 | n19417 ;
  assign n19419 = n19260 ^ n14099 ^ 1'b0 ;
  assign n19420 = n19419 ^ n8583 ^ 1'b0 ;
  assign n19421 = ~n19418 & n19420 ;
  assign n19422 = n10664 ^ n5909 ^ 1'b0 ;
  assign n19423 = n11611 & ~n19422 ;
  assign n19424 = n19423 ^ n1393 ^ 1'b0 ;
  assign n19425 = n9380 & ~n19424 ;
  assign n19426 = n5144 & n9208 ;
  assign n19427 = n9411 | n10127 ;
  assign n19428 = n756 & ~n19427 ;
  assign n19429 = n19426 | n19428 ;
  assign n19430 = n19425 | n19429 ;
  assign n19431 = n19430 ^ n14061 ^ 1'b0 ;
  assign n19432 = n7741 & ~n10203 ;
  assign n19433 = ~n7741 & n19432 ;
  assign n19434 = n19433 ^ n2931 ^ 1'b0 ;
  assign n19435 = n6188 & n8572 ;
  assign n19436 = n2838 & n19435 ;
  assign n19437 = n15042 | n16898 ;
  assign n19438 = n19436 & ~n19437 ;
  assign n19439 = n9686 & n12251 ;
  assign n19440 = ~n17385 & n19439 ;
  assign n19441 = ( n397 & n9129 ) | ( n397 & ~n19047 ) | ( n9129 & ~n19047 ) ;
  assign n19442 = ( n2853 & n17585 ) | ( n2853 & ~n19119 ) | ( n17585 & ~n19119 ) ;
  assign n19443 = n10779 & ~n17970 ;
  assign n19444 = n9100 ^ n1444 ^ 1'b0 ;
  assign n19445 = n19443 | n19444 ;
  assign n19446 = n16968 ^ n11274 ^ 1'b0 ;
  assign n19447 = ~n9650 & n16942 ;
  assign n19448 = n19447 ^ n9886 ^ 1'b0 ;
  assign n19449 = n12970 ^ n503 ^ 1'b0 ;
  assign n19450 = n5592 & n19449 ;
  assign n19451 = n19257 & n19450 ;
  assign n19452 = n6441 & n19451 ;
  assign n19453 = n17266 ^ n16249 ^ n5684 ;
  assign n19454 = n11699 ^ n6459 ^ 1'b0 ;
  assign n19455 = n5285 | n15928 ;
  assign n19456 = ~n4373 & n12309 ;
  assign n19457 = n19456 ^ n8989 ^ 1'b0 ;
  assign n19461 = n8962 & n13204 ;
  assign n19462 = n19461 ^ n5015 ^ 1'b0 ;
  assign n19458 = n1204 & ~n4295 ;
  assign n19459 = n19458 ^ n2765 ^ 1'b0 ;
  assign n19460 = ~n17059 & n19459 ;
  assign n19463 = n19462 ^ n19460 ^ 1'b0 ;
  assign n19464 = n527 | n1947 ;
  assign n19465 = n3055 & ~n19263 ;
  assign n19467 = n2466 & n3748 ;
  assign n19466 = n6790 & ~n12340 ;
  assign n19468 = n19467 ^ n19466 ^ 1'b0 ;
  assign n19469 = ~n2428 & n17320 ;
  assign n19470 = n19469 ^ n10136 ^ 1'b0 ;
  assign n19471 = n19470 ^ n14486 ^ 1'b0 ;
  assign n19472 = n17811 ^ n5403 ^ 1'b0 ;
  assign n19473 = n12091 ^ n9953 ^ 1'b0 ;
  assign n19474 = n604 & ~n19473 ;
  assign n19475 = n5850 | n18856 ;
  assign n19476 = n3011 ^ n2312 ^ 1'b0 ;
  assign n19477 = n15584 & n19476 ;
  assign n19478 = n19477 ^ n8779 ^ n5085 ;
  assign n19479 = n2862 & ~n14190 ;
  assign n19480 = n19479 ^ n6932 ^ 1'b0 ;
  assign n19481 = n3460 | n6630 ;
  assign n19482 = n874 | n19481 ;
  assign n19483 = ~n1560 & n8142 ;
  assign n19484 = n19483 ^ n12762 ^ 1'b0 ;
  assign n19485 = ( n4705 & ~n8449 ) | ( n4705 & n19484 ) | ( ~n8449 & n19484 ) ;
  assign n19486 = n10482 ^ n1479 ^ n1077 ;
  assign n19487 = ~n13734 & n19486 ;
  assign n19488 = ( n796 & n1970 ) | ( n796 & n12096 ) | ( n1970 & n12096 ) ;
  assign n19489 = n5695 & n18898 ;
  assign n19490 = n19488 & ~n19489 ;
  assign n19491 = n8260 & n19490 ;
  assign n19492 = n17064 ^ n1778 ^ 1'b0 ;
  assign n19493 = n14480 & ~n19492 ;
  assign n19494 = n8833 ^ n4013 ^ 1'b0 ;
  assign n19495 = n3988 | n19494 ;
  assign n19496 = n1629 | n10479 ;
  assign n19497 = n17861 | n19496 ;
  assign n19498 = n1881 & ~n9629 ;
  assign n19499 = n19498 ^ n12030 ^ n8630 ;
  assign n19500 = ~n11275 & n13070 ;
  assign n19501 = n19500 ^ n10530 ^ 1'b0 ;
  assign n19502 = n10602 | n12583 ;
  assign n19503 = n10130 & ~n15633 ;
  assign n19506 = n6376 ^ n3209 ^ 1'b0 ;
  assign n19507 = n5422 & ~n19506 ;
  assign n19504 = n10754 ^ n2898 ^ 1'b0 ;
  assign n19505 = ~n9732 & n19504 ;
  assign n19508 = n19507 ^ n19505 ^ n1355 ;
  assign n19509 = n19508 ^ n13017 ^ n8577 ;
  assign n19510 = n553 & n11391 ;
  assign n19511 = ~n2423 & n2553 ;
  assign n19512 = n19511 ^ n14553 ^ 1'b0 ;
  assign n19515 = n244 | n299 ;
  assign n19516 = n19515 ^ n7504 ^ 1'b0 ;
  assign n19517 = n4556 & n7934 ;
  assign n19518 = n1978 & n19517 ;
  assign n19519 = n17133 | n19518 ;
  assign n19520 = n19519 ^ n2305 ^ 1'b0 ;
  assign n19521 = n19516 & n19520 ;
  assign n19514 = n2176 & n9804 ;
  assign n19513 = n6855 & ~n8106 ;
  assign n19522 = n19521 ^ n19514 ^ n19513 ;
  assign n19523 = n2121 & ~n7575 ;
  assign n19524 = n17259 & n19523 ;
  assign n19525 = n6356 | n18377 ;
  assign n19526 = n1308 ^ x56 ^ 1'b0 ;
  assign n19527 = n4451 & n19526 ;
  assign n19528 = n13040 | n14696 ;
  assign n19529 = n19527 | n19528 ;
  assign n19530 = ( ~n732 & n7736 ) | ( ~n732 & n16457 ) | ( n7736 & n16457 ) ;
  assign n19531 = n1569 & ~n9286 ;
  assign n19536 = n2561 & n10054 ;
  assign n19537 = ~n10775 & n19536 ;
  assign n19532 = ~n9051 & n14108 ;
  assign n19533 = n12247 ^ n5805 ^ n1295 ;
  assign n19534 = n14619 | n19533 ;
  assign n19535 = n19532 | n19534 ;
  assign n19538 = n19537 ^ n19535 ^ 1'b0 ;
  assign n19539 = n3837 & ~n10061 ;
  assign n19540 = ~n9530 & n19539 ;
  assign n19541 = n3903 | n19540 ;
  assign n19542 = n13810 & ~n19541 ;
  assign n19543 = n4669 ^ n3649 ^ 1'b0 ;
  assign n19544 = ~n8508 & n15964 ;
  assign n19545 = n3921 & n4793 ;
  assign n19546 = n19545 ^ n8552 ^ 1'b0 ;
  assign n19547 = ~n18382 & n19546 ;
  assign n19551 = n283 & ~n8844 ;
  assign n19552 = n4883 | n19551 ;
  assign n19548 = n5448 ^ n5093 ^ 1'b0 ;
  assign n19549 = n4978 | n19548 ;
  assign n19550 = n11603 | n19549 ;
  assign n19553 = n19552 ^ n19550 ^ 1'b0 ;
  assign n19554 = n4942 & n9717 ;
  assign n19555 = n9570 & ~n19554 ;
  assign n19556 = ~n2280 & n12994 ;
  assign n19557 = n591 & n3319 ;
  assign n19558 = n11202 ^ n3253 ^ 1'b0 ;
  assign n19559 = n1793 & ~n8595 ;
  assign n19560 = n17489 ^ n12837 ^ 1'b0 ;
  assign n19561 = ( n1133 & ~n7659 ) | ( n1133 & n19560 ) | ( ~n7659 & n19560 ) ;
  assign n19562 = n15310 ^ n4611 ^ 1'b0 ;
  assign n19563 = n19561 & ~n19562 ;
  assign n19564 = n6949 & n10550 ;
  assign n19565 = n19564 ^ n14801 ^ 1'b0 ;
  assign n19566 = ~n1386 & n5608 ;
  assign n19567 = n19566 ^ n9236 ^ 1'b0 ;
  assign n19568 = n11419 | n19567 ;
  assign n19569 = n19565 | n19568 ;
  assign n19570 = n3655 | n6017 ;
  assign n19571 = n12249 ^ n6327 ^ 1'b0 ;
  assign n19572 = n1962 & ~n19571 ;
  assign n19573 = n7765 & ~n16573 ;
  assign n19574 = n19573 ^ n10133 ^ 1'b0 ;
  assign n19575 = n19574 ^ n3483 ^ 1'b0 ;
  assign n19576 = n19575 ^ n134 ^ 1'b0 ;
  assign n19577 = n12150 & ~n19576 ;
  assign n19578 = n19577 ^ x79 ^ 1'b0 ;
  assign n19579 = n19572 & ~n19578 ;
  assign n19580 = n14468 ^ n11945 ^ n229 ;
  assign n19581 = n1637 | n6252 ;
  assign n19582 = n4334 & ~n19581 ;
  assign n19583 = n19582 ^ n15784 ^ 1'b0 ;
  assign n19584 = n3233 | n6545 ;
  assign n19585 = ~n7337 & n9765 ;
  assign n19586 = n19584 & n19585 ;
  assign n19587 = n14573 ^ n10190 ^ n4633 ;
  assign n19588 = n19587 ^ n6618 ^ 1'b0 ;
  assign n19589 = n5219 & n19588 ;
  assign n19590 = n14643 ^ n553 ^ 1'b0 ;
  assign n19591 = n12409 ^ n5363 ^ x119 ;
  assign n19592 = n19591 ^ n2262 ^ n417 ;
  assign n19593 = n16186 & ~n19592 ;
  assign n19594 = n19593 ^ n8016 ^ 1'b0 ;
  assign n19595 = ~n4095 & n19594 ;
  assign n19599 = n1676 & n2153 ;
  assign n19597 = ~n1231 & n7577 ;
  assign n19598 = n930 & n19597 ;
  assign n19600 = n19599 ^ n19598 ^ 1'b0 ;
  assign n19596 = n6818 & ~n7033 ;
  assign n19601 = n19600 ^ n19596 ^ n14610 ;
  assign n19603 = n11241 ^ n7690 ^ 1'b0 ;
  assign n19604 = n5957 | n19603 ;
  assign n19602 = n1527 & ~n9385 ;
  assign n19605 = n19604 ^ n19602 ^ n10050 ;
  assign n19606 = n2392 | n9367 ;
  assign n19607 = n19605 & ~n19606 ;
  assign n19608 = ~n2344 & n3953 ;
  assign n19609 = n10161 & ~n15464 ;
  assign n19610 = n11983 ^ n669 ^ 1'b0 ;
  assign n19611 = n1200 & n19610 ;
  assign n19612 = n1011 | n6120 ;
  assign n19613 = n19612 ^ n12226 ^ 1'b0 ;
  assign n19614 = n7764 & ~n14333 ;
  assign n19615 = n16521 & n19614 ;
  assign n19616 = n9092 & ~n19615 ;
  assign n19617 = n16956 ^ n2678 ^ 1'b0 ;
  assign n19618 = n9722 | n19617 ;
  assign n19619 = n5546 & n19618 ;
  assign n19620 = n1248 | n19619 ;
  assign n19621 = n15618 & ~n19620 ;
  assign n19622 = n15731 ^ n1937 ^ 1'b0 ;
  assign n19623 = n10728 & n11117 ;
  assign n19624 = n19583 ^ n5733 ^ 1'b0 ;
  assign n19625 = n13384 | n16643 ;
  assign n19626 = n1300 & ~n4411 ;
  assign n19627 = ( n1224 & n1772 ) | ( n1224 & ~n3414 ) | ( n1772 & ~n3414 ) ;
  assign n19628 = n19627 ^ n17850 ^ 1'b0 ;
  assign n19629 = n19626 | n19628 ;
  assign n19630 = n4747 | n16314 ;
  assign n19631 = x45 & n17547 ;
  assign n19632 = n19631 ^ n3737 ^ n1831 ;
  assign n19633 = n19630 | n19632 ;
  assign n19634 = n7451 | n10418 ;
  assign n19635 = n7137 | n19634 ;
  assign n19636 = n19633 | n19635 ;
  assign n19637 = n5693 & ~n9759 ;
  assign n19638 = n19637 ^ n5463 ^ 1'b0 ;
  assign n19639 = n19638 ^ n6050 ^ 1'b0 ;
  assign n19640 = n16056 & n19639 ;
  assign n19641 = n19640 ^ n18759 ^ n12129 ;
  assign n19642 = n11891 & n16323 ;
  assign n19643 = n471 & n7730 ;
  assign n19644 = ~n13465 & n19643 ;
  assign n19645 = n19644 ^ n7698 ^ 1'b0 ;
  assign n19646 = n12188 & ~n13521 ;
  assign n19647 = ~n2823 & n19646 ;
  assign n19648 = n12260 & ~n13854 ;
  assign n19649 = ~n2563 & n2904 ;
  assign n19650 = n589 & n767 ;
  assign n19651 = ~n589 & n19650 ;
  assign n19652 = n10734 & ~n19651 ;
  assign n19653 = ~n8089 & n19652 ;
  assign n19654 = ~n19652 & n19653 ;
  assign n19655 = ( n1195 & n17301 ) | ( n1195 & n19654 ) | ( n17301 & n19654 ) ;
  assign n19656 = n14655 ^ n5667 ^ n2826 ;
  assign n19657 = ~n8803 & n19656 ;
  assign n19658 = n3099 ^ n1911 ^ 1'b0 ;
  assign n19659 = ~n1750 & n19658 ;
  assign n19660 = n6432 ^ n468 ^ 1'b0 ;
  assign n19661 = n1070 ^ n787 ^ n525 ;
  assign n19662 = n19661 ^ n7698 ^ n3514 ;
  assign n19663 = ~n5471 & n13443 ;
  assign n19664 = n19663 ^ n3055 ^ 1'b0 ;
  assign n19665 = n15024 | n19664 ;
  assign n19669 = n180 & n3025 ;
  assign n19670 = ~n180 & n19669 ;
  assign n19671 = n10831 | n14561 ;
  assign n19672 = n1259 & ~n19671 ;
  assign n19673 = n19671 & n19672 ;
  assign n19674 = n19670 | n19673 ;
  assign n19666 = n11300 ^ n3792 ^ 1'b0 ;
  assign n19667 = n824 & ~n19666 ;
  assign n19668 = ~n824 & n19667 ;
  assign n19675 = n19674 ^ n19668 ^ 1'b0 ;
  assign n19676 = ~n11767 & n19675 ;
  assign n19677 = n13176 & n16778 ;
  assign n19678 = n3504 ^ n3004 ^ 1'b0 ;
  assign n19679 = n1028 | n19678 ;
  assign n19680 = ~n19677 & n19679 ;
  assign n19681 = n3873 & ~n19680 ;
  assign n19682 = n741 | n4547 ;
  assign n19683 = n6472 & ~n19682 ;
  assign n19684 = n13803 ^ n5676 ^ 1'b0 ;
  assign n19685 = n13900 ^ n2580 ^ 1'b0 ;
  assign n19686 = ~n19684 & n19685 ;
  assign n19687 = n7110 ^ n5176 ^ 1'b0 ;
  assign n19688 = n14957 | n19687 ;
  assign n19689 = n3556 ^ n3021 ^ 1'b0 ;
  assign n19690 = ~n755 & n19689 ;
  assign n19691 = ~n19688 & n19690 ;
  assign n19692 = n821 & n12674 ;
  assign n19693 = ~n3708 & n5228 ;
  assign n19694 = ~n3654 & n15929 ;
  assign n19695 = ~n4408 & n6946 ;
  assign n19696 = n15213 & n19695 ;
  assign n19697 = ~n4430 & n10728 ;
  assign n19698 = n5181 & ~n5523 ;
  assign n19699 = n377 | n19698 ;
  assign n19700 = n19699 ^ n19494 ^ n1908 ;
  assign n19701 = n3795 & ~n9017 ;
  assign n19702 = ~n1689 & n19701 ;
  assign n19703 = n6828 | n15683 ;
  assign n19704 = n4781 & n18928 ;
  assign n19705 = n6323 ^ n5419 ^ 1'b0 ;
  assign n19706 = ~n9703 & n19705 ;
  assign n19707 = n4428 & ~n7612 ;
  assign n19708 = ~n19706 & n19707 ;
  assign n19709 = n6327 ^ n1527 ^ 1'b0 ;
  assign n19710 = n5687 & n13005 ;
  assign n19711 = ( n2075 & n19709 ) | ( n2075 & ~n19710 ) | ( n19709 & ~n19710 ) ;
  assign n19712 = n10722 ^ n3491 ^ 1'b0 ;
  assign n19713 = n13551 & ~n13917 ;
  assign n19714 = n8657 & ~n9984 ;
  assign n19715 = n13373 & n19714 ;
  assign n19716 = n2626 & n6069 ;
  assign n19717 = ~n336 & n19716 ;
  assign n19718 = n5807 | n9937 ;
  assign n19719 = ~n19717 & n19718 ;
  assign n19720 = n9462 & ~n15951 ;
  assign n19721 = n12043 & ~n18965 ;
  assign n19722 = n17350 & n19721 ;
  assign n19723 = n5183 | n16643 ;
  assign n19724 = n19723 ^ n8684 ^ 1'b0 ;
  assign n19725 = n2351 ^ n808 ^ 1'b0 ;
  assign n19726 = n3474 & n15629 ;
  assign n19727 = n11753 & n19726 ;
  assign n19728 = ~n6584 & n19727 ;
  assign n19729 = n4901 ^ n3858 ^ 1'b0 ;
  assign n19730 = ~n4561 & n19729 ;
  assign n19731 = ~x0 & n2053 ;
  assign n19732 = n19731 ^ n11962 ^ 1'b0 ;
  assign n19733 = n4337 & n19732 ;
  assign n19734 = ~n19730 & n19733 ;
  assign n19735 = n11981 ^ n3907 ^ 1'b0 ;
  assign n19736 = n10011 ^ n1975 ^ 1'b0 ;
  assign n19737 = ~n1213 & n1597 ;
  assign n19738 = n15163 & ~n16852 ;
  assign n19739 = ~n6893 & n19738 ;
  assign n19740 = ~n2189 & n9097 ;
  assign n19741 = n11084 ^ n4808 ^ 1'b0 ;
  assign n19742 = ~n15176 & n19741 ;
  assign n19743 = n13114 ^ n2067 ^ 1'b0 ;
  assign n19744 = ~n5770 & n19743 ;
  assign n19745 = n5109 | n19744 ;
  assign n19746 = ( ~n4893 & n7075 ) | ( ~n4893 & n19745 ) | ( n7075 & n19745 ) ;
  assign n19747 = n14434 & ~n19746 ;
  assign n19748 = n4630 & ~n8787 ;
  assign n19749 = n12391 & n19748 ;
  assign n19750 = ~n10627 & n16260 ;
  assign n19751 = ~n4998 & n19750 ;
  assign n19752 = n1851 & ~n4893 ;
  assign n19753 = n19752 ^ n3738 ^ 1'b0 ;
  assign n19754 = ( n1765 & ~n6407 ) | ( n1765 & n10511 ) | ( ~n6407 & n10511 ) ;
  assign n19755 = n12612 ^ n8797 ^ 1'b0 ;
  assign n19756 = n19754 & ~n19755 ;
  assign n19757 = ~n11957 & n17888 ;
  assign n19758 = n6049 ^ n1740 ^ 1'b0 ;
  assign n19759 = ( ~n5240 & n17120 ) | ( ~n5240 & n19758 ) | ( n17120 & n19758 ) ;
  assign n19760 = n7687 & n17555 ;
  assign n19761 = n19760 ^ n4305 ^ 1'b0 ;
  assign n19762 = n5774 & n17056 ;
  assign n19763 = n19762 ^ n12588 ^ 1'b0 ;
  assign n19764 = n14641 ^ n879 ^ 1'b0 ;
  assign n19765 = ~n994 & n19764 ;
  assign n19766 = n3601 ^ n3111 ^ 1'b0 ;
  assign n19767 = ~n456 & n5955 ;
  assign n19768 = n19766 & n19767 ;
  assign n19769 = n6503 | n12856 ;
  assign n19770 = ~n9345 & n15051 ;
  assign n19771 = n2340 & n19770 ;
  assign n19772 = n2382 & n8187 ;
  assign n19773 = n19772 ^ n7173 ^ 1'b0 ;
  assign n19774 = ~n4555 & n15410 ;
  assign n19775 = n19774 ^ n9942 ^ 1'b0 ;
  assign n19776 = n7858 ^ n145 ^ 1'b0 ;
  assign n19777 = n13981 ^ n6940 ^ 1'b0 ;
  assign n19778 = n19776 & ~n19777 ;
  assign n19779 = ~n476 & n11529 ;
  assign n19780 = n19779 ^ n5583 ^ 1'b0 ;
  assign n19781 = n3505 & ~n6534 ;
  assign n19782 = n19781 ^ n11664 ^ 1'b0 ;
  assign n19783 = n6989 & n19782 ;
  assign n19784 = n19783 ^ n4647 ^ 1'b0 ;
  assign n19785 = n3498 ^ n400 ^ 1'b0 ;
  assign n19786 = n556 & ~n19785 ;
  assign n19787 = n19786 ^ n1882 ^ 1'b0 ;
  assign n19788 = n10086 ^ n9898 ^ n7528 ;
  assign n19789 = n842 & n6457 ;
  assign n19790 = ~n19788 & n19789 ;
  assign n19791 = n6852 & n19790 ;
  assign n19792 = ( n973 & ~n8921 ) | ( n973 & n14995 ) | ( ~n8921 & n14995 ) ;
  assign n19793 = n19792 ^ n12208 ^ 1'b0 ;
  assign n19794 = n16438 & ~n19793 ;
  assign n19795 = n16456 ^ n7532 ^ 1'b0 ;
  assign n19796 = ~n2937 & n12161 ;
  assign n19797 = ~n1404 & n19796 ;
  assign n19798 = ~n18753 & n19797 ;
  assign n19799 = n12587 & ~n19798 ;
  assign n19800 = n9348 & n19799 ;
  assign n19801 = n6041 ^ n331 ^ 1'b0 ;
  assign n19802 = x86 | n2300 ;
  assign n19803 = n4036 & n19802 ;
  assign n19804 = ~n5022 & n19803 ;
  assign n19805 = ( ~n5823 & n19801 ) | ( ~n5823 & n19804 ) | ( n19801 & n19804 ) ;
  assign n19806 = n10323 | n19805 ;
  assign n19807 = ~n7329 & n9694 ;
  assign n19808 = n19807 ^ n2905 ^ 1'b0 ;
  assign n19809 = n10580 ^ n10075 ^ n9768 ;
  assign n19810 = n19809 ^ n8075 ^ 1'b0 ;
  assign n19811 = ~n19808 & n19810 ;
  assign n19812 = ~n5546 & n8097 ;
  assign n19813 = n19812 ^ n7143 ^ 1'b0 ;
  assign n19814 = n13663 & n19813 ;
  assign n19815 = n19812 ^ n5500 ^ n2102 ;
  assign n19816 = n1089 | n6348 ;
  assign n19817 = n19816 ^ x23 ^ 1'b0 ;
  assign n19818 = n2984 | n14460 ;
  assign n19819 = ( n1230 & ~n1439 ) | ( n1230 & n19818 ) | ( ~n1439 & n19818 ) ;
  assign n19820 = n9136 | n19819 ;
  assign n19821 = ~n13452 & n19820 ;
  assign n19822 = ~n19817 & n19821 ;
  assign n19823 = n2920 & n18256 ;
  assign n19824 = n19123 ^ n1392 ^ 1'b0 ;
  assign n19825 = ~n2936 & n3850 ;
  assign n19826 = ~n4467 & n19825 ;
  assign n19827 = ~n9604 & n19826 ;
  assign n19828 = n3505 | n19245 ;
  assign n19829 = n10472 ^ n4734 ^ 1'b0 ;
  assign n19830 = n4123 & ~n12602 ;
  assign n19831 = n19830 ^ n10823 ^ 1'b0 ;
  assign n19832 = n5605 | n9994 ;
  assign n19833 = n17547 | n19832 ;
  assign n19834 = n3887 & ~n15002 ;
  assign n19835 = n1275 & n19834 ;
  assign n19836 = n1552 & n3567 ;
  assign n19837 = n15431 & n19836 ;
  assign n19838 = n5995 & n10045 ;
  assign n19839 = ( ~n4793 & n6731 ) | ( ~n4793 & n19838 ) | ( n6731 & n19838 ) ;
  assign n19840 = n9060 & ~n13878 ;
  assign n19841 = n10695 ^ n2914 ^ 1'b0 ;
  assign n19842 = ~n1761 & n19841 ;
  assign n19843 = ~n903 & n19842 ;
  assign n19844 = n19843 ^ n1838 ^ 1'b0 ;
  assign n19845 = n7959 & n19844 ;
  assign n19846 = n9888 & ~n19845 ;
  assign n19847 = n4708 ^ n3799 ^ 1'b0 ;
  assign n19848 = n6167 & ~n19847 ;
  assign n19849 = n12000 & ~n16054 ;
  assign n19850 = n7609 ^ n5074 ^ 1'b0 ;
  assign n19851 = n9950 ^ n2525 ^ 1'b0 ;
  assign n19852 = ~n19850 & n19851 ;
  assign n19853 = ~n3348 & n10204 ;
  assign n19854 = n12962 & n19853 ;
  assign n19855 = n2312 | n8185 ;
  assign n19856 = n661 & n19855 ;
  assign n19857 = n8746 ^ n4555 ^ n814 ;
  assign n19858 = n278 | n13599 ;
  assign n19859 = n19858 ^ n3336 ^ 1'b0 ;
  assign n19860 = n3109 | n13919 ;
  assign n19861 = n11013 ^ n1897 ^ 1'b0 ;
  assign n19862 = n18623 & ~n19861 ;
  assign n19863 = ~n8809 & n19862 ;
  assign n19864 = n19860 & n19863 ;
  assign n19865 = n832 | n1150 ;
  assign n19866 = n15030 & ~n19865 ;
  assign n19867 = n16683 ^ n15491 ^ 1'b0 ;
  assign n19868 = n3693 & ~n3879 ;
  assign n19869 = n18343 & n19868 ;
  assign n19870 = n8810 | n19869 ;
  assign n19871 = n4555 & ~n15823 ;
  assign n19872 = n19871 ^ n12480 ^ 1'b0 ;
  assign n19873 = n2940 & ~n5214 ;
  assign n19874 = n19872 & n19873 ;
  assign n19875 = n19874 ^ n10019 ^ n6871 ;
  assign n19876 = n12508 ^ n511 ^ 1'b0 ;
  assign n19877 = ~n5351 & n16234 ;
  assign n19878 = n19877 ^ n19129 ^ 1'b0 ;
  assign n19879 = n13942 ^ n7380 ^ 1'b0 ;
  assign n19880 = n1697 & ~n16200 ;
  assign n19881 = n18468 & n19880 ;
  assign n19882 = n8353 & ~n10501 ;
  assign n19883 = n8723 ^ n588 ^ 1'b0 ;
  assign n19884 = n15488 & n19883 ;
  assign n19885 = n6399 & n19884 ;
  assign n19886 = n6821 ^ n1086 ^ 1'b0 ;
  assign n19887 = ( n5650 & ~n11839 ) | ( n5650 & n19886 ) | ( ~n11839 & n19886 ) ;
  assign n19888 = n17904 ^ n9845 ^ 1'b0 ;
  assign n19889 = n4261 & n6585 ;
  assign n19890 = n9000 & n19889 ;
  assign n19891 = n2127 ^ n208 ^ 1'b0 ;
  assign n19892 = ~n11187 & n19891 ;
  assign n19893 = n585 & ~n6105 ;
  assign n19894 = n12677 & n19893 ;
  assign n19895 = n3543 | n7210 ;
  assign n19896 = n19895 ^ n1479 ^ 1'b0 ;
  assign n19897 = n19896 ^ n13476 ^ 1'b0 ;
  assign n19898 = n5605 | n19897 ;
  assign n19899 = n17218 ^ n10530 ^ 1'b0 ;
  assign n19903 = n8240 & n18467 ;
  assign n19901 = n3824 ^ n1670 ^ 1'b0 ;
  assign n19900 = ~n506 & n2234 ;
  assign n19902 = n19901 ^ n19900 ^ 1'b0 ;
  assign n19904 = n19903 ^ n19902 ^ n11332 ;
  assign n19905 = n16057 & n19904 ;
  assign n19906 = n18351 ^ n5112 ^ 1'b0 ;
  assign n19907 = n13500 | n19906 ;
  assign n19908 = n9041 & ~n19907 ;
  assign n19909 = n16931 ^ n3895 ^ 1'b0 ;
  assign n19910 = n2740 ^ n2048 ^ 1'b0 ;
  assign n19911 = n15802 ^ n11146 ^ 1'b0 ;
  assign n19912 = n19910 & n19911 ;
  assign n19913 = n19912 ^ n12662 ^ n8996 ;
  assign n19914 = ~n2737 & n8423 ;
  assign n19915 = n19914 ^ n6292 ^ 1'b0 ;
  assign n19916 = n19751 | n19915 ;
  assign n19917 = n7942 & ~n19916 ;
  assign n19918 = n6839 ^ n3354 ^ 1'b0 ;
  assign n19919 = ~n19917 & n19918 ;
  assign n19920 = n6436 & n19875 ;
  assign n19921 = n6629 & n19920 ;
  assign n19922 = n1155 & n16762 ;
  assign n19923 = n9445 & n19922 ;
  assign n19924 = n4380 & n19923 ;
  assign n19926 = n11990 ^ n10417 ^ 1'b0 ;
  assign n19927 = n8679 | n19926 ;
  assign n19925 = n517 | n2235 ;
  assign n19928 = n19927 ^ n19925 ^ n11056 ;
  assign n19929 = ~n1038 & n5358 ;
  assign n19930 = ~n3205 & n19929 ;
  assign n19931 = n10547 & n19930 ;
  assign n19932 = n5726 | n16975 ;
  assign n19933 = n19932 ^ n3574 ^ 1'b0 ;
  assign n19934 = n4275 & ~n7920 ;
  assign n19935 = n2533 & n9245 ;
  assign n19936 = n19934 & n19935 ;
  assign n19937 = n2053 & n8282 ;
  assign n19938 = n19937 ^ n7637 ^ 1'b0 ;
  assign n19939 = n838 & ~n19938 ;
  assign n19940 = n13235 & ~n19939 ;
  assign n19941 = ~n19936 & n19940 ;
  assign n19942 = n19941 ^ n5086 ^ 1'b0 ;
  assign n19943 = ~n11123 & n15844 ;
  assign n19944 = n12670 ^ n10106 ^ 1'b0 ;
  assign n19945 = ~n881 & n7619 ;
  assign n19946 = n19945 ^ n9273 ^ 1'b0 ;
  assign n19947 = n16497 ^ n16374 ^ n10954 ;
  assign n19948 = n8429 & n16276 ;
  assign n19949 = n19948 ^ n11738 ^ 1'b0 ;
  assign n19950 = ~n17511 & n19949 ;
  assign n19951 = n5907 & n16267 ;
  assign n19952 = n19951 ^ x41 ^ 1'b0 ;
  assign n19953 = ~n6120 & n14456 ;
  assign n19954 = ~n8943 & n19953 ;
  assign n19955 = n7878 ^ n5279 ^ n5080 ;
  assign n19956 = n16668 & ~n19955 ;
  assign n19957 = n971 & ~n5324 ;
  assign n19958 = n19957 ^ n4362 ^ 1'b0 ;
  assign n19959 = n9394 | n19958 ;
  assign n19960 = ~n1015 & n11784 ;
  assign n19961 = n19959 & n19960 ;
  assign n19962 = ( n4467 & ~n15503 ) | ( n4467 & n19961 ) | ( ~n15503 & n19961 ) ;
  assign n19963 = ~n1138 & n7457 ;
  assign n19964 = n19963 ^ n5300 ^ 1'b0 ;
  assign n19965 = n3331 ^ n368 ^ 1'b0 ;
  assign n19966 = n5830 & n19965 ;
  assign n19967 = n8590 | n13346 ;
  assign n19968 = n14075 ^ n8287 ^ 1'b0 ;
  assign n19969 = n3202 | n6132 ;
  assign n19970 = n6132 & ~n19969 ;
  assign n19971 = n6529 ^ n2321 ^ 1'b0 ;
  assign n19972 = n16957 & ~n19971 ;
  assign n19973 = n19972 ^ n13732 ^ n10818 ;
  assign n19974 = ( n11863 & n19970 ) | ( n11863 & n19973 ) | ( n19970 & n19973 ) ;
  assign n19975 = n19380 & ~n19974 ;
  assign n19976 = n19975 ^ n6006 ^ 1'b0 ;
  assign n19977 = n2869 ^ n892 ^ 1'b0 ;
  assign n19978 = ~n16988 & n19977 ;
  assign n19979 = n10176 ^ n6817 ^ 1'b0 ;
  assign n19980 = n6376 & n9229 ;
  assign n19981 = n5102 ^ n562 ^ 1'b0 ;
  assign n19982 = n11190 ^ n1348 ^ n600 ;
  assign n19983 = n4578 & ~n14456 ;
  assign n19984 = ~n1483 & n19983 ;
  assign n19985 = n243 & n3331 ;
  assign n19986 = x116 & ~n8619 ;
  assign n19987 = ~n19985 & n19986 ;
  assign n19988 = n8931 ^ n5505 ^ n4327 ;
  assign n19989 = ~n14998 & n19988 ;
  assign n19990 = ~n10577 & n19989 ;
  assign n19991 = n4568 ^ n2525 ^ 1'b0 ;
  assign n19992 = n16105 ^ n9613 ^ n6472 ;
  assign n19993 = n19991 & n19992 ;
  assign n19994 = n19990 | n19993 ;
  assign n19995 = n351 | n4600 ;
  assign n19996 = n1572 ^ n1439 ^ 1'b0 ;
  assign n19997 = n9978 | n19996 ;
  assign n19998 = n19995 & ~n19997 ;
  assign n20007 = n3761 ^ n3524 ^ n3460 ;
  assign n19999 = n11110 & n15800 ;
  assign n20000 = n7141 ^ n2671 ^ 1'b0 ;
  assign n20001 = n5413 & n20000 ;
  assign n20002 = n6105 | n20001 ;
  assign n20003 = n667 & ~n20002 ;
  assign n20004 = n20003 ^ n1201 ^ 1'b0 ;
  assign n20005 = n19999 & ~n20004 ;
  assign n20006 = ~n3215 & n20005 ;
  assign n20008 = n20007 ^ n20006 ^ 1'b0 ;
  assign n20009 = n959 & ~n13962 ;
  assign n20010 = n2605 | n6277 ;
  assign n20011 = n5040 ^ n2837 ^ 1'b0 ;
  assign n20012 = n5608 | n13675 ;
  assign n20013 = n13475 | n20012 ;
  assign n20014 = n20013 ^ n14448 ^ n13790 ;
  assign n20015 = n4829 & ~n11910 ;
  assign n20016 = n8688 | n20015 ;
  assign n20017 = n20015 & ~n20016 ;
  assign n20018 = n3491 ^ n1159 ^ n854 ;
  assign n20019 = ~n3968 & n20018 ;
  assign n20020 = ~n20018 & n20019 ;
  assign n20021 = n10759 & n20020 ;
  assign n20022 = ~n12457 & n20021 ;
  assign n20023 = ~n20021 & n20022 ;
  assign n20024 = n1304 | n8314 ;
  assign n20025 = n20024 ^ n2026 ^ 1'b0 ;
  assign n20026 = ~n2701 & n20025 ;
  assign n20027 = ~n20025 & n20026 ;
  assign n20028 = n5593 & ~n20027 ;
  assign n20029 = ~n5593 & n20028 ;
  assign n20030 = n20029 ^ n10541 ^ n7876 ;
  assign n20031 = n8992 & ~n20030 ;
  assign n20032 = ~n20023 & n20031 ;
  assign n20033 = n20032 ^ n3304 ^ 1'b0 ;
  assign n20034 = ( n3716 & n20017 ) | ( n3716 & ~n20033 ) | ( n20017 & ~n20033 ) ;
  assign n20035 = n10632 ^ n2676 ^ 1'b0 ;
  assign n20036 = n15211 ^ n1701 ^ 1'b0 ;
  assign n20037 = n2723 & n4639 ;
  assign n20038 = n20036 & n20037 ;
  assign n20039 = n6623 ^ n297 ^ 1'b0 ;
  assign n20040 = n11324 & n20039 ;
  assign n20041 = ~n4273 & n20040 ;
  assign n20042 = n7936 & n11307 ;
  assign n20043 = n4344 & n15595 ;
  assign n20044 = n19129 ^ n2492 ^ 1'b0 ;
  assign n20045 = n1172 & ~n4212 ;
  assign n20046 = n20045 ^ n10344 ^ 1'b0 ;
  assign n20047 = n19807 | n20046 ;
  assign n20048 = n14049 ^ n10460 ^ 1'b0 ;
  assign n20049 = ~n15985 & n20048 ;
  assign n20050 = n9148 | n19518 ;
  assign n20051 = n20050 ^ n11615 ^ 1'b0 ;
  assign n20052 = n17316 ^ n6021 ^ 1'b0 ;
  assign n20053 = n4424 | n6675 ;
  assign n20054 = n20053 ^ n3851 ^ x1 ;
  assign n20055 = n3389 | n8561 ;
  assign n20056 = n20054 & ~n20055 ;
  assign n20057 = n10152 & n13580 ;
  assign n20058 = n2624 & ~n17122 ;
  assign n20059 = n20058 ^ n12215 ^ 1'b0 ;
  assign n20060 = n5219 ^ n3400 ^ 1'b0 ;
  assign n20061 = n4468 | n4924 ;
  assign n20062 = n14372 & ~n20061 ;
  assign n20063 = n12214 ^ n7145 ^ 1'b0 ;
  assign n20064 = n8332 ^ n1526 ^ 1'b0 ;
  assign n20065 = ( ~n3820 & n9971 ) | ( ~n3820 & n20064 ) | ( n9971 & n20064 ) ;
  assign n20066 = n7711 | n20065 ;
  assign n20067 = n7501 & n12880 ;
  assign n20068 = ~n5914 & n20067 ;
  assign n20069 = n1190 & n8226 ;
  assign n20070 = ~n10878 & n15257 ;
  assign n20071 = n1372 & n20070 ;
  assign n20072 = n11259 ^ n7578 ^ n3318 ;
  assign n20073 = n11449 | n20072 ;
  assign n20074 = n20073 ^ n6105 ^ 1'b0 ;
  assign n20075 = n14608 ^ n11620 ^ 1'b0 ;
  assign n20076 = ( n1319 & n4953 ) | ( n1319 & ~n20075 ) | ( n4953 & ~n20075 ) ;
  assign n20077 = n8840 ^ n6539 ^ 1'b0 ;
  assign n20078 = n7995 | n16535 ;
  assign n20079 = n10831 & ~n20078 ;
  assign n20080 = n16981 & ~n18373 ;
  assign n20081 = ~n2125 & n20080 ;
  assign n20082 = n8791 ^ n2928 ^ 1'b0 ;
  assign n20083 = n1541 | n3408 ;
  assign n20084 = n20083 ^ n1834 ^ 1'b0 ;
  assign n20085 = n2235 & ~n20084 ;
  assign n20086 = n20085 ^ n15942 ^ n14560 ;
  assign n20087 = n4099 ^ n2075 ^ 1'b0 ;
  assign n20088 = n5477 & ~n20087 ;
  assign n20089 = n20088 ^ n9763 ^ 1'b0 ;
  assign n20090 = n8656 | n14446 ;
  assign n20091 = ~n2559 & n20090 ;
  assign n20092 = n20091 ^ n9505 ^ 1'b0 ;
  assign n20093 = ~n16612 & n17900 ;
  assign n20094 = n8590 & ~n20093 ;
  assign n20095 = n1408 & ~n9621 ;
  assign n20096 = n9229 ^ n5283 ^ n4766 ;
  assign n20097 = n294 | n20096 ;
  assign n20098 = n1200 | n13680 ;
  assign n20099 = n15598 & n16376 ;
  assign n20100 = ( n801 & n1336 ) | ( n801 & ~n8062 ) | ( n1336 & ~n8062 ) ;
  assign n20101 = n20100 ^ n8819 ^ 1'b0 ;
  assign n20102 = n10311 | n20101 ;
  assign n20103 = n20102 ^ n8938 ^ n4528 ;
  assign n20104 = n20103 ^ n7226 ^ 1'b0 ;
  assign n20105 = n8651 | n20104 ;
  assign n20106 = n17859 ^ n1180 ^ 1'b0 ;
  assign n20107 = n10152 ^ n4605 ^ 1'b0 ;
  assign n20108 = n9837 & ~n20107 ;
  assign n20109 = n4174 & ~n4963 ;
  assign n20110 = ~n6999 & n9706 ;
  assign n20111 = ~n20109 & n20110 ;
  assign n20112 = n2170 ^ n496 ^ 1'b0 ;
  assign n20113 = n19143 | n20112 ;
  assign n20114 = n20113 ^ n8425 ^ 1'b0 ;
  assign n20115 = n632 & n7136 ;
  assign n20116 = ~n4215 & n20115 ;
  assign n20117 = n4387 & ~n20116 ;
  assign n20118 = n20117 ^ n4639 ^ 1'b0 ;
  assign n20119 = n444 | n20118 ;
  assign n20120 = n20119 ^ n19838 ^ 1'b0 ;
  assign n20121 = n13448 ^ n7030 ^ 1'b0 ;
  assign n20122 = n16476 ^ n4534 ^ 1'b0 ;
  assign n20123 = n5647 | n18341 ;
  assign n20124 = n5842 ^ n5360 ^ n3799 ;
  assign n20125 = n13487 | n20124 ;
  assign n20126 = n16230 ^ n13292 ^ 1'b0 ;
  assign n20127 = n10361 & ~n20126 ;
  assign n20128 = n3205 ^ n2390 ^ 1'b0 ;
  assign n20129 = n20128 ^ n2132 ^ n699 ;
  assign n20130 = n4536 | n14663 ;
  assign n20131 = n5518 | n20130 ;
  assign n20132 = n12935 & ~n20131 ;
  assign n20133 = n20132 ^ n8226 ^ 1'b0 ;
  assign n20134 = n20129 | n20133 ;
  assign n20135 = ( n18008 & n20127 ) | ( n18008 & n20134 ) | ( n20127 & n20134 ) ;
  assign n20136 = ~n10516 & n13521 ;
  assign n20137 = n6124 | n16150 ;
  assign n20138 = n11840 ^ n10858 ^ 1'b0 ;
  assign n20139 = n20137 & ~n20138 ;
  assign n20140 = n20139 ^ n4201 ^ x106 ;
  assign n20141 = n6801 & ~n8809 ;
  assign n20142 = n5751 ^ n5243 ^ n2333 ;
  assign n20143 = ( n19774 & n20141 ) | ( n19774 & ~n20142 ) | ( n20141 & ~n20142 ) ;
  assign n20144 = ~n7075 & n19392 ;
  assign n20145 = n20143 & n20144 ;
  assign n20146 = n7908 & n11308 ;
  assign n20147 = n2824 & n18817 ;
  assign n20148 = ~n2824 & n20147 ;
  assign n20149 = n20148 ^ n5453 ^ 1'b0 ;
  assign n20150 = ~n20146 & n20149 ;
  assign n20151 = n5550 & ~n5822 ;
  assign n20152 = n5822 & n20151 ;
  assign n20153 = n20150 & ~n20152 ;
  assign n20154 = ~n20150 & n20153 ;
  assign n20155 = n20154 ^ n3029 ^ 1'b0 ;
  assign n20156 = n17284 & n20155 ;
  assign n20157 = n6059 & n7258 ;
  assign n20158 = ( n1861 & n9085 ) | ( n1861 & ~n20157 ) | ( n9085 & ~n20157 ) ;
  assign n20159 = ~n852 & n985 ;
  assign n20160 = ~n767 & n20159 ;
  assign n20161 = n16162 | n20160 ;
  assign n20162 = n20158 & ~n20161 ;
  assign n20163 = n4757 ^ n973 ^ 1'b0 ;
  assign n20164 = n9172 ^ n6428 ^ 1'b0 ;
  assign n20165 = n4793 & n20164 ;
  assign n20166 = n3481 ^ n2510 ^ 1'b0 ;
  assign n20167 = n6212 & ~n20166 ;
  assign n20168 = ~n12780 & n15378 ;
  assign n20169 = ~n13758 & n15045 ;
  assign n20170 = n20169 ^ n16433 ^ 1'b0 ;
  assign n20172 = n904 ^ n480 ^ 1'b0 ;
  assign n20171 = n9978 ^ n1329 ^ 1'b0 ;
  assign n20173 = n20172 ^ n20171 ^ n12662 ;
  assign n20174 = n4090 & ~n19725 ;
  assign n20176 = n1031 & ~n2339 ;
  assign n20175 = n1578 | n5324 ;
  assign n20177 = n20176 ^ n20175 ^ 1'b0 ;
  assign n20179 = n2750 & ~n4065 ;
  assign n20178 = ( n1251 & n1651 ) | ( n1251 & n10529 ) | ( n1651 & n10529 ) ;
  assign n20180 = n20179 ^ n20178 ^ 1'b0 ;
  assign n20181 = n11717 | n20180 ;
  assign n20182 = n2232 & ~n13268 ;
  assign n20183 = n20182 ^ n13080 ^ 1'b0 ;
  assign n20184 = n20183 ^ n10408 ^ 1'b0 ;
  assign n20185 = n1211 | n18736 ;
  assign n20186 = n13976 ^ n11637 ^ 1'b0 ;
  assign n20187 = ( n3869 & n7558 ) | ( n3869 & ~n20186 ) | ( n7558 & ~n20186 ) ;
  assign n20188 = n12071 | n13329 ;
  assign n20189 = n20188 ^ n16308 ^ 1'b0 ;
  assign n20191 = n9343 ^ n5613 ^ 1'b0 ;
  assign n20192 = n17384 | n20191 ;
  assign n20193 = n20192 ^ n15148 ^ 1'b0 ;
  assign n20190 = n4304 & ~n19489 ;
  assign n20194 = n20193 ^ n20190 ^ 1'b0 ;
  assign n20196 = n4053 | n16181 ;
  assign n20195 = n13057 & n17768 ;
  assign n20197 = n20196 ^ n20195 ^ 1'b0 ;
  assign n20198 = n17214 ^ n2596 ^ 1'b0 ;
  assign n20199 = n10450 ^ n3395 ^ 1'b0 ;
  assign n20200 = n13981 ^ n5381 ^ 1'b0 ;
  assign n20201 = ~n6869 & n7677 ;
  assign n20202 = n16206 & ~n19118 ;
  assign n20203 = ~n15528 & n20202 ;
  assign n20204 = ~n14499 & n20203 ;
  assign n20205 = n14642 ^ n8803 ^ 1'b0 ;
  assign n20206 = ~n5336 & n18210 ;
  assign n20207 = n14296 | n16179 ;
  assign n20208 = n10284 | n20207 ;
  assign n20209 = n2832 ^ n157 ^ 1'b0 ;
  assign n20210 = n2222 & ~n20209 ;
  assign n20211 = n20210 ^ x86 ^ 1'b0 ;
  assign n20212 = n2882 & ~n20211 ;
  assign n20213 = ~n616 & n20212 ;
  assign n20214 = n15834 ^ n6232 ^ 1'b0 ;
  assign n20215 = n5557 & n7542 ;
  assign n20216 = n20215 ^ n2748 ^ 1'b0 ;
  assign n20217 = n1212 & n1359 ;
  assign n20218 = n20217 ^ n13043 ^ 1'b0 ;
  assign n20219 = n12537 | n20218 ;
  assign n20220 = n13340 ^ n9383 ^ n3963 ;
  assign n20221 = ( n5894 & n8855 ) | ( n5894 & ~n16728 ) | ( n8855 & ~n16728 ) ;
  assign n20222 = n6074 & ~n19557 ;
  assign n20223 = n16357 ^ n8319 ^ 1'b0 ;
  assign n20224 = n9924 | n16945 ;
  assign n20225 = n7263 ^ n6137 ^ 1'b0 ;
  assign n20226 = n9151 ^ n4766 ^ 1'b0 ;
  assign n20227 = n20225 & n20226 ;
  assign n20228 = n13223 | n20227 ;
  assign n20229 = ~n6440 & n8475 ;
  assign n20230 = n6440 & n20229 ;
  assign n20235 = n3424 & ~n3639 ;
  assign n20236 = ~n3424 & n20235 ;
  assign n20231 = n475 & ~n487 ;
  assign n20232 = n487 & n20231 ;
  assign n20233 = n1222 & ~n20232 ;
  assign n20234 = ~n1222 & n20233 ;
  assign n20237 = n20236 ^ n20234 ^ 1'b0 ;
  assign n20238 = n20230 | n20237 ;
  assign n20239 = n20230 & ~n20238 ;
  assign n20240 = n20239 ^ n14303 ^ 1'b0 ;
  assign n20241 = n18958 ^ n14091 ^ 1'b0 ;
  assign n20242 = ~n20240 & n20241 ;
  assign n20243 = ~n5497 & n12395 ;
  assign n20244 = n18386 ^ n2009 ^ 1'b0 ;
  assign n20245 = n9800 | n20244 ;
  assign n20246 = n5862 & n20245 ;
  assign n20247 = n16629 ^ n5711 ^ 1'b0 ;
  assign n20248 = n18271 ^ n17385 ^ 1'b0 ;
  assign n20249 = n19321 ^ n16172 ^ n3816 ;
  assign n20252 = n672 & n17566 ;
  assign n20250 = n6610 | n16113 ;
  assign n20251 = n16768 | n20250 ;
  assign n20253 = n20252 ^ n20251 ^ 1'b0 ;
  assign n20254 = n13082 ^ n4551 ^ 1'b0 ;
  assign n20255 = ~n1711 & n5066 ;
  assign n20256 = n20254 & n20255 ;
  assign n20257 = n1097 ^ n678 ^ 1'b0 ;
  assign n20258 = n20256 | n20257 ;
  assign n20259 = n1465 | n1991 ;
  assign n20260 = n10080 | n20259 ;
  assign n20261 = n20260 ^ n1821 ^ 1'b0 ;
  assign n20262 = n16158 & n20261 ;
  assign n20263 = n3787 | n5514 ;
  assign n20264 = x37 & ~n7353 ;
  assign n20265 = n9156 ^ n4811 ^ 1'b0 ;
  assign n20266 = n3860 & ~n20265 ;
  assign n20267 = n6864 | n9439 ;
  assign n20268 = n12902 & ~n20267 ;
  assign n20269 = n8005 ^ n6843 ^ n6484 ;
  assign n20270 = n901 & n7096 ;
  assign n20271 = n20270 ^ n8592 ^ 1'b0 ;
  assign n20272 = n20269 & ~n20271 ;
  assign n20273 = n16150 ^ n15804 ^ 1'b0 ;
  assign n20274 = n14599 ^ n11322 ^ 1'b0 ;
  assign n20275 = n13066 ^ n10952 ^ 1'b0 ;
  assign n20276 = n20274 | n20275 ;
  assign n20277 = n14913 & ~n18062 ;
  assign n20278 = n18079 | n20277 ;
  assign n20279 = n20278 ^ n4892 ^ 1'b0 ;
  assign n20280 = n18295 ^ n10664 ^ 1'b0 ;
  assign n20281 = ~n1275 & n20280 ;
  assign n20282 = n8274 & n20281 ;
  assign n20283 = ~n3789 & n20282 ;
  assign n20284 = n4183 | n18569 ;
  assign n20285 = n20284 ^ n19397 ^ 1'b0 ;
  assign n20286 = ~n4325 & n19430 ;
  assign n20287 = n20286 ^ n6613 ^ 1'b0 ;
  assign n20288 = n15197 ^ n6148 ^ 1'b0 ;
  assign n20289 = n20288 ^ n9918 ^ 1'b0 ;
  assign n20290 = n676 & n10242 ;
  assign n20291 = n16375 ^ n4355 ^ 1'b0 ;
  assign n20292 = n9899 ^ n826 ^ 1'b0 ;
  assign n20293 = n20292 ^ n11000 ^ 1'b0 ;
  assign n20294 = n20291 & n20293 ;
  assign n20295 = n20294 ^ n6935 ^ n1481 ;
  assign n20296 = n14505 ^ n6155 ^ n3850 ;
  assign n20297 = n8273 & ~n18411 ;
  assign n20298 = n17261 & n20297 ;
  assign n20299 = n11699 ^ n6187 ^ 1'b0 ;
  assign n20300 = n2113 | n3715 ;
  assign n20301 = n20300 ^ n1865 ^ 1'b0 ;
  assign n20302 = n2730 & n6932 ;
  assign n20303 = n20301 & ~n20302 ;
  assign n20306 = n10307 | n13878 ;
  assign n20304 = ~n5022 & n10201 ;
  assign n20305 = n5693 & ~n20304 ;
  assign n20307 = n20306 ^ n20305 ^ 1'b0 ;
  assign n20308 = n4255 & n5458 ;
  assign n20309 = n17790 ^ n11593 ^ 1'b0 ;
  assign n20310 = x116 & n11948 ;
  assign n20311 = ~n3294 & n20310 ;
  assign n20312 = n15020 & n20311 ;
  assign n20313 = n5492 ^ n4172 ^ n1532 ;
  assign n20314 = n8510 ^ n4452 ^ 1'b0 ;
  assign n20315 = n8363 & n20314 ;
  assign n20316 = n13137 ^ n13114 ^ 1'b0 ;
  assign n20317 = n5849 & n20316 ;
  assign n20318 = ~n15557 & n20317 ;
  assign n20319 = n7990 & n20318 ;
  assign n20320 = ~n20315 & n20319 ;
  assign n20323 = n15406 ^ x3 ^ 1'b0 ;
  assign n20324 = n3313 & n20323 ;
  assign n20321 = n2102 & ~n9141 ;
  assign n20322 = n20321 ^ n7203 ^ 1'b0 ;
  assign n20325 = n20324 ^ n20322 ^ 1'b0 ;
  assign n20326 = n4800 ^ n4028 ^ 1'b0 ;
  assign n20327 = n7866 & n19078 ;
  assign n20328 = ( n3869 & ~n8048 ) | ( n3869 & n20327 ) | ( ~n8048 & n20327 ) ;
  assign n20329 = n542 | n1645 ;
  assign n20330 = n6391 & ~n20329 ;
  assign n20331 = n8109 ^ n3352 ^ 1'b0 ;
  assign n20332 = n20330 | n20331 ;
  assign n20333 = n20332 ^ n12736 ^ 1'b0 ;
  assign n20334 = n1406 & ~n6342 ;
  assign n20335 = ~n10431 & n20247 ;
  assign n20336 = ~n20334 & n20335 ;
  assign n20337 = n3128 & n3190 ;
  assign n20338 = n14769 & n20337 ;
  assign n20339 = n6693 & ~n20338 ;
  assign n20340 = ~n3539 & n20339 ;
  assign n20341 = n9732 ^ n8571 ^ 1'b0 ;
  assign n20342 = n20341 ^ n12792 ^ 1'b0 ;
  assign n20343 = n2938 ^ n1903 ^ 1'b0 ;
  assign n20346 = n5556 | n6563 ;
  assign n20347 = n6594 & ~n20346 ;
  assign n20344 = n815 | n1401 ;
  assign n20345 = n16787 & ~n20344 ;
  assign n20348 = n20347 ^ n20345 ^ 1'b0 ;
  assign n20349 = ~n3276 & n10897 ;
  assign n20350 = n1283 & n20349 ;
  assign n20353 = n10540 ^ n1733 ^ n993 ;
  assign n20354 = x39 | n20353 ;
  assign n20351 = n10619 ^ n1481 ^ 1'b0 ;
  assign n20352 = n13682 | n20351 ;
  assign n20355 = n20354 ^ n20352 ^ 1'b0 ;
  assign n20356 = n1830 ^ x13 ^ 1'b0 ;
  assign n20357 = n7087 & ~n18111 ;
  assign n20358 = n2030 | n5466 ;
  assign n20359 = n20357 & ~n20358 ;
  assign n20360 = n20359 ^ n3546 ^ 1'b0 ;
  assign n20361 = n20356 | n20360 ;
  assign n20367 = ~n2529 & n2638 ;
  assign n20362 = n4992 ^ n628 ^ 1'b0 ;
  assign n20363 = n20362 ^ n18764 ^ 1'b0 ;
  assign n20364 = ~n5841 & n20363 ;
  assign n20365 = ~n13167 & n20364 ;
  assign n20366 = n7213 & n20365 ;
  assign n20368 = n20367 ^ n20366 ^ 1'b0 ;
  assign n20369 = n203 | n14663 ;
  assign n20370 = n4161 ^ n4037 ^ 1'b0 ;
  assign n20371 = n5357 | n20370 ;
  assign n20372 = n16185 ^ n2637 ^ 1'b0 ;
  assign n20373 = x104 & n20372 ;
  assign n20374 = n6520 ^ n1735 ^ 1'b0 ;
  assign n20375 = n20373 & ~n20374 ;
  assign n20376 = n421 & n12202 ;
  assign n20377 = n14589 ^ n13002 ^ 1'b0 ;
  assign n20378 = n12148 & n15013 ;
  assign n20379 = n9829 & ~n20378 ;
  assign n20380 = n11484 & n20379 ;
  assign n20381 = ( n8203 & n10512 ) | ( n8203 & ~n10993 ) | ( n10512 & ~n10993 ) ;
  assign n20382 = n20381 ^ n15250 ^ 1'b0 ;
  assign n20383 = n13775 ^ n11235 ^ n6827 ;
  assign n20384 = n20383 ^ n4382 ^ 1'b0 ;
  assign n20385 = n9616 | n17930 ;
  assign n20386 = n14441 ^ n344 ^ 1'b0 ;
  assign n20387 = ~n2153 & n20386 ;
  assign n20388 = ~n1219 & n3846 ;
  assign n20389 = n18403 & ~n20388 ;
  assign n20390 = n5910 | n15203 ;
  assign n20391 = n8257 ^ n4134 ^ n708 ;
  assign n20392 = n7992 ^ n1578 ^ 1'b0 ;
  assign n20393 = n565 | n20392 ;
  assign n20394 = n20393 ^ n11600 ^ 1'b0 ;
  assign n20395 = n8096 ^ n4632 ^ 1'b0 ;
  assign n20396 = n574 & ~n8897 ;
  assign n20397 = ~n15197 & n20396 ;
  assign n20398 = n14493 & n20397 ;
  assign n20399 = ~n12537 & n18954 ;
  assign n20400 = n6942 & n20399 ;
  assign n20401 = n246 & ~n20175 ;
  assign n20402 = n7164 | n12023 ;
  assign n20404 = ( n400 & n1133 ) | ( n400 & n2778 ) | ( n1133 & n2778 ) ;
  assign n20403 = n2742 & ~n2802 ;
  assign n20405 = n20404 ^ n20403 ^ 1'b0 ;
  assign n20406 = n15566 ^ n14242 ^ 1'b0 ;
  assign n20407 = ~n5754 & n20406 ;
  assign n20408 = n11519 ^ n6940 ^ 1'b0 ;
  assign n20409 = n4007 | n20408 ;
  assign n20410 = n18554 ^ n14166 ^ 1'b0 ;
  assign n20411 = n5707 ^ n3251 ^ 1'b0 ;
  assign n20412 = ~n20410 & n20411 ;
  assign n20413 = n12040 ^ n695 ^ 1'b0 ;
  assign n20414 = n8756 & ~n10124 ;
  assign n20415 = n20414 ^ n17532 ^ 1'b0 ;
  assign n20416 = ~n16304 & n16479 ;
  assign n20417 = n20416 ^ n8106 ^ 1'b0 ;
  assign n20418 = ~n3314 & n20417 ;
  assign n20419 = ~n20415 & n20418 ;
  assign n20420 = n20413 | n20419 ;
  assign n20421 = n20420 ^ n14495 ^ 1'b0 ;
  assign n20422 = ( n231 & n1963 ) | ( n231 & n2462 ) | ( n1963 & n2462 ) ;
  assign n20423 = ~n2928 & n10732 ;
  assign n20424 = n556 & n19552 ;
  assign n20425 = n20423 & n20424 ;
  assign n20426 = n13315 ^ n5524 ^ 1'b0 ;
  assign n20427 = n276 & n12549 ;
  assign n20428 = n10012 & ~n20427 ;
  assign n20429 = n16206 & n17425 ;
  assign n20430 = n15378 ^ n8282 ^ 1'b0 ;
  assign n20431 = n3214 | n4510 ;
  assign n20432 = n20431 ^ x94 ^ 1'b0 ;
  assign n20433 = n20430 & n20432 ;
  assign n20434 = n6322 & n12219 ;
  assign n20435 = n5863 & n5967 ;
  assign n20436 = n20435 ^ n12446 ^ n1606 ;
  assign n20437 = n12853 ^ n3671 ^ n3032 ;
  assign n20438 = ( ~n2816 & n5131 ) | ( ~n2816 & n20437 ) | ( n5131 & n20437 ) ;
  assign n20439 = n3550 & ~n10357 ;
  assign n20440 = ~n9749 & n20439 ;
  assign n20441 = n14832 & ~n20440 ;
  assign n20442 = n20441 ^ n4299 ^ 1'b0 ;
  assign n20443 = ~n6623 & n20442 ;
  assign n20444 = n1109 | n10652 ;
  assign n20445 = n7760 | n8236 ;
  assign n20446 = n10278 ^ x52 ^ 1'b0 ;
  assign n20447 = n6802 | n20446 ;
  assign n20448 = n9199 & n20447 ;
  assign n20449 = ( ~n6278 & n10357 ) | ( ~n6278 & n12692 ) | ( n10357 & n12692 ) ;
  assign n20450 = n20449 ^ n12248 ^ 1'b0 ;
  assign n20451 = n11324 & n20450 ;
  assign n20452 = n13636 | n20451 ;
  assign n20453 = n8957 ^ n6415 ^ 1'b0 ;
  assign n20454 = n15854 & n20453 ;
  assign n20455 = n19805 ^ n4048 ^ 1'b0 ;
  assign n20456 = n15564 & ~n16037 ;
  assign n20458 = n2235 ^ n1068 ^ 1'b0 ;
  assign n20459 = n20458 ^ n8306 ^ 1'b0 ;
  assign n20460 = ~n677 & n20459 ;
  assign n20457 = n15949 ^ n11040 ^ n3879 ;
  assign n20461 = n20460 ^ n20457 ^ n5457 ;
  assign n20462 = n18854 ^ n14267 ^ 1'b0 ;
  assign n20463 = n5634 | n12897 ;
  assign n20464 = n5577 ^ n3855 ^ 1'b0 ;
  assign n20465 = n13031 & ~n20464 ;
  assign n20466 = n20465 ^ n9154 ^ 1'b0 ;
  assign n20467 = n404 & ~n20466 ;
  assign n20468 = n1632 | n17264 ;
  assign n20469 = n20468 ^ n6720 ^ 1'b0 ;
  assign n20470 = n4647 ^ n400 ^ 1'b0 ;
  assign n20471 = ~n3266 & n20470 ;
  assign n20472 = n10571 | n12436 ;
  assign n20473 = n18399 ^ n17033 ^ n16678 ;
  assign n20474 = n16431 ^ n1102 ^ 1'b0 ;
  assign n20475 = n10485 | n20474 ;
  assign n20476 = n9055 ^ n4150 ^ 1'b0 ;
  assign n20477 = n15164 ^ n8830 ^ n2402 ;
  assign n20478 = n7190 ^ n2364 ^ 1'b0 ;
  assign n20479 = ~n18670 & n20478 ;
  assign n20480 = ~n2021 & n5584 ;
  assign n20481 = n20480 ^ n6574 ^ 1'b0 ;
  assign n20482 = n5692 & n9462 ;
  assign n20483 = n8768 & n10791 ;
  assign n20484 = n20483 ^ n13084 ^ 1'b0 ;
  assign n20485 = n8056 & n9959 ;
  assign n20486 = n20485 ^ n5495 ^ 1'b0 ;
  assign n20487 = n3528 | n4897 ;
  assign n20488 = ~n3090 & n20487 ;
  assign n20489 = ~n6289 & n6753 ;
  assign n20490 = ~n6959 & n20489 ;
  assign n20491 = n10479 | n20490 ;
  assign n20492 = n1244 ^ x17 ^ 1'b0 ;
  assign n20493 = n4827 & n6594 ;
  assign n20494 = n20493 ^ n2899 ^ 1'b0 ;
  assign n20495 = n6103 & ~n8741 ;
  assign n20496 = n17353 & n20495 ;
  assign n20497 = n20496 ^ n19632 ^ 1'b0 ;
  assign n20498 = n20494 & ~n20497 ;
  assign n20499 = n12635 & ~n15290 ;
  assign n20500 = n20499 ^ n19855 ^ 1'b0 ;
  assign n20501 = n15878 ^ n4804 ^ 1'b0 ;
  assign n20502 = n4995 & n14095 ;
  assign n20503 = n20502 ^ n9850 ^ 1'b0 ;
  assign n20504 = n2562 & ~n8331 ;
  assign n20505 = ~n12552 & n20504 ;
  assign n20506 = n20505 ^ n9962 ^ 1'b0 ;
  assign n20507 = n12871 & ~n16584 ;
  assign n20508 = n1901 & ~n10512 ;
  assign n20510 = n6821 ^ n4438 ^ n2170 ;
  assign n20509 = n10851 & n17552 ;
  assign n20511 = n20510 ^ n20509 ^ 1'b0 ;
  assign n20512 = n20004 | n20511 ;
  assign n20513 = n6398 ^ x117 ^ 1'b0 ;
  assign n20514 = n13992 | n20513 ;
  assign n20515 = ~n3613 & n9071 ;
  assign n20516 = n12421 ^ n6271 ^ 1'b0 ;
  assign n20517 = ~n5561 & n9003 ;
  assign n20518 = n1661 | n10969 ;
  assign n20519 = n10985 & ~n13755 ;
  assign n20520 = n7198 | n14592 ;
  assign n20521 = ~n7377 & n10475 ;
  assign n20522 = n4712 & n20521 ;
  assign n20523 = ( n4581 & ~n20520 ) | ( n4581 & n20522 ) | ( ~n20520 & n20522 ) ;
  assign n20524 = n7234 ^ n5678 ^ 1'b0 ;
  assign n20525 = ~n7674 & n20524 ;
  assign n20526 = ( n1209 & ~n8315 ) | ( n1209 & n20525 ) | ( ~n8315 & n20525 ) ;
  assign n20527 = n3894 ^ n1377 ^ 1'b0 ;
  assign n20528 = x69 & n20527 ;
  assign n20529 = n18383 ^ n10608 ^ 1'b0 ;
  assign n20530 = n20528 & ~n20529 ;
  assign n20531 = ~n10064 & n12721 ;
  assign n20532 = n20531 ^ n709 ^ 1'b0 ;
  assign n20533 = ~n208 & n15218 ;
  assign n20534 = n20533 ^ n2050 ^ 1'b0 ;
  assign n20535 = ~n9763 & n18424 ;
  assign n20536 = n3800 ^ n2121 ^ 1'b0 ;
  assign n20537 = ~n909 & n9350 ;
  assign n20538 = n16979 | n20537 ;
  assign n20539 = n2501 & n13955 ;
  assign n20540 = n20539 ^ n15402 ^ 1'b0 ;
  assign n20541 = n20540 ^ n13315 ^ n1831 ;
  assign n20542 = n419 | n4613 ;
  assign n20543 = n1399 ^ x50 ^ 1'b0 ;
  assign n20544 = n308 & n20543 ;
  assign n20545 = n7636 & ~n20544 ;
  assign n20546 = ~n14795 & n15986 ;
  assign n20547 = n20546 ^ n8477 ^ 1'b0 ;
  assign n20548 = n14271 ^ n6606 ^ 1'b0 ;
  assign n20549 = n12705 | n15176 ;
  assign n20550 = n20549 ^ n4010 ^ 1'b0 ;
  assign n20551 = n20550 ^ n2562 ^ n2131 ;
  assign n20552 = ~n2462 & n18136 ;
  assign n20555 = ~n1143 & n1295 ;
  assign n20556 = n580 & ~n9460 ;
  assign n20557 = n20555 & n20556 ;
  assign n20554 = n3414 & ~n9435 ;
  assign n20558 = n20557 ^ n20554 ^ 1'b0 ;
  assign n20553 = n1899 & ~n7036 ;
  assign n20559 = n20558 ^ n20553 ^ 1'b0 ;
  assign n20560 = n1448 | n3467 ;
  assign n20561 = n11767 | n20560 ;
  assign n20562 = n15749 & ~n17576 ;
  assign n20563 = n10236 & n20562 ;
  assign n20564 = n11713 ^ n1659 ^ 1'b0 ;
  assign n20565 = ~n9676 & n20564 ;
  assign n20566 = n3974 & ~n11568 ;
  assign n20567 = n20566 ^ n578 ^ 1'b0 ;
  assign n20568 = ~n4287 & n20567 ;
  assign n20569 = ( n11550 & n13128 ) | ( n11550 & ~n17136 ) | ( n13128 & ~n17136 ) ;
  assign n20573 = ~n18736 & n20388 ;
  assign n20574 = ~n8816 & n20573 ;
  assign n20570 = n4569 ^ x39 ^ 1'b0 ;
  assign n20571 = n5290 | n20570 ;
  assign n20572 = n1254 & ~n20571 ;
  assign n20575 = n20574 ^ n20572 ^ 1'b0 ;
  assign n20576 = n9125 ^ n2170 ^ 1'b0 ;
  assign n20577 = n744 & n20576 ;
  assign n20578 = n4893 ^ n2136 ^ 1'b0 ;
  assign n20579 = n9288 | n20578 ;
  assign n20580 = ~n4884 & n19988 ;
  assign n20581 = ~n3869 & n6599 ;
  assign n20582 = ( n7800 & ~n17146 ) | ( n7800 & n20581 ) | ( ~n17146 & n20581 ) ;
  assign n20583 = n2783 | n6122 ;
  assign n20584 = n11324 | n20583 ;
  assign n20585 = n1296 | n7324 ;
  assign n20586 = n555 | n7787 ;
  assign n20587 = n464 & ~n20586 ;
  assign n20588 = n20585 | n20587 ;
  assign n20589 = n3020 ^ n1863 ^ 1'b0 ;
  assign n20590 = n3528 & n20589 ;
  assign n20592 = n11902 ^ n722 ^ 1'b0 ;
  assign n20591 = n9154 ^ n4102 ^ 1'b0 ;
  assign n20593 = n20592 ^ n20591 ^ n7110 ;
  assign n20594 = n18064 ^ n15454 ^ 1'b0 ;
  assign n20595 = n13994 ^ n2953 ^ 1'b0 ;
  assign n20596 = n20595 ^ n3937 ^ 1'b0 ;
  assign n20597 = n9265 & n9297 ;
  assign n20598 = n2354 & n20597 ;
  assign n20599 = ~n7744 & n19891 ;
  assign n20600 = n20599 ^ n7368 ^ 1'b0 ;
  assign n20601 = n8399 & n20600 ;
  assign n20602 = ( n203 & n3370 ) | ( n203 & ~n11660 ) | ( n3370 & ~n11660 ) ;
  assign n20603 = ~n3114 & n20602 ;
  assign n20604 = n760 | n4705 ;
  assign n20605 = n20604 ^ n4171 ^ 1'b0 ;
  assign n20606 = n11018 & n20605 ;
  assign n20607 = n14889 | n17105 ;
  assign n20608 = n20607 ^ n16190 ^ 1'b0 ;
  assign n20609 = n14713 ^ x102 ^ 1'b0 ;
  assign n20610 = n5561 | n20609 ;
  assign n20611 = n20610 ^ n423 ^ 1'b0 ;
  assign n20612 = n506 & ~n12882 ;
  assign n20613 = n148 & n20612 ;
  assign n20614 = n16793 ^ n15045 ^ 1'b0 ;
  assign n20615 = n10382 ^ n7221 ^ 1'b0 ;
  assign n20616 = ~n5219 & n10772 ;
  assign n20617 = n20616 ^ n16723 ^ 1'b0 ;
  assign n20618 = ( n1491 & ~n3381 ) | ( n1491 & n20617 ) | ( ~n3381 & n20617 ) ;
  assign n20619 = n8309 | n8575 ;
  assign n20620 = n18988 ^ n10496 ^ 1'b0 ;
  assign n20621 = n5519 ^ n1084 ^ 1'b0 ;
  assign n20622 = n3399 | n20621 ;
  assign n20623 = n14596 & ~n20622 ;
  assign n20624 = ~n5450 & n16264 ;
  assign n20625 = n1758 | n7624 ;
  assign n20626 = n10100 & n20625 ;
  assign n20627 = n1190 | n19263 ;
  assign n20628 = n13924 & ~n20302 ;
  assign n20629 = ( n4502 & n4556 ) | ( n4502 & ~n13871 ) | ( n4556 & ~n13871 ) ;
  assign n20630 = ~n1324 & n18995 ;
  assign n20631 = n10647 ^ n5193 ^ 1'b0 ;
  assign n20632 = ~n10402 & n10673 ;
  assign n20633 = n5374 & n20632 ;
  assign n20634 = n14456 ^ n2585 ^ 1'b0 ;
  assign n20635 = n941 & n8722 ;
  assign n20636 = n10107 ^ n9524 ^ 1'b0 ;
  assign n20637 = n5989 ^ n3844 ^ 1'b0 ;
  assign n20638 = n3300 | n20637 ;
  assign n20639 = n20638 ^ n15142 ^ 1'b0 ;
  assign n20640 = n4613 & n20639 ;
  assign n20641 = n10331 | n10535 ;
  assign n20642 = n3758 & n18513 ;
  assign n20643 = n20642 ^ n9802 ^ 1'b0 ;
  assign n20644 = n9327 ^ n8466 ^ 1'b0 ;
  assign n20645 = n9604 | n20644 ;
  assign n20646 = n4875 | n12438 ;
  assign n20647 = n7319 & ~n20646 ;
  assign n20648 = n14048 ^ n9495 ^ 1'b0 ;
  assign n20650 = n2243 | n19872 ;
  assign n20649 = n8224 | n17557 ;
  assign n20651 = n20650 ^ n20649 ^ n9897 ;
  assign n20652 = n6201 ^ n2585 ^ 1'b0 ;
  assign n20653 = n3215 | n20652 ;
  assign n20654 = n20653 ^ n4831 ^ 1'b0 ;
  assign n20655 = ( n1068 & ~n4323 ) | ( n1068 & n5011 ) | ( ~n4323 & n5011 ) ;
  assign n20656 = ( n9796 & n16788 ) | ( n9796 & ~n20655 ) | ( n16788 & ~n20655 ) ;
  assign n20658 = n3564 ^ n3372 ^ 1'b0 ;
  assign n20659 = n10904 | n20658 ;
  assign n20657 = n7953 ^ n5951 ^ 1'b0 ;
  assign n20660 = n20659 ^ n20657 ^ 1'b0 ;
  assign n20661 = ~n7102 & n20660 ;
  assign n20662 = n20656 & n20661 ;
  assign n20663 = n18190 ^ n15010 ^ 1'b0 ;
  assign n20664 = n2948 | n20663 ;
  assign n20665 = n3870 | n6671 ;
  assign n20666 = n20665 ^ n10770 ^ 1'b0 ;
  assign n20667 = n17024 ^ n15399 ^ 1'b0 ;
  assign n20668 = n20666 & ~n20667 ;
  assign n20669 = n3041 | n16287 ;
  assign n20670 = n3246 | n20669 ;
  assign n20671 = ( n4987 & n6050 ) | ( n4987 & ~n20670 ) | ( n6050 & ~n20670 ) ;
  assign n20672 = n2987 | n4307 ;
  assign n20673 = n20672 ^ n437 ^ 1'b0 ;
  assign n20674 = n12302 ^ n942 ^ 1'b0 ;
  assign n20675 = n7998 & ~n20674 ;
  assign n20676 = n3988 | n5129 ;
  assign n20677 = n10161 | n20676 ;
  assign n20678 = n7602 & n20546 ;
  assign n20679 = ~n2135 & n12520 ;
  assign n20680 = n11632 & n20679 ;
  assign n20681 = n11365 & ~n20680 ;
  assign n20682 = n20681 ^ n6432 ^ 1'b0 ;
  assign n20683 = n17566 ^ n4694 ^ 1'b0 ;
  assign n20684 = n11215 | n13439 ;
  assign n20685 = n1285 & n20684 ;
  assign n20686 = n20685 ^ n9242 ^ 1'b0 ;
  assign n20687 = n1585 | n15499 ;
  assign n20688 = n20687 ^ n17082 ^ 1'b0 ;
  assign n20689 = n16940 & n20688 ;
  assign n20690 = n182 & n16618 ;
  assign n20691 = n20690 ^ n4927 ^ 1'b0 ;
  assign n20692 = n12946 ^ n567 ^ 1'b0 ;
  assign n20693 = n2146 & n8045 ;
  assign n20694 = n808 & ~n9645 ;
  assign n20695 = n20694 ^ n2752 ^ 1'b0 ;
  assign n20696 = n18185 ^ n11635 ^ x67 ;
  assign n20697 = x46 & ~n4522 ;
  assign n20698 = n2648 | n18168 ;
  assign n20699 = n2170 & n20698 ;
  assign n20700 = ~n1062 & n8710 ;
  assign n20701 = n20700 ^ n10061 ^ 1'b0 ;
  assign n20702 = n2622 | n7245 ;
  assign n20703 = n1361 | n6093 ;
  assign n20704 = n920 & ~n20703 ;
  assign n20705 = n9598 & n20704 ;
  assign n20706 = n20702 & n20705 ;
  assign n20707 = ~n336 & n2782 ;
  assign n20708 = x89 & ~n5810 ;
  assign n20709 = n20708 ^ n8058 ^ n6801 ;
  assign n20710 = n1271 & n5383 ;
  assign n20711 = ~n6448 & n8520 ;
  assign n20712 = n20711 ^ n6451 ^ 1'b0 ;
  assign n20713 = ~n12170 & n20712 ;
  assign n20714 = n20713 ^ n13099 ^ 1'b0 ;
  assign n20715 = n20714 ^ n7344 ^ 1'b0 ;
  assign n20716 = n19129 ^ n1599 ^ 1'b0 ;
  assign n20717 = ~n12129 & n20716 ;
  assign n20718 = n9585 & n15195 ;
  assign n20719 = n12670 & ~n15898 ;
  assign n20720 = n7297 & n11709 ;
  assign n20721 = n5191 ^ n2931 ^ 1'b0 ;
  assign n20722 = n10615 | n20721 ;
  assign n20723 = n11837 ^ n5942 ^ 1'b0 ;
  assign n20724 = ~n3269 & n18324 ;
  assign n20725 = n13042 & ~n13048 ;
  assign n20726 = n18869 ^ n13345 ^ n4542 ;
  assign n20727 = ~n16304 & n20726 ;
  assign n20728 = ~n5092 & n6137 ;
  assign n20729 = n20727 & ~n20728 ;
  assign n20730 = ~n1367 & n7577 ;
  assign n20731 = n6370 & ~n14629 ;
  assign n20732 = n16712 & n20731 ;
  assign n20733 = n9255 | n20732 ;
  assign n20734 = n20730 | n20733 ;
  assign n20735 = ~n2321 & n6322 ;
  assign n20736 = n20735 ^ n9273 ^ n4586 ;
  assign n20737 = n14394 ^ n11743 ^ n8342 ;
  assign n20738 = n2645 | n2931 ;
  assign n20739 = n8774 | n9121 ;
  assign n20740 = n10336 ^ n9880 ^ 1'b0 ;
  assign n20741 = n11410 | n20740 ;
  assign n20742 = ( ~n2113 & n7828 ) | ( ~n2113 & n12746 ) | ( n7828 & n12746 ) ;
  assign n20743 = n20742 ^ n11010 ^ n866 ;
  assign n20744 = n3339 & ~n20743 ;
  assign n20745 = n20744 ^ n16483 ^ 1'b0 ;
  assign n20746 = n756 ^ x47 ^ 1'b0 ;
  assign n20747 = n20440 ^ n11826 ^ 1'b0 ;
  assign n20748 = n20746 | n20747 ;
  assign n20749 = n3924 | n9319 ;
  assign n20750 = n1817 | n14854 ;
  assign n20751 = n20750 ^ n3261 ^ 1'b0 ;
  assign n20752 = n11438 & ~n20211 ;
  assign n20753 = n20752 ^ n9191 ^ 1'b0 ;
  assign n20754 = n14573 ^ n9412 ^ 1'b0 ;
  assign n20755 = ~n2370 & n20754 ;
  assign n20756 = n494 & n20755 ;
  assign n20757 = n20756 ^ n11034 ^ 1'b0 ;
  assign n20758 = ( n1761 & ~n7382 ) | ( n1761 & n20364 ) | ( ~n7382 & n20364 ) ;
  assign n20759 = n1945 & n20758 ;
  assign n20760 = ( n6397 & n7881 ) | ( n6397 & n12591 ) | ( n7881 & n12591 ) ;
  assign n20761 = n20760 ^ n4030 ^ 1'b0 ;
  assign n20762 = ~n8344 & n20761 ;
  assign n20763 = ~n4516 & n20191 ;
  assign n20764 = n4745 & n12308 ;
  assign n20765 = n20764 ^ n3877 ^ n1939 ;
  assign n20766 = n16559 ^ n5500 ^ 1'b0 ;
  assign n20768 = ~n4175 & n18518 ;
  assign n20767 = n6093 & ~n11990 ;
  assign n20769 = n20768 ^ n20767 ^ 1'b0 ;
  assign n20770 = n20769 ^ n7594 ^ 1'b0 ;
  assign n20771 = n6290 & n20770 ;
  assign n20773 = ~n4775 & n10736 ;
  assign n20774 = n13593 & n20773 ;
  assign n20772 = n6803 ^ n5243 ^ 1'b0 ;
  assign n20775 = n20774 ^ n20772 ^ 1'b0 ;
  assign n20776 = ~n2085 & n9163 ;
  assign n20777 = n20776 ^ n11910 ^ 1'b0 ;
  assign n20778 = n8954 ^ n3547 ^ 1'b0 ;
  assign n20779 = n6768 ^ n3629 ^ 1'b0 ;
  assign n20780 = n632 & ~n20779 ;
  assign n20781 = n20780 ^ n20362 ^ n11632 ;
  assign n20782 = n3359 & n7998 ;
  assign n20783 = n20782 ^ n19345 ^ 1'b0 ;
  assign n20784 = n20783 ^ n18968 ^ 1'b0 ;
  assign n20785 = n5952 | n7777 ;
  assign n20786 = n8849 ^ n5157 ^ 1'b0 ;
  assign n20787 = n19493 & ~n20786 ;
  assign n20788 = ~n6921 & n7690 ;
  assign n20789 = ~n4065 & n20788 ;
  assign n20790 = n3268 & ~n9616 ;
  assign n20791 = ( n2814 & n5490 ) | ( n2814 & n14378 ) | ( n5490 & n14378 ) ;
  assign n20792 = n18181 ^ n15479 ^ 1'b0 ;
  assign n20793 = ~n2303 & n2961 ;
  assign n20794 = n5267 & n20793 ;
  assign n20795 = n20794 ^ n14652 ^ 1'b0 ;
  assign n20796 = n13274 ^ n11269 ^ 1'b0 ;
  assign n20797 = n5755 | n20796 ;
  assign n20798 = n20797 ^ n2436 ^ 1'b0 ;
  assign n20799 = n6538 & ~n20798 ;
  assign n20800 = n18595 ^ n4164 ^ n4106 ;
  assign n20801 = n17674 ^ n5693 ^ n4109 ;
  assign n20802 = n8916 ^ n4418 ^ n175 ;
  assign n20803 = n2474 & ~n17862 ;
  assign n20804 = n18814 & ~n20803 ;
  assign n20805 = ~n20802 & n20804 ;
  assign n20806 = n6653 | n8247 ;
  assign n20807 = n7794 ^ n6579 ^ 1'b0 ;
  assign n20808 = n20807 ^ n2735 ^ 1'b0 ;
  assign n20809 = ~n171 & n10370 ;
  assign n20810 = n20809 ^ n6176 ^ 1'b0 ;
  assign n20811 = n11740 & ~n20810 ;
  assign n20812 = n3010 & ~n3373 ;
  assign n20813 = n5649 & ~n12866 ;
  assign n20814 = n9987 & ~n16242 ;
  assign n20815 = n4082 & ~n4514 ;
  assign n20816 = n6771 & ~n20815 ;
  assign n20817 = ~n2830 & n20816 ;
  assign n20818 = n11131 | n18424 ;
  assign n20819 = n1107 & ~n20818 ;
  assign n20820 = n14724 ^ n637 ^ 1'b0 ;
  assign n20821 = n18817 ^ n6050 ^ 1'b0 ;
  assign n20822 = n5969 & ~n20821 ;
  assign n20823 = n8368 & n20822 ;
  assign n20824 = n20823 ^ n832 ^ 1'b0 ;
  assign n20825 = n7043 & n20824 ;
  assign n20826 = n3376 & ~n14555 ;
  assign n20827 = n5321 & n5394 ;
  assign n20828 = ~n19545 & n20827 ;
  assign n20829 = n8910 & n11823 ;
  assign n20830 = n857 & n2174 ;
  assign n20831 = n12511 ^ n11544 ^ n6580 ;
  assign n20832 = n11274 ^ n9022 ^ 1'b0 ;
  assign n20833 = n1738 & ~n20832 ;
  assign n20834 = n11034 & n14679 ;
  assign n20835 = n7689 & n20834 ;
  assign n20836 = n1756 | n20835 ;
  assign n20837 = n20836 ^ n1892 ^ 1'b0 ;
  assign n20838 = n20833 & n20837 ;
  assign n20839 = ( n531 & n2564 ) | ( n531 & ~n6863 ) | ( n2564 & ~n6863 ) ;
  assign n20841 = ( ~n1003 & n19061 ) | ( ~n1003 & n19661 ) | ( n19061 & n19661 ) ;
  assign n20840 = n13636 ^ n6550 ^ 1'b0 ;
  assign n20842 = n20841 ^ n20840 ^ n14930 ;
  assign n20843 = ~n13634 & n20170 ;
  assign n20844 = n18125 & n20843 ;
  assign n20845 = n3903 | n9660 ;
  assign n20846 = n20845 ^ n9865 ^ 1'b0 ;
  assign n20847 = ~n1287 & n4530 ;
  assign n20848 = n20847 ^ n13215 ^ 1'b0 ;
  assign n20849 = n4333 & ~n12754 ;
  assign n20850 = n1835 & n20849 ;
  assign n20851 = n13021 & ~n20850 ;
  assign n20852 = n7228 ^ n5315 ^ 1'b0 ;
  assign n20853 = ( ~n2922 & n7532 ) | ( ~n2922 & n20852 ) | ( n7532 & n20852 ) ;
  assign n20854 = ( n20848 & n20851 ) | ( n20848 & ~n20853 ) | ( n20851 & ~n20853 ) ;
  assign n20855 = ( ~n6415 & n8158 ) | ( ~n6415 & n9127 ) | ( n8158 & n9127 ) ;
  assign n20856 = ~n13758 & n20855 ;
  assign n20857 = n11797 & ~n14336 ;
  assign n20858 = n20857 ^ n3520 ^ 1'b0 ;
  assign n20859 = n20858 ^ n469 ^ 1'b0 ;
  assign n20862 = n3270 ^ n1231 ^ 1'b0 ;
  assign n20863 = n868 | n20862 ;
  assign n20860 = n2249 | n8531 ;
  assign n20861 = ~n11026 & n20860 ;
  assign n20864 = n20863 ^ n20861 ^ 1'b0 ;
  assign n20865 = n1201 ^ n859 ^ 1'b0 ;
  assign n20866 = ~n19648 & n20865 ;
  assign n20867 = n1200 & n8788 ;
  assign n20868 = n15759 & n20867 ;
  assign n20869 = n14014 ^ n6789 ^ 1'b0 ;
  assign n20870 = n4033 & n6658 ;
  assign n20871 = n20870 ^ n9266 ^ 1'b0 ;
  assign n20872 = n20869 & ~n20871 ;
  assign n20873 = n4002 | n9613 ;
  assign n20874 = n2915 | n20873 ;
  assign n20875 = ( n6060 & n8210 ) | ( n6060 & ~n20874 ) | ( n8210 & ~n20874 ) ;
  assign n20876 = n9273 & ~n18782 ;
  assign n20877 = ~n12853 & n20876 ;
  assign n20878 = n9601 | n20877 ;
  assign n20879 = n12727 ^ n2053 ^ 1'b0 ;
  assign n20880 = ~n1402 & n20879 ;
  assign n20881 = n6437 ^ n5043 ^ 1'b0 ;
  assign n20882 = ~n9880 & n20881 ;
  assign n20883 = n17862 ^ n13035 ^ 1'b0 ;
  assign n20884 = n9421 & ~n20883 ;
  assign n20885 = ~n5351 & n5787 ;
  assign n20886 = n20885 ^ n4273 ^ 1'b0 ;
  assign n20887 = n10850 ^ n8452 ^ n3942 ;
  assign n20888 = n4994 ^ n1865 ^ 1'b0 ;
  assign n20889 = n12443 ^ n1467 ^ n618 ;
  assign n20890 = ~n3564 & n20889 ;
  assign n20891 = n1133 & ~n19544 ;
  assign n20892 = ~n141 & n852 ;
  assign n20893 = n14846 ^ n13648 ^ 1'b0 ;
  assign n20894 = n16152 ^ n10017 ^ n2684 ;
  assign n20895 = n10485 ^ n5304 ^ 1'b0 ;
  assign n20896 = ~n5598 & n20895 ;
  assign n20897 = ~n12092 & n20896 ;
  assign n20898 = n20897 ^ n2103 ^ n1049 ;
  assign n20899 = n16179 ^ n4776 ^ 1'b0 ;
  assign n20900 = n5291 & ~n20899 ;
  assign n20901 = n20900 ^ n6334 ^ 1'b0 ;
  assign n20902 = ~n12778 & n12896 ;
  assign n20903 = n1909 & n20902 ;
  assign n20904 = ~n1419 & n5373 ;
  assign n20905 = ~n5020 & n8413 ;
  assign n20906 = n20905 ^ n5358 ^ 1'b0 ;
  assign n20907 = n20906 ^ n307 ^ 1'b0 ;
  assign n20908 = ~n4493 & n20907 ;
  assign n20909 = n6940 & ~n12071 ;
  assign n20910 = ( n560 & n11071 ) | ( n560 & ~n20909 ) | ( n11071 & ~n20909 ) ;
  assign n20914 = n487 | n3075 ;
  assign n20911 = n625 & ~n1796 ;
  assign n20912 = n20911 ^ n7842 ^ 1'b0 ;
  assign n20913 = ~n13516 & n20912 ;
  assign n20915 = n20914 ^ n20913 ^ 1'b0 ;
  assign n20916 = n3792 & n6954 ;
  assign n20917 = n198 & n20916 ;
  assign n20918 = n3238 & ~n20917 ;
  assign n20919 = n12684 ^ n789 ^ 1'b0 ;
  assign n20920 = n1868 & ~n20919 ;
  assign n20921 = n1627 | n3757 ;
  assign n20922 = n20921 ^ n3124 ^ 1'b0 ;
  assign n20923 = n20922 ^ n10084 ^ 1'b0 ;
  assign n20924 = n6652 ^ n3027 ^ 1'b0 ;
  assign n20925 = n20923 | n20924 ;
  assign n20926 = n14847 ^ n7822 ^ 1'b0 ;
  assign n20927 = n8794 & ~n14877 ;
  assign n20928 = ~n4565 & n20927 ;
  assign n20929 = n1157 | n20928 ;
  assign n20930 = n11154 & n15222 ;
  assign n20931 = n15147 ^ n13082 ^ n2224 ;
  assign n20932 = n20931 ^ n17746 ^ 1'b0 ;
  assign n20933 = ~n504 & n10643 ;
  assign n20934 = n20933 ^ n16863 ^ 1'b0 ;
  assign n20935 = n4423 & n20934 ;
  assign n20936 = n4666 & ~n6426 ;
  assign n20937 = n2758 & n20936 ;
  assign n20938 = ~n875 & n20937 ;
  assign n20939 = n9290 | n12782 ;
  assign n20940 = n6547 & ~n20939 ;
  assign n20941 = n6930 & ~n9005 ;
  assign n20942 = n3286 & n20941 ;
  assign n20943 = n10520 | n12081 ;
  assign n20944 = n17638 | n20943 ;
  assign n20945 = n20944 ^ n1620 ^ 1'b0 ;
  assign n20946 = n7568 ^ n4115 ^ n2280 ;
  assign n20947 = ~n7878 & n8100 ;
  assign n20948 = n20947 ^ n453 ^ 1'b0 ;
  assign n20949 = n18026 & n20948 ;
  assign n20950 = n20949 ^ n5374 ^ 1'b0 ;
  assign n20954 = n8868 & ~n11968 ;
  assign n20955 = n2233 & n4472 ;
  assign n20956 = n20955 ^ n6511 ^ 1'b0 ;
  assign n20957 = n20956 ^ n13133 ^ 1'b0 ;
  assign n20958 = n20954 & ~n20957 ;
  assign n20951 = n339 & n2919 ;
  assign n20952 = n19614 & n20951 ;
  assign n20953 = n20952 ^ n10755 ^ 1'b0 ;
  assign n20959 = n20958 ^ n20953 ^ 1'b0 ;
  assign n20960 = n13392 ^ n842 ^ 1'b0 ;
  assign n20961 = ~n623 & n3498 ;
  assign n20962 = n3740 & n20961 ;
  assign n20963 = n4648 | n15822 ;
  assign n20964 = n20963 ^ n6139 ^ n811 ;
  assign n20965 = ~n1916 & n2308 ;
  assign n20966 = ~n292 & n20965 ;
  assign n20967 = n20966 ^ n7384 ^ n971 ;
  assign n20968 = n10046 ^ n2635 ^ 1'b0 ;
  assign n20969 = ~n15833 & n18813 ;
  assign n20970 = n20969 ^ n3482 ^ 1'b0 ;
  assign n20971 = n6458 & n20970 ;
  assign n20972 = x93 & ~n5834 ;
  assign n20973 = n2823 | n3403 ;
  assign n20974 = n14142 | n20973 ;
  assign n20975 = n20974 ^ n19293 ^ 1'b0 ;
  assign n20976 = n10528 & ~n19184 ;
  assign n20977 = n20976 ^ n12902 ^ 1'b0 ;
  assign n20978 = n3286 ^ n3164 ^ 1'b0 ;
  assign n20979 = n997 & ~n20978 ;
  assign n20980 = n18365 ^ n5930 ^ 1'b0 ;
  assign n20981 = ( ~n7532 & n20979 ) | ( ~n7532 & n20980 ) | ( n20979 & n20980 ) ;
  assign n20982 = n17953 ^ n3065 ^ n2899 ;
  assign n20983 = n2332 | n4190 ;
  assign n20984 = n18558 | n20983 ;
  assign n20985 = n20984 ^ n7866 ^ 1'b0 ;
  assign n20986 = n6216 | n11277 ;
  assign n20987 = n20986 ^ n4430 ^ 1'b0 ;
  assign n20988 = ~n1079 & n7349 ;
  assign n20989 = n2366 & n20988 ;
  assign n20990 = n468 | n20989 ;
  assign n20991 = n10054 & ~n14995 ;
  assign n20992 = ~n2942 & n8854 ;
  assign n20993 = n632 & n20992 ;
  assign n20994 = n8061 ^ x79 ^ 1'b0 ;
  assign n20995 = n1619 | n5906 ;
  assign n20996 = n562 | n20995 ;
  assign n20997 = ( n309 & n10887 ) | ( n309 & ~n19533 ) | ( n10887 & ~n19533 ) ;
  assign n20998 = n13621 ^ x1 ^ 1'b0 ;
  assign n20999 = n438 & ~n20998 ;
  assign n21000 = ~n5301 & n20999 ;
  assign n21001 = ( ~n1281 & n11778 ) | ( ~n1281 & n21000 ) | ( n11778 & n21000 ) ;
  assign n21002 = n6550 & n19644 ;
  assign n21003 = n1126 | n6961 ;
  assign n21004 = x102 | n21003 ;
  assign n21005 = ~n15554 & n15609 ;
  assign n21006 = n14313 & n21005 ;
  assign n21007 = n21006 ^ n14929 ^ 1'b0 ;
  assign n21008 = n21004 & n21007 ;
  assign n21009 = ~n4268 & n9441 ;
  assign n21010 = ~n3740 & n21009 ;
  assign n21011 = n21010 ^ n8738 ^ 1'b0 ;
  assign n21012 = n965 & ~n21011 ;
  assign n21013 = n15387 | n18631 ;
  assign n21014 = n21013 ^ n6263 ^ 1'b0 ;
  assign n21015 = n4611 | n21014 ;
  assign n21016 = n1450 & n3746 ;
  assign n21017 = n21016 ^ n7866 ^ 1'b0 ;
  assign n21018 = n17438 ^ n8913 ^ x41 ;
  assign n21019 = n14841 & ~n21018 ;
  assign n21020 = n10909 & n13601 ;
  assign n21021 = n11473 ^ n2137 ^ 1'b0 ;
  assign n21022 = n7222 & ~n19009 ;
  assign n21023 = n21022 ^ n6384 ^ 1'b0 ;
  assign n21024 = ( n269 & ~n388 ) | ( n269 & n10977 ) | ( ~n388 & n10977 ) ;
  assign n21025 = n1948 & n15269 ;
  assign n21026 = n9625 & n21025 ;
  assign n21027 = ~n2463 & n21026 ;
  assign n21028 = n13082 ^ n10806 ^ n3501 ;
  assign n21029 = n21028 ^ n2444 ^ 1'b0 ;
  assign n21030 = n15769 ^ n12031 ^ 1'b0 ;
  assign n21031 = ~n7794 & n21030 ;
  assign n21032 = ~n8395 & n15012 ;
  assign n21033 = n7526 & n21032 ;
  assign n21035 = n1411 | n5002 ;
  assign n21034 = n3961 ^ n2830 ^ 1'b0 ;
  assign n21036 = n21035 ^ n21034 ^ 1'b0 ;
  assign n21037 = ( n6659 & n8476 ) | ( n6659 & n10389 ) | ( n8476 & n10389 ) ;
  assign n21038 = n1821 & ~n6744 ;
  assign n21039 = n3105 | n11666 ;
  assign n21040 = n21038 | n21039 ;
  assign n21041 = n1030 | n7902 ;
  assign n21042 = n21041 ^ n621 ^ 1'b0 ;
  assign n21043 = n4235 | n15046 ;
  assign n21044 = n21043 ^ n14632 ^ 1'b0 ;
  assign n21045 = n17818 | n21044 ;
  assign n21046 = n3773 & ~n4308 ;
  assign n21047 = n21046 ^ n6421 ^ 1'b0 ;
  assign n21048 = ( n2983 & n11366 ) | ( n2983 & n21047 ) | ( n11366 & n21047 ) ;
  assign n21049 = ( n3604 & ~n8129 ) | ( n3604 & n10842 ) | ( ~n8129 & n10842 ) ;
  assign n21053 = n7807 | n11253 ;
  assign n21050 = n2827 | n4979 ;
  assign n21051 = ~n4771 & n21050 ;
  assign n21052 = n586 & n21051 ;
  assign n21054 = n21053 ^ n21052 ^ 1'b0 ;
  assign n21055 = n2694 ^ n2215 ^ 1'b0 ;
  assign n21056 = ~n476 & n21055 ;
  assign n21057 = n2070 | n21056 ;
  assign n21058 = n13021 & ~n21057 ;
  assign n21059 = n14615 ^ n225 ^ 1'b0 ;
  assign n21060 = ~n3564 & n8595 ;
  assign n21061 = ~n12774 & n21060 ;
  assign n21062 = n7711 ^ n371 ^ 1'b0 ;
  assign n21063 = ~n1797 & n3344 ;
  assign n21064 = n6015 & n21063 ;
  assign n21065 = ( n12455 & ~n21062 ) | ( n12455 & n21064 ) | ( ~n21062 & n21064 ) ;
  assign n21066 = n3820 ^ n1526 ^ 1'b0 ;
  assign n21067 = ~n2670 & n21066 ;
  assign n21068 = n4588 | n10463 ;
  assign n21069 = n21067 | n21068 ;
  assign n21070 = n21069 ^ n16081 ^ 1'b0 ;
  assign n21071 = n21070 ^ n20934 ^ n16062 ;
  assign n21072 = ( n1166 & n1271 ) | ( n1166 & n7705 ) | ( n1271 & n7705 ) ;
  assign n21073 = n5046 ^ n788 ^ 1'b0 ;
  assign n21074 = n15043 & n21073 ;
  assign n21075 = n21072 & n21074 ;
  assign n21076 = n14614 ^ n8878 ^ 1'b0 ;
  assign n21077 = n11882 ^ n9802 ^ 1'b0 ;
  assign n21078 = n3510 ^ n1747 ^ 1'b0 ;
  assign n21079 = n9211 ^ n357 ^ 1'b0 ;
  assign n21080 = n5430 & ~n12712 ;
  assign n21081 = ~n14267 & n21080 ;
  assign n21082 = n4786 & ~n21081 ;
  assign n21083 = n1676 & ~n17006 ;
  assign n21084 = n21083 ^ n867 ^ 1'b0 ;
  assign n21087 = n7877 ^ n1418 ^ 1'b0 ;
  assign n21088 = n3139 | n21087 ;
  assign n21085 = n1011 | n16222 ;
  assign n21086 = n21085 ^ n6809 ^ 1'b0 ;
  assign n21089 = n21088 ^ n21086 ^ n13683 ;
  assign n21090 = ( ~n6764 & n10551 ) | ( ~n6764 & n16134 ) | ( n10551 & n16134 ) ;
  assign n21091 = ~n11029 & n11842 ;
  assign n21092 = n21091 ^ n1317 ^ 1'b0 ;
  assign n21093 = n2738 ^ n1774 ^ 1'b0 ;
  assign n21094 = n15164 & n21093 ;
  assign n21095 = n795 & n15341 ;
  assign n21096 = n21095 ^ n10307 ^ 1'b0 ;
  assign n21097 = n21096 ^ n13926 ^ 1'b0 ;
  assign n21098 = n6946 & ~n8873 ;
  assign n21099 = n1192 | n16518 ;
  assign n21100 = n21099 ^ n13623 ^ n5063 ;
  assign n21101 = n962 | n21100 ;
  assign n21102 = ~n5050 & n13172 ;
  assign n21103 = ~n8760 & n21102 ;
  assign n21104 = n21103 ^ n10064 ^ 1'b0 ;
  assign n21105 = n19797 ^ n2213 ^ 1'b0 ;
  assign n21106 = n3061 | n21105 ;
  assign n21107 = n8826 & ~n21106 ;
  assign n21108 = n6210 & n21107 ;
  assign n21109 = n14769 | n21108 ;
  assign n21110 = n8671 ^ n8491 ^ 1'b0 ;
  assign n21111 = n21110 ^ n18784 ^ n3744 ;
  assign n21112 = n5069 & n12215 ;
  assign n21113 = n15983 ^ n8695 ^ 1'b0 ;
  assign n21114 = n17138 & n21113 ;
  assign n21115 = n13659 ^ n12555 ^ n10162 ;
  assign n21116 = n9920 & n16559 ;
  assign n21117 = ~n21115 & n21116 ;
  assign n21118 = n20292 ^ n13439 ^ n11554 ;
  assign n21119 = n4797 & ~n10035 ;
  assign n21120 = n5189 & ~n6728 ;
  assign n21121 = n6519 & n8827 ;
  assign n21122 = n9812 ^ n3848 ^ 1'b0 ;
  assign n21123 = n6277 | n21122 ;
  assign n21125 = n2289 & n12445 ;
  assign n21124 = n981 & n1803 ;
  assign n21126 = n21125 ^ n21124 ^ 1'b0 ;
  assign n21127 = n3488 | n17708 ;
  assign n21128 = n21127 ^ n6665 ^ 1'b0 ;
  assign n21129 = n20703 ^ n6488 ^ n905 ;
  assign n21130 = ~n8801 & n12577 ;
  assign n21131 = n21130 ^ n3773 ^ n941 ;
  assign n21132 = n3401 & n16297 ;
  assign n21133 = n18113 ^ n6242 ^ 1'b0 ;
  assign n21134 = n4148 ^ n2656 ^ 1'b0 ;
  assign n21135 = n17598 ^ n6559 ^ 1'b0 ;
  assign n21136 = n14171 & ~n21135 ;
  assign n21137 = n6571 ^ n4542 ^ 1'b0 ;
  assign n21138 = n1394 & n21137 ;
  assign n21139 = n19102 | n21138 ;
  assign n21140 = n3655 | n10075 ;
  assign n21141 = n16881 | n21140 ;
  assign n21142 = n3367 & ~n15789 ;
  assign n21143 = ~n1766 & n21142 ;
  assign n21144 = n21062 | n21143 ;
  assign n21145 = n14045 ^ n630 ^ 1'b0 ;
  assign n21146 = ( n5152 & n18425 ) | ( n5152 & n19602 ) | ( n18425 & n19602 ) ;
  assign n21147 = n21146 ^ n7244 ^ 1'b0 ;
  assign n21148 = n6758 & ~n10039 ;
  assign n21149 = n10039 & n21148 ;
  assign n21150 = n20378 ^ n15068 ^ 1'b0 ;
  assign n21151 = n8420 ^ n694 ^ 1'b0 ;
  assign n21152 = n165 | n21151 ;
  assign n21153 = n220 | n3524 ;
  assign n21154 = n9342 | n21153 ;
  assign n21155 = n17677 ^ n12565 ^ 1'b0 ;
  assign n21156 = n18396 ^ n8514 ^ 1'b0 ;
  assign n21157 = n17325 & ~n21156 ;
  assign n21158 = n21157 ^ n5634 ^ 1'b0 ;
  assign n21159 = n18014 ^ n4700 ^ 1'b0 ;
  assign n21160 = n8458 & ~n19737 ;
  assign n21161 = n21160 ^ n4147 ^ 1'b0 ;
  assign n21163 = n5062 | n11723 ;
  assign n21162 = n425 & n12044 ;
  assign n21164 = n21163 ^ n21162 ^ 1'b0 ;
  assign n21165 = n18973 ^ x79 ^ 1'b0 ;
  assign n21166 = ~n19233 & n21165 ;
  assign n21167 = n9998 ^ n1012 ^ 1'b0 ;
  assign n21168 = n2417 & ~n15489 ;
  assign n21169 = n21168 ^ n6318 ^ 1'b0 ;
  assign n21170 = ~n2033 & n5584 ;
  assign n21171 = n1163 & ~n21170 ;
  assign n21172 = n9472 ^ n3503 ^ 1'b0 ;
  assign n21173 = n21171 & ~n21172 ;
  assign n21174 = n6140 & n13788 ;
  assign n21175 = ~n21173 & n21174 ;
  assign n21176 = n8323 ^ n8097 ^ 1'b0 ;
  assign n21180 = n5446 & ~n9022 ;
  assign n21178 = n8265 ^ n163 ^ 1'b0 ;
  assign n21179 = n5014 & ~n21178 ;
  assign n21177 = n11715 ^ n10729 ^ n1464 ;
  assign n21181 = n21180 ^ n21179 ^ n21177 ;
  assign n21182 = n17941 ^ n14149 ^ 1'b0 ;
  assign n21184 = n13057 ^ n11275 ^ n5127 ;
  assign n21183 = n9139 & n20807 ;
  assign n21185 = n21184 ^ n21183 ^ 1'b0 ;
  assign n21186 = n3210 ^ n1096 ^ 1'b0 ;
  assign n21187 = n4774 & n21186 ;
  assign n21188 = n21187 ^ n4443 ^ 1'b0 ;
  assign n21190 = n2529 & n3399 ;
  assign n21189 = n6037 & n14172 ;
  assign n21191 = n21190 ^ n21189 ^ n1505 ;
  assign n21192 = n10606 ^ n335 ^ 1'b0 ;
  assign n21193 = n1295 & ~n6263 ;
  assign n21194 = n4224 & ~n8172 ;
  assign n21195 = ~n6565 & n21194 ;
  assign n21196 = ( ~n1221 & n10105 ) | ( ~n1221 & n21195 ) | ( n10105 & n21195 ) ;
  assign n21197 = n14243 | n21196 ;
  assign n21198 = n21193 | n21197 ;
  assign n21199 = n3795 | n4440 ;
  assign n21200 = n6201 ^ n5046 ^ n4849 ;
  assign n21201 = n11933 & ~n20145 ;
  assign n21202 = ~n6442 & n21201 ;
  assign n21203 = ( ~n555 & n1374 ) | ( ~n555 & n2861 ) | ( n1374 & n2861 ) ;
  assign n21204 = ( n5074 & n10232 ) | ( n5074 & n21203 ) | ( n10232 & n21203 ) ;
  assign n21205 = n14990 & ~n16136 ;
  assign n21206 = ~n1990 & n21205 ;
  assign n21207 = n21206 ^ n3133 ^ 1'b0 ;
  assign n21208 = n11882 | n21207 ;
  assign n21209 = n15502 | n21208 ;
  assign n21210 = n8237 | n21209 ;
  assign n21211 = n3367 ^ x23 ^ 1'b0 ;
  assign n21212 = ( n440 & ~n2168 ) | ( n440 & n3515 ) | ( ~n2168 & n3515 ) ;
  assign n21213 = n2513 & n3390 ;
  assign n21214 = ~n15246 & n21213 ;
  assign n21215 = n832 & n6347 ;
  assign n21216 = n13777 ^ n3968 ^ 1'b0 ;
  assign n21217 = n1586 | n21216 ;
  assign n21218 = n4997 ^ x69 ^ 1'b0 ;
  assign n21219 = ~n21217 & n21218 ;
  assign n21220 = n12812 ^ n7687 ^ n6111 ;
  assign n21221 = n21220 ^ n16768 ^ 1'b0 ;
  assign n21222 = ~x17 & n2280 ;
  assign n21223 = n2508 ^ n551 ^ 1'b0 ;
  assign n21224 = n13991 & n21223 ;
  assign n21225 = ~n10535 & n17787 ;
  assign n21226 = ~x34 & n11863 ;
  assign n21227 = n17344 ^ n13227 ^ 1'b0 ;
  assign n21228 = ~n7493 & n21227 ;
  assign n21229 = n5283 & ~n11680 ;
  assign n21230 = n21229 ^ n16670 ^ 1'b0 ;
  assign n21231 = n14471 ^ n1670 ^ 1'b0 ;
  assign n21232 = n16108 & ~n16344 ;
  assign n21233 = n3041 ^ n2684 ^ n1348 ;
  assign n21234 = ~n4073 & n7547 ;
  assign n21235 = ( n1432 & ~n3222 ) | ( n1432 & n6264 ) | ( ~n3222 & n6264 ) ;
  assign n21236 = n3413 | n7851 ;
  assign n21237 = n21235 | n21236 ;
  assign n21238 = n21237 ^ n6652 ^ 1'b0 ;
  assign n21239 = n11315 & n16511 ;
  assign n21240 = n21239 ^ n6240 ^ 1'b0 ;
  assign n21241 = n7002 & n14939 ;
  assign n21242 = ~n8446 & n10941 ;
  assign n21243 = n4967 ^ n3761 ^ 1'b0 ;
  assign n21244 = n19461 ^ n16689 ^ 1'b0 ;
  assign n21245 = n9522 ^ n4881 ^ 1'b0 ;
  assign n21246 = n7002 & n21245 ;
  assign n21247 = n21246 ^ n10862 ^ 1'b0 ;
  assign n21248 = n503 & ~n5894 ;
  assign n21249 = n21248 ^ n506 ^ 1'b0 ;
  assign n21250 = n500 & n21249 ;
  assign n21251 = n21250 ^ n4432 ^ 1'b0 ;
  assign n21252 = n1599 & n21251 ;
  assign n21253 = n14108 | n14609 ;
  assign n21254 = n14381 | n21253 ;
  assign n21255 = n4216 & ~n9473 ;
  assign n21256 = n2221 & n21255 ;
  assign n21257 = n21256 ^ n3033 ^ 1'b0 ;
  assign n21258 = n21254 & n21257 ;
  assign n21259 = n10198 | n14761 ;
  assign n21260 = ~n10311 & n18378 ;
  assign n21261 = ( n10657 & n11251 ) | ( n10657 & ~n12915 ) | ( n11251 & ~n12915 ) ;
  assign n21262 = n4766 | n21261 ;
  assign n21263 = n21262 ^ n10224 ^ 1'b0 ;
  assign n21264 = n3215 | n21263 ;
  assign n21265 = n2211 | n7880 ;
  assign n21266 = n1204 | n21265 ;
  assign n21267 = ~n9236 & n15410 ;
  assign n21268 = ~n14801 & n18435 ;
  assign n21269 = n591 & n21268 ;
  assign n21270 = n21269 ^ n5868 ^ 1'b0 ;
  assign n21271 = n3790 & n10128 ;
  assign n21272 = ~n625 & n2333 ;
  assign n21273 = n13656 ^ n4697 ^ 1'b0 ;
  assign n21274 = ~n21272 & n21273 ;
  assign n21275 = n17082 & ~n21274 ;
  assign n21276 = n2270 & ~n5881 ;
  assign n21277 = ~n11760 & n21276 ;
  assign n21278 = n21277 ^ n6109 ^ 1'b0 ;
  assign n21279 = ~n1635 & n4547 ;
  assign n21280 = n3724 & n21279 ;
  assign n21281 = n8231 | n21280 ;
  assign n21282 = n21281 ^ n9366 ^ 1'b0 ;
  assign n21283 = n21282 ^ n16150 ^ n7755 ;
  assign n21284 = ~n2756 & n10433 ;
  assign n21285 = n12302 & ~n19797 ;
  assign n21286 = n21285 ^ n8599 ^ 1'b0 ;
  assign n21287 = ~n6099 & n21286 ;
  assign n21288 = n21287 ^ n3606 ^ 1'b0 ;
  assign n21289 = ~n4777 & n15649 ;
  assign n21290 = n21024 ^ n19382 ^ 1'b0 ;
  assign n21297 = n1120 | n17931 ;
  assign n21291 = ~n4333 & n14561 ;
  assign n21292 = ~n1950 & n3303 ;
  assign n21293 = n21291 & n21292 ;
  assign n21294 = n4412 ^ n2030 ^ 1'b0 ;
  assign n21295 = n9758 & ~n21294 ;
  assign n21296 = ~n21293 & n21295 ;
  assign n21298 = n21297 ^ n21296 ^ 1'b0 ;
  assign n21299 = n5559 & ~n21298 ;
  assign n21300 = n18780 & n21299 ;
  assign n21301 = n137 | n12706 ;
  assign n21302 = n21301 ^ n1150 ^ 1'b0 ;
  assign n21303 = ~n3378 & n12896 ;
  assign n21304 = n21303 ^ n2676 ^ 1'b0 ;
  assign n21305 = n21302 | n21304 ;
  assign n21306 = n192 & ~n859 ;
  assign n21307 = ~n192 & n21306 ;
  assign n21308 = ~n623 & n982 ;
  assign n21309 = n623 & n21308 ;
  assign n21310 = n21309 ^ n1761 ^ 1'b0 ;
  assign n21311 = ~n21307 & n21310 ;
  assign n21312 = n4199 & n21311 ;
  assign n21313 = n732 & n21312 ;
  assign n21314 = n7481 | n21313 ;
  assign n21315 = n21314 ^ n13031 ^ n8023 ;
  assign n21316 = n6626 | n7235 ;
  assign n21317 = n21316 ^ n147 ^ 1'b0 ;
  assign n21318 = n2416 & ~n16296 ;
  assign n21319 = n10345 | n19138 ;
  assign n21325 = n5927 & ~n7942 ;
  assign n21320 = n3442 | n5443 ;
  assign n21321 = n3442 & ~n21320 ;
  assign n21322 = n666 | n21321 ;
  assign n21323 = n666 & ~n21322 ;
  assign n21324 = n6669 & ~n21323 ;
  assign n21326 = n21325 ^ n21324 ^ 1'b0 ;
  assign n21327 = n792 & ~n21326 ;
  assign n21328 = ~n3122 & n5398 ;
  assign n21329 = n642 & n8709 ;
  assign n21330 = n21329 ^ n1464 ^ 1'b0 ;
  assign n21331 = n19399 ^ n5958 ^ 1'b0 ;
  assign n21332 = n11099 ^ n971 ^ 1'b0 ;
  assign n21333 = ~n4978 & n21332 ;
  assign n21334 = n21333 ^ n486 ^ 1'b0 ;
  assign n21335 = n2076 & ~n5015 ;
  assign n21336 = n6923 | n19634 ;
  assign n21337 = n5256 | n21336 ;
  assign n21338 = n7325 & ~n8121 ;
  assign n21339 = n14339 ^ n2497 ^ 1'b0 ;
  assign n21340 = n12014 ^ n2797 ^ 1'b0 ;
  assign n21341 = n15433 | n21340 ;
  assign n21342 = ( n21338 & ~n21339 ) | ( n21338 & n21341 ) | ( ~n21339 & n21341 ) ;
  assign n21343 = ~n741 & n2289 ;
  assign n21344 = n21343 ^ n1180 ^ 1'b0 ;
  assign n21345 = n11877 & n21344 ;
  assign n21346 = ~n4271 & n16088 ;
  assign n21347 = ~n21325 & n21346 ;
  assign n21348 = n16115 ^ n2893 ^ 1'b0 ;
  assign n21349 = n21347 | n21348 ;
  assign n21350 = n6046 & n13982 ;
  assign n21351 = n5124 | n10072 ;
  assign n21352 = n5492 | n21351 ;
  assign n21353 = n1300 & n16767 ;
  assign n21354 = n3558 & n21353 ;
  assign n21355 = n13131 | n21354 ;
  assign n21356 = n21352 & ~n21355 ;
  assign n21357 = ~n882 & n11739 ;
  assign n21358 = n21357 ^ n4176 ^ 1'b0 ;
  assign n21359 = n5203 & ~n21358 ;
  assign n21360 = ~n874 & n7610 ;
  assign n21361 = n14811 & ~n19446 ;
  assign n21362 = n1165 & ~n3694 ;
  assign n21363 = n14149 | n17208 ;
  assign n21364 = n8262 & ~n19367 ;
  assign n21365 = n21364 ^ n13137 ^ 1'b0 ;
  assign n21366 = n3401 ^ n1804 ^ 1'b0 ;
  assign n21367 = n8434 & ~n21366 ;
  assign n21368 = ~n19192 & n21367 ;
  assign n21369 = ( ~n694 & n14878 ) | ( ~n694 & n16013 ) | ( n14878 & n16013 ) ;
  assign n21370 = n3615 & ~n12561 ;
  assign n21371 = n869 & n21370 ;
  assign n21372 = n11406 ^ n8368 ^ 1'b0 ;
  assign n21373 = n13048 ^ n666 ^ 1'b0 ;
  assign n21374 = ~n1545 & n21373 ;
  assign n21375 = ~n3209 & n6508 ;
  assign n21376 = n7158 ^ n1124 ^ 1'b0 ;
  assign n21377 = ~n21375 & n21376 ;
  assign n21380 = n7673 ^ n4302 ^ 1'b0 ;
  assign n21381 = n9256 & ~n21380 ;
  assign n21382 = ~n1785 & n2740 ;
  assign n21383 = ~n4082 & n21382 ;
  assign n21384 = ( n4359 & ~n6879 ) | ( n4359 & n21383 ) | ( ~n6879 & n21383 ) ;
  assign n21385 = ( ~n13293 & n21381 ) | ( ~n13293 & n21384 ) | ( n21381 & n21384 ) ;
  assign n21379 = ~n9344 & n13426 ;
  assign n21386 = n21385 ^ n21379 ^ 1'b0 ;
  assign n21378 = ~n3542 & n8112 ;
  assign n21387 = n21386 ^ n21378 ^ 1'b0 ;
  assign n21388 = n11758 & ~n20797 ;
  assign n21389 = n3908 & ~n13757 ;
  assign n21390 = ~n1545 & n16196 ;
  assign n21391 = n2529 & ~n2866 ;
  assign n21392 = n21391 ^ n10312 ^ 1'b0 ;
  assign n21393 = n5061 & n21392 ;
  assign n21394 = n6074 ^ n3046 ^ 1'b0 ;
  assign n21395 = n10222 & ~n21394 ;
  assign n21396 = n1959 & n14652 ;
  assign n21397 = n2546 & n11635 ;
  assign n21398 = n18452 ^ n10889 ^ n8339 ;
  assign n21401 = ( ~n1030 & n3130 ) | ( ~n1030 & n7951 ) | ( n3130 & n7951 ) ;
  assign n21402 = n21401 ^ n13064 ^ 1'b0 ;
  assign n21403 = n1565 & n21402 ;
  assign n21399 = ( n368 & n2473 ) | ( n368 & n4872 ) | ( n2473 & n4872 ) ;
  assign n21400 = n21399 ^ n9117 ^ 1'b0 ;
  assign n21404 = n21403 ^ n21400 ^ n11559 ;
  assign n21405 = n767 & n9186 ;
  assign n21406 = n4775 & n11665 ;
  assign n21407 = n6292 ^ n6055 ^ 1'b0 ;
  assign n21408 = n2658 & ~n21407 ;
  assign n21409 = n12069 ^ n3212 ^ 1'b0 ;
  assign n21410 = n16300 ^ n13775 ^ 1'b0 ;
  assign n21411 = n21409 | n21410 ;
  assign n21412 = n7753 & n16931 ;
  assign n21413 = n13425 & n18843 ;
  assign n21414 = ( n1845 & ~n15769 ) | ( n1845 & n21413 ) | ( ~n15769 & n21413 ) ;
  assign n21420 = x6 & n12569 ;
  assign n21421 = ~n6987 & n21420 ;
  assign n21415 = n20007 ^ n11410 ^ 1'b0 ;
  assign n21416 = n9363 | n13921 ;
  assign n21417 = n4037 & ~n21416 ;
  assign n21418 = n6886 & ~n21417 ;
  assign n21419 = ~n21415 & n21418 ;
  assign n21422 = n21421 ^ n21419 ^ n3246 ;
  assign n21423 = n4793 & n5613 ;
  assign n21424 = ~n5618 & n16640 ;
  assign n21425 = n3825 | n10346 ;
  assign n21426 = n14290 | n21425 ;
  assign n21427 = n8820 & n21426 ;
  assign n21429 = n150 & ~n1708 ;
  assign n21428 = n14086 | n17638 ;
  assign n21430 = n21429 ^ n21428 ^ 1'b0 ;
  assign n21431 = n4516 | n13602 ;
  assign n21432 = n12478 ^ n8451 ^ 1'b0 ;
  assign n21433 = n560 & n3800 ;
  assign n21434 = n4069 & n9984 ;
  assign n21435 = n16624 ^ n7713 ^ 1'b0 ;
  assign n21436 = n21434 | n21435 ;
  assign n21437 = n4843 & ~n20688 ;
  assign n21438 = n21437 ^ n4076 ^ 1'b0 ;
  assign n21439 = n3289 | n3292 ;
  assign n21440 = n161 & ~n9865 ;
  assign n21441 = n21439 & n21440 ;
  assign n21442 = n18445 ^ n5727 ^ n5176 ;
  assign n21443 = ( n3594 & n6419 ) | ( n3594 & n8167 ) | ( n6419 & n8167 ) ;
  assign n21444 = n21443 ^ n18790 ^ 1'b0 ;
  assign n21446 = n11512 ^ n240 ^ 1'b0 ;
  assign n21447 = ~n19549 & n21446 ;
  assign n21445 = n3074 | n8934 ;
  assign n21448 = n21447 ^ n21445 ^ 1'b0 ;
  assign n21449 = n12205 & ~n21448 ;
  assign n21450 = ( n15964 & n17107 ) | ( n15964 & n20914 ) | ( n17107 & n20914 ) ;
  assign n21451 = n21450 ^ n19766 ^ 1'b0 ;
  assign n21452 = n21451 ^ n12452 ^ 1'b0 ;
  assign n21453 = n8443 ^ n5492 ^ n2074 ;
  assign n21454 = n12391 ^ n7039 ^ 1'b0 ;
  assign n21455 = x23 | n21454 ;
  assign n21456 = n4396 & n17532 ;
  assign n21458 = n14372 ^ n10497 ^ 1'b0 ;
  assign n21459 = n10081 & ~n21458 ;
  assign n21460 = ~n417 & n1333 ;
  assign n21461 = ~n21459 & n21460 ;
  assign n21457 = n5062 & n14575 ;
  assign n21462 = n21461 ^ n21457 ^ 1'b0 ;
  assign n21463 = n6488 ^ n5654 ^ 1'b0 ;
  assign n21464 = n7941 & n21463 ;
  assign n21465 = ~n15479 & n21067 ;
  assign n21467 = ~n4292 & n9662 ;
  assign n21468 = ~n2020 & n21467 ;
  assign n21466 = n2790 ^ n1651 ^ 1'b0 ;
  assign n21469 = n21468 ^ n21466 ^ 1'b0 ;
  assign n21470 = ~n21465 & n21469 ;
  assign n21474 = n13832 ^ n10127 ^ 1'b0 ;
  assign n21471 = n1914 & ~n2800 ;
  assign n21472 = n7385 & n21471 ;
  assign n21473 = n1972 & ~n21472 ;
  assign n21475 = n21474 ^ n21473 ^ 1'b0 ;
  assign n21476 = n6659 ^ x120 ^ 1'b0 ;
  assign n21477 = ~n4293 & n21476 ;
  assign n21478 = n19247 ^ n8903 ^ n2370 ;
  assign n21479 = n13224 ^ n10527 ^ 1'b0 ;
  assign n21480 = n14094 | n21479 ;
  assign n21481 = n5580 ^ n3635 ^ n3336 ;
  assign n21482 = n573 & ~n9799 ;
  assign n21483 = n21482 ^ n9657 ^ 1'b0 ;
  assign n21484 = n12799 ^ n4350 ^ 1'b0 ;
  assign n21485 = n3479 ^ n1315 ^ 1'b0 ;
  assign n21486 = n17801 ^ n3744 ^ 1'b0 ;
  assign n21487 = n1774 | n21486 ;
  assign n21489 = ( ~n147 & n299 ) | ( ~n147 & n2931 ) | ( n299 & n2931 ) ;
  assign n21488 = n2680 & n17968 ;
  assign n21490 = n21489 ^ n21488 ^ 1'b0 ;
  assign n21491 = n17050 ^ n4601 ^ n3389 ;
  assign n21492 = n10715 | n21491 ;
  assign n21493 = n21492 ^ n13046 ^ 1'b0 ;
  assign n21494 = ~n12716 & n21493 ;
  assign n21495 = n8764 & ~n19258 ;
  assign n21496 = n3075 & ~n5801 ;
  assign n21497 = n1545 | n8247 ;
  assign n21498 = n8247 & ~n21497 ;
  assign n21499 = n373 | n21498 ;
  assign n21500 = n21498 & ~n21499 ;
  assign n21501 = n1562 | n21500 ;
  assign n21502 = n1562 & ~n21501 ;
  assign n21503 = n6474 | n21502 ;
  assign n21504 = n6474 & ~n21503 ;
  assign n21505 = n6340 ^ n3483 ^ 1'b0 ;
  assign n21506 = n3828 & n21505 ;
  assign n21507 = n959 & n3085 ;
  assign n21508 = ~n2455 & n21507 ;
  assign n21509 = n21508 ^ n4045 ^ 1'b0 ;
  assign n21510 = n21506 & ~n21509 ;
  assign n21511 = n21510 ^ n2405 ^ 1'b0 ;
  assign n21513 = ~n7731 & n12315 ;
  assign n21514 = n437 & n5064 ;
  assign n21515 = n3866 & n21514 ;
  assign n21516 = n21513 & n21515 ;
  assign n21512 = n7984 & ~n9973 ;
  assign n21517 = n21516 ^ n21512 ^ 1'b0 ;
  assign n21518 = ~n186 & n11406 ;
  assign n21519 = n4921 & n10244 ;
  assign n21520 = n2101 & n3326 ;
  assign n21521 = n7146 ^ n147 ^ 1'b0 ;
  assign n21522 = n3376 & ~n21521 ;
  assign n21523 = n3289 & ~n21522 ;
  assign n21524 = n21523 ^ n1965 ^ 1'b0 ;
  assign n21525 = n5814 & ~n21524 ;
  assign n21526 = n7006 ^ n5650 ^ 1'b0 ;
  assign n21527 = n21525 & n21526 ;
  assign n21528 = n12391 ^ n4769 ^ 1'b0 ;
  assign n21529 = ~n5156 & n13842 ;
  assign n21530 = n21528 & n21529 ;
  assign n21531 = n3452 | n3896 ;
  assign n21532 = n5208 & ~n21531 ;
  assign n21533 = n21532 ^ n964 ^ 1'b0 ;
  assign n21534 = n7039 | n21533 ;
  assign n21535 = ( n521 & n11072 ) | ( n521 & ~n15437 ) | ( n11072 & ~n15437 ) ;
  assign n21536 = n14419 | n14804 ;
  assign n21537 = n1951 & ~n6459 ;
  assign n21538 = n9351 & n21537 ;
  assign n21539 = n777 & ~n1619 ;
  assign n21540 = n19855 ^ n10997 ^ 1'b0 ;
  assign n21541 = n12394 | n21540 ;
  assign n21542 = n21541 ^ n15425 ^ 1'b0 ;
  assign n21543 = n4536 | n21542 ;
  assign n21544 = n13469 ^ n6488 ^ n1505 ;
  assign n21545 = n9376 ^ n175 ^ 1'b0 ;
  assign n21546 = n21544 | n21545 ;
  assign n21547 = n5012 | n21546 ;
  assign n21549 = ( n849 & n2906 ) | ( n849 & n3660 ) | ( n2906 & n3660 ) ;
  assign n21548 = n531 & n4065 ;
  assign n21550 = n21549 ^ n21548 ^ 1'b0 ;
  assign n21551 = n6940 ^ n6667 ^ 1'b0 ;
  assign n21552 = n21551 ^ n11224 ^ 1'b0 ;
  assign n21553 = n21550 & n21552 ;
  assign n21554 = n21298 ^ n351 ^ 1'b0 ;
  assign n21555 = n4156 | n18378 ;
  assign n21556 = n8355 | n12052 ;
  assign n21557 = ( n1899 & ~n10763 ) | ( n1899 & n16141 ) | ( ~n10763 & n16141 ) ;
  assign n21558 = n14591 ^ n4204 ^ 1'b0 ;
  assign n21559 = n7447 & ~n20544 ;
  assign n21560 = n18085 ^ n9666 ^ 1'b0 ;
  assign n21561 = ~n20850 & n21560 ;
  assign n21562 = n5797 & n14585 ;
  assign n21563 = n16032 ^ n3998 ^ 1'b0 ;
  assign n21564 = n21562 & n21563 ;
  assign n21565 = n16782 | n21564 ;
  assign n21566 = n5486 ^ n4859 ^ 1'b0 ;
  assign n21567 = n1597 & ~n5424 ;
  assign n21568 = n21567 ^ n9888 ^ 1'b0 ;
  assign n21569 = n11584 ^ n7449 ^ 1'b0 ;
  assign n21570 = n1103 | n21569 ;
  assign n21571 = n17095 & ~n21570 ;
  assign n21572 = n13930 ^ n11937 ^ 1'b0 ;
  assign n21573 = n14419 & n21572 ;
  assign n21574 = n13863 ^ n12573 ^ 1'b0 ;
  assign n21575 = ~n6620 & n21574 ;
  assign n21576 = n21575 ^ n11071 ^ 1'b0 ;
  assign n21578 = n12623 | n19826 ;
  assign n21577 = n5015 | n9678 ;
  assign n21579 = n21578 ^ n21577 ^ 1'b0 ;
  assign n21580 = n462 & n17445 ;
  assign n21581 = n19393 ^ n9587 ^ 1'b0 ;
  assign n21582 = n11596 ^ n8835 ^ 1'b0 ;
  assign n21583 = n19648 ^ n4434 ^ 1'b0 ;
  assign n21584 = n7282 & ~n11284 ;
  assign n21585 = n10851 & n21584 ;
  assign n21586 = n13849 ^ n2405 ^ 1'b0 ;
  assign n21587 = n14333 ^ n3390 ^ 1'b0 ;
  assign n21588 = n17541 ^ n1638 ^ 1'b0 ;
  assign n21589 = n2569 | n3544 ;
  assign n21590 = ~n12080 & n18931 ;
  assign n21591 = n21590 ^ n5301 ^ 1'b0 ;
  assign n21592 = n2235 & ~n10244 ;
  assign n21593 = n21591 & n21592 ;
  assign n21594 = n17457 ^ n16681 ^ 1'b0 ;
  assign n21596 = ~n3505 & n12532 ;
  assign n21595 = n7775 | n9525 ;
  assign n21597 = n21596 ^ n21595 ^ 1'b0 ;
  assign n21598 = n19575 ^ n3058 ^ 1'b0 ;
  assign n21599 = n6439 & ~n21598 ;
  assign n21600 = n5590 & ~n21599 ;
  assign n21601 = n5579 & n15391 ;
  assign n21602 = n4892 & n20491 ;
  assign n21603 = n11740 & ~n20141 ;
  assign n21604 = x105 & n14831 ;
  assign n21605 = ~n1919 & n21604 ;
  assign n21606 = n17426 ^ n3719 ^ n2168 ;
  assign n21607 = n11482 | n21606 ;
  assign n21608 = ~n14296 & n21607 ;
  assign n21609 = n1186 & ~n21608 ;
  assign n21610 = n179 & n3528 ;
  assign n21611 = n21610 ^ n2159 ^ 1'b0 ;
  assign n21612 = n6037 | n21611 ;
  assign n21613 = ( x114 & ~n10148 ) | ( x114 & n15229 ) | ( ~n10148 & n15229 ) ;
  assign n21614 = ~n3350 & n5193 ;
  assign n21615 = n4125 ^ n2396 ^ 1'b0 ;
  assign n21616 = n674 & ~n21615 ;
  assign n21617 = n21616 ^ n14049 ^ 1'b0 ;
  assign n21618 = ( n11241 & n21614 ) | ( n11241 & n21617 ) | ( n21614 & n21617 ) ;
  assign n21619 = ~n12465 & n13070 ;
  assign n21620 = ~n10363 & n21619 ;
  assign n21621 = n5524 & ~n8299 ;
  assign n21622 = n3095 | n3995 ;
  assign n21623 = n21621 | n21622 ;
  assign n21624 = n6327 | n12640 ;
  assign n21625 = n21623 | n21624 ;
  assign n21626 = ~n5923 & n21625 ;
  assign n21627 = ( n1898 & n19419 ) | ( n1898 & n21261 ) | ( n19419 & n21261 ) ;
  assign n21628 = n6050 & n9015 ;
  assign n21629 = n21628 ^ n6002 ^ 1'b0 ;
  assign n21630 = n676 & n21629 ;
  assign n21631 = ~n21627 & n21630 ;
  assign n21632 = n15429 ^ n5389 ^ 1'b0 ;
  assign n21633 = ~n9624 & n12367 ;
  assign n21634 = n1899 & n6147 ;
  assign n21635 = n5062 & n17838 ;
  assign n21636 = n21635 ^ n19934 ^ n6763 ;
  assign n21637 = ~n1907 & n20885 ;
  assign n21638 = ~n16289 & n21637 ;
  assign n21639 = n21203 ^ n3452 ^ 1'b0 ;
  assign n21640 = ( n2787 & ~n12499 ) | ( n2787 & n14825 ) | ( ~n12499 & n14825 ) ;
  assign n21641 = n21640 ^ n3279 ^ 1'b0 ;
  assign n21642 = ~n18869 & n21641 ;
  assign n21643 = ~n6817 & n13761 ;
  assign n21644 = n9990 & n21643 ;
  assign n21645 = n1536 & ~n5548 ;
  assign n21646 = n1421 & n21645 ;
  assign n21647 = n21646 ^ n5846 ^ 1'b0 ;
  assign n21648 = n1710 & ~n21647 ;
  assign n21649 = n2333 | n3542 ;
  assign n21650 = n2916 & ~n21649 ;
  assign n21651 = ~n10564 & n21650 ;
  assign n21652 = n21651 ^ n3964 ^ 1'b0 ;
  assign n21653 = n21648 & ~n21652 ;
  assign n21654 = n11510 & n21653 ;
  assign n21655 = n7033 ^ n315 ^ 1'b0 ;
  assign n21656 = n17672 & ~n21655 ;
  assign n21657 = n18498 ^ n13937 ^ n11559 ;
  assign n21658 = n6337 & ~n6727 ;
  assign n21659 = n9911 | n10579 ;
  assign n21660 = ~n18871 & n21659 ;
  assign n21661 = n1790 & n7532 ;
  assign n21662 = n21661 ^ n17636 ^ 1'b0 ;
  assign n21663 = n10435 & n16186 ;
  assign n21664 = n21662 & n21663 ;
  assign n21665 = n18150 ^ n361 ^ 1'b0 ;
  assign n21666 = n21664 | n21665 ;
  assign n21667 = n6821 & ~n7367 ;
  assign n21668 = ~n11403 & n21667 ;
  assign n21669 = n13955 & ~n21668 ;
  assign n21670 = n21669 ^ n6362 ^ 1'b0 ;
  assign n21671 = n4782 & n6323 ;
  assign n21672 = ~n6933 & n21671 ;
  assign n21673 = n224 & n20460 ;
  assign n21674 = ~n16640 & n21673 ;
  assign n21675 = n1200 | n19229 ;
  assign n21676 = n21674 & ~n21675 ;
  assign n21677 = n21676 ^ n224 ^ 1'b0 ;
  assign n21678 = n12088 | n21677 ;
  assign n21679 = n21678 ^ n10087 ^ 1'b0 ;
  assign n21680 = ~n21672 & n21679 ;
  assign n21681 = ( ~n8555 & n11985 ) | ( ~n8555 & n12882 ) | ( n11985 & n12882 ) ;
  assign n21682 = n15516 | n21681 ;
  assign n21683 = n7524 | n21682 ;
  assign n21684 = n12999 ^ n9396 ^ 1'b0 ;
  assign n21685 = n14850 | n21684 ;
  assign n21686 = ~n2013 & n2481 ;
  assign n21687 = n21686 ^ n4314 ^ 1'b0 ;
  assign n21688 = n21687 ^ n15778 ^ 1'b0 ;
  assign n21689 = n585 | n19644 ;
  assign n21690 = n21689 ^ n4408 ^ n2302 ;
  assign n21691 = n5625 ^ n4235 ^ 1'b0 ;
  assign n21692 = n7274 & ~n21691 ;
  assign n21693 = n13341 & n21692 ;
  assign n21694 = n16570 ^ n1884 ^ 1'b0 ;
  assign n21695 = n21694 ^ n19538 ^ 1'b0 ;
  assign n21696 = ~n14540 & n14954 ;
  assign n21697 = n21696 ^ n5787 ^ 1'b0 ;
  assign n21698 = n21697 ^ n11191 ^ 1'b0 ;
  assign n21699 = n7057 & ~n21698 ;
  assign n21700 = n5654 & n6545 ;
  assign n21701 = n9064 ^ n1810 ^ 1'b0 ;
  assign n21702 = n10318 | n21701 ;
  assign n21703 = n16732 ^ n5720 ^ 1'b0 ;
  assign n21704 = n14901 | n21703 ;
  assign n21705 = n5000 | n6268 ;
  assign n21706 = ~n15527 & n21705 ;
  assign n21707 = n21706 ^ n3768 ^ 1'b0 ;
  assign n21708 = n6836 & ~n13373 ;
  assign n21709 = n21708 ^ n8927 ^ 1'b0 ;
  assign n21710 = ( n7692 & n9586 ) | ( n7692 & n21709 ) | ( n9586 & n21709 ) ;
  assign n21711 = n15341 ^ n2062 ^ 1'b0 ;
  assign n21712 = n13414 ^ n5031 ^ 1'b0 ;
  assign n21713 = n2566 & ~n21712 ;
  assign n21714 = n12812 | n14248 ;
  assign n21715 = n722 & ~n21714 ;
  assign n21716 = n677 & ~n6476 ;
  assign n21717 = n21716 ^ n7629 ^ 1'b0 ;
  assign n21718 = n16283 ^ n14957 ^ n13487 ;
  assign n21719 = ( ~n549 & n20143 ) | ( ~n549 & n21718 ) | ( n20143 & n21718 ) ;
  assign n21720 = x78 | n7207 ;
  assign n21721 = n376 & ~n6529 ;
  assign n21722 = ( n12549 & n21720 ) | ( n12549 & n21721 ) | ( n21720 & n21721 ) ;
  assign n21728 = n1532 & n1570 ;
  assign n21729 = ~n1532 & n21728 ;
  assign n21730 = x52 | n21729 ;
  assign n21723 = ~n5547 & n17413 ;
  assign n21724 = n5547 & n21723 ;
  assign n21725 = n3532 & n21724 ;
  assign n21726 = ~n7430 & n21725 ;
  assign n21727 = n7751 & n21726 ;
  assign n21731 = n21730 ^ n21727 ^ n9926 ;
  assign n21732 = n21731 ^ n18838 ^ 1'b0 ;
  assign n21734 = n4044 & ~n6943 ;
  assign n21733 = n7925 | n10106 ;
  assign n21735 = n21734 ^ n21733 ^ 1'b0 ;
  assign n21736 = n21476 ^ n3853 ^ 1'b0 ;
  assign n21737 = n21735 & n21736 ;
  assign n21738 = n14704 ^ n14280 ^ 1'b0 ;
  assign n21739 = n7925 & ~n11255 ;
  assign n21740 = n2603 & n21739 ;
  assign n21741 = n11647 | n18386 ;
  assign n21742 = ~n10298 & n16138 ;
  assign n21743 = n21742 ^ n11053 ^ 1'b0 ;
  assign n21744 = ~n11826 & n16298 ;
  assign n21745 = n13028 ^ n556 ^ 1'b0 ;
  assign n21746 = n9592 & n21745 ;
  assign n21747 = n15171 ^ n3399 ^ 1'b0 ;
  assign n21748 = n21746 & ~n21747 ;
  assign n21749 = n8909 ^ n753 ^ 1'b0 ;
  assign n21750 = n5445 & ~n21749 ;
  assign n21751 = ~n709 & n21750 ;
  assign n21752 = ~n21748 & n21751 ;
  assign n21753 = n1376 & n19112 ;
  assign n21754 = n10549 ^ n10529 ^ 1'b0 ;
  assign n21755 = n1632 & n14784 ;
  assign n21756 = n18458 ^ n11745 ^ 1'b0 ;
  assign n21757 = n853 & ~n1991 ;
  assign n21759 = n2462 | n2624 ;
  assign n21758 = ~n607 & n1966 ;
  assign n21760 = n21759 ^ n21758 ^ 1'b0 ;
  assign n21761 = ~n5273 & n21760 ;
  assign n21762 = n21761 ^ n1645 ^ 1'b0 ;
  assign n21763 = n1552 & n7941 ;
  assign n21764 = ~n9116 & n11859 ;
  assign n21765 = n21763 & n21764 ;
  assign n21766 = n18123 ^ n11998 ^ n1950 ;
  assign n21767 = n9429 ^ n2328 ^ 1'b0 ;
  assign n21768 = n4524 | n21767 ;
  assign n21769 = n1457 ^ n1219 ^ 1'b0 ;
  assign n21770 = ~n14507 & n21769 ;
  assign n21771 = n3761 | n21770 ;
  assign n21772 = ~n3757 & n18985 ;
  assign n21773 = ~n4728 & n21772 ;
  assign n21774 = n11154 ^ n7014 ^ 1'b0 ;
  assign n21775 = n2673 & n21774 ;
  assign n21776 = ~n855 & n21775 ;
  assign n21777 = n15614 & n21776 ;
  assign n21778 = n7525 & n21777 ;
  assign n21779 = n180 & n7164 ;
  assign n21780 = ( n2889 & n3511 ) | ( n2889 & n21779 ) | ( n3511 & n21779 ) ;
  assign n21781 = ( n2131 & ~n16712 ) | ( n2131 & n21780 ) | ( ~n16712 & n21780 ) ;
  assign n21782 = ~n10579 & n19162 ;
  assign n21783 = n6396 & ~n11110 ;
  assign n21784 = n21783 ^ n19887 ^ 1'b0 ;
  assign n21785 = n8247 ^ n156 ^ 1'b0 ;
  assign n21786 = ~n17384 & n21785 ;
  assign n21787 = n6138 & n21786 ;
  assign n21788 = n21787 ^ n10712 ^ 1'b0 ;
  assign n21789 = n21788 ^ n4746 ^ n2709 ;
  assign n21790 = ~n16054 & n21789 ;
  assign n21791 = n20047 ^ n17955 ^ 1'b0 ;
  assign n21792 = n12948 ^ n1463 ^ 1'b0 ;
  assign n21793 = n13564 ^ n7137 ^ 1'b0 ;
  assign n21794 = n8552 | n21793 ;
  assign n21795 = n11538 & n21794 ;
  assign n21796 = n2783 | n10318 ;
  assign n21797 = n1555 & ~n2322 ;
  assign n21798 = n7571 & ~n19145 ;
  assign n21799 = n6891 & n12347 ;
  assign n21800 = ( n1836 & n2389 ) | ( n1836 & ~n4069 ) | ( n2389 & ~n4069 ) ;
  assign n21801 = n21800 ^ n20137 ^ 1'b0 ;
  assign n21802 = n1242 & n21801 ;
  assign n21803 = n560 | n8219 ;
  assign n21804 = n8931 | n10295 ;
  assign n21805 = n21804 ^ n4152 ^ 1'b0 ;
  assign n21806 = n16731 ^ n1939 ^ 1'b0 ;
  assign n21807 = n8703 & ~n21806 ;
  assign n21808 = n11649 ^ n1867 ^ n1785 ;
  assign n21809 = n791 & n6148 ;
  assign n21810 = n17186 ^ n9077 ^ 1'b0 ;
  assign n21811 = n4723 & ~n17549 ;
  assign n21812 = n7341 & ~n19017 ;
  assign n21813 = ~n5381 & n21812 ;
  assign n21814 = ( n308 & n3641 ) | ( n308 & n5678 ) | ( n3641 & n5678 ) ;
  assign n21815 = n21814 ^ n21143 ^ n587 ;
  assign n21816 = n3217 & n4906 ;
  assign n21817 = n21816 ^ n6440 ^ 1'b0 ;
  assign n21818 = n3757 ^ x21 ^ 1'b0 ;
  assign n21819 = n10602 ^ n1997 ^ 1'b0 ;
  assign n21820 = ~n7778 & n21819 ;
  assign n21821 = n11054 ^ n10530 ^ 1'b0 ;
  assign n21822 = n210 & ~n12887 ;
  assign n21823 = n14313 & n21822 ;
  assign n21824 = n12195 ^ n10861 ^ n8460 ;
  assign n21825 = ( n5576 & ~n7781 ) | ( n5576 & n21824 ) | ( ~n7781 & n21824 ) ;
  assign n21826 = n6875 ^ n5100 ^ 1'b0 ;
  assign n21827 = n3558 | n21826 ;
  assign n21828 = n21827 ^ n6943 ^ n6398 ;
  assign n21829 = n4151 | n4657 ;
  assign n21830 = n2718 & ~n21829 ;
  assign n21831 = n11320 ^ n881 ^ 1'b0 ;
  assign n21832 = n21830 | n21831 ;
  assign n21833 = n6421 & n21832 ;
  assign n21834 = n3572 & n20557 ;
  assign n21835 = ( ~x29 & n1545 ) | ( ~x29 & n10840 ) | ( n1545 & n10840 ) ;
  assign n21836 = n258 & n3404 ;
  assign n21837 = n227 & n18867 ;
  assign n21838 = n11753 & n21837 ;
  assign n21839 = n17581 & n17768 ;
  assign n21840 = n1686 | n1909 ;
  assign n21841 = n21840 ^ n20423 ^ 1'b0 ;
  assign n21842 = n8092 | n8854 ;
  assign n21843 = n21842 ^ n1922 ^ 1'b0 ;
  assign n21844 = n17721 & n21843 ;
  assign n21845 = n8704 ^ n1237 ^ 1'b0 ;
  assign n21846 = n15755 ^ n11178 ^ 1'b0 ;
  assign n21847 = n2381 & ~n21846 ;
  assign n21848 = n17291 ^ n11861 ^ n8801 ;
  assign n21849 = ~n16428 & n21848 ;
  assign n21850 = n4583 ^ n634 ^ 1'b0 ;
  assign n21851 = n7871 & ~n9846 ;
  assign n21852 = x26 & ~n5109 ;
  assign n21853 = n21852 ^ n9568 ^ 1'b0 ;
  assign n21854 = ( ~n20315 & n21851 ) | ( ~n20315 & n21853 ) | ( n21851 & n21853 ) ;
  assign n21855 = ( n2222 & n4380 ) | ( n2222 & ~n4848 ) | ( n4380 & ~n4848 ) ;
  assign n21857 = n14505 ^ n2758 ^ 1'b0 ;
  assign n21856 = n6594 & ~n15213 ;
  assign n21858 = n21857 ^ n21856 ^ 1'b0 ;
  assign n21859 = n4237 & ~n4424 ;
  assign n21860 = n21859 ^ n14428 ^ 1'b0 ;
  assign n21861 = n6807 | n21860 ;
  assign n21862 = n2146 | n21861 ;
  assign n21863 = n5446 & n12614 ;
  assign n21864 = ~n1303 & n21863 ;
  assign n21865 = n9703 & ~n21864 ;
  assign n21866 = n12229 ^ n5240 ^ 1'b0 ;
  assign n21867 = n15430 ^ n10657 ^ n2463 ;
  assign n21868 = n13757 ^ x25 ^ 1'b0 ;
  assign n21869 = n3364 | n21868 ;
  assign n21870 = n7478 & ~n21869 ;
  assign n21871 = n2564 & n21870 ;
  assign n21872 = n10149 ^ n6101 ^ 1'b0 ;
  assign n21873 = n21872 ^ n12460 ^ n2953 ;
  assign n21874 = n21873 ^ n3595 ^ 1'b0 ;
  assign n21875 = n3194 | n10732 ;
  assign n21876 = n7160 & ~n21875 ;
  assign n21877 = ( n11474 & n13006 ) | ( n11474 & n16165 ) | ( n13006 & n16165 ) ;
  assign n21878 = n713 | n10024 ;
  assign n21879 = ( n3027 & ~n5837 ) | ( n3027 & n19263 ) | ( ~n5837 & n19263 ) ;
  assign n21882 = n1324 | n15237 ;
  assign n21883 = n21882 ^ n9570 ^ 1'b0 ;
  assign n21880 = n7373 ^ n1908 ^ 1'b0 ;
  assign n21881 = n8653 & n21880 ;
  assign n21884 = n21883 ^ n21881 ^ n529 ;
  assign n21885 = n20170 ^ n19731 ^ 1'b0 ;
  assign n21886 = ~x63 & n261 ;
  assign n21887 = n21886 ^ n10327 ^ n5834 ;
  assign n21888 = ( n5092 & ~n9790 ) | ( n5092 & n19661 ) | ( ~n9790 & n19661 ) ;
  assign n21889 = n8321 | n9265 ;
  assign n21890 = n8379 ^ n5715 ^ 1'b0 ;
  assign n21891 = ~n7637 & n21890 ;
  assign n21892 = n15009 | n17984 ;
  assign n21893 = n6661 & n8101 ;
  assign n21895 = n2626 & n7259 ;
  assign n21896 = ~n3224 & n21895 ;
  assign n21894 = n3851 | n20394 ;
  assign n21897 = n21896 ^ n21894 ^ 1'b0 ;
  assign n21898 = n5747 | n10971 ;
  assign n21899 = n342 | n21898 ;
  assign n21900 = n21899 ^ n8405 ^ 1'b0 ;
  assign n21901 = n21900 ^ n2389 ^ 1'b0 ;
  assign n21902 = n16053 ^ n5231 ^ 1'b0 ;
  assign n21903 = n17023 ^ n1838 ^ 1'b0 ;
  assign n21904 = n10426 & ~n15746 ;
  assign n21905 = n21904 ^ x37 ^ 1'b0 ;
  assign n21906 = n577 & ~n21905 ;
  assign n21907 = ( ~n4942 & n18026 ) | ( ~n4942 & n21906 ) | ( n18026 & n21906 ) ;
  assign n21908 = n3230 ^ n788 ^ 1'b0 ;
  assign n21909 = n2300 | n11000 ;
  assign n21910 = n21909 ^ n4085 ^ 1'b0 ;
  assign n21911 = n6131 & ~n10825 ;
  assign n21912 = n21911 ^ n9685 ^ 1'b0 ;
  assign n21913 = n888 & ~n5181 ;
  assign n21914 = ~n2476 & n21913 ;
  assign n21915 = n20794 & n21914 ;
  assign n21916 = n792 & ~n5020 ;
  assign n21917 = ~n6037 & n21916 ;
  assign n21918 = ~n11811 & n12549 ;
  assign n21919 = n9411 | n15388 ;
  assign n21920 = n21918 & ~n21919 ;
  assign n21921 = n7356 & ~n20989 ;
  assign n21922 = ~n12561 & n21396 ;
  assign n21923 = n3087 & n10487 ;
  assign n21924 = n21923 ^ n13109 ^ 1'b0 ;
  assign n21925 = n20046 & n21924 ;
  assign n21926 = n1510 | n19233 ;
  assign n21927 = n21926 ^ n11137 ^ 1'b0 ;
  assign n21928 = n8832 ^ n1654 ^ 1'b0 ;
  assign n21929 = n9988 & n21928 ;
  assign n21930 = x25 & n6323 ;
  assign n21931 = n10826 & n21930 ;
  assign n21932 = n9494 & ~n11292 ;
  assign n21933 = n21932 ^ n939 ^ 1'b0 ;
  assign n21934 = n7141 | n21933 ;
  assign n21935 = n7847 & ~n15103 ;
  assign n21936 = n21935 ^ n9446 ^ 1'b0 ;
  assign n21937 = n21934 | n21936 ;
  assign n21938 = n21937 ^ n6631 ^ 1'b0 ;
  assign n21939 = n6455 ^ n4710 ^ 1'b0 ;
  assign n21940 = n758 & ~n21939 ;
  assign n21941 = n789 & n21940 ;
  assign n21942 = n21941 ^ n13786 ^ 1'b0 ;
  assign n21943 = n1338 & n1766 ;
  assign n21944 = ~n1766 & n21943 ;
  assign n21945 = ~n1117 & n1361 ;
  assign n21946 = n21944 & n21945 ;
  assign n21947 = n1289 & n21946 ;
  assign n21948 = n21947 ^ n8509 ^ 1'b0 ;
  assign n21949 = ~n5757 & n21948 ;
  assign n21950 = n5757 & n21949 ;
  assign n21951 = ( n3401 & n11893 ) | ( n3401 & ~n21950 ) | ( n11893 & ~n21950 ) ;
  assign n21952 = n21951 ^ n2589 ^ n2319 ;
  assign n21958 = n21491 ^ n2433 ^ 1'b0 ;
  assign n21959 = n3295 ^ n2816 ^ 1'b0 ;
  assign n21960 = ~n21958 & n21959 ;
  assign n21956 = n21399 ^ n519 ^ 1'b0 ;
  assign n21957 = n3885 | n21956 ;
  assign n21954 = n5642 ^ n1172 ^ 1'b0 ;
  assign n21953 = ~n8627 & n11938 ;
  assign n21955 = n21954 ^ n21953 ^ 1'b0 ;
  assign n21961 = n21960 ^ n21957 ^ n21955 ;
  assign n21962 = n907 ^ n559 ^ 1'b0 ;
  assign n21963 = n11777 | n21962 ;
  assign n21964 = ( n3179 & ~n5040 ) | ( n3179 & n7815 ) | ( ~n5040 & n7815 ) ;
  assign n21965 = n21964 ^ n8812 ^ 1'b0 ;
  assign n21966 = n19877 & n21965 ;
  assign n21967 = ~n1884 & n21700 ;
  assign n21968 = n4759 & n5775 ;
  assign n21969 = n19775 ^ n11845 ^ 1'b0 ;
  assign n21970 = ~n4897 & n11253 ;
  assign n21971 = n21877 & n21970 ;
  assign n21972 = n440 | n1793 ;
  assign n21973 = n4798 & ~n11246 ;
  assign n21974 = n17301 ^ n12593 ^ 1'b0 ;
  assign n21975 = n384 | n1505 ;
  assign n21976 = n5374 & n21975 ;
  assign n21977 = n17650 ^ n4177 ^ 1'b0 ;
  assign n21978 = n7057 & ~n21977 ;
  assign n21979 = n11284 | n11917 ;
  assign n21980 = ( n9754 & n21578 ) | ( n9754 & ~n21979 ) | ( n21578 & ~n21979 ) ;
  assign n21981 = n8470 | n10987 ;
  assign n21982 = n21981 ^ n6094 ^ 1'b0 ;
  assign n21983 = n3517 ^ n2198 ^ 1'b0 ;
  assign n21984 = n20561 ^ n4611 ^ 1'b0 ;
  assign n21985 = n21983 & n21984 ;
  assign n21986 = n3190 & n14770 ;
  assign n21988 = ~n5652 & n10301 ;
  assign n21987 = ~n6787 & n11293 ;
  assign n21989 = n21988 ^ n21987 ^ 1'b0 ;
  assign n21990 = ~n8472 & n19718 ;
  assign n21991 = n4784 & ~n15566 ;
  assign n21992 = n215 & n21991 ;
  assign n21993 = n1588 | n12555 ;
  assign n21994 = n21993 ^ n1438 ^ 1'b0 ;
  assign n21995 = n21994 ^ n16573 ^ n15873 ;
  assign n21996 = n437 & ~n13241 ;
  assign n21997 = ~n1481 & n4514 ;
  assign n21998 = n21997 ^ n525 ^ 1'b0 ;
  assign n21999 = n5965 & ~n14418 ;
  assign n22000 = n4119 ^ n616 ^ 1'b0 ;
  assign n22001 = ~n21999 & n22000 ;
  assign n22002 = n22001 ^ n10728 ^ n6158 ;
  assign n22003 = n1823 & n21325 ;
  assign n22004 = ~n20368 & n22003 ;
  assign n22005 = n157 & n11598 ;
  assign n22006 = n5094 & n22005 ;
  assign n22007 = n2899 & n22006 ;
  assign n22008 = n22007 ^ n17746 ^ 1'b0 ;
  assign n22009 = ~n9590 & n9802 ;
  assign n22010 = n22009 ^ n9940 ^ 1'b0 ;
  assign n22011 = n8398 | n16626 ;
  assign n22012 = n22011 ^ n2217 ^ 1'b0 ;
  assign n22013 = n17266 ^ n12547 ^ n879 ;
  assign n22014 = n22013 ^ n12391 ^ 1'b0 ;
  assign n22015 = n2931 | n14937 ;
  assign n22016 = n14495 | n22015 ;
  assign n22017 = n22016 ^ n456 ^ 1'b0 ;
  assign n22018 = ~n10889 & n12695 ;
  assign n22019 = n22018 ^ n896 ^ 1'b0 ;
  assign n22020 = ~n7439 & n17019 ;
  assign n22021 = ~n1473 & n22020 ;
  assign n22022 = n3124 & n8943 ;
  assign n22023 = n15327 | n22022 ;
  assign n22024 = n829 & ~n15612 ;
  assign n22025 = n22023 & n22024 ;
  assign n22026 = n4434 | n9846 ;
  assign n22027 = n11279 & ~n22026 ;
  assign n22028 = n17085 ^ n10787 ^ 1'b0 ;
  assign n22029 = n15352 ^ n4398 ^ 1'b0 ;
  assign n22032 = n4123 & ~n9481 ;
  assign n22033 = n14561 | n22032 ;
  assign n22030 = n9476 & ~n13802 ;
  assign n22031 = ~n5508 & n22030 ;
  assign n22034 = n22033 ^ n22031 ^ 1'b0 ;
  assign n22035 = n19131 & ~n19567 ;
  assign n22036 = n22035 ^ n7654 ^ 1'b0 ;
  assign n22037 = n1931 & ~n5206 ;
  assign n22038 = ~n12493 & n22037 ;
  assign n22039 = n8705 & n11537 ;
  assign n22040 = n1461 & ~n5244 ;
  assign n22041 = ~n12747 & n22040 ;
  assign n22042 = n22041 ^ n8946 ^ 1'b0 ;
  assign n22043 = n11107 | n15876 ;
  assign n22044 = n9608 & ~n14190 ;
  assign n22045 = n21286 ^ n20727 ^ 1'b0 ;
  assign n22046 = ~n18222 & n19532 ;
  assign n22047 = n1726 ^ n1361 ^ 1'b0 ;
  assign n22048 = n15290 ^ n4009 ^ 1'b0 ;
  assign n22049 = ~n22047 & n22048 ;
  assign n22050 = n10087 ^ n6124 ^ 1'b0 ;
  assign n22051 = n12071 | n22050 ;
  assign n22052 = n13877 ^ n5642 ^ 1'b0 ;
  assign n22053 = x108 & ~n22052 ;
  assign n22054 = n15854 & ~n21587 ;
  assign n22055 = n1491 & n6167 ;
  assign n22056 = ~n12027 & n22055 ;
  assign n22057 = n3274 & ~n22056 ;
  assign n22058 = n22057 ^ n3313 ^ 1'b0 ;
  assign n22059 = ~n7282 & n16411 ;
  assign n22060 = n22059 ^ n1981 ^ 1'b0 ;
  assign n22061 = n2412 | n15563 ;
  assign n22063 = n14446 & ~n18782 ;
  assign n22064 = n4290 & n22063 ;
  assign n22062 = n10715 | n13689 ;
  assign n22065 = n22064 ^ n22062 ^ 1'b0 ;
  assign n22066 = ~n13252 & n19062 ;
  assign n22067 = n9023 | n16479 ;
  assign n22068 = n18818 ^ n9847 ^ 1'b0 ;
  assign n22069 = n10612 ^ n4310 ^ 1'b0 ;
  assign n22070 = n1534 | n2328 ;
  assign n22071 = n4575 | n22070 ;
  assign n22072 = ( n302 & ~n1685 ) | ( n302 & n22071 ) | ( ~n1685 & n22071 ) ;
  assign n22073 = n1143 & n14256 ;
  assign n22074 = n9245 & n17120 ;
  assign n22075 = ~n22073 & n22074 ;
  assign n22076 = ~n3295 & n6006 ;
  assign n22077 = n22076 ^ n11732 ^ 1'b0 ;
  assign n22078 = n22077 ^ n12140 ^ 1'b0 ;
  assign n22080 = n17224 & n19322 ;
  assign n22079 = n16934 | n18847 ;
  assign n22081 = n22080 ^ n22079 ^ 1'b0 ;
  assign n22082 = n581 & n19244 ;
  assign n22083 = n4759 & ~n4944 ;
  assign n22084 = n22083 ^ n4405 ^ 1'b0 ;
  assign n22085 = n10398 ^ n2080 ^ 1'b0 ;
  assign n22086 = n20458 & n22085 ;
  assign n22087 = ( n8170 & n11511 ) | ( n8170 & ~n17405 ) | ( n11511 & ~n17405 ) ;
  assign n22088 = n22086 & ~n22087 ;
  assign n22089 = n5052 ^ n3025 ^ n1169 ;
  assign n22090 = n1680 & ~n10885 ;
  assign n22091 = n3925 & n4575 ;
  assign n22092 = n13257 ^ n4619 ^ 1'b0 ;
  assign n22093 = n6366 & ~n14319 ;
  assign n22094 = n8746 ^ n5836 ^ 1'b0 ;
  assign n22095 = n16234 & n22094 ;
  assign n22096 = n22095 ^ n12420 ^ 1'b0 ;
  assign n22097 = n901 | n15260 ;
  assign n22098 = ( ~n4373 & n16853 ) | ( ~n4373 & n22097 ) | ( n16853 & n22097 ) ;
  assign n22099 = ~n881 & n21888 ;
  assign n22100 = n22099 ^ n4186 ^ 1'b0 ;
  assign n22101 = ~n5351 & n14838 ;
  assign n22102 = x57 & n1334 ;
  assign n22103 = n22101 & n22102 ;
  assign n22104 = n14446 | n22103 ;
  assign n22105 = n1444 & n2494 ;
  assign n22106 = n22105 ^ n5692 ^ 1'b0 ;
  assign n22107 = x38 & ~n5009 ;
  assign n22108 = n22106 & n22107 ;
  assign n22109 = n9061 ^ n8343 ^ 1'b0 ;
  assign n22110 = n9258 | n22109 ;
  assign n22111 = n2227 ^ n1774 ^ 1'b0 ;
  assign n22112 = n4259 & ~n7075 ;
  assign n22113 = n5930 ^ n5796 ^ 1'b0 ;
  assign n22114 = n7054 & ~n22113 ;
  assign n22115 = n4204 & n22114 ;
  assign n22116 = n22115 ^ n6716 ^ 1'b0 ;
  assign n22117 = n14230 ^ n5810 ^ 1'b0 ;
  assign n22118 = ~n22116 & n22117 ;
  assign n22119 = n6940 | n12915 ;
  assign n22120 = n21544 & ~n22119 ;
  assign n22125 = n8418 ^ n3737 ^ 1'b0 ;
  assign n22121 = n6090 & n16564 ;
  assign n22122 = n22121 ^ n6279 ^ 1'b0 ;
  assign n22123 = n2198 | n22122 ;
  assign n22124 = ~n14099 & n22123 ;
  assign n22126 = n22125 ^ n22124 ^ 1'b0 ;
  assign n22127 = n22126 ^ n13223 ^ 1'b0 ;
  assign n22128 = n12087 ^ n10072 ^ 1'b0 ;
  assign n22129 = n1597 & n14331 ;
  assign n22130 = n19565 ^ n11458 ^ 1'b0 ;
  assign n22131 = n5497 | n17288 ;
  assign n22132 = n13589 | n18208 ;
  assign n22133 = n22132 ^ n9116 ^ 1'b0 ;
  assign n22134 = n13455 & ~n22133 ;
  assign n22135 = n3489 & n22134 ;
  assign n22136 = n8496 ^ n6759 ^ n4132 ;
  assign n22137 = n10956 | n11768 ;
  assign n22138 = n22137 ^ n4482 ^ 1'b0 ;
  assign n22139 = ~n344 & n17850 ;
  assign n22140 = n6261 & n22139 ;
  assign n22141 = n22140 ^ n732 ^ 1'b0 ;
  assign n22142 = n16887 ^ n13249 ^ n7291 ;
  assign n22143 = n13057 & ~n18799 ;
  assign n22144 = ~n892 & n22143 ;
  assign n22145 = n3770 & n8965 ;
  assign n22146 = n1495 & n22145 ;
  assign n22147 = n4377 ^ n2142 ^ 1'b0 ;
  assign n22148 = ~n12889 & n22147 ;
  assign n22149 = n18259 & n22148 ;
  assign n22150 = ~n13907 & n22149 ;
  assign n22151 = n4798 & n11732 ;
  assign n22152 = n8071 | n22151 ;
  assign n22153 = n22152 ^ n4104 ^ 1'b0 ;
  assign n22156 = ~n1579 & n2334 ;
  assign n22157 = n841 & n22156 ;
  assign n22158 = n2805 & ~n22157 ;
  assign n22159 = n22158 ^ n16824 ^ 1'b0 ;
  assign n22160 = ( n13298 & n19869 ) | ( n13298 & ~n22159 ) | ( n19869 & ~n22159 ) ;
  assign n22154 = ~n8033 & n18043 ;
  assign n22155 = n1503 & n22154 ;
  assign n22161 = n22160 ^ n22155 ^ 1'b0 ;
  assign n22162 = ~n531 & n6720 ;
  assign n22163 = n13910 ^ n903 ^ 1'b0 ;
  assign n22164 = n17056 & ~n22163 ;
  assign n22165 = n9105 ^ n4793 ^ 1'b0 ;
  assign n22166 = n6759 | n22165 ;
  assign n22167 = ~n2036 & n2249 ;
  assign n22168 = n22167 ^ n1219 ^ 1'b0 ;
  assign n22169 = n8926 & n15729 ;
  assign n22170 = n21280 & n22169 ;
  assign n22171 = n10778 ^ n2341 ^ n1114 ;
  assign n22172 = n14150 & n17615 ;
  assign n22173 = n22172 ^ n4947 ^ 1'b0 ;
  assign n22174 = n14014 ^ n3873 ^ 1'b0 ;
  assign n22175 = n14072 ^ n2637 ^ 1'b0 ;
  assign n22176 = ~n22174 & n22175 ;
  assign n22177 = n9009 & n22176 ;
  assign n22178 = n22177 ^ x6 ^ 1'b0 ;
  assign n22179 = n5954 & ~n12783 ;
  assign n22180 = n22179 ^ n3920 ^ 1'b0 ;
  assign n22181 = n4976 ^ n548 ^ x95 ;
  assign n22182 = ~n1315 & n21171 ;
  assign n22183 = n22181 & n22182 ;
  assign n22184 = n13924 ^ n2268 ^ 1'b0 ;
  assign n22185 = n10275 | n22184 ;
  assign n22186 = n11293 | n22185 ;
  assign n22188 = n11555 ^ n7755 ^ 1'b0 ;
  assign n22187 = n8158 | n9573 ;
  assign n22189 = n22188 ^ n22187 ^ 1'b0 ;
  assign n22190 = n1756 | n8292 ;
  assign n22191 = n8292 & ~n22190 ;
  assign n22192 = n630 | n10526 ;
  assign n22193 = n630 & ~n22192 ;
  assign n22194 = n3497 | n22193 ;
  assign n22195 = n22193 & ~n22194 ;
  assign n22196 = n3431 ^ n1419 ^ 1'b0 ;
  assign n22197 = n12758 | n22196 ;
  assign n22198 = n12758 & ~n22197 ;
  assign n22199 = n22195 | n22198 ;
  assign n22200 = n22191 & ~n22199 ;
  assign n22201 = n7512 & n12593 ;
  assign n22202 = n22200 & n22201 ;
  assign n22203 = ~n1659 & n8854 ;
  assign n22204 = n22203 ^ n12046 ^ 1'b0 ;
  assign n22205 = n6020 & ~n22204 ;
  assign n22206 = n22205 ^ n1592 ^ 1'b0 ;
  assign n22207 = ~n4316 & n19205 ;
  assign n22208 = ~n5154 & n22207 ;
  assign n22209 = n22208 ^ n14954 ^ 1'b0 ;
  assign n22210 = n22209 ^ n9971 ^ n5129 ;
  assign n22211 = n12583 ^ n10370 ^ 1'b0 ;
  assign n22212 = n2176 & ~n22211 ;
  assign n22213 = n3022 & ~n18295 ;
  assign n22214 = n22213 ^ n6013 ^ 1'b0 ;
  assign n22215 = n10934 & ~n22214 ;
  assign n22216 = n22215 ^ n4797 ^ 1'b0 ;
  assign n22217 = n16824 ^ n11770 ^ 1'b0 ;
  assign n22218 = n6244 & n22217 ;
  assign n22219 = n14002 ^ n651 ^ 1'b0 ;
  assign n22220 = ~n18154 & n22219 ;
  assign n22221 = n21996 & ~n22220 ;
  assign n22222 = n3450 & ~n9476 ;
  assign n22223 = ~n3595 & n22222 ;
  assign n22224 = n13976 ^ n243 ^ 1'b0 ;
  assign n22225 = n3481 | n22224 ;
  assign n22226 = n19291 & ~n22225 ;
  assign n22227 = n22223 & n22226 ;
  assign n22228 = n13179 | n15065 ;
  assign n22229 = ( n17337 & n17457 ) | ( n17337 & n22228 ) | ( n17457 & n22228 ) ;
  assign n22230 = x46 & n6046 ;
  assign n22231 = n5713 & n22230 ;
  assign n22232 = n6171 & ~n8503 ;
  assign n22233 = n22232 ^ n2448 ^ 1'b0 ;
  assign n22234 = n11775 & n22233 ;
  assign n22235 = n4150 | n22234 ;
  assign n22236 = ( n3289 & n22231 ) | ( n3289 & n22235 ) | ( n22231 & n22235 ) ;
  assign n22237 = n5220 ^ n4496 ^ n680 ;
  assign n22238 = n22237 ^ n1543 ^ 1'b0 ;
  assign n22239 = n2093 | n22238 ;
  assign n22240 = ( n950 & n5410 ) | ( n950 & ~n22239 ) | ( n5410 & ~n22239 ) ;
  assign n22241 = n9141 & n22240 ;
  assign n22242 = x32 & ~n986 ;
  assign n22243 = n12900 ^ n4118 ^ 1'b0 ;
  assign n22244 = n3122 & n13013 ;
  assign n22245 = n22244 ^ n9004 ^ 1'b0 ;
  assign n22246 = n2298 & n8996 ;
  assign n22247 = n22246 ^ n7362 ^ 1'b0 ;
  assign n22248 = n13031 & n13666 ;
  assign n22249 = ~n22247 & n22248 ;
  assign n22250 = n14279 ^ n8232 ^ 1'b0 ;
  assign n22251 = n7154 ^ n922 ^ 1'b0 ;
  assign n22252 = n4066 | n22251 ;
  assign n22253 = n5741 | n22252 ;
  assign n22254 = ~n22250 & n22253 ;
  assign n22255 = n12797 ^ n3666 ^ 1'b0 ;
  assign n22259 = n5274 ^ n1881 ^ 1'b0 ;
  assign n22256 = n3530 | n19519 ;
  assign n22257 = n437 | n22256 ;
  assign n22258 = ~n3214 & n22257 ;
  assign n22260 = n22259 ^ n22258 ^ 1'b0 ;
  assign n22261 = n3343 ^ n897 ^ 1'b0 ;
  assign n22262 = n1393 | n21088 ;
  assign n22263 = n2043 & ~n22262 ;
  assign n22264 = n5176 ^ n4352 ^ 1'b0 ;
  assign n22265 = n6416 | n22264 ;
  assign n22266 = n22265 ^ n12716 ^ n357 ;
  assign n22267 = ~n14553 & n22266 ;
  assign n22268 = n3287 ^ n1816 ^ 1'b0 ;
  assign n22269 = n22268 ^ n14702 ^ n1615 ;
  assign n22270 = n13340 ^ n5652 ^ 1'b0 ;
  assign n22271 = n9657 & ~n22270 ;
  assign n22272 = n294 & n12627 ;
  assign n22273 = n11518 ^ n9412 ^ 1'b0 ;
  assign n22274 = ( n9460 & n12880 ) | ( n9460 & ~n19198 ) | ( n12880 & ~n19198 ) ;
  assign n22275 = ( ~n6631 & n14187 ) | ( ~n6631 & n20413 ) | ( n14187 & n20413 ) ;
  assign n22276 = n21930 ^ n2501 ^ 1'b0 ;
  assign n22277 = ~n3264 & n4903 ;
  assign n22278 = n8948 & n21050 ;
  assign n22279 = x109 & n3058 ;
  assign n22280 = n22279 ^ n10301 ^ 1'b0 ;
  assign n22281 = n4861 & ~n22280 ;
  assign n22282 = n22281 ^ n10310 ^ 1'b0 ;
  assign n22283 = n19050 ^ n3620 ^ 1'b0 ;
  assign n22284 = n19844 & n22283 ;
  assign n22285 = ~n1378 & n5191 ;
  assign n22286 = ~n3135 & n22285 ;
  assign n22287 = n3974 & ~n22286 ;
  assign n22288 = n17835 & n22287 ;
  assign n22289 = n2771 ^ n2763 ^ 1'b0 ;
  assign n22290 = n1956 | n4506 ;
  assign n22291 = n22290 ^ n16150 ^ 1'b0 ;
  assign n22292 = n12315 & n18256 ;
  assign n22293 = n14554 & n19230 ;
  assign n22294 = ~n2513 & n22293 ;
  assign n22296 = n19464 ^ n1128 ^ 1'b0 ;
  assign n22297 = n397 & ~n22296 ;
  assign n22295 = n5820 & ~n9154 ;
  assign n22298 = n22297 ^ n22295 ^ 1'b0 ;
  assign n22299 = n1586 | n8301 ;
  assign n22300 = n21676 & ~n22299 ;
  assign n22301 = ~n5735 & n16359 ;
  assign n22302 = n22301 ^ n6116 ^ 1'b0 ;
  assign n22303 = ~n1128 & n15807 ;
  assign n22304 = n1275 ^ n152 ^ 1'b0 ;
  assign n22305 = ~n224 & n22304 ;
  assign n22306 = n22305 ^ n13992 ^ 1'b0 ;
  assign n22307 = n22306 ^ n1092 ^ 1'b0 ;
  assign n22308 = n5265 | n17306 ;
  assign n22309 = n5640 ^ n2228 ^ 1'b0 ;
  assign n22310 = n22308 & n22309 ;
  assign n22311 = x68 & n13377 ;
  assign n22312 = n19390 & n22311 ;
  assign n22313 = n892 | n22312 ;
  assign n22314 = n8403 & n16885 ;
  assign n22315 = n17792 ^ n11065 ^ n2090 ;
  assign n22316 = n4345 | n22315 ;
  assign n22317 = n22314 | n22316 ;
  assign n22318 = ~n3795 & n6347 ;
  assign n22319 = n22318 ^ n8176 ^ 1'b0 ;
  assign n22320 = n2090 & ~n10318 ;
  assign n22321 = n22320 ^ n22231 ^ 1'b0 ;
  assign n22322 = n13999 & n22321 ;
  assign n22323 = n3145 & n13368 ;
  assign n22324 = n10312 ^ n7274 ^ 1'b0 ;
  assign n22325 = ~n6354 & n22324 ;
  assign n22326 = ( ~x4 & n10564 ) | ( ~x4 & n22325 ) | ( n10564 & n22325 ) ;
  assign n22327 = ( n4738 & n7055 ) | ( n4738 & ~n12152 ) | ( n7055 & ~n12152 ) ;
  assign n22328 = ~n17465 & n21464 ;
  assign n22329 = n22328 ^ n14342 ^ 1'b0 ;
  assign n22330 = n814 & ~n11295 ;
  assign n22331 = n3025 & ~n21081 ;
  assign n22332 = ~n19838 & n22331 ;
  assign n22333 = n4605 ^ x71 ^ 1'b0 ;
  assign n22334 = n4794 | n22333 ;
  assign n22335 = ( n985 & ~n3987 ) | ( n985 & n22334 ) | ( ~n3987 & n22334 ) ;
  assign n22336 = n256 | n22335 ;
  assign n22337 = n22336 ^ n2556 ^ 1'b0 ;
  assign n22338 = ~n8476 & n22337 ;
  assign n22339 = n4481 & ~n22338 ;
  assign n22340 = ~n2810 & n4143 ;
  assign n22341 = n22340 ^ n10769 ^ 1'b0 ;
  assign n22342 = n7453 ^ n1635 ^ 1'b0 ;
  assign n22343 = n3897 | n22342 ;
  assign n22344 = n2234 | n5389 ;
  assign n22345 = n22344 ^ n2450 ^ 1'b0 ;
  assign n22346 = n468 & n22345 ;
  assign n22347 = n3649 & ~n10715 ;
  assign n22348 = n973 & ~n10019 ;
  assign n22349 = ~n12253 & n14229 ;
  assign n22350 = ~n4542 & n4836 ;
  assign n22351 = n9211 | n22350 ;
  assign n22352 = ~n468 & n4429 ;
  assign n22353 = n1656 & n8710 ;
  assign n22354 = n21734 ^ n16981 ^ 1'b0 ;
  assign n22355 = n16151 & ~n22354 ;
  assign n22356 = n2963 | n14657 ;
  assign n22357 = ( n1031 & n12969 ) | ( n1031 & n22356 ) | ( n12969 & n22356 ) ;
  assign n22358 = n11577 & ~n22357 ;
  assign n22359 = n6454 ^ n4973 ^ n4813 ;
  assign n22360 = n22359 ^ n10527 ^ n3550 ;
  assign n22361 = n14767 ^ x124 ^ 1'b0 ;
  assign n22362 = n7914 & n22361 ;
  assign n22363 = n11333 ^ n8993 ^ 1'b0 ;
  assign n22364 = n4058 | n11575 ;
  assign n22365 = ~n22363 & n22364 ;
  assign n22366 = n15423 ^ n12782 ^ 1'b0 ;
  assign n22369 = n18753 ^ n17476 ^ 1'b0 ;
  assign n22367 = n822 & n8101 ;
  assign n22368 = n13087 & n22367 ;
  assign n22370 = n22369 ^ n22368 ^ n16700 ;
  assign n22371 = n7453 & ~n14344 ;
  assign n22372 = n5281 & ~n6932 ;
  assign n22373 = ~n15240 & n22372 ;
  assign n22374 = n5145 & n13242 ;
  assign n22375 = n22374 ^ n15840 ^ 1'b0 ;
  assign n22376 = n7729 ^ n4262 ^ 1'b0 ;
  assign n22377 = ( ~n1745 & n2629 ) | ( ~n1745 & n3204 ) | ( n2629 & n3204 ) ;
  assign n22378 = n13343 ^ n3528 ^ 1'b0 ;
  assign n22379 = n5826 | n6882 ;
  assign n22380 = n14284 | n22379 ;
  assign n22381 = n8666 | n22380 ;
  assign n22382 = n7039 & ~n8322 ;
  assign n22383 = ~n14135 & n22382 ;
  assign n22384 = n22383 ^ n4292 ^ 1'b0 ;
  assign n22385 = n12349 & n22384 ;
  assign n22386 = n2228 & n15372 ;
  assign n22387 = ~n1124 & n22386 ;
  assign n22388 = n22387 ^ n12677 ^ 1'b0 ;
  assign n22389 = ~n13082 & n22388 ;
  assign n22390 = ~n209 & n2537 ;
  assign n22391 = n22390 ^ n6604 ^ 1'b0 ;
  assign n22392 = n16020 | n22391 ;
  assign n22393 = n22392 ^ n20178 ^ 1'b0 ;
  assign n22394 = n2476 | n22393 ;
  assign n22395 = n3162 | n10814 ;
  assign n22396 = n22394 & ~n22395 ;
  assign n22397 = ~n15814 & n17136 ;
  assign n22398 = n22397 ^ x102 ^ 1'b0 ;
  assign n22399 = ( n697 & ~n8343 ) | ( n697 & n12520 ) | ( ~n8343 & n12520 ) ;
  assign n22400 = n2330 ^ n2238 ^ n258 ;
  assign n22401 = ~n858 & n12813 ;
  assign n22402 = n22401 ^ n6080 ^ 1'b0 ;
  assign n22406 = ~n2809 & n6356 ;
  assign n22407 = ~n8520 & n22406 ;
  assign n22403 = ~n8317 & n21954 ;
  assign n22404 = n6686 | n14254 ;
  assign n22405 = ( n13080 & n22403 ) | ( n13080 & ~n22404 ) | ( n22403 & ~n22404 ) ;
  assign n22408 = n22407 ^ n22405 ^ 1'b0 ;
  assign n22409 = n7678 & ~n22408 ;
  assign n22410 = n17475 ^ n3424 ^ 1'b0 ;
  assign n22411 = n21786 & ~n22410 ;
  assign n22412 = n5297 & ~n9672 ;
  assign n22413 = n8829 & n22412 ;
  assign n22414 = n7874 ^ n7391 ^ 1'b0 ;
  assign n22415 = ~n22413 & n22414 ;
  assign n22416 = n11783 ^ n464 ^ 1'b0 ;
  assign n22417 = ( n645 & ~n749 ) | ( n645 & n1853 ) | ( ~n749 & n1853 ) ;
  assign n22418 = n4237 & n22417 ;
  assign n22419 = n19671 ^ n15148 ^ 1'b0 ;
  assign n22420 = n14908 ^ n4523 ^ 1'b0 ;
  assign n22421 = n4264 & ~n6101 ;
  assign n22422 = n22421 ^ n675 ^ n562 ;
  assign n22423 = n8405 | n22422 ;
  assign n22424 = n8710 | n22423 ;
  assign n22425 = n22424 ^ n12609 ^ 1'b0 ;
  assign n22426 = n18692 & n22425 ;
  assign n22427 = ( n12993 & ~n18400 ) | ( n12993 & n22334 ) | ( ~n18400 & n22334 ) ;
  assign n22428 = n2593 ^ n678 ^ n204 ;
  assign n22429 = ( n7053 & n12588 ) | ( n7053 & ~n22428 ) | ( n12588 & ~n22428 ) ;
  assign n22430 = n14777 ^ n6108 ^ n5088 ;
  assign n22431 = n1333 & ~n22430 ;
  assign n22432 = n22431 ^ n6009 ^ 1'b0 ;
  assign n22433 = n22116 ^ n18380 ^ 1'b0 ;
  assign n22434 = n9758 & ~n22433 ;
  assign n22435 = n15106 ^ n2665 ^ 1'b0 ;
  assign n22436 = n14995 & ~n22435 ;
  assign n22437 = ~n916 & n17244 ;
  assign n22438 = ~n22436 & n22437 ;
  assign n22439 = n21979 & ~n22438 ;
  assign n22440 = n11976 & ~n15920 ;
  assign n22441 = n11251 ^ n5967 ^ 1'b0 ;
  assign n22442 = n3142 | n22441 ;
  assign n22443 = n12076 | n22442 ;
  assign n22444 = n3231 & ~n7525 ;
  assign n22445 = n4874 & n22444 ;
  assign n22446 = n586 | n8006 ;
  assign n22447 = x34 & n22446 ;
  assign n22448 = ~n3552 & n22447 ;
  assign n22449 = ~n874 & n10053 ;
  assign n22450 = n2062 | n15645 ;
  assign n22451 = n22450 ^ n9604 ^ 1'b0 ;
  assign n22452 = n22449 & ~n22451 ;
  assign n22453 = n166 | n2085 ;
  assign n22454 = n7188 & ~n22453 ;
  assign n22455 = n14499 & n22454 ;
  assign n22456 = ~n468 & n3729 ;
  assign n22457 = n6675 & ~n22456 ;
  assign n22458 = n22457 ^ n21177 ^ n6626 ;
  assign n22459 = ~n1053 & n6090 ;
  assign n22460 = ~n6090 & n22459 ;
  assign n22461 = n21095 ^ n9994 ^ 1'b0 ;
  assign n22462 = ~n10644 & n22461 ;
  assign n22463 = n22460 & n22462 ;
  assign n22464 = n3745 ^ n2617 ^ 1'b0 ;
  assign n22465 = n22464 ^ n12677 ^ 1'b0 ;
  assign n22466 = n2331 & n22465 ;
  assign n22467 = n4055 & n22466 ;
  assign n22468 = n468 & n7746 ;
  assign n22469 = ~n468 & n22468 ;
  assign n22470 = ~n3842 & n4456 ;
  assign n22471 = n10544 & n22470 ;
  assign n22472 = n17476 | n22471 ;
  assign n22473 = n22471 & ~n22472 ;
  assign n22474 = ( n6218 & n22469 ) | ( n6218 & ~n22473 ) | ( n22469 & ~n22473 ) ;
  assign n22475 = ( n2131 & ~n20659 ) | ( n2131 & n22474 ) | ( ~n20659 & n22474 ) ;
  assign n22476 = ~n1115 & n2605 ;
  assign n22477 = n13648 & n22112 ;
  assign n22479 = ~n6049 & n7710 ;
  assign n22478 = n14592 | n18544 ;
  assign n22480 = n22479 ^ n22478 ^ 1'b0 ;
  assign n22482 = ~n7742 & n9071 ;
  assign n22481 = n5614 & ~n20613 ;
  assign n22483 = n22482 ^ n22481 ^ 1'b0 ;
  assign n22484 = ~n5836 & n22403 ;
  assign n22485 = n1083 | n7549 ;
  assign n22486 = n833 & n19493 ;
  assign n22487 = n22485 & n22486 ;
  assign n22488 = n12877 ^ n3601 ^ n657 ;
  assign n22489 = n22488 ^ n21610 ^ 1'b0 ;
  assign n22490 = ~n6392 & n15781 ;
  assign n22491 = n7851 & ~n22490 ;
  assign n22492 = ~n6958 & n22491 ;
  assign n22493 = n5423 & n6714 ;
  assign n22494 = n22493 ^ x24 ^ 1'b0 ;
  assign n22495 = n4389 & ~n22494 ;
  assign n22496 = n22495 ^ n4246 ^ 1'b0 ;
  assign n22497 = n6901 ^ n1633 ^ 1'b0 ;
  assign n22498 = n1601 & n5916 ;
  assign n22499 = n8602 & n22498 ;
  assign n22500 = ~n3481 & n15210 ;
  assign n22501 = n6094 & n22500 ;
  assign n22502 = n22501 ^ n5573 ^ 1'b0 ;
  assign n22504 = n476 & n21648 ;
  assign n22503 = n7548 | n10265 ;
  assign n22505 = n22504 ^ n22503 ^ 1'b0 ;
  assign n22506 = n22505 ^ n6071 ^ 1'b0 ;
  assign n22507 = n17206 ^ n2726 ^ 1'b0 ;
  assign n22508 = ~n13183 & n22507 ;
  assign n22509 = ~n1745 & n3729 ;
  assign n22510 = n22509 ^ n7688 ^ 1'b0 ;
  assign n22511 = n1124 & ~n22510 ;
  assign n22512 = n12554 ^ n2153 ^ 1'b0 ;
  assign n22513 = n2935 | n9703 ;
  assign n22514 = n22513 ^ n9026 ^ 1'b0 ;
  assign n22515 = ~n3510 & n22514 ;
  assign n22516 = n18265 ^ n4437 ^ 1'b0 ;
  assign n22517 = ~n6612 & n15995 ;
  assign n22519 = x56 & ~n12227 ;
  assign n22518 = n3287 & n14801 ;
  assign n22520 = n22519 ^ n22518 ^ 1'b0 ;
  assign n22521 = n5863 | n22407 ;
  assign n22522 = n11300 & ~n16252 ;
  assign n22523 = n13301 ^ n6497 ^ 1'b0 ;
  assign n22524 = n14341 & n20833 ;
  assign n22525 = ~n22523 & n22524 ;
  assign n22526 = n9862 ^ n2044 ^ 1'b0 ;
  assign n22527 = n10445 | n16317 ;
  assign n22528 = ( n5470 & n6169 ) | ( n5470 & ~n22527 ) | ( n6169 & ~n22527 ) ;
  assign n22529 = n6062 ^ n2176 ^ 1'b0 ;
  assign n22530 = n14994 ^ n14856 ^ 1'b0 ;
  assign n22531 = n4295 & ~n19280 ;
  assign n22532 = ( n5262 & n10039 ) | ( n5262 & ~n14159 ) | ( n10039 & ~n14159 ) ;
  assign n22533 = n22532 ^ n15948 ^ 1'b0 ;
  assign n22535 = ( n1001 & ~n21827 ) | ( n1001 & n22509 ) | ( ~n21827 & n22509 ) ;
  assign n22534 = n3694 & ~n6354 ;
  assign n22536 = n22535 ^ n22534 ^ 1'b0 ;
  assign n22537 = n7958 ^ n5996 ^ n2402 ;
  assign n22538 = n9471 & ~n22537 ;
  assign n22539 = n19078 ^ n7645 ^ 1'b0 ;
  assign n22540 = n1416 | n22539 ;
  assign n22541 = n20688 ^ n6411 ^ 1'b0 ;
  assign n22542 = n456 | n14828 ;
  assign n22543 = n1143 | n22542 ;
  assign n22544 = n6075 & ~n8992 ;
  assign n22545 = ~n2070 & n10416 ;
  assign n22546 = n6671 & n22545 ;
  assign n22547 = n2856 ^ n2684 ^ 1'b0 ;
  assign n22548 = n7219 | n22547 ;
  assign n22549 = n15757 ^ n9994 ^ 1'b0 ;
  assign n22550 = ~n14217 & n22549 ;
  assign n22551 = n2170 | n5249 ;
  assign n22552 = ~n2213 & n11617 ;
  assign n22553 = n22551 & n22552 ;
  assign n22554 = ~n6598 & n14786 ;
  assign n22555 = n10568 & n22554 ;
  assign n22556 = n10825 & n22555 ;
  assign n22557 = n22556 ^ n7253 ^ 1'b0 ;
  assign n22558 = n13869 ^ n11531 ^ 1'b0 ;
  assign n22559 = n1999 | n6279 ;
  assign n22560 = n4195 & ~n22559 ;
  assign n22563 = n7038 ^ n3811 ^ 1'b0 ;
  assign n22564 = n22563 ^ n10825 ^ 1'b0 ;
  assign n22565 = n7155 ^ n4315 ^ 1'b0 ;
  assign n22566 = n9868 & n22565 ;
  assign n22567 = n22566 ^ n5459 ^ 1'b0 ;
  assign n22568 = ( ~n3411 & n22564 ) | ( ~n3411 & n22567 ) | ( n22564 & n22567 ) ;
  assign n22561 = x69 & n22209 ;
  assign n22562 = ~n677 & n22561 ;
  assign n22569 = n22568 ^ n22562 ^ 1'b0 ;
  assign n22570 = n20172 ^ n3860 ^ n1641 ;
  assign n22571 = n14847 ^ n8063 ^ 1'b0 ;
  assign n22572 = n4665 & n22571 ;
  assign n22573 = ~n1531 & n5354 ;
  assign n22574 = n22573 ^ n3814 ^ 1'b0 ;
  assign n22575 = ( ~n1130 & n8185 ) | ( ~n1130 & n10053 ) | ( n8185 & n10053 ) ;
  assign n22576 = n13979 & ~n22575 ;
  assign n22582 = n2438 & n2892 ;
  assign n22583 = ~n11831 & n22582 ;
  assign n22577 = ~n2689 & n9046 ;
  assign n22578 = n22577 ^ n4077 ^ 1'b0 ;
  assign n22579 = ~n6432 & n22578 ;
  assign n22580 = n10013 ^ n366 ^ 1'b0 ;
  assign n22581 = n22579 & ~n22580 ;
  assign n22584 = n22583 ^ n22581 ^ n17228 ;
  assign n22585 = n1413 & ~n7157 ;
  assign n22586 = ~n7865 & n22585 ;
  assign n22587 = n22586 ^ n20069 ^ n851 ;
  assign n22588 = ( n543 & n1166 ) | ( n543 & ~n4159 ) | ( n1166 & ~n4159 ) ;
  assign n22589 = n13942 & n22588 ;
  assign n22590 = n22589 ^ n8702 ^ 1'b0 ;
  assign n22591 = n10070 | n22590 ;
  assign n22592 = n22591 ^ n8124 ^ 1'b0 ;
  assign n22593 = n357 | n534 ;
  assign n22594 = n3927 & ~n22593 ;
  assign n22595 = ~n4490 & n22594 ;
  assign n22596 = n14870 ^ n6591 ^ 1'b0 ;
  assign n22598 = n4555 & n4973 ;
  assign n22597 = ( n3938 & n4819 ) | ( n3938 & ~n9996 ) | ( n4819 & ~n9996 ) ;
  assign n22599 = n22598 ^ n22597 ^ 1'b0 ;
  assign n22600 = n5206 ^ n2418 ^ 1'b0 ;
  assign n22601 = n20334 ^ n2497 ^ n645 ;
  assign n22602 = n10905 | n22335 ;
  assign n22603 = n22602 ^ n14607 ^ 1'b0 ;
  assign n22604 = n22603 ^ n8770 ^ n2539 ;
  assign n22605 = n7125 | n22166 ;
  assign n22606 = n22605 ^ n4364 ^ 1'b0 ;
  assign n22607 = n853 & n21799 ;
  assign n22608 = ~n21746 & n22607 ;
  assign n22609 = n16364 & ~n17146 ;
  assign n22610 = n7105 & n8242 ;
  assign n22611 = n22610 ^ n5031 ^ 1'b0 ;
  assign n22612 = n331 & n5165 ;
  assign n22613 = n22612 ^ n9863 ^ 1'b0 ;
  assign n22614 = n8622 & n12716 ;
  assign n22615 = n3287 & ~n5958 ;
  assign n22616 = ~n5448 & n10193 ;
  assign n22617 = n287 | n13747 ;
  assign n22618 = n17489 | n22617 ;
  assign n22619 = n3140 & n19413 ;
  assign n22620 = ~n8752 & n22619 ;
  assign n22622 = n15347 ^ n6126 ^ 1'b0 ;
  assign n22623 = n3097 | n22622 ;
  assign n22621 = ~n8608 & n15971 ;
  assign n22624 = n22623 ^ n22621 ^ 1'b0 ;
  assign n22625 = n3006 & ~n17541 ;
  assign n22626 = n22625 ^ n17077 ^ x28 ;
  assign n22627 = n15334 ^ n12626 ^ n8679 ;
  assign n22628 = n5958 ^ n3226 ^ 1'b0 ;
  assign n22629 = n1897 & n22628 ;
  assign n22630 = n18438 ^ n16576 ^ 1'b0 ;
  assign n22631 = n3629 & ~n22630 ;
  assign n22632 = n3474 & n22631 ;
  assign n22633 = ~n22629 & n22632 ;
  assign n22634 = n10937 ^ n9202 ^ 1'b0 ;
  assign n22635 = n11000 ^ n540 ^ 1'b0 ;
  assign n22636 = n22635 ^ n3374 ^ 1'b0 ;
  assign n22637 = n4579 | n11609 ;
  assign n22638 = n22637 ^ n16458 ^ 1'b0 ;
  assign n22639 = n11231 & ~n14228 ;
  assign n22640 = n14001 | n17543 ;
  assign n22641 = n2179 & n4382 ;
  assign n22642 = n22641 ^ n143 ^ 1'b0 ;
  assign n22643 = n22642 ^ n6486 ^ 1'b0 ;
  assign n22644 = n3240 | n7881 ;
  assign n22645 = n1590 & n4923 ;
  assign n22646 = ~n2407 & n3530 ;
  assign n22647 = n20686 | n21545 ;
  assign n22648 = n22646 & ~n22647 ;
  assign n22649 = n11431 ^ n2892 ^ 1'b0 ;
  assign n22650 = n4440 & n22649 ;
  assign n22651 = n4963 | n22650 ;
  assign n22652 = ~n1077 & n14479 ;
  assign n22653 = n14813 ^ n1831 ^ 1'b0 ;
  assign n22658 = ~n854 & n1427 ;
  assign n22659 = ~n3839 & n22658 ;
  assign n22654 = n1457 ^ n301 ^ 1'b0 ;
  assign n22655 = n5986 | n22654 ;
  assign n22656 = n7673 | n9242 ;
  assign n22657 = n22655 & ~n22656 ;
  assign n22660 = n22659 ^ n22657 ^ 1'b0 ;
  assign n22661 = n22660 ^ n5457 ^ 1'b0 ;
  assign n22662 = n1778 | n22661 ;
  assign n22663 = ( n1402 & n22653 ) | ( n1402 & n22662 ) | ( n22653 & n22662 ) ;
  assign n22664 = n8284 ^ n1252 ^ 1'b0 ;
  assign n22665 = n5345 & n7048 ;
  assign n22666 = ~n22664 & n22665 ;
  assign n22667 = n16824 ^ x6 ^ 1'b0 ;
  assign n22668 = n16923 & ~n22667 ;
  assign n22669 = n5479 & ~n9831 ;
  assign n22670 = ~n8713 & n22669 ;
  assign n22671 = ~n7705 & n22670 ;
  assign n22672 = n22668 & ~n22671 ;
  assign n22673 = n19765 & n22672 ;
  assign n22674 = ~n5052 & n18227 ;
  assign n22675 = n6437 ^ n2667 ^ n1639 ;
  assign n22676 = n6938 | n22675 ;
  assign n22677 = n22674 | n22676 ;
  assign n22678 = n9084 ^ n5074 ^ n2290 ;
  assign n22679 = ( n377 & n1174 ) | ( n377 & n22678 ) | ( n1174 & n22678 ) ;
  assign n22680 = ( n6565 & n8284 ) | ( n6565 & n15684 ) | ( n8284 & n15684 ) ;
  assign n22681 = n7527 ^ n7105 ^ 1'b0 ;
  assign n22682 = n5274 & n16728 ;
  assign n22683 = n15384 & n22682 ;
  assign n22684 = n10896 & ~n22683 ;
  assign n22685 = ~n22681 & n22684 ;
  assign n22687 = n20458 ^ n250 ^ 1'b0 ;
  assign n22688 = n19999 | n22687 ;
  assign n22686 = ~n3336 & n17082 ;
  assign n22689 = n22688 ^ n22686 ^ 1'b0 ;
  assign n22690 = n8052 ^ n4456 ^ 1'b0 ;
  assign n22691 = ~n934 & n6504 ;
  assign n22692 = n489 | n5694 ;
  assign n22693 = n3115 & ~n22692 ;
  assign n22694 = n19614 & n22693 ;
  assign n22695 = n16222 ^ n1350 ^ 1'b0 ;
  assign n22697 = n3104 & ~n8418 ;
  assign n22696 = n2596 & n2802 ;
  assign n22698 = n22697 ^ n22696 ^ 1'b0 ;
  assign n22699 = ~n5792 & n16456 ;
  assign n22700 = n977 & n22699 ;
  assign n22701 = n11865 ^ n9009 ^ 1'b0 ;
  assign n22702 = n20224 | n22701 ;
  assign n22703 = n5580 | n11026 ;
  assign n22704 = n22703 ^ n2409 ^ 1'b0 ;
  assign n22705 = ~x75 & n22704 ;
  assign n22706 = ~n3595 & n22705 ;
  assign n22707 = n20853 | n22706 ;
  assign n22708 = n22707 ^ n18893 ^ 1'b0 ;
  assign n22709 = n7423 & ~n15623 ;
  assign n22710 = ~n7920 & n22709 ;
  assign n22711 = n22708 & n22710 ;
  assign n22712 = n4436 | n16312 ;
  assign n22713 = n22712 ^ n147 ^ 1'b0 ;
  assign n22714 = n22713 ^ n786 ^ n556 ;
  assign n22715 = n488 | n13004 ;
  assign n22716 = n15384 ^ n1327 ^ 1'b0 ;
  assign n22717 = n2103 & n22716 ;
  assign n22718 = n20749 ^ n13463 ^ 1'b0 ;
  assign n22719 = n835 | n22718 ;
  assign n22720 = n13326 ^ n4093 ^ n2445 ;
  assign n22721 = n22720 ^ n5669 ^ n5521 ;
  assign n22722 = x35 & ~n2167 ;
  assign n22723 = n10124 & n22722 ;
  assign n22724 = n875 | n13229 ;
  assign n22725 = n22723 & ~n22724 ;
  assign n22726 = n3072 | n19644 ;
  assign n22727 = ( n18236 & n22725 ) | ( n18236 & ~n22726 ) | ( n22725 & ~n22726 ) ;
  assign n22728 = n1681 & ~n2978 ;
  assign n22729 = n1115 & n22728 ;
  assign n22730 = n11891 ^ n2235 ^ 1'b0 ;
  assign n22731 = n3384 | n4759 ;
  assign n22732 = n22731 ^ n1426 ^ 1'b0 ;
  assign n22733 = n11036 | n16636 ;
  assign n22734 = n22732 | n22733 ;
  assign n22735 = n3062 & n21574 ;
  assign n22736 = n22735 ^ n5220 ^ 1'b0 ;
  assign n22737 = n8587 ^ n6358 ^ 1'b0 ;
  assign n22738 = n8448 & n22737 ;
  assign n22739 = n10782 & n22738 ;
  assign n22740 = n1311 & ~n16113 ;
  assign n22741 = ~n16667 & n22740 ;
  assign n22742 = n20281 | n22741 ;
  assign n22743 = ~n3741 & n17442 ;
  assign n22744 = n2917 & n22743 ;
  assign n22745 = n8859 ^ n2804 ^ 1'b0 ;
  assign n22746 = ~n541 & n2254 ;
  assign n22747 = n7389 | n22746 ;
  assign n22748 = n19717 ^ n697 ^ 1'b0 ;
  assign n22749 = n13207 ^ n4856 ^ 1'b0 ;
  assign n22750 = n20090 ^ n19203 ^ n15078 ;
  assign n22751 = n16141 ^ n15240 ^ 1'b0 ;
  assign n22752 = n14534 ^ n5992 ^ 1'b0 ;
  assign n22753 = ~n13343 & n14724 ;
  assign n22754 = n8167 | n11475 ;
  assign n22755 = n12345 & ~n22754 ;
  assign n22756 = ~n17745 & n22755 ;
  assign n22757 = n3290 | n9117 ;
  assign n22758 = n681 | n4268 ;
  assign n22759 = n22758 ^ n9904 ^ 1'b0 ;
  assign n22760 = ( n8888 & n14906 ) | ( n8888 & n15905 ) | ( n14906 & n15905 ) ;
  assign n22761 = ~n17527 & n22760 ;
  assign n22762 = n22761 ^ n5223 ^ 1'b0 ;
  assign n22763 = n10868 & n20723 ;
  assign n22764 = n3239 ^ n2718 ^ 1'b0 ;
  assign n22765 = n3605 ^ n362 ^ 1'b0 ;
  assign n22766 = n22764 & ~n22765 ;
  assign n22767 = n20860 ^ n4664 ^ 1'b0 ;
  assign n22768 = n6124 & ~n22767 ;
  assign n22769 = x83 & n13625 ;
  assign n22770 = n15843 ^ n462 ^ 1'b0 ;
  assign n22771 = n11267 ^ n2096 ^ 1'b0 ;
  assign n22772 = n398 | n22771 ;
  assign n22773 = n18480 ^ n17851 ^ 1'b0 ;
  assign n22774 = n8352 & n22773 ;
  assign n22775 = ~n9051 & n22774 ;
  assign n22776 = n22772 & n22775 ;
  assign n22777 = n2338 & ~n9481 ;
  assign n22778 = n22777 ^ n10248 ^ 1'b0 ;
  assign n22779 = n3859 & n9888 ;
  assign n22780 = n5644 & ~n5711 ;
  assign n22781 = n12464 | n22780 ;
  assign n22782 = ( n2763 & ~n3899 ) | ( n2763 & n22456 ) | ( ~n3899 & n22456 ) ;
  assign n22783 = ( ~n5634 & n22781 ) | ( ~n5634 & n22782 ) | ( n22781 & n22782 ) ;
  assign n22784 = n3027 | n9689 ;
  assign n22785 = n22784 ^ n16324 ^ 1'b0 ;
  assign n22786 = ( ~x97 & n7453 ) | ( ~x97 & n22785 ) | ( n7453 & n22785 ) ;
  assign n22787 = ~n4994 & n5088 ;
  assign n22788 = n22787 ^ n16301 ^ 1'b0 ;
  assign n22789 = n7353 | n14923 ;
  assign n22790 = n22789 ^ n6758 ^ 1'b0 ;
  assign n22791 = ( ~n222 & n21649 ) | ( ~n222 & n22790 ) | ( n21649 & n22790 ) ;
  assign n22792 = n22791 ^ n7496 ^ 1'b0 ;
  assign n22793 = n1567 & n22792 ;
  assign n22794 = n6486 ^ n2938 ^ 1'b0 ;
  assign n22795 = ~n13245 & n22794 ;
  assign n22796 = n7235 | n17970 ;
  assign n22797 = n11282 & ~n22796 ;
  assign n22798 = n3880 & n5963 ;
  assign n22799 = n22798 ^ n10301 ^ 1'b0 ;
  assign n22800 = n9675 & ~n22799 ;
  assign n22801 = ~n15240 & n21889 ;
  assign n22802 = n22490 ^ n4081 ^ 1'b0 ;
  assign n22804 = ( n336 & n553 ) | ( n336 & n6151 ) | ( n553 & n6151 ) ;
  assign n22803 = n9106 & n12890 ;
  assign n22805 = n22804 ^ n22803 ^ 1'b0 ;
  assign n22806 = n11368 ^ n7854 ^ 1'b0 ;
  assign n22807 = n22806 ^ n17962 ^ n2545 ;
  assign n22808 = n7636 ^ n1038 ^ 1'b0 ;
  assign n22809 = n11162 & ~n18081 ;
  assign n22810 = n4052 | n8080 ;
  assign n22811 = n22810 ^ n17850 ^ 1'b0 ;
  assign n22812 = n2928 | n9473 ;
  assign n22813 = n22812 ^ n3384 ^ 1'b0 ;
  assign n22814 = n3533 ^ n1211 ^ n344 ;
  assign n22815 = n22814 ^ n13686 ^ x63 ;
  assign n22817 = ~n480 & n12083 ;
  assign n22816 = n5028 & ~n16756 ;
  assign n22818 = n22817 ^ n22816 ^ n6153 ;
  assign n22819 = n3251 | n5876 ;
  assign n22820 = n13345 | n22819 ;
  assign n22821 = ~n1498 & n14205 ;
  assign n22822 = ~n22820 & n22821 ;
  assign n22823 = n7032 ^ n1199 ^ 1'b0 ;
  assign n22824 = ~n8563 & n9696 ;
  assign n22825 = ~n17927 & n22824 ;
  assign n22826 = n2634 | n22825 ;
  assign n22827 = n20142 & ~n22826 ;
  assign n22828 = n15090 ^ n12251 ^ 1'b0 ;
  assign n22829 = ~n6555 & n22828 ;
  assign n22830 = ~n6840 & n6990 ;
  assign n22831 = ~n6917 & n22830 ;
  assign n22832 = n22831 ^ n16386 ^ 1'b0 ;
  assign n22833 = n22829 & ~n22832 ;
  assign n22834 = n10150 ^ x11 ^ 1'b0 ;
  assign n22835 = n3973 ^ n3960 ^ 1'b0 ;
  assign n22836 = n17833 ^ n208 ^ 1'b0 ;
  assign n22837 = n3429 ^ x15 ^ 1'b0 ;
  assign n22838 = n11842 | n22837 ;
  assign n22839 = n13299 ^ n11292 ^ 1'b0 ;
  assign n22840 = n13341 & n22839 ;
  assign n22841 = n2956 & ~n17890 ;
  assign n22842 = n2826 | n10889 ;
  assign n22843 = n15917 | n22842 ;
  assign n22844 = ~n14674 & n16378 ;
  assign n22845 = n22844 ^ n8339 ^ 1'b0 ;
  assign n22846 = n7607 ^ n3162 ^ 1'b0 ;
  assign n22847 = ( n249 & n1835 ) | ( n249 & ~n4041 ) | ( n1835 & ~n4041 ) ;
  assign n22848 = n3740 & n22847 ;
  assign n22849 = n10304 | n22815 ;
  assign n22850 = n22849 ^ n7652 ^ 1'b0 ;
  assign n22851 = n2605 & n18731 ;
  assign n22852 = ~n6387 & n22851 ;
  assign n22853 = n11404 ^ n10216 ^ 1'b0 ;
  assign n22854 = ~n22852 & n22853 ;
  assign n22856 = n1689 | n10820 ;
  assign n22857 = n4547 & ~n22856 ;
  assign n22855 = n12240 ^ n11181 ^ 1'b0 ;
  assign n22858 = n22857 ^ n22855 ^ 1'b0 ;
  assign n22859 = n5486 | n10600 ;
  assign n22860 = n22859 ^ n18949 ^ 1'b0 ;
  assign n22861 = n16714 ^ n4012 ^ 1'b0 ;
  assign n22862 = n7330 & ~n22861 ;
  assign n22863 = ~n15634 & n22862 ;
  assign n22864 = n12996 & n14610 ;
  assign n22865 = n2737 & n22864 ;
  assign n22866 = ~n2154 & n10903 ;
  assign n22868 = ~n13075 & n16056 ;
  assign n22867 = n6712 | n13544 ;
  assign n22869 = n22868 ^ n22867 ^ 1'b0 ;
  assign n22870 = n22869 ^ x16 ^ 1'b0 ;
  assign n22871 = n2814 ^ n224 ^ 1'b0 ;
  assign n22872 = n14336 ^ n1552 ^ 1'b0 ;
  assign n22873 = n20721 | n22872 ;
  assign n22874 = n586 | n4107 ;
  assign n22876 = x69 & n6140 ;
  assign n22875 = n4510 & n15769 ;
  assign n22877 = n22876 ^ n22875 ^ 1'b0 ;
  assign n22878 = n7906 & ~n22877 ;
  assign n22879 = n22878 ^ n3897 ^ 1'b0 ;
  assign n22880 = n15618 ^ n4482 ^ 1'b0 ;
  assign n22881 = n6148 & ~n8829 ;
  assign n22882 = n22881 ^ n6370 ^ 1'b0 ;
  assign n22883 = n22882 ^ n15806 ^ 1'b0 ;
  assign n22884 = ~n8853 & n22883 ;
  assign n22885 = n1463 | n11014 ;
  assign n22886 = x6 & ~n22885 ;
  assign n22887 = ~n22884 & n22886 ;
  assign n22888 = n6529 & n22738 ;
  assign n22889 = n6775 & n22888 ;
  assign n22890 = n22889 ^ n17461 ^ 1'b0 ;
  assign n22891 = n5374 & ~n11872 ;
  assign n22892 = n4324 & n22891 ;
  assign n22893 = n9923 ^ x48 ^ 1'b0 ;
  assign n22894 = n9276 | n9348 ;
  assign n22895 = n22894 ^ n6727 ^ 1'b0 ;
  assign n22896 = n8535 | n22895 ;
  assign n22897 = n1697 | n8489 ;
  assign n22898 = n15289 & n22897 ;
  assign n22899 = n1681 & n22898 ;
  assign n22900 = ~n3839 & n20283 ;
  assign n22901 = ( ~n147 & n8080 ) | ( ~n147 & n10356 ) | ( n8080 & n10356 ) ;
  assign n22902 = n11416 ^ n10506 ^ 1'b0 ;
  assign n22903 = n3171 & ~n22902 ;
  assign n22904 = ~n22901 & n22903 ;
  assign n22905 = ~n351 & n22904 ;
  assign n22906 = n5462 & n9885 ;
  assign n22907 = ~n21102 & n22906 ;
  assign n22908 = n22907 ^ n1819 ^ 1'b0 ;
  assign n22909 = n16456 & n22908 ;
  assign n22910 = n7600 ^ n3278 ^ 1'b0 ;
  assign n22911 = n19626 ^ n16287 ^ 1'b0 ;
  assign n22912 = n2235 & n7347 ;
  assign n22913 = n22912 ^ n3439 ^ 1'b0 ;
  assign n22914 = n152 & ~n22913 ;
  assign n22915 = n20341 ^ n154 ^ 1'b0 ;
  assign n22916 = n18048 & ~n22915 ;
  assign n22917 = n5594 ^ n3188 ^ 1'b0 ;
  assign n22918 = n11165 ^ n5329 ^ 1'b0 ;
  assign n22919 = ~n1270 & n18843 ;
  assign n22920 = n22919 ^ n2091 ^ 1'b0 ;
  assign n22921 = n12724 ^ n6092 ^ 1'b0 ;
  assign n22922 = ~n4551 & n22921 ;
  assign n22923 = n4093 ^ n1399 ^ 1'b0 ;
  assign n22924 = n11758 ^ n11269 ^ 1'b0 ;
  assign n22925 = n17017 | n22924 ;
  assign n22926 = n1970 & n13326 ;
  assign n22927 = n5716 ^ n5074 ^ 1'b0 ;
  assign n22928 = n4355 | n7778 ;
  assign n22929 = n22928 ^ n1879 ^ 1'b0 ;
  assign n22930 = x51 & ~n22929 ;
  assign n22931 = ~n11961 & n22930 ;
  assign n22932 = n22931 ^ n14314 ^ 1'b0 ;
  assign n22933 = n8702 & n15002 ;
  assign n22934 = n12921 & n19304 ;
  assign n22935 = n6820 & n22934 ;
  assign n22936 = n2207 ^ n1495 ^ 1'b0 ;
  assign n22937 = n22936 ^ n4134 ^ 1'b0 ;
  assign n22938 = x32 & n18374 ;
  assign n22939 = n2905 & ~n22938 ;
  assign n22940 = ~n1710 & n8005 ;
  assign n22941 = n19887 ^ n13757 ^ 1'b0 ;
  assign n22942 = n11063 & ~n13669 ;
  assign n22943 = n22942 ^ n3116 ^ 1'b0 ;
  assign n22944 = ~n15617 & n22943 ;
  assign n22945 = n849 & n22944 ;
  assign n22946 = n6900 & n14328 ;
  assign n22947 = n22946 ^ n4418 ^ 1'b0 ;
  assign n22948 = ~n8651 & n10695 ;
  assign n22949 = ( n3968 & ~n6416 ) | ( n3968 & n8527 ) | ( ~n6416 & n8527 ) ;
  assign n22950 = n17006 ^ n9416 ^ n2414 ;
  assign n22951 = n22950 ^ n6230 ^ 1'b0 ;
  assign n22952 = n680 | n12334 ;
  assign n22953 = n22952 ^ n15921 ^ 1'b0 ;
  assign n22954 = n5738 ^ n3233 ^ 1'b0 ;
  assign n22955 = n14526 & n22954 ;
  assign n22956 = n8920 & n21173 ;
  assign n22957 = n19552 ^ n7905 ^ 1'b0 ;
  assign n22958 = n15740 ^ n1898 ^ 1'b0 ;
  assign n22959 = n8583 ^ n7781 ^ 1'b0 ;
  assign n22960 = n6720 & ~n10532 ;
  assign n22961 = n18344 & n22960 ;
  assign n22962 = n10784 & n19300 ;
  assign n22963 = ~n5135 & n5974 ;
  assign n22964 = n12919 & n22963 ;
  assign n22965 = n6575 & ~n10891 ;
  assign n22966 = n2146 ^ n1450 ^ 1'b0 ;
  assign n22967 = n5297 & n22966 ;
  assign n22968 = n6665 | n22967 ;
  assign n22969 = n22968 ^ n6953 ^ 1'b0 ;
  assign n22970 = n22969 ^ n8737 ^ n2804 ;
  assign n22971 = n1535 | n20211 ;
  assign n22972 = n22971 ^ n6237 ^ 1'b0 ;
  assign n22973 = n12240 ^ n9158 ^ 1'b0 ;
  assign n22974 = n22972 & ~n22973 ;
  assign n22975 = n6174 ^ x71 ^ 1'b0 ;
  assign n22976 = n19058 | n19117 ;
  assign n22977 = n22976 ^ n13521 ^ 1'b0 ;
  assign n22978 = n2802 ^ n254 ^ 1'b0 ;
  assign n22979 = ~n20783 & n22978 ;
  assign n22980 = n4329 & ~n7360 ;
  assign n22981 = ( n1103 & ~n5200 ) | ( n1103 & n22980 ) | ( ~n5200 & n22980 ) ;
  assign n22982 = ~n10208 & n15202 ;
  assign n22983 = n22982 ^ n13397 ^ 1'b0 ;
  assign n22984 = n15113 | n15486 ;
  assign n22985 = n4766 & ~n22984 ;
  assign n22986 = n1377 & n2382 ;
  assign n22987 = n18081 ^ n15171 ^ 1'b0 ;
  assign n22988 = n10941 | n22987 ;
  assign n22989 = n15840 ^ n361 ^ 1'b0 ;
  assign n22990 = n17970 ^ n17504 ^ 1'b0 ;
  assign n22991 = n3576 & ~n19930 ;
  assign n22992 = n20619 | n22991 ;
  assign n22993 = n16755 ^ n3951 ^ 1'b0 ;
  assign n22994 = n17072 | n22993 ;
  assign n22995 = n3788 & n4881 ;
  assign n22996 = n22995 ^ n11550 ^ 1'b0 ;
  assign n22997 = ~n17651 & n22996 ;
  assign n22998 = ~n14313 & n14952 ;
  assign n22999 = ( n16354 & n22997 ) | ( n16354 & n22998 ) | ( n22997 & n22998 ) ;
  assign n23000 = n1121 & ~n6619 ;
  assign n23001 = n23000 ^ n2882 ^ 1'b0 ;
  assign n23003 = n11938 ^ n10885 ^ 1'b0 ;
  assign n23002 = n2440 | n13734 ;
  assign n23004 = n23003 ^ n23002 ^ 1'b0 ;
  assign n23005 = n4976 | n14251 ;
  assign n23006 = n23004 & ~n23005 ;
  assign n23007 = n3206 | n20228 ;
  assign n23008 = n23007 ^ n3738 ^ 1'b0 ;
  assign n23009 = n17314 | n22953 ;
  assign n23010 = n4844 ^ n2638 ^ 1'b0 ;
  assign n23011 = n9668 ^ n9071 ^ 1'b0 ;
  assign n23012 = n4073 | n13097 ;
  assign n23013 = n23012 ^ n6493 ^ 1'b0 ;
  assign n23014 = n1856 & ~n2167 ;
  assign n23015 = n980 & n23014 ;
  assign n23016 = n2561 & ~n23015 ;
  assign n23017 = n23016 ^ n8224 ^ 1'b0 ;
  assign n23018 = n2401 & ~n2531 ;
  assign n23019 = n19257 & n20015 ;
  assign n23020 = n6592 ^ n3520 ^ 1'b0 ;
  assign n23021 = n9027 & n23020 ;
  assign n23022 = n12906 | n23021 ;
  assign n23023 = n23022 ^ n9540 ^ 1'b0 ;
  assign n23024 = n9438 | n23023 ;
  assign n23026 = ~n2630 & n7535 ;
  assign n23025 = ~n4318 & n9693 ;
  assign n23027 = n23026 ^ n23025 ^ 1'b0 ;
  assign n23028 = n11995 ^ n5178 ^ 1'b0 ;
  assign n23029 = n1157 | n1880 ;
  assign n23030 = n9269 & ~n23029 ;
  assign n23031 = n23030 ^ n283 ^ 1'b0 ;
  assign n23032 = n6110 & ~n15249 ;
  assign n23033 = ~n23031 & n23032 ;
  assign n23034 = n9616 | n11366 ;
  assign n23035 = ( n2410 & n16020 ) | ( n2410 & n18002 ) | ( n16020 & n18002 ) ;
  assign n23036 = n7194 & n7641 ;
  assign n23037 = ( n466 & ~n21734 ) | ( n466 & n23036 ) | ( ~n21734 & n23036 ) ;
  assign n23038 = n7030 | n11049 ;
  assign n23039 = n23038 ^ n4443 ^ 1'b0 ;
  assign n23040 = n7986 | n15777 ;
  assign n23041 = n23040 ^ n21314 ^ 1'b0 ;
  assign n23042 = n12762 ^ n548 ^ 1'b0 ;
  assign n23043 = n204 | n23042 ;
  assign n23044 = n4447 ^ n1524 ^ 1'b0 ;
  assign n23045 = ~n6936 & n9578 ;
  assign n23046 = ~n23044 & n23045 ;
  assign n23047 = n9001 & ~n17537 ;
  assign n23048 = n7590 & n17824 ;
  assign n23049 = n11485 & ~n23048 ;
  assign n23050 = n3145 & n11912 ;
  assign n23051 = n14969 ^ n13413 ^ n9023 ;
  assign n23052 = n19002 ^ n12262 ^ 1'b0 ;
  assign n23053 = n1719 & n3420 ;
  assign n23054 = ~n10222 & n23053 ;
  assign n23056 = n6273 & n7736 ;
  assign n23057 = n23056 ^ n1046 ^ 1'b0 ;
  assign n23055 = n2868 | n12088 ;
  assign n23058 = n23057 ^ n23055 ^ 1'b0 ;
  assign n23059 = n774 | n19055 ;
  assign n23062 = n3968 | n11416 ;
  assign n23063 = n6762 | n23062 ;
  assign n23060 = n10507 & ~n20130 ;
  assign n23061 = n23060 ^ n719 ^ 1'b0 ;
  assign n23064 = n23063 ^ n23061 ^ 1'b0 ;
  assign n23065 = ~n1939 & n11364 ;
  assign n23066 = n23065 ^ n4769 ^ 1'b0 ;
  assign n23067 = n10990 ^ n4549 ^ 1'b0 ;
  assign n23068 = n15383 ^ n3546 ^ 1'b0 ;
  assign n23069 = n12842 ^ n10274 ^ 1'b0 ;
  assign n23070 = n23068 | n23069 ;
  assign n23071 = ~n10039 & n11687 ;
  assign n23072 = n2156 & ~n23071 ;
  assign n23073 = n23072 ^ n7643 ^ 1'b0 ;
  assign n23074 = ~n23070 & n23073 ;
  assign n23075 = n12883 ^ n9712 ^ n4710 ;
  assign n23076 = n5935 ^ n4675 ^ 1'b0 ;
  assign n23077 = n4671 | n23076 ;
  assign n23078 = n16150 ^ n6249 ^ 1'b0 ;
  assign n23079 = n5931 & n23078 ;
  assign n23080 = n23077 & n23079 ;
  assign n23081 = ( n6108 & n21069 ) | ( n6108 & ~n23080 ) | ( n21069 & ~n23080 ) ;
  assign n23082 = n8306 & n9998 ;
  assign n23083 = n11605 & n23082 ;
  assign n23084 = n22027 | n23083 ;
  assign n23085 = n23084 ^ n16433 ^ 1'b0 ;
  assign n23086 = n8889 ^ n3699 ^ 1'b0 ;
  assign n23087 = n8711 | n15548 ;
  assign n23088 = n4357 & ~n23087 ;
  assign n23089 = n5840 & n6133 ;
  assign n23090 = ~n10615 & n23089 ;
  assign n23091 = n23090 ^ n20519 ^ n9015 ;
  assign n23092 = n23091 ^ n5050 ^ 1'b0 ;
  assign n23093 = n5614 & ~n23092 ;
  assign n23094 = n2235 | n18279 ;
  assign n23095 = n1113 & n6029 ;
  assign n23096 = ( ~n3565 & n21347 ) | ( ~n3565 & n23095 ) | ( n21347 & n23095 ) ;
  assign n23097 = n12481 ^ n2694 ^ 1'b0 ;
  assign n23098 = n2103 & ~n10161 ;
  assign n23099 = n8845 ^ n6474 ^ 1'b0 ;
  assign n23100 = n23098 & ~n23099 ;
  assign n23101 = n23097 & n23100 ;
  assign n23102 = n4014 & n14559 ;
  assign n23103 = n23102 ^ n17082 ^ 1'b0 ;
  assign n23104 = n9191 & ~n23103 ;
  assign n23105 = n23104 ^ n13692 ^ 1'b0 ;
  assign n23106 = n17470 ^ n3973 ^ 1'b0 ;
  assign n23107 = n2204 | n3888 ;
  assign n23108 = n23107 ^ n489 ^ 1'b0 ;
  assign n23109 = ~n4411 & n23108 ;
  assign n23110 = n19814 ^ n7527 ^ 1'b0 ;
  assign n23111 = n17970 & ~n23110 ;
  assign n23112 = n16658 ^ n5970 ^ 1'b0 ;
  assign n23113 = n20211 & n23112 ;
  assign n23114 = n22136 ^ n583 ^ 1'b0 ;
  assign n23115 = n1869 & ~n23114 ;
  assign n23116 = n23115 ^ x124 ^ 1'b0 ;
  assign n23117 = n5356 & ~n19677 ;
  assign n23118 = n3165 & ~n5614 ;
  assign n23119 = n1365 & ~n13505 ;
  assign n23120 = n6565 & n23119 ;
  assign n23121 = n10165 ^ n9837 ^ 1'b0 ;
  assign n23122 = n16196 & ~n23121 ;
  assign n23123 = ( n6717 & ~n11734 ) | ( n6717 & n21900 ) | ( ~n11734 & n21900 ) ;
  assign n23128 = n14610 ^ n4472 ^ 1'b0 ;
  assign n23124 = ~n466 & n4506 ;
  assign n23125 = n18964 ^ n15195 ^ 1'b0 ;
  assign n23126 = x35 & ~n23125 ;
  assign n23127 = n23124 & n23126 ;
  assign n23129 = n23128 ^ n23127 ^ 1'b0 ;
  assign n23130 = n718 | n8773 ;
  assign n23131 = n23130 ^ n3866 ^ 1'b0 ;
  assign n23132 = n12935 & ~n14771 ;
  assign n23133 = n23132 ^ n1429 ^ 1'b0 ;
  assign n23134 = n3085 & ~n23133 ;
  assign n23135 = n12476 ^ n10063 ^ 1'b0 ;
  assign n23136 = n14243 ^ n4843 ^ 1'b0 ;
  assign n23137 = ~n391 & n9528 ;
  assign n23138 = n23137 ^ n19298 ^ 1'b0 ;
  assign n23143 = n3999 | n8118 ;
  assign n23144 = n13637 & ~n23143 ;
  assign n23145 = n3536 & ~n23144 ;
  assign n23146 = n23145 ^ n10217 ^ 1'b0 ;
  assign n23139 = n4784 ^ n2960 ^ 1'b0 ;
  assign n23140 = n10345 | n23139 ;
  assign n23141 = n23140 ^ n2963 ^ 1'b0 ;
  assign n23142 = n3726 & ~n23141 ;
  assign n23147 = n23146 ^ n23142 ^ 1'b0 ;
  assign n23148 = n7942 & ~n17576 ;
  assign n23149 = n15479 & n23148 ;
  assign n23150 = n5623 | n18271 ;
  assign n23151 = n14869 ^ n3404 ^ 1'b0 ;
  assign n23152 = n3465 | n23151 ;
  assign n23153 = n17675 ^ n2337 ^ 1'b0 ;
  assign n23154 = ~n19973 & n23153 ;
  assign n23156 = n2189 ^ n843 ^ 1'b0 ;
  assign n23157 = n7110 & ~n23156 ;
  assign n23158 = n4853 | n9831 ;
  assign n23159 = n23157 | n23158 ;
  assign n23155 = n3319 | n15177 ;
  assign n23160 = n23159 ^ n23155 ^ 1'b0 ;
  assign n23163 = n240 & ~n1224 ;
  assign n23164 = n15925 & n23163 ;
  assign n23161 = ~n735 & n1867 ;
  assign n23162 = ~n5623 & n23161 ;
  assign n23165 = n23164 ^ n23162 ^ 1'b0 ;
  assign n23166 = ( n1083 & n1232 ) | ( n1083 & ~n3336 ) | ( n1232 & ~n3336 ) ;
  assign n23167 = ~n1329 & n23166 ;
  assign n23168 = ~n2948 & n23167 ;
  assign n23169 = n11942 ^ n6277 ^ 1'b0 ;
  assign n23170 = n2330 & n23169 ;
  assign n23171 = ~n9931 & n23170 ;
  assign n23172 = ~n16618 & n23171 ;
  assign n23173 = ~n3167 & n3589 ;
  assign n23174 = n709 & n23173 ;
  assign n23175 = n15544 & n20057 ;
  assign n23176 = n18448 ^ n18383 ^ 1'b0 ;
  assign n23177 = n5203 | n14237 ;
  assign n23178 = n10321 ^ n9528 ^ 1'b0 ;
  assign n23179 = ~n1893 & n23178 ;
  assign n23185 = n8862 ^ n4717 ^ 1'b0 ;
  assign n23180 = n311 & ~n779 ;
  assign n23181 = ~n311 & n23180 ;
  assign n23182 = n14251 | n23181 ;
  assign n23183 = n23181 & ~n23182 ;
  assign n23184 = n17021 | n23183 ;
  assign n23186 = n23185 ^ n23184 ^ 1'b0 ;
  assign n23187 = n11714 ^ n1646 ^ 1'b0 ;
  assign n23188 = ~n7024 & n21143 ;
  assign n23189 = n23188 ^ n2802 ^ 1'b0 ;
  assign n23190 = n2250 & ~n3413 ;
  assign n23191 = n23190 ^ n1664 ^ 1'b0 ;
  assign n23192 = n22783 ^ n15037 ^ 1'b0 ;
  assign n23193 = n4906 & ~n23192 ;
  assign n23194 = n2382 & ~n20721 ;
  assign n23195 = n23194 ^ n349 ^ 1'b0 ;
  assign n23196 = ( n1861 & ~n2608 ) | ( n1861 & n5154 ) | ( ~n2608 & n5154 ) ;
  assign n23197 = n7362 | n23196 ;
  assign n23198 = n23197 ^ n1821 ^ 1'b0 ;
  assign n23199 = n8582 ^ n3470 ^ 1'b0 ;
  assign n23200 = n9882 ^ n9169 ^ 1'b0 ;
  assign n23201 = ~n23199 & n23200 ;
  assign n23202 = n16181 | n23201 ;
  assign n23203 = ~n10352 & n11190 ;
  assign n23204 = n23203 ^ n15632 ^ n6568 ;
  assign n23205 = n17441 ^ n5918 ^ 1'b0 ;
  assign n23206 = n17557 ^ n581 ^ 1'b0 ;
  assign n23207 = n23206 ^ n2109 ^ 1'b0 ;
  assign n23208 = n9022 ^ n2671 ^ 1'b0 ;
  assign n23209 = n8416 ^ n3944 ^ 1'b0 ;
  assign n23210 = n6994 & ~n11990 ;
  assign n23211 = ~n340 & n23210 ;
  assign n23212 = n23211 ^ n4940 ^ 1'b0 ;
  assign n23213 = n23209 | n23212 ;
  assign n23214 = n11990 ^ n4120 ^ 1'b0 ;
  assign n23215 = ~n2804 & n23214 ;
  assign n23216 = n18898 ^ n13612 ^ 1'b0 ;
  assign n23217 = n16195 ^ n3921 ^ 1'b0 ;
  assign n23218 = ~n14929 & n21466 ;
  assign n23219 = ~n1011 & n13987 ;
  assign n23220 = n2020 & n23219 ;
  assign n23221 = n16141 ^ x75 ^ 1'b0 ;
  assign n23224 = n5787 ^ n2582 ^ 1'b0 ;
  assign n23222 = ( ~n468 & n5645 ) | ( ~n468 & n5904 ) | ( n5645 & n5904 ) ;
  assign n23223 = n23222 ^ n17085 ^ n3986 ;
  assign n23225 = n23224 ^ n23223 ^ 1'b0 ;
  assign n23226 = n19991 & ~n23225 ;
  assign n23227 = n11965 ^ n3626 ^ 1'b0 ;
  assign n23228 = n6244 ^ n1863 ^ 1'b0 ;
  assign n23229 = ~n2949 & n16714 ;
  assign n23230 = n22151 | n23229 ;
  assign n23231 = n5544 & n23230 ;
  assign n23232 = n9733 & ~n23231 ;
  assign n23233 = n23232 ^ n723 ^ 1'b0 ;
  assign n23234 = ~n7134 & n23233 ;
  assign n23235 = n8078 ^ n3674 ^ 1'b0 ;
  assign n23237 = n5249 | n10183 ;
  assign n23238 = n23237 ^ n11178 ^ 1'b0 ;
  assign n23239 = n2952 & ~n23238 ;
  assign n23240 = n23239 ^ n9664 ^ 1'b0 ;
  assign n23236 = n14702 & ~n23206 ;
  assign n23241 = n23240 ^ n23236 ^ 1'b0 ;
  assign n23243 = ~n4368 & n9265 ;
  assign n23242 = n8654 | n10307 ;
  assign n23244 = n23243 ^ n23242 ^ 1'b0 ;
  assign n23245 = n9923 & n13114 ;
  assign n23246 = ~n874 & n23245 ;
  assign n23247 = ~n4520 & n17662 ;
  assign n23248 = n4867 & n23247 ;
  assign n23250 = ( n2861 & n8641 ) | ( n2861 & n17606 ) | ( n8641 & n17606 ) ;
  assign n23249 = n747 & n10343 ;
  assign n23251 = n23250 ^ n23249 ^ 1'b0 ;
  assign n23252 = n4776 ^ n141 ^ 1'b0 ;
  assign n23253 = n1568 & ~n23252 ;
  assign n23254 = ~n5332 & n23253 ;
  assign n23255 = n5854 & ~n23254 ;
  assign n23256 = n12799 & n23255 ;
  assign n23257 = n20600 ^ n11478 ^ 1'b0 ;
  assign n23258 = n16188 & ~n23257 ;
  assign n23259 = n11611 ^ n6981 ^ 1'b0 ;
  assign n23260 = n23259 ^ n12031 ^ n10527 ;
  assign n23262 = n1742 | n4252 ;
  assign n23263 = n23262 ^ n4877 ^ 1'b0 ;
  assign n23261 = ~n5468 & n16050 ;
  assign n23264 = n23263 ^ n23261 ^ n10072 ;
  assign n23265 = n21439 ^ n9613 ^ 1'b0 ;
  assign n23266 = ~n7305 & n23265 ;
  assign n23267 = n1300 & ~n20969 ;
  assign n23268 = n9163 ^ n3298 ^ 1'b0 ;
  assign n23269 = n7536 & n23268 ;
  assign n23270 = n15369 ^ n10237 ^ 1'b0 ;
  assign n23271 = n15137 ^ n11948 ^ 1'b0 ;
  assign n23272 = ( n5088 & ~n5408 ) | ( n5088 & n10274 ) | ( ~n5408 & n10274 ) ;
  assign n23273 = ~n6022 & n23272 ;
  assign n23274 = ( n6807 & ~n16468 ) | ( n6807 & n19949 ) | ( ~n16468 & n19949 ) ;
  assign n23275 = n23274 ^ n6468 ^ 1'b0 ;
  assign n23276 = n1495 | n23275 ;
  assign n23277 = ( ~n4733 & n7857 ) | ( ~n4733 & n12088 ) | ( n7857 & n12088 ) ;
  assign n23278 = n8855 & ~n16934 ;
  assign n23279 = ~n23277 & n23278 ;
  assign n23280 = n6640 ^ n472 ^ 1'b0 ;
  assign n23281 = n3636 & ~n23280 ;
  assign n23282 = ~n2444 & n23281 ;
  assign n23283 = n11797 ^ n3804 ^ 1'b0 ;
  assign n23284 = n4820 & ~n23283 ;
  assign n23285 = ~n4604 & n23284 ;
  assign n23286 = n5154 & n23285 ;
  assign n23287 = n4077 ^ n1189 ^ 1'b0 ;
  assign n23288 = ~n419 & n3255 ;
  assign n23289 = n23288 ^ n15429 ^ 1'b0 ;
  assign n23290 = ~n1406 & n23289 ;
  assign n23291 = n503 & ~n14579 ;
  assign n23292 = n464 | n13343 ;
  assign n23293 = n23292 ^ n17736 ^ 1'b0 ;
  assign n23294 = n10971 | n12621 ;
  assign n23295 = n23294 ^ n8269 ^ 1'b0 ;
  assign n23296 = n14151 & ~n14248 ;
  assign n23297 = n299 & n21381 ;
  assign n23298 = n9383 ^ n2038 ^ 1'b0 ;
  assign n23299 = n15279 & ~n23298 ;
  assign n23300 = n19792 ^ n13032 ^ 1'b0 ;
  assign n23301 = n3286 | n10947 ;
  assign n23302 = n19532 | n23301 ;
  assign n23303 = ~n11883 & n18533 ;
  assign n23304 = n12580 ^ n3411 ^ 1'b0 ;
  assign n23305 = x75 & ~n13576 ;
  assign n23306 = n23305 ^ n20694 ^ 1'b0 ;
  assign n23307 = n5385 & ~n8388 ;
  assign n23308 = n23307 ^ n16956 ^ 1'b0 ;
  assign n23309 = n1529 & n11175 ;
  assign n23310 = ~n1801 & n23309 ;
  assign n23311 = n8906 | n23310 ;
  assign n23312 = n14592 & ~n23311 ;
  assign n23313 = n3481 & ~n15093 ;
  assign n23314 = n7194 ^ n5265 ^ 1'b0 ;
  assign n23315 = n17991 & ~n23314 ;
  assign n23316 = x54 | n1247 ;
  assign n23317 = ~n9484 & n23316 ;
  assign n23318 = n12420 & n23317 ;
  assign n23319 = n829 & n12996 ;
  assign n23320 = ~n15836 & n23319 ;
  assign n23321 = n9768 & n15712 ;
  assign n23322 = ( ~n4808 & n5613 ) | ( ~n4808 & n9130 ) | ( n5613 & n9130 ) ;
  assign n23323 = n22337 ^ n12059 ^ 1'b0 ;
  assign n23324 = n7713 & n23323 ;
  assign n23325 = ( n1413 & n23322 ) | ( n1413 & ~n23324 ) | ( n23322 & ~n23324 ) ;
  assign n23326 = n11457 | n19906 ;
  assign n23327 = n23326 ^ n1422 ^ 1'b0 ;
  assign n23328 = n4251 ^ n2558 ^ 1'b0 ;
  assign n23329 = n3459 | n23328 ;
  assign n23330 = n15929 & ~n22797 ;
  assign n23331 = n23330 ^ n18782 ^ 1'b0 ;
  assign n23332 = n8659 ^ n7488 ^ 1'b0 ;
  assign n23333 = n3115 & ~n6177 ;
  assign n23334 = n14804 & n23333 ;
  assign n23335 = ~n8684 & n9645 ;
  assign n23336 = ~n23334 & n23335 ;
  assign n23337 = n4433 & ~n9527 ;
  assign n23338 = n12623 & n23337 ;
  assign n23339 = ~n4526 & n10808 ;
  assign n23340 = n23339 ^ n17988 ^ 1'b0 ;
  assign n23341 = n11993 | n19584 ;
  assign n23342 = n12332 ^ n6078 ^ 1'b0 ;
  assign n23343 = n2405 & n15638 ;
  assign n23344 = n23343 ^ n12087 ^ 1'b0 ;
  assign n23345 = n513 | n23344 ;
  assign n23346 = n9134 | n11807 ;
  assign n23347 = n17031 ^ n12131 ^ 1'b0 ;
  assign n23348 = n10740 & n23347 ;
  assign n23349 = n3910 | n5958 ;
  assign n23350 = n10201 & ~n12092 ;
  assign n23351 = n12197 ^ n156 ^ 1'b0 ;
  assign n23354 = n1189 & n2213 ;
  assign n23355 = n23354 ^ n9756 ^ 1'b0 ;
  assign n23352 = n13680 ^ n3495 ^ 1'b0 ;
  assign n23353 = n10204 & n23352 ;
  assign n23356 = n23355 ^ n23353 ^ n10689 ;
  assign n23357 = n13972 ^ n1773 ^ 1'b0 ;
  assign n23358 = n14784 ^ n4260 ^ 1'b0 ;
  assign n23359 = n3991 & ~n23358 ;
  assign n23360 = ~n12692 & n18788 ;
  assign n23361 = n4536 & n23360 ;
  assign n23362 = n11401 ^ n297 ^ 1'b0 ;
  assign n23363 = n13114 & ~n23362 ;
  assign n23364 = ~n12963 & n23363 ;
  assign n23365 = n23364 ^ n15548 ^ 1'b0 ;
  assign n23366 = n5667 & n14664 ;
  assign n23367 = ~n17934 & n23366 ;
  assign n23368 = n10804 | n12011 ;
  assign n23369 = n23368 ^ n978 ^ 1'b0 ;
  assign n23370 = n14966 & n23369 ;
  assign n23371 = n10183 ^ n4355 ^ 1'b0 ;
  assign n23372 = n23371 ^ n12816 ^ n6478 ;
  assign n23373 = ~n9656 & n13402 ;
  assign n23374 = n9164 & n14614 ;
  assign n23375 = n23374 ^ n1819 ^ 1'b0 ;
  assign n23376 = n8776 & ~n23375 ;
  assign n23377 = n6990 & ~n7100 ;
  assign n23378 = ~n4287 & n5637 ;
  assign n23379 = n23378 ^ n11025 ^ 1'b0 ;
  assign n23380 = n20638 | n23379 ;
  assign n23381 = ~n10320 & n22122 ;
  assign n23382 = n16188 ^ n2818 ^ 1'b0 ;
  assign n23383 = n23382 ^ n13583 ^ n9009 ;
  assign n23384 = n17552 ^ n9225 ^ 1'b0 ;
  assign n23385 = n504 ^ n148 ^ 1'b0 ;
  assign n23386 = n23385 ^ n4630 ^ 1'b0 ;
  assign n23387 = n5179 | n23012 ;
  assign n23388 = n23387 ^ n4217 ^ 1'b0 ;
  assign n23389 = ~n11889 & n18817 ;
  assign n23390 = n23389 ^ n1821 ^ 1'b0 ;
  assign n23391 = n5262 & n10585 ;
  assign n23392 = n7678 & ~n18823 ;
  assign n23393 = n23392 ^ n14968 ^ 1'b0 ;
  assign n23394 = n23393 ^ n1011 ^ 1'b0 ;
  assign n23395 = n4865 & n11056 ;
  assign n23396 = n17725 ^ n13622 ^ 1'b0 ;
  assign n23397 = n7727 ^ n1588 ^ 1'b0 ;
  assign n23398 = n23397 ^ n11606 ^ n3764 ;
  assign n23399 = n23398 ^ n3198 ^ 1'b0 ;
  assign n23400 = n23399 ^ n14463 ^ 1'b0 ;
  assign n23401 = n1635 | n23400 ;
  assign n23402 = n6189 & n7054 ;
  assign n23403 = n3547 & ~n5655 ;
  assign n23404 = n23403 ^ n9610 ^ 1'b0 ;
  assign n23405 = n13937 & ~n20295 ;
  assign n23406 = n23405 ^ n3853 ^ 1'b0 ;
  assign n23407 = ~n1597 & n20657 ;
  assign n23408 = n9290 | n11111 ;
  assign n23409 = ~n4033 & n4420 ;
  assign n23410 = n4005 & n22368 ;
  assign n23411 = n23410 ^ n6511 ^ n5250 ;
  assign n23412 = ~n11127 & n14556 ;
  assign n23413 = n23412 ^ n4387 ^ 1'b0 ;
  assign n23414 = n16595 ^ n1254 ^ 1'b0 ;
  assign n23415 = n23413 | n23414 ;
  assign n23416 = n4759 | n16725 ;
  assign n23417 = n4551 | n6473 ;
  assign n23418 = n2366 & ~n23417 ;
  assign n23419 = n137 & ~n8781 ;
  assign n23420 = n7649 | n23419 ;
  assign n23421 = n2272 & n19925 ;
  assign n23422 = n4292 | n22563 ;
  assign n23423 = n4113 ^ n1162 ^ 1'b0 ;
  assign n23424 = n4084 & n23423 ;
  assign n23425 = ~n4512 & n13965 ;
  assign n23426 = n23425 ^ n275 ^ 1'b0 ;
  assign n23427 = ~n5301 & n7071 ;
  assign n23428 = n6019 & n7297 ;
  assign n23429 = n23428 ^ n14507 ^ 1'b0 ;
  assign n23430 = ~n8744 & n11798 ;
  assign n23431 = ~n23429 & n23430 ;
  assign n23432 = n14260 & n21143 ;
  assign n23433 = n692 | n6704 ;
  assign n23434 = n5980 ^ n3746 ^ 1'b0 ;
  assign n23435 = ( n9504 & ~n23107 ) | ( n9504 & n23434 ) | ( ~n23107 & n23434 ) ;
  assign n23436 = n14022 & n18968 ;
  assign n23437 = n1906 & n23436 ;
  assign n23438 = n4250 & n4782 ;
  assign n23439 = n23438 ^ n7449 ^ 1'b0 ;
  assign n23440 = n4921 ^ n795 ^ 1'b0 ;
  assign n23441 = n23439 | n23440 ;
  assign n23442 = n6415 & ~n23048 ;
  assign n23443 = ~n2851 & n3799 ;
  assign n23444 = n23443 ^ n13596 ^ 1'b0 ;
  assign n23445 = n12903 & n21555 ;
  assign n23446 = ~n23444 & n23445 ;
  assign n23447 = n5889 | n12194 ;
  assign n23448 = n4292 | n23447 ;
  assign n23449 = n23448 ^ n255 ^ 1'b0 ;
  assign n23450 = n14846 & ~n23449 ;
  assign n23451 = ( ~n13204 & n15223 ) | ( ~n13204 & n19877 ) | ( n15223 & n19877 ) ;
  assign n23452 = n5102 & ~n19223 ;
  assign n23453 = x108 & ~n4309 ;
  assign n23454 = n16714 ^ n3381 ^ 1'b0 ;
  assign n23455 = n16169 | n23454 ;
  assign n23456 = n16775 ^ n11413 ^ 1'b0 ;
  assign n23457 = ( ~n8723 & n14229 ) | ( ~n8723 & n23456 ) | ( n14229 & n23456 ) ;
  assign n23458 = n7695 ^ n4371 ^ 1'b0 ;
  assign n23459 = n3594 & ~n5183 ;
  assign n23460 = n1348 & n23459 ;
  assign n23461 = n23460 ^ n275 ^ 1'b0 ;
  assign n23462 = n13713 ^ n1920 ^ 1'b0 ;
  assign n23463 = n10985 & ~n23462 ;
  assign n23464 = n14698 ^ n3015 ^ 1'b0 ;
  assign n23465 = n19985 & ~n23464 ;
  assign n23466 = n15953 & n23465 ;
  assign n23467 = ~n13810 & n13869 ;
  assign n23468 = ~n799 & n23467 ;
  assign n23469 = n11972 ^ n9628 ^ 1'b0 ;
  assign n23470 = n6051 | n23469 ;
  assign n23471 = n23470 ^ n2530 ^ 1'b0 ;
  assign n23472 = n11105 & ~n23471 ;
  assign n23473 = n6246 ^ n758 ^ 1'b0 ;
  assign n23474 = n23472 & n23473 ;
  assign n23475 = n23474 ^ n13777 ^ 1'b0 ;
  assign n23476 = n6680 ^ n1681 ^ 1'b0 ;
  assign n23477 = ~n10683 & n20200 ;
  assign n23478 = n23477 ^ n22901 ^ 1'b0 ;
  assign n23479 = n9758 & ~n20217 ;
  assign n23480 = n2341 | n4739 ;
  assign n23482 = n16276 ^ n10633 ^ n353 ;
  assign n23481 = x118 & n1639 ;
  assign n23483 = n23482 ^ n23481 ^ 1'b0 ;
  assign n23484 = n19574 ^ n4148 ^ 1'b0 ;
  assign n23485 = n4141 & ~n23127 ;
  assign n23486 = n7408 & ~n11928 ;
  assign n23487 = ~n475 & n11121 ;
  assign n23488 = n17790 | n23487 ;
  assign n23489 = n2842 | n20828 ;
  assign n23490 = n23489 ^ n20180 ^ 1'b0 ;
  assign n23491 = ~n6568 & n9847 ;
  assign n23492 = n10361 ^ n7164 ^ 1'b0 ;
  assign n23500 = n13282 ^ n1385 ^ 1'b0 ;
  assign n23501 = n21912 & n23500 ;
  assign n23493 = n6090 ^ n4888 ^ n208 ;
  assign n23494 = n5462 & ~n23493 ;
  assign n23495 = n3733 ^ n1937 ^ 1'b0 ;
  assign n23496 = n10983 & n23495 ;
  assign n23497 = ~n1396 & n23496 ;
  assign n23498 = ~n23494 & n23497 ;
  assign n23499 = n3286 | n23498 ;
  assign n23502 = n23501 ^ n23499 ^ 1'b0 ;
  assign n23503 = n23443 ^ n17200 ^ 1'b0 ;
  assign n23504 = n23503 ^ n10757 ^ 1'b0 ;
  assign n23505 = n20989 ^ n2458 ^ 1'b0 ;
  assign n23506 = n16795 & n23505 ;
  assign n23508 = ~n218 & n9525 ;
  assign n23509 = n23508 ^ n2802 ^ 1'b0 ;
  assign n23507 = ~n391 & n1507 ;
  assign n23510 = n23509 ^ n23507 ^ n16434 ;
  assign n23511 = n19363 ^ n18971 ^ 1'b0 ;
  assign n23512 = n6269 ^ n1021 ^ 1'b0 ;
  assign n23513 = n23512 ^ n1213 ^ 1'b0 ;
  assign n23514 = n4750 ^ n1361 ^ 1'b0 ;
  assign n23515 = n4463 & n15219 ;
  assign n23516 = n23515 ^ n20666 ^ 1'b0 ;
  assign n23517 = ~n2489 & n5787 ;
  assign n23518 = n23517 ^ n8491 ^ 1'b0 ;
  assign n23519 = n4441 & n20712 ;
  assign n23520 = ~n19597 & n23519 ;
  assign n23521 = ~n7707 & n8854 ;
  assign n23522 = n23521 ^ n10046 ^ 1'b0 ;
  assign n23523 = ( n23518 & n23520 ) | ( n23518 & n23522 ) | ( n23520 & n23522 ) ;
  assign n23524 = n8023 ^ n2650 ^ 1'b0 ;
  assign n23525 = ~n585 & n15681 ;
  assign n23526 = ( x51 & ~n1927 ) | ( x51 & n5104 ) | ( ~n1927 & n5104 ) ;
  assign n23527 = n11586 & n23526 ;
  assign n23528 = n23527 ^ n1103 ^ 1'b0 ;
  assign n23529 = ~n9846 & n10950 ;
  assign n23530 = n7876 ^ n477 ^ 1'b0 ;
  assign n23531 = n3478 & n23530 ;
  assign n23532 = n14527 ^ n4159 ^ 1'b0 ;
  assign n23533 = n16667 & ~n23532 ;
  assign n23534 = n22396 ^ n1168 ^ 1'b0 ;
  assign n23535 = n15491 & ~n23534 ;
  assign n23536 = n23385 ^ n3744 ^ 1'b0 ;
  assign n23539 = n17729 ^ n15213 ^ 1'b0 ;
  assign n23537 = n922 & ~n8299 ;
  assign n23538 = n20415 & ~n23537 ;
  assign n23540 = n23539 ^ n23538 ^ 1'b0 ;
  assign n23541 = n13919 ^ n9664 ^ 1'b0 ;
  assign n23542 = n15706 & ~n23541 ;
  assign n23543 = n9262 & n19284 ;
  assign n23544 = n23543 ^ n5149 ^ 1'b0 ;
  assign n23545 = n5109 | n6476 ;
  assign n23546 = n23545 ^ n8691 ^ 1'b0 ;
  assign n23548 = n8619 ^ n2463 ^ 1'b0 ;
  assign n23547 = n3344 & n20362 ;
  assign n23549 = n23548 ^ n23547 ^ n6449 ;
  assign n23550 = n4686 ^ n2685 ^ 1'b0 ;
  assign n23551 = n23550 ^ n18894 ^ x84 ;
  assign n23552 = n18096 ^ n8684 ^ 1'b0 ;
  assign n23553 = n7317 ^ n1398 ^ 1'b0 ;
  assign n23554 = n4596 & ~n23553 ;
  assign n23555 = n12849 ^ n3973 ^ 1'b0 ;
  assign n23556 = ~n9837 & n23555 ;
  assign n23557 = ~n18549 & n23556 ;
  assign n23558 = n438 | n8309 ;
  assign n23559 = n7190 & ~n11559 ;
  assign n23560 = ~n23558 & n23559 ;
  assign n23561 = n4987 | n5705 ;
  assign n23562 = n7528 | n23561 ;
  assign n23563 = n21687 | n23562 ;
  assign n23564 = n15602 ^ n13430 ^ 1'b0 ;
  assign n23565 = n18367 ^ n391 ^ 1'b0 ;
  assign n23566 = n23564 & n23565 ;
  assign n23567 = n23566 ^ n2596 ^ 1'b0 ;
  assign n23568 = n7930 & ~n23567 ;
  assign n23569 = n1695 | n15076 ;
  assign n23570 = n4036 & n23569 ;
  assign n23571 = n23570 ^ n1962 ^ 1'b0 ;
  assign n23572 = n23571 ^ n3143 ^ 1'b0 ;
  assign n23573 = n23568 & n23572 ;
  assign n23574 = n4548 & ~n12030 ;
  assign n23575 = n8548 & n23574 ;
  assign n23576 = ~n10039 & n22614 ;
  assign n23577 = n23575 & n23576 ;
  assign n23578 = n20288 ^ n17768 ^ n11252 ;
  assign n23579 = n23230 ^ n21507 ^ 1'b0 ;
  assign n23580 = n8595 ^ n2067 ^ 1'b0 ;
  assign n23581 = n12071 | n23580 ;
  assign n23582 = ~n23512 & n23581 ;
  assign n23583 = ~n388 & n14510 ;
  assign n23584 = n2953 & n23583 ;
  assign n23585 = n5759 & ~n23584 ;
  assign n23586 = n18323 ^ n15884 ^ x126 ;
  assign n23587 = n13179 & n17457 ;
  assign n23588 = n7590 & n23587 ;
  assign n23589 = n1552 | n5492 ;
  assign n23590 = n16678 & ~n23589 ;
  assign n23591 = n23590 ^ n16918 ^ 1'b0 ;
  assign n23592 = n6985 ^ n6040 ^ 1'b0 ;
  assign n23593 = ( n5881 & n6946 ) | ( n5881 & n23592 ) | ( n6946 & n23592 ) ;
  assign n23594 = n3842 | n5791 ;
  assign n23595 = n23594 ^ n7802 ^ 1'b0 ;
  assign n23596 = n23595 ^ n2192 ^ 1'b0 ;
  assign n23597 = n4395 & ~n23596 ;
  assign n23598 = n22247 ^ n13005 ^ n6034 ;
  assign n23599 = n23598 ^ n21653 ^ 1'b0 ;
  assign n23600 = n1396 | n22364 ;
  assign n23601 = n23600 ^ n12717 ^ 1'b0 ;
  assign n23602 = n17915 ^ n15935 ^ 1'b0 ;
  assign n23605 = n4331 ^ x108 ^ 1'b0 ;
  assign n23606 = n15830 & n23605 ;
  assign n23603 = n3869 & ~n11853 ;
  assign n23604 = ( n5086 & ~n17208 ) | ( n5086 & n23603 ) | ( ~n17208 & n23603 ) ;
  assign n23607 = n23606 ^ n23604 ^ n17484 ;
  assign n23608 = n1370 & n9721 ;
  assign n23609 = n23608 ^ n12153 ^ n10798 ;
  assign n23610 = ~n2827 & n23609 ;
  assign n23611 = n12712 & n23610 ;
  assign n23612 = n6928 | n7816 ;
  assign n23613 = n3404 ^ n469 ^ 1'b0 ;
  assign n23614 = n8413 & ~n23613 ;
  assign n23615 = n12583 ^ n3215 ^ 1'b0 ;
  assign n23616 = n23614 & ~n23615 ;
  assign n23617 = n5962 & n23616 ;
  assign n23618 = ~n2257 & n6437 ;
  assign n23619 = n23618 ^ n20202 ^ 1'b0 ;
  assign n23620 = n20671 ^ n20116 ^ 1'b0 ;
  assign n23621 = n8288 & ~n23620 ;
  assign n23622 = n14710 ^ n11606 ^ 1'b0 ;
  assign n23623 = n12355 ^ n6907 ^ 1'b0 ;
  assign n23624 = n6124 | n23623 ;
  assign n23625 = n17209 ^ n17040 ^ 1'b0 ;
  assign n23626 = n13710 | n23625 ;
  assign n23627 = ( n10148 & ~n23624 ) | ( n10148 & n23626 ) | ( ~n23624 & n23626 ) ;
  assign n23628 = n4785 | n8911 ;
  assign n23629 = n23628 ^ n17144 ^ n3987 ;
  assign n23632 = ( n1680 & n9066 ) | ( n1680 & n11607 ) | ( n9066 & n11607 ) ;
  assign n23633 = n7308 & ~n7696 ;
  assign n23634 = n23632 & n23633 ;
  assign n23630 = n19886 ^ n19245 ^ 1'b0 ;
  assign n23631 = n13731 & n23630 ;
  assign n23635 = n23634 ^ n23631 ^ 1'b0 ;
  assign n23636 = n742 & n9813 ;
  assign n23637 = ( ~n377 & n9623 ) | ( ~n377 & n10730 ) | ( n9623 & n10730 ) ;
  assign n23638 = ~n11660 & n17456 ;
  assign n23639 = ~n23637 & n23638 ;
  assign n23640 = n1862 | n23639 ;
  assign n23641 = n14980 ^ n1541 ^ 1'b0 ;
  assign n23642 = ~n17451 & n21750 ;
  assign n23643 = n23642 ^ n4698 ^ 1'b0 ;
  assign n23644 = n2779 & ~n23643 ;
  assign n23645 = n12948 ^ n4180 ^ 1'b0 ;
  assign n23646 = n3212 & ~n23645 ;
  assign n23647 = n23646 ^ n3556 ^ n1761 ;
  assign n23648 = ~n2054 & n16511 ;
  assign n23649 = ~n853 & n3245 ;
  assign n23650 = n11957 ^ n8038 ^ 1'b0 ;
  assign n23651 = n12476 & ~n23650 ;
  assign n23652 = n21264 ^ n9913 ^ 1'b0 ;
  assign n23653 = n11473 ^ n8938 ^ 1'b0 ;
  assign n23654 = n2908 & n23653 ;
  assign n23655 = n2746 | n13798 ;
  assign n23656 = ( n2172 & n15096 ) | ( n2172 & ~n23655 ) | ( n15096 & ~n23655 ) ;
  assign n23657 = n3066 ^ n1167 ^ 1'b0 ;
  assign n23658 = ~n11291 & n16032 ;
  assign n23659 = n23658 ^ n4566 ^ 1'b0 ;
  assign n23660 = n12421 ^ n8236 ^ 1'b0 ;
  assign n23661 = n23659 & n23660 ;
  assign n23663 = x62 | n7305 ;
  assign n23662 = n172 & n10392 ;
  assign n23664 = n23663 ^ n23662 ^ 1'b0 ;
  assign n23665 = n10130 ^ n1616 ^ 1'b0 ;
  assign n23666 = n12422 & n23665 ;
  assign n23667 = n11677 ^ n4416 ^ n2863 ;
  assign n23668 = n5960 | n23667 ;
  assign n23669 = n10304 & n14931 ;
  assign n23670 = n23669 ^ n20388 ^ n11768 ;
  assign n23671 = n23668 & ~n23670 ;
  assign n23672 = ~n8212 & n13857 ;
  assign n23673 = n23672 ^ n11391 ^ 1'b0 ;
  assign n23674 = ~n22697 & n23673 ;
  assign n23675 = n13013 ^ n9408 ^ n3605 ;
  assign n23676 = n23674 | n23675 ;
  assign n23680 = n4906 & n6073 ;
  assign n23677 = ~n6135 & n7713 ;
  assign n23678 = n12025 & n23677 ;
  assign n23679 = ~n2563 & n23678 ;
  assign n23681 = n23680 ^ n23679 ^ 1'b0 ;
  assign n23682 = ( n2394 & ~n5203 ) | ( n2394 & n10791 ) | ( ~n5203 & n10791 ) ;
  assign n23683 = n8171 ^ n7887 ^ 1'b0 ;
  assign n23684 = ~n23682 & n23683 ;
  assign n23685 = n15793 ^ n292 ^ 1'b0 ;
  assign n23686 = n672 | n23685 ;
  assign n23687 = n2969 & ~n19934 ;
  assign n23688 = n23687 ^ n21673 ^ 1'b0 ;
  assign n23689 = n23688 ^ n2958 ^ 1'b0 ;
  assign n23690 = ~n23686 & n23689 ;
  assign n23691 = n1933 | n5389 ;
  assign n23692 = ~n815 & n23691 ;
  assign n23693 = n16924 ^ n4013 ^ 1'b0 ;
  assign n23694 = n3997 ^ n1787 ^ 1'b0 ;
  assign n23695 = n20655 & n23694 ;
  assign n23697 = ~n11756 & n13325 ;
  assign n23698 = n12458 ^ n2670 ^ 1'b0 ;
  assign n23699 = n23697 | n23698 ;
  assign n23700 = n11488 | n23699 ;
  assign n23696 = n3450 & ~n16629 ;
  assign n23701 = n23700 ^ n23696 ^ 1'b0 ;
  assign n23702 = n17981 ^ n1390 ^ 1'b0 ;
  assign n23703 = n21653 ^ n16291 ^ 1'b0 ;
  assign n23704 = n3478 & ~n8702 ;
  assign n23705 = ~n10834 & n23704 ;
  assign n23706 = n23705 ^ n6698 ^ 1'b0 ;
  assign n23707 = n23706 ^ n6437 ^ n2839 ;
  assign n23708 = n10526 | n21833 ;
  assign n23709 = n9628 & ~n23708 ;
  assign n23710 = n1412 | n23709 ;
  assign n23711 = n332 | n23710 ;
  assign n23712 = n6391 | n9046 ;
  assign n23713 = ~n4345 & n9269 ;
  assign n23714 = n3700 & ~n10806 ;
  assign n23715 = ~n4678 & n23714 ;
  assign n23716 = n2088 | n11571 ;
  assign n23717 = n19306 | n23716 ;
  assign n23719 = n2591 | n8119 ;
  assign n23718 = n4076 & n6073 ;
  assign n23720 = n23719 ^ n23718 ^ 1'b0 ;
  assign n23721 = n23720 ^ n3724 ^ 1'b0 ;
  assign n23722 = n23717 & ~n23721 ;
  assign n23723 = ( ~x102 & n4488 ) | ( ~x102 & n9167 ) | ( n4488 & n9167 ) ;
  assign n23724 = n2289 | n2399 ;
  assign n23725 = n23724 ^ n9768 ^ n7305 ;
  assign n23726 = n6310 & n18790 ;
  assign n23727 = n2874 & ~n3613 ;
  assign n23728 = n471 & n14685 ;
  assign n23729 = n23728 ^ x63 ^ 1'b0 ;
  assign n23730 = n23729 ^ n5133 ^ 1'b0 ;
  assign n23731 = n3610 & n23730 ;
  assign n23732 = ~n17821 & n23731 ;
  assign n23733 = ~n632 & n4244 ;
  assign n23734 = ~n12412 & n23733 ;
  assign n23735 = n23734 ^ n3930 ^ 1'b0 ;
  assign n23736 = n1973 | n22359 ;
  assign n23737 = n23736 ^ n4681 ^ 1'b0 ;
  assign n23738 = ~n7285 & n15962 ;
  assign n23739 = n23738 ^ n11665 ^ n11435 ;
  assign n23740 = n182 | n13919 ;
  assign n23741 = n16344 & ~n23740 ;
  assign n23742 = n21203 ^ n6640 ^ 1'b0 ;
  assign n23743 = n17342 | n23742 ;
  assign n23744 = n5462 | n23743 ;
  assign n23745 = n10363 & n23605 ;
  assign n23746 = n23745 ^ n6902 ^ 1'b0 ;
  assign n23747 = n2372 & ~n6006 ;
  assign n23748 = n6378 ^ n2078 ^ 1'b0 ;
  assign n23749 = n23748 ^ n17639 ^ n1863 ;
  assign n23750 = n4513 & n6626 ;
  assign n23751 = ~n5979 & n23750 ;
  assign n23752 = n1303 & n1920 ;
  assign n23753 = n23752 ^ n17264 ^ 1'b0 ;
  assign n23754 = n6053 | n9319 ;
  assign n23755 = ~n23753 & n23754 ;
  assign n23756 = n20287 ^ n13904 ^ 1'b0 ;
  assign n23757 = n4574 & n23756 ;
  assign n23758 = n15276 & n18238 ;
  assign n23759 = n16133 ^ n371 ^ 1'b0 ;
  assign n23760 = n13718 & n23759 ;
  assign n23763 = n8637 & ~n9841 ;
  assign n23764 = n11738 ^ n4216 ^ 1'b0 ;
  assign n23765 = n23763 & ~n23764 ;
  assign n23761 = n15588 & n23448 ;
  assign n23762 = n23761 ^ n4530 ^ 1'b0 ;
  assign n23766 = n23765 ^ n23762 ^ n143 ;
  assign n23767 = n16054 | n19165 ;
  assign n23768 = n23766 | n23767 ;
  assign n23769 = n22664 & ~n23768 ;
  assign n23771 = n5015 | n5646 ;
  assign n23772 = n672 | n23771 ;
  assign n23770 = n20746 | n22432 ;
  assign n23773 = n23772 ^ n23770 ^ 1'b0 ;
  assign n23774 = ( ~n1078 & n1512 ) | ( ~n1078 & n13766 ) | ( n1512 & n13766 ) ;
  assign n23776 = n768 ^ n475 ^ 1'b0 ;
  assign n23777 = n7472 & n23776 ;
  assign n23775 = n12215 & ~n17223 ;
  assign n23778 = n23777 ^ n23775 ^ 1'b0 ;
  assign n23779 = n23778 ^ n16428 ^ 1'b0 ;
  assign n23780 = n4216 ^ n2340 ^ 1'b0 ;
  assign n23781 = ~n6043 & n11736 ;
  assign n23782 = n23781 ^ n11674 ^ 1'b0 ;
  assign n23783 = ~n969 & n6300 ;
  assign n23784 = n5054 & ~n7704 ;
  assign n23785 = n23784 ^ n1155 ^ 1'b0 ;
  assign n23786 = ~n789 & n17930 ;
  assign n23787 = ~n15210 & n23786 ;
  assign n23788 = n9169 | n15260 ;
  assign n23789 = n14935 & n23788 ;
  assign n23790 = n23789 ^ n20703 ^ 1'b0 ;
  assign n23791 = n3331 ^ n444 ^ 1'b0 ;
  assign n23792 = ~n9671 & n17024 ;
  assign n23793 = n8582 ^ x50 ^ 1'b0 ;
  assign n23794 = n23793 ^ n23284 ^ n5812 ;
  assign n23795 = n12887 ^ n7086 ^ 1'b0 ;
  assign n23796 = n2283 & ~n19995 ;
  assign n23797 = n3992 & ~n23796 ;
  assign n23798 = n13087 & n23797 ;
  assign n23799 = n3700 & ~n6584 ;
  assign n23800 = n23799 ^ n13722 ^ 1'b0 ;
  assign n23801 = n5899 & ~n12291 ;
  assign n23802 = n22464 & n23801 ;
  assign n23803 = n23802 ^ n6171 ^ 1'b0 ;
  assign n23804 = n23800 | n23803 ;
  assign n23805 = n20850 ^ n7133 ^ 1'b0 ;
  assign n23806 = n1489 & n23805 ;
  assign n23807 = n12335 ^ n8485 ^ 1'b0 ;
  assign n23808 = ( n6633 & n15286 ) | ( n6633 & n19058 ) | ( n15286 & n19058 ) ;
  assign n23809 = n2969 | n23808 ;
  assign n23810 = ( ~n3647 & n7645 ) | ( ~n3647 & n23809 ) | ( n7645 & n23809 ) ;
  assign n23811 = n4353 & n19883 ;
  assign n23812 = n9103 & n23811 ;
  assign n23813 = n2204 & ~n14219 ;
  assign n23814 = n23813 ^ n11711 ^ 1'b0 ;
  assign n23815 = n10084 ^ n973 ^ 1'b0 ;
  assign n23816 = n22335 | n23815 ;
  assign n23817 = n12271 | n19461 ;
  assign n23818 = n20943 & ~n23817 ;
  assign n23819 = n10072 | n11054 ;
  assign n23820 = n412 & ~n23819 ;
  assign n23821 = n23820 ^ n6850 ^ n1659 ;
  assign n23822 = n21722 ^ n19644 ^ n17721 ;
  assign n23823 = ~n922 & n1497 ;
  assign n23825 = n3768 & ~n5028 ;
  assign n23826 = n23825 ^ n3615 ^ 1'b0 ;
  assign n23824 = n16689 | n19725 ;
  assign n23827 = n23826 ^ n23824 ^ 1'b0 ;
  assign n23828 = n12129 ^ n5245 ^ 1'b0 ;
  assign n23829 = ~n2561 & n3245 ;
  assign n23830 = n19623 ^ n19108 ^ 1'b0 ;
  assign n23831 = n10271 | n11053 ;
  assign n23832 = ~n5832 & n23831 ;
  assign n23833 = n23503 ^ n4068 ^ 1'b0 ;
  assign n23834 = n4194 ^ n1458 ^ 1'b0 ;
  assign n23835 = n21930 | n23834 ;
  assign n23836 = n11410 | n21659 ;
  assign n23837 = n3636 | n6550 ;
  assign n23838 = n8058 & ~n23837 ;
  assign n23839 = ~n7948 & n10990 ;
  assign n23840 = n23839 ^ n9823 ^ n3212 ;
  assign n23841 = n7076 | n15099 ;
  assign n23842 = n23840 | n23841 ;
  assign n23843 = n5419 ^ n1761 ^ 1'b0 ;
  assign n23844 = n18637 | n23843 ;
  assign n23845 = ( n15554 & n16834 ) | ( n15554 & n23844 ) | ( n16834 & n23844 ) ;
  assign n23846 = n1440 | n23845 ;
  assign n23847 = n6361 & ~n23846 ;
  assign n23848 = n2885 & ~n23847 ;
  assign n23849 = n23848 ^ n12622 ^ 1'b0 ;
  assign n23850 = n9651 ^ n7403 ^ 1'b0 ;
  assign n23851 = n10564 & ~n23850 ;
  assign n23852 = n560 & ~n4113 ;
  assign n23853 = ~n8296 & n23852 ;
  assign n23854 = ~n3948 & n23853 ;
  assign n23855 = n3571 | n4212 ;
  assign n23856 = n23855 ^ n3405 ^ 1'b0 ;
  assign n23857 = n2103 | n16416 ;
  assign n23858 = n23857 ^ n19011 ^ n9071 ;
  assign n23859 = ~n1711 & n18077 ;
  assign n23860 = n23859 ^ n6273 ^ 1'b0 ;
  assign n23861 = n5439 | n5904 ;
  assign n23862 = n23860 & ~n23861 ;
  assign n23863 = n11340 & ~n23862 ;
  assign n23864 = ~n19839 & n23863 ;
  assign n23865 = n1703 & ~n18096 ;
  assign n23866 = n23865 ^ n20069 ^ 1'b0 ;
  assign n23867 = n20208 & ~n23866 ;
  assign n23868 = n1279 & ~n19775 ;
  assign n23869 = ~n3518 & n7876 ;
  assign n23870 = n14134 ^ n8164 ^ 1'b0 ;
  assign n23871 = ( ~n10331 & n13712 ) | ( ~n10331 & n13713 ) | ( n13712 & n13713 ) ;
  assign n23872 = ~n2730 & n16413 ;
  assign n23873 = n7377 | n10884 ;
  assign n23874 = n18971 | n23873 ;
  assign n23875 = n930 & ~n18685 ;
  assign n23877 = n14154 ^ n8472 ^ 1'b0 ;
  assign n23878 = n2120 | n23877 ;
  assign n23876 = n21421 ^ n16498 ^ n15410 ;
  assign n23879 = n23878 ^ n23876 ^ 1'b0 ;
  assign n23880 = n23879 ^ n4204 ^ 1'b0 ;
  assign n23881 = n16095 & ~n16490 ;
  assign n23882 = n23881 ^ n2751 ^ 1'b0 ;
  assign n23883 = n2930 & ~n7412 ;
  assign n23884 = n23883 ^ n530 ^ 1'b0 ;
  assign n23885 = n18619 ^ n13766 ^ 1'b0 ;
  assign n23886 = ~n9779 & n23885 ;
  assign n23887 = n23884 & n23886 ;
  assign n23888 = n15223 ^ n7154 ^ 1'b0 ;
  assign n23889 = n2967 ^ n1433 ^ 1'b0 ;
  assign n23890 = n8691 & n16969 ;
  assign n23891 = n10265 & n23890 ;
  assign n23892 = n10677 & n23891 ;
  assign n23893 = n5897 & n21451 ;
  assign n23894 = n14969 & ~n23893 ;
  assign n23895 = n5277 & n23894 ;
  assign n23896 = n23895 ^ n5042 ^ 1'b0 ;
  assign n23897 = n6910 & n14554 ;
  assign n23898 = ~n5437 & n23897 ;
  assign n23899 = ( n2160 & n9200 ) | ( n2160 & ~n17945 ) | ( n9200 & ~n17945 ) ;
  assign n23900 = ~n8931 & n23899 ;
  assign n23901 = n19294 ^ n8948 ^ n3683 ;
  assign n23902 = n18843 ^ n8966 ^ 1'b0 ;
  assign n23903 = n978 & n1758 ;
  assign n23904 = ~n857 & n23903 ;
  assign n23905 = ~n3430 & n13780 ;
  assign n23906 = n6183 & n23905 ;
  assign n23907 = n6372 | n23906 ;
  assign n23908 = n23904 & ~n23907 ;
  assign n23909 = n18821 ^ n2450 ^ 1'b0 ;
  assign n23910 = ~n7800 & n19660 ;
  assign n23911 = n4450 & ~n21130 ;
  assign n23912 = n23911 ^ n4989 ^ 1'b0 ;
  assign n23913 = n14782 & ~n23912 ;
  assign n23914 = n20364 ^ n15347 ^ 1'b0 ;
  assign n23915 = n3790 & n9187 ;
  assign n23916 = n23915 ^ n5863 ^ 1'b0 ;
  assign n23917 = n4455 & ~n23916 ;
  assign n23918 = n13317 ^ n9127 ^ 1'b0 ;
  assign n23919 = ~n17855 & n23918 ;
  assign n23920 = ~n12414 & n22122 ;
  assign n23921 = n23920 ^ n507 ^ 1'b0 ;
  assign n23922 = n1714 | n8147 ;
  assign n23923 = n10732 & ~n23922 ;
  assign n23924 = n6088 & ~n23923 ;
  assign n23925 = n1076 & n23924 ;
  assign n23926 = n1481 & n4927 ;
  assign n23927 = n15299 & n23926 ;
  assign n23928 = n23925 & n23927 ;
  assign n23929 = n236 | n9416 ;
  assign n23930 = n23929 ^ n14001 ^ 1'b0 ;
  assign n23931 = n23930 ^ n4168 ^ 1'b0 ;
  assign n23932 = ~n2281 & n9353 ;
  assign n23933 = n23932 ^ n9703 ^ 1'b0 ;
  assign n23934 = n12313 ^ n4884 ^ 1'b0 ;
  assign n23935 = ~n15647 & n23934 ;
  assign n23936 = ~n9182 & n12077 ;
  assign n23939 = n5893 ^ n3248 ^ 1'b0 ;
  assign n23937 = n3698 & n5955 ;
  assign n23938 = ~n3393 & n23937 ;
  assign n23940 = n23939 ^ n23938 ^ n2014 ;
  assign n23941 = ~n3203 & n9037 ;
  assign n23942 = n15698 ^ n272 ^ 1'b0 ;
  assign n23943 = n10384 & ~n23942 ;
  assign n23944 = n1470 & ~n4628 ;
  assign n23945 = ~n15698 & n23944 ;
  assign n23946 = n3078 & ~n23427 ;
  assign n23947 = n11116 ^ n5744 ^ 1'b0 ;
  assign n23948 = n8984 & ~n23947 ;
  assign n23949 = n9089 & n23948 ;
  assign n23950 = n13798 ^ n937 ^ 1'b0 ;
  assign n23951 = n7951 | n23950 ;
  assign n23952 = n18517 ^ n9418 ^ 1'b0 ;
  assign n23953 = ~n3719 & n5511 ;
  assign n23954 = n4323 & n23953 ;
  assign n23955 = ~n11291 & n23954 ;
  assign n23956 = n23952 & n23955 ;
  assign n23957 = x25 & n2156 ;
  assign n23958 = ~n569 & n11290 ;
  assign n23959 = ~n3401 & n23958 ;
  assign n23960 = n19839 & ~n23959 ;
  assign n23961 = n23960 ^ n17325 ^ 1'b0 ;
  assign n23962 = n10951 ^ n2910 ^ 1'b0 ;
  assign n23963 = n1568 & ~n15217 ;
  assign n23964 = n1136 & ~n12057 ;
  assign n23965 = ~n1909 & n11324 ;
  assign n23966 = n21302 & n23965 ;
  assign n23967 = n10988 ^ n10985 ^ 1'b0 ;
  assign n23968 = n17434 | n23967 ;
  assign n23969 = n1270 & ~n23968 ;
  assign n23970 = n4216 & ~n4592 ;
  assign n23971 = n5057 & n8242 ;
  assign n23972 = ( n18663 & n23440 ) | ( n18663 & n23971 ) | ( n23440 & n23971 ) ;
  assign n23973 = n4204 ^ n3083 ^ 1'b0 ;
  assign n23974 = n4319 & n23973 ;
  assign n23975 = n18729 | n23974 ;
  assign n23976 = n137 | n1392 ;
  assign n23977 = n23976 ^ n11292 ^ 1'b0 ;
  assign n23978 = n4382 & n4824 ;
  assign n23979 = ~n5106 & n23978 ;
  assign n23980 = n18401 & ~n23979 ;
  assign n23981 = ~n1735 & n23980 ;
  assign n23982 = n773 & n23981 ;
  assign n23983 = n2331 & n9975 ;
  assign n23984 = n23983 ^ n1904 ^ 1'b0 ;
  assign n23985 = n4305 ^ n3972 ^ 1'b0 ;
  assign n23986 = ( ~n2714 & n12642 ) | ( ~n2714 & n14777 ) | ( n12642 & n14777 ) ;
  assign n23987 = ( n4966 & ~n10775 ) | ( n4966 & n23986 ) | ( ~n10775 & n23986 ) ;
  assign n23988 = ~n12420 & n19324 ;
  assign n23989 = n10665 & n11811 ;
  assign n23990 = n23989 ^ n15479 ^ n3204 ;
  assign n23991 = ( n11010 & n23988 ) | ( n11010 & n23990 ) | ( n23988 & n23990 ) ;
  assign n23992 = n7050 ^ n5486 ^ 1'b0 ;
  assign n23993 = n5119 & n23992 ;
  assign n23994 = n16300 | n23993 ;
  assign n23995 = n7643 & n12049 ;
  assign n23996 = n3202 & n23995 ;
  assign n23997 = n2948 & ~n18253 ;
  assign n23998 = ( ~n3861 & n4315 ) | ( ~n3861 & n19080 ) | ( n4315 & n19080 ) ;
  assign n23999 = n23998 ^ n8331 ^ 1'b0 ;
  assign n24000 = ~n222 & n23999 ;
  assign n24001 = n10216 ^ n9006 ^ 1'b0 ;
  assign n24002 = n10011 | n24001 ;
  assign n24003 = n20726 | n24002 ;
  assign n24004 = n1509 | n11942 ;
  assign n24005 = n24004 ^ n14995 ^ 1'b0 ;
  assign n24006 = n10271 & ~n19944 ;
  assign n24007 = n24006 ^ n7644 ^ 1'b0 ;
  assign n24008 = n8227 & ~n10780 ;
  assign n24009 = n15467 & n24008 ;
  assign n24010 = n24009 ^ n18799 ^ 1'b0 ;
  assign n24011 = n389 | n16539 ;
  assign n24012 = n14512 & n24011 ;
  assign n24013 = n18326 ^ n2031 ^ 1'b0 ;
  assign n24014 = n14028 & n24013 ;
  assign n24015 = n1970 & ~n3270 ;
  assign n24016 = n24015 ^ n14263 ^ 1'b0 ;
  assign n24017 = ~n833 & n4145 ;
  assign n24018 = n1761 & n14808 ;
  assign n24019 = n24018 ^ n11609 ^ 1'b0 ;
  assign n24020 = ~n19256 & n24019 ;
  assign n24021 = n855 & n24020 ;
  assign n24023 = n9186 & ~n13337 ;
  assign n24024 = n17060 & n24023 ;
  assign n24022 = ~n12658 & n14414 ;
  assign n24025 = n24024 ^ n24022 ^ 1'b0 ;
  assign n24026 = ~n4227 & n10547 ;
  assign n24027 = n16468 & n24026 ;
  assign n24028 = n24027 ^ n15917 ^ 1'b0 ;
  assign n24029 = n13450 ^ n12505 ^ n6386 ;
  assign n24030 = n7809 | n12410 ;
  assign n24032 = n2302 & ~n2615 ;
  assign n24033 = ( ~n22001 & n23012 ) | ( ~n22001 & n24032 ) | ( n23012 & n24032 ) ;
  assign n24031 = n5402 & n10204 ;
  assign n24034 = n24033 ^ n24031 ^ 1'b0 ;
  assign n24035 = n6529 & ~n23116 ;
  assign n24036 = n1128 & n4304 ;
  assign n24037 = n24036 ^ n17444 ^ 1'b0 ;
  assign n24038 = n10499 ^ n6850 ^ 1'b0 ;
  assign n24039 = n1757 & n24038 ;
  assign n24040 = n24039 ^ n2108 ^ 1'b0 ;
  assign n24041 = n3616 & ~n24040 ;
  assign n24042 = n3420 & n19820 ;
  assign n24043 = n4493 & n24042 ;
  assign n24044 = ~n2414 & n8061 ;
  assign n24045 = n24044 ^ n7297 ^ 1'b0 ;
  assign n24046 = ( n2948 & n7980 ) | ( n2948 & n24045 ) | ( n7980 & n24045 ) ;
  assign n24047 = n9458 ^ n598 ^ 1'b0 ;
  assign n24048 = n3465 | n10463 ;
  assign n24049 = n2361 | n24048 ;
  assign n24050 = n11228 | n22439 ;
  assign n24051 = n994 | n3376 ;
  assign n24052 = n12475 & ~n24051 ;
  assign n24053 = n2575 | n23748 ;
  assign n24054 = n24052 & ~n24053 ;
  assign n24055 = n2031 & n4722 ;
  assign n24056 = ~n468 & n24055 ;
  assign n24057 = n8852 | n24056 ;
  assign n24058 = n1793 | n24057 ;
  assign n24059 = n23132 ^ n2759 ^ n1192 ;
  assign n24060 = n1248 | n13982 ;
  assign n24061 = n7542 & n21456 ;
  assign n24062 = n13238 & n19419 ;
  assign n24063 = n24062 ^ n23284 ^ 1'b0 ;
  assign n24064 = ~n8452 & n11272 ;
  assign n24065 = n188 | n2494 ;
  assign n24066 = n24065 ^ n21479 ^ 1'b0 ;
  assign n24067 = n5390 & n8106 ;
  assign n24069 = n17155 ^ n13788 ^ n10739 ;
  assign n24070 = n5466 | n8956 ;
  assign n24071 = n24069 | n24070 ;
  assign n24068 = n15822 | n22184 ;
  assign n24072 = n24071 ^ n24068 ^ 1'b0 ;
  assign n24073 = n5510 | n24072 ;
  assign n24074 = n11010 & ~n24073 ;
  assign n24075 = n10545 ^ n9796 ^ 1'b0 ;
  assign n24076 = n11067 ^ n4683 ^ n1816 ;
  assign n24077 = n8996 & ~n11750 ;
  assign n24078 = ~n4919 & n11638 ;
  assign n24079 = n24078 ^ n16428 ^ 1'b0 ;
  assign n24080 = n21824 & ~n24079 ;
  assign n24081 = n9460 | n21912 ;
  assign n24082 = ~n1701 & n3659 ;
  assign n24083 = n24082 ^ n5974 ^ 1'b0 ;
  assign n24084 = ~n2412 & n24073 ;
  assign n24085 = n1788 & ~n4887 ;
  assign n24086 = n14413 ^ n3226 ^ 1'b0 ;
  assign n24087 = n1680 | n2812 ;
  assign n24088 = n24087 ^ n10046 ^ 1'b0 ;
  assign n24089 = ~n24086 & n24088 ;
  assign n24090 = n23537 ^ n14877 ^ 1'b0 ;
  assign n24091 = n7920 | n9066 ;
  assign n24092 = ( ~n14551 & n15621 ) | ( ~n14551 & n23449 ) | ( n15621 & n23449 ) ;
  assign n24093 = n1003 & n1431 ;
  assign n24094 = n4295 & ~n15099 ;
  assign n24095 = n24094 ^ n23638 ^ 1'b0 ;
  assign n24096 = n9446 ^ n9046 ^ 1'b0 ;
  assign n24097 = n1500 | n16285 ;
  assign n24098 = n24096 & ~n24097 ;
  assign n24101 = ~n9649 & n13670 ;
  assign n24102 = n5911 & n24101 ;
  assign n24099 = n5507 ^ x126 ^ 1'b0 ;
  assign n24100 = ~n21900 & n24099 ;
  assign n24103 = n24102 ^ n24100 ^ 1'b0 ;
  assign n24104 = n573 | n24103 ;
  assign n24105 = n13654 ^ n9008 ^ 1'b0 ;
  assign n24106 = n16449 ^ n11711 ^ 1'b0 ;
  assign n24107 = n3289 | n24106 ;
  assign n24108 = n24107 ^ n11719 ^ 1'b0 ;
  assign n24109 = n24105 | n24108 ;
  assign n24110 = n3605 & n15943 ;
  assign n24111 = n4912 & n22913 ;
  assign n24112 = n24111 ^ n10100 ^ 1'b0 ;
  assign n24113 = n5843 & ~n6718 ;
  assign n24114 = n24113 ^ n15615 ^ 1'b0 ;
  assign n24115 = n24112 & ~n24114 ;
  assign n24116 = n227 & ~n23894 ;
  assign n24117 = n15303 ^ n12402 ^ 1'b0 ;
  assign n24118 = n17194 & n24117 ;
  assign n24119 = n23163 | n24118 ;
  assign n24120 = n8543 ^ n4917 ^ 1'b0 ;
  assign n24121 = n2172 ^ n838 ^ 1'b0 ;
  assign n24122 = ~n6520 & n15602 ;
  assign n24123 = n11750 ^ n8910 ^ 1'b0 ;
  assign n24124 = n24122 & n24123 ;
  assign n24125 = n6340 & n10024 ;
  assign n24126 = n24125 ^ n18450 ^ n5715 ;
  assign n24128 = ~n4969 & n18637 ;
  assign n24127 = n2174 & n2889 ;
  assign n24129 = n24128 ^ n24127 ^ 1'b0 ;
  assign n24130 = ~n16768 & n24129 ;
  assign n24131 = ~n2756 & n10632 ;
  assign n24132 = ~n374 & n24131 ;
  assign n24133 = n1287 | n2859 ;
  assign n24134 = n24133 ^ n16729 ^ 1'b0 ;
  assign n24135 = n17778 ^ n16075 ^ n11318 ;
  assign n24136 = n240 & ~n11798 ;
  assign n24137 = n24136 ^ n3193 ^ 1'b0 ;
  assign n24138 = n24135 & n24137 ;
  assign n24139 = n3222 | n12289 ;
  assign n24140 = ~n364 & n4604 ;
  assign n24141 = n13819 ^ n5642 ^ 1'b0 ;
  assign n24142 = ~n19626 & n24141 ;
  assign n24143 = n1600 & n19253 ;
  assign n24144 = n1535 & n24143 ;
  assign n24145 = n19903 & n24144 ;
  assign n24146 = n7052 & ~n18116 ;
  assign n24147 = n7393 | n18247 ;
  assign n24148 = n24147 ^ n2228 ^ 1'b0 ;
  assign n24149 = n9498 & ~n11952 ;
  assign n24150 = ~n24148 & n24149 ;
  assign n24151 = n4892 ^ n3386 ^ 1'b0 ;
  assign n24152 = n14781 & n24151 ;
  assign n24153 = n15793 ^ n2928 ^ 1'b0 ;
  assign n24154 = ~n12799 & n24153 ;
  assign n24155 = n1959 & n3284 ;
  assign n24156 = n24155 ^ n23334 ^ 1'b0 ;
  assign n24157 = ~n12561 & n22420 ;
  assign n24158 = n24157 ^ n22171 ^ 1'b0 ;
  assign n24160 = n17120 ^ n16587 ^ n10683 ;
  assign n24159 = n5669 & n12998 ;
  assign n24161 = n24160 ^ n24159 ^ 1'b0 ;
  assign n24162 = n21964 ^ n3290 ^ 1'b0 ;
  assign n24163 = n19203 & n24162 ;
  assign n24164 = n24163 ^ n22322 ^ 1'b0 ;
  assign n24165 = n8840 & ~n24164 ;
  assign n24166 = ~n4596 & n20404 ;
  assign n24167 = n14520 ^ n10522 ^ n8982 ;
  assign n24170 = n1476 | n2769 ;
  assign n24171 = n4395 | n24170 ;
  assign n24168 = n11993 & n17615 ;
  assign n24169 = ~n4319 & n24168 ;
  assign n24172 = n24171 ^ n24169 ^ 1'b0 ;
  assign n24173 = n1511 & n2195 ;
  assign n24174 = ~n2445 & n24173 ;
  assign n24175 = n11561 | n17895 ;
  assign n24176 = n13475 & n14865 ;
  assign n24177 = n10300 ^ n1331 ^ 1'b0 ;
  assign n24178 = n1512 & ~n24177 ;
  assign n24179 = n24178 ^ n3131 ^ 1'b0 ;
  assign n24180 = n2351 & ~n9358 ;
  assign n24181 = n3537 & n24180 ;
  assign n24182 = n24181 ^ n3130 ^ 1'b0 ;
  assign n24183 = n24182 ^ n23556 ^ n8908 ;
  assign n24184 = ~n266 & n14038 ;
  assign n24185 = ~n11382 & n24184 ;
  assign n24186 = n17824 & n24185 ;
  assign n24187 = n10499 ^ n6551 ^ 1'b0 ;
  assign n24188 = n19143 | n24187 ;
  assign n24189 = n24188 ^ n18344 ^ 1'b0 ;
  assign n24190 = n24189 ^ n20969 ^ 1'b0 ;
  assign n24191 = n11348 | n14382 ;
  assign n24192 = n9632 | n22893 ;
  assign n24193 = n9942 ^ n7777 ^ 1'b0 ;
  assign n24194 = ~n17085 & n24193 ;
  assign n24195 = n4653 | n5048 ;
  assign n24196 = n14126 & ~n24195 ;
  assign n24197 = n24196 ^ n20015 ^ 1'b0 ;
  assign n24198 = n24197 ^ n4403 ^ 1'b0 ;
  assign n24199 = n18729 | n18753 ;
  assign n24200 = n8630 & ~n19013 ;
  assign n24201 = ~n14085 & n24200 ;
  assign n24202 = n19805 ^ n1666 ^ 1'b0 ;
  assign n24203 = n134 & n4056 ;
  assign n24206 = n10136 & ~n12344 ;
  assign n24207 = n24206 ^ n20672 ^ 1'b0 ;
  assign n24204 = n7716 | n18470 ;
  assign n24205 = n24204 ^ n175 ^ 1'b0 ;
  assign n24208 = n24207 ^ n24205 ^ 1'b0 ;
  assign n24210 = n6062 ^ n5804 ^ 1'b0 ;
  assign n24211 = n1325 | n24210 ;
  assign n24209 = n5787 & ~n8556 ;
  assign n24212 = n24211 ^ n24209 ^ 1'b0 ;
  assign n24213 = n18517 ^ n4468 ^ 1'b0 ;
  assign n24214 = n9882 | n22744 ;
  assign n24215 = n18906 | n24214 ;
  assign n24216 = n560 & n8077 ;
  assign n24217 = ~n17547 & n24216 ;
  assign n24218 = n4334 & n14160 ;
  assign n24219 = ~n455 & n11191 ;
  assign n24220 = n24219 ^ n18663 ^ 1'b0 ;
  assign n24221 = ~n20223 & n24220 ;
  assign n24222 = n24221 ^ n15847 ^ 1'b0 ;
  assign n24223 = n5079 & ~n9253 ;
  assign n24224 = n10808 & n24223 ;
  assign n24225 = n2436 ^ n2386 ^ 1'b0 ;
  assign n24226 = n24224 | n24225 ;
  assign n24227 = n6036 & ~n24226 ;
  assign n24228 = n10685 ^ n3219 ^ 1'b0 ;
  assign n24229 = ~n1805 & n24228 ;
  assign n24230 = n5170 ^ n2951 ^ 1'b0 ;
  assign n24231 = n5517 & ~n24230 ;
  assign n24232 = ( n10758 & ~n17405 ) | ( n10758 & n24231 ) | ( ~n17405 & n24231 ) ;
  assign n24233 = n5220 & ~n8146 ;
  assign n24234 = n8146 & n24233 ;
  assign n24235 = n7617 & ~n24234 ;
  assign n24236 = n14610 | n24235 ;
  assign n24237 = n24236 ^ n13840 ^ 1'b0 ;
  assign n24238 = n5439 | n7959 ;
  assign n24239 = n24238 ^ n12816 ^ 1'b0 ;
  assign n24240 = ~n637 & n22371 ;
  assign n24241 = n24240 ^ n1907 ^ 1'b0 ;
  assign n24242 = n22007 ^ n1190 ^ 1'b0 ;
  assign n24243 = n23427 | n24242 ;
  assign n24244 = n24243 ^ n1143 ^ 1'b0 ;
  assign n24245 = n5531 | n8430 ;
  assign n24246 = n152 | n7037 ;
  assign n24247 = n24246 ^ n22447 ^ 1'b0 ;
  assign n24248 = n21663 ^ n8092 ^ 1'b0 ;
  assign n24249 = n8584 & n9299 ;
  assign n24250 = n24249 ^ n7057 ^ 1'b0 ;
  assign n24251 = x6 & n24250 ;
  assign n24252 = ~n1237 & n2920 ;
  assign n24253 = n24252 ^ n6891 ^ 1'b0 ;
  assign n24254 = n23857 & n24253 ;
  assign n24255 = n3702 ^ n1761 ^ 1'b0 ;
  assign n24256 = ( n5345 & n12880 ) | ( n5345 & ~n24255 ) | ( n12880 & ~n24255 ) ;
  assign n24257 = n14680 ^ n14048 ^ n13274 ;
  assign n24258 = n13596 ^ n6455 ^ 1'b0 ;
  assign n24259 = n4917 & n24258 ;
  assign n24260 = n1769 | n18790 ;
  assign n24261 = n24260 ^ n15085 ^ 1'b0 ;
  assign n24262 = n1172 & ~n24261 ;
  assign n24263 = n24262 ^ n860 ^ 1'b0 ;
  assign n24264 = x115 & ~n7279 ;
  assign n24265 = n24264 ^ n849 ^ 1'b0 ;
  assign n24266 = n702 & n11740 ;
  assign n24267 = n24266 ^ n9428 ^ 1'b0 ;
  assign n24268 = n24265 | n24267 ;
  assign n24269 = n17007 ^ n6899 ^ 1'b0 ;
  assign n24270 = ~n7649 & n13846 ;
  assign n24271 = n24270 ^ n198 ^ 1'b0 ;
  assign n24272 = n24271 ^ n22969 ^ n2349 ;
  assign n24273 = ( n9950 & n10320 ) | ( n9950 & ~n10321 ) | ( n10320 & ~n10321 ) ;
  assign n24274 = ~n490 & n13460 ;
  assign n24275 = n12866 ^ n2577 ^ 1'b0 ;
  assign n24276 = n24274 & n24275 ;
  assign n24277 = ( n7556 & n9190 ) | ( n7556 & ~n12564 ) | ( n9190 & ~n12564 ) ;
  assign n24278 = n24277 ^ n19735 ^ 1'b0 ;
  assign n24279 = n22576 & ~n24278 ;
  assign n24280 = n7469 & n24279 ;
  assign n24281 = n21562 ^ n16244 ^ 1'b0 ;
  assign n24282 = ~n20330 & n24281 ;
  assign n24283 = n4601 & ~n15024 ;
  assign n24284 = n24283 ^ n5764 ^ 1'b0 ;
  assign n24285 = n2527 & ~n14237 ;
  assign n24286 = n6773 & n13709 ;
  assign n24287 = n9671 & n15769 ;
  assign n24288 = n24287 ^ n21718 ^ n9527 ;
  assign n24289 = n18535 ^ n4201 ^ 1'b0 ;
  assign n24292 = ~n2029 & n2561 ;
  assign n24293 = n24292 ^ n2227 ^ 1'b0 ;
  assign n24290 = n1252 & n16166 ;
  assign n24291 = n24290 ^ n3246 ^ 1'b0 ;
  assign n24294 = n24293 ^ n24291 ^ 1'b0 ;
  assign n24295 = ~n21383 & n22979 ;
  assign n24296 = n24295 ^ n6252 ^ 1'b0 ;
  assign n24297 = n5398 ^ n3830 ^ 1'b0 ;
  assign n24298 = ~n15508 & n24297 ;
  assign n24299 = n4623 | n23808 ;
  assign n24301 = n11890 ^ n4428 ^ 1'b0 ;
  assign n24302 = ( ~n676 & n1611 ) | ( ~n676 & n24301 ) | ( n1611 & n24301 ) ;
  assign n24300 = n22434 & ~n24027 ;
  assign n24303 = n24302 ^ n24300 ^ 1'b0 ;
  assign n24305 = n19321 ^ n7595 ^ 1'b0 ;
  assign n24304 = n2882 & ~n8297 ;
  assign n24306 = n24305 ^ n24304 ^ 1'b0 ;
  assign n24307 = n1028 & ~n24306 ;
  assign n24308 = n14489 ^ n4208 ^ 1'b0 ;
  assign n24309 = n2778 & ~n24308 ;
  assign n24310 = n8020 & n24309 ;
  assign n24311 = ( n2365 & n10186 ) | ( n2365 & n24310 ) | ( n10186 & n24310 ) ;
  assign n24315 = n6568 ^ n4887 ^ n3734 ;
  assign n24313 = n9349 ^ n993 ^ 1'b0 ;
  assign n24314 = n324 | n24313 ;
  assign n24316 = n24315 ^ n24314 ^ 1'b0 ;
  assign n24312 = ( n13298 & ~n15229 ) | ( n13298 & n19540 ) | ( ~n15229 & n19540 ) ;
  assign n24317 = n24316 ^ n24312 ^ 1'b0 ;
  assign n24318 = n5657 & n10161 ;
  assign n24319 = n12281 | n24318 ;
  assign n24320 = n5537 | n24319 ;
  assign n24321 = n3778 | n14833 ;
  assign n24322 = n3745 & ~n24321 ;
  assign n24323 = n4423 & n5828 ;
  assign n24324 = n3778 & n24323 ;
  assign n24325 = n24324 ^ n12260 ^ 1'b0 ;
  assign n24326 = n1291 & n24325 ;
  assign n24327 = n15400 & ~n20743 ;
  assign n24328 = n21674 ^ x1 ^ 1'b0 ;
  assign n24329 = n901 & n6396 ;
  assign n24330 = n24329 ^ n2956 ^ 1'b0 ;
  assign n24331 = n2266 & ~n24330 ;
  assign n24332 = ~n7185 & n22490 ;
  assign y0 = x2 ;
  assign y1 = x5 ;
  assign y2 = x6 ;
  assign y3 = x8 ;
  assign y4 = x9 ;
  assign y5 = x11 ;
  assign y6 = x13 ;
  assign y7 = x20 ;
  assign y8 = x26 ;
  assign y9 = x30 ;
  assign y10 = x31 ;
  assign y11 = x32 ;
  assign y12 = x37 ;
  assign y13 = x43 ;
  assign y14 = x44 ;
  assign y15 = x47 ;
  assign y16 = x49 ;
  assign y17 = x51 ;
  assign y18 = x57 ;
  assign y19 = x61 ;
  assign y20 = x70 ;
  assign y21 = x71 ;
  assign y22 = x75 ;
  assign y23 = x76 ;
  assign y24 = x78 ;
  assign y25 = x80 ;
  assign y26 = x81 ;
  assign y27 = x85 ;
  assign y28 = x88 ;
  assign y29 = x91 ;
  assign y30 = x92 ;
  assign y31 = x97 ;
  assign y32 = x98 ;
  assign y33 = x105 ;
  assign y34 = x108 ;
  assign y35 = x110 ;
  assign y36 = x111 ;
  assign y37 = x113 ;
  assign y38 = x116 ;
  assign y39 = x117 ;
  assign y40 = x118 ;
  assign y41 = x121 ;
  assign y42 = x123 ;
  assign y43 = x125 ;
  assign y44 = n129 ;
  assign y45 = ~n131 ;
  assign y46 = ~1'b0 ;
  assign y47 = n133 ;
  assign y48 = n134 ;
  assign y49 = ~1'b0 ;
  assign y50 = n138 ;
  assign y51 = n139 ;
  assign y52 = ~n141 ;
  assign y53 = ~1'b0 ;
  assign y54 = n144 ;
  assign y55 = ~n145 ;
  assign y56 = ~n147 ;
  assign y57 = ~n150 ;
  assign y58 = ~n154 ;
  assign y59 = n157 ;
  assign y60 = ~n159 ;
  assign y61 = n161 ;
  assign y62 = n163 ;
  assign y63 = ~n166 ;
  assign y64 = ~1'b0 ;
  assign y65 = ~n174 ;
  assign y66 = ~n177 ;
  assign y67 = ~n182 ;
  assign y68 = ~n184 ;
  assign y69 = ~n188 ;
  assign y70 = n190 ;
  assign y71 = ~n194 ;
  assign y72 = n195 ;
  assign y73 = ~1'b0 ;
  assign y74 = n196 ;
  assign y75 = ~n202 ;
  assign y76 = n205 ;
  assign y77 = n210 ;
  assign y78 = ~n218 ;
  assign y79 = ~n220 ;
  assign y80 = ~1'b0 ;
  assign y81 = ~1'b0 ;
  assign y82 = ~n224 ;
  assign y83 = ~1'b0 ;
  assign y84 = n225 ;
  assign y85 = n227 ;
  assign y86 = n231 ;
  assign y87 = ~n236 ;
  assign y88 = ~n238 ;
  assign y89 = ~1'b0 ;
  assign y90 = n246 ;
  assign y91 = ~n250 ;
  assign y92 = ~n252 ;
  assign y93 = ~1'b0 ;
  assign y94 = n255 ;
  assign y95 = ~n256 ;
  assign y96 = ~1'b0 ;
  assign y97 = n257 ;
  assign y98 = ~n260 ;
  assign y99 = ~1'b0 ;
  assign y100 = n261 ;
  assign y101 = n276 ;
  assign y102 = n277 ;
  assign y103 = ~n283 ;
  assign y104 = ~1'b0 ;
  assign y105 = ~n285 ;
  assign y106 = ~1'b0 ;
  assign y107 = ~1'b0 ;
  assign y108 = ~n287 ;
  assign y109 = n288 ;
  assign y110 = ~n293 ;
  assign y111 = n294 ;
  assign y112 = ~1'b0 ;
  assign y113 = n297 ;
  assign y114 = ~n301 ;
  assign y115 = ~n307 ;
  assign y116 = ~n313 ;
  assign y117 = ~1'b0 ;
  assign y118 = n321 ;
  assign y119 = ~n326 ;
  assign y120 = n331 ;
  assign y121 = n334 ;
  assign y122 = n336 ;
  assign y123 = n339 ;
  assign y124 = ~1'b0 ;
  assign y125 = ~1'b0 ;
  assign y126 = ~n344 ;
  assign y127 = ~n345 ;
  assign y128 = ~n351 ;
  assign y129 = ~n358 ;
  assign y130 = ~1'b0 ;
  assign y131 = n359 ;
  assign y132 = ~n361 ;
  assign y133 = ~n363 ;
  assign y134 = ~1'b0 ;
  assign y135 = ~n368 ;
  assign y136 = ~n369 ;
  assign y137 = n371 ;
  assign y138 = n374 ;
  assign y139 = n379 ;
  assign y140 = ~1'b0 ;
  assign y141 = ~n386 ;
  assign y142 = ~1'b0 ;
  assign y143 = ~n388 ;
  assign y144 = n392 ;
  assign y145 = n393 ;
  assign y146 = ~n398 ;
  assign y147 = n403 ;
  assign y148 = ~n404 ;
  assign y149 = n407 ;
  assign y150 = ~n414 ;
  assign y151 = ~n415 ;
  assign y152 = ~n417 ;
  assign y153 = ~n421 ;
  assign y154 = ~1'b0 ;
  assign y155 = n425 ;
  assign y156 = n428 ;
  assign y157 = n175 ;
  assign y158 = n438 ;
  assign y159 = ~n444 ;
  assign y160 = ~1'b0 ;
  assign y161 = n445 ;
  assign y162 = ~n448 ;
  assign y163 = 1'b0 ;
  assign y164 = ~n455 ;
  assign y165 = ~n456 ;
  assign y166 = ~1'b0 ;
  assign y167 = ~1'b0 ;
  assign y168 = n458 ;
  assign y169 = ~1'b0 ;
  assign y170 = ~1'b0 ;
  assign y171 = ~1'b0 ;
  assign y172 = ~n461 ;
  assign y173 = ~n468 ;
  assign y174 = ~n472 ;
  assign y175 = ~n476 ;
  assign y176 = n479 ;
  assign y177 = ~n481 ;
  assign y178 = ~n483 ;
  assign y179 = n486 ;
  assign y180 = ~n487 ;
  assign y181 = n489 ;
  assign y182 = n494 ;
  assign y183 = n496 ;
  assign y184 = n500 ;
  assign y185 = ~1'b0 ;
  assign y186 = ~1'b0 ;
  assign y187 = ~1'b0 ;
  assign y188 = n501 ;
  assign y189 = ~n504 ;
  assign y190 = n506 ;
  assign y191 = n519 ;
  assign y192 = ~1'b0 ;
  assign y193 = n527 ;
  assign y194 = ~1'b0 ;
  assign y195 = ~n531 ;
  assign y196 = ~1'b0 ;
  assign y197 = x1 ;
  assign y198 = ~1'b0 ;
  assign y199 = ~n533 ;
  assign y200 = ~n534 ;
  assign y201 = n538 ;
  assign y202 = ~1'b0 ;
  assign y203 = x6 ;
  assign y204 = ~n539 ;
  assign y205 = ~1'b0 ;
  assign y206 = n540 ;
  assign y207 = ~n541 ;
  assign y208 = ~n542 ;
  assign y209 = ~n545 ;
  assign y210 = ~n548 ;
  assign y211 = ~n551 ;
  assign y212 = n557 ;
  assign y213 = n489 ;
  assign y214 = n571 ;
  assign y215 = ~n577 ;
  assign y216 = ~1'b0 ;
  assign y217 = n578 ;
  assign y218 = n580 ;
  assign y219 = ~1'b0 ;
  assign y220 = n583 ;
  assign y221 = ~1'b0 ;
  assign y222 = n585 ;
  assign y223 = n591 ;
  assign y224 = ~n593 ;
  assign y225 = n597 ;
  assign y226 = ~n605 ;
  assign y227 = n612 ;
  assign y228 = ~n615 ;
  assign y229 = n616 ;
  assign y230 = ~1'b0 ;
  assign y231 = ~n623 ;
  assign y232 = ~1'b0 ;
  assign y233 = n627 ;
  assign y234 = n628 ;
  assign y235 = ~1'b0 ;
  assign y236 = ~1'b0 ;
  assign y237 = ~n630 ;
  assign y238 = n632 ;
  assign y239 = n634 ;
  assign y240 = ~1'b0 ;
  assign y241 = n636 ;
  assign y242 = ~1'b0 ;
  assign y243 = ~n641 ;
  assign y244 = ~n400 ;
  assign y245 = ~1'b0 ;
  assign y246 = n642 ;
  assign y247 = n649 ;
  assign y248 = ~n656 ;
  assign y249 = ~n660 ;
  assign y250 = ~n662 ;
  assign y251 = n632 ;
  assign y252 = n664 ;
  assign y253 = x70 ;
  assign y254 = ~1'b0 ;
  assign y255 = n163 ;
  assign y256 = n667 ;
  assign y257 = n671 ;
  assign y258 = n672 ;
  assign y259 = n674 ;
  assign y260 = ~1'b0 ;
  assign y261 = n675 ;
  assign y262 = ~n677 ;
  assign y263 = n678 ;
  assign y264 = ~n679 ;
  assign y265 = ~1'b0 ;
  assign y266 = ~n680 ;
  assign y267 = ~n683 ;
  assign y268 = ~n687 ;
  assign y269 = n676 ;
  assign y270 = n692 ;
  assign y271 = ~1'b0 ;
  assign y272 = n697 ;
  assign y273 = ~n701 ;
  assign y274 = n708 ;
  assign y275 = ~n710 ;
  assign y276 = n714 ;
  assign y277 = ~n718 ;
  assign y278 = n722 ;
  assign y279 = ~x6 ;
  assign y280 = ~1'b0 ;
  assign y281 = n725 ;
  assign y282 = ~1'b0 ;
  assign y283 = ~n726 ;
  assign y284 = n730 ;
  assign y285 = ~n732 ;
  assign y286 = ~1'b0 ;
  assign y287 = ~n737 ;
  assign y288 = ~1'b0 ;
  assign y289 = n738 ;
  assign y290 = n722 ;
  assign y291 = n741 ;
  assign y292 = n742 ;
  assign y293 = ~n745 ;
  assign y294 = ~n746 ;
  assign y295 = n747 ;
  assign y296 = ~1'b0 ;
  assign y297 = ~n751 ;
  assign y298 = ~n754 ;
  assign y299 = ~1'b0 ;
  assign y300 = n758 ;
  assign y301 = n762 ;
  assign y302 = ~1'b0 ;
  assign y303 = ~n766 ;
  assign y304 = n768 ;
  assign y305 = ~1'b0 ;
  assign y306 = n769 ;
  assign y307 = ~n770 ;
  assign y308 = n771 ;
  assign y309 = ~n777 ;
  assign y310 = ~1'b0 ;
  assign y311 = ~n779 ;
  assign y312 = ~1'b0 ;
  assign y313 = n781 ;
  assign y314 = ~n789 ;
  assign y315 = ~x98 ;
  assign y316 = ~1'b0 ;
  assign y317 = ~n796 ;
  assign y318 = 1'b0 ;
  assign y319 = n797 ;
  assign y320 = ~n802 ;
  assign y321 = n808 ;
  assign y322 = n809 ;
  assign y323 = n810 ;
  assign y324 = ~n811 ;
  assign y325 = ~n815 ;
  assign y326 = ~n816 ;
  assign y327 = n821 ;
  assign y328 = n822 ;
  assign y329 = n825 ;
  assign y330 = ~1'b0 ;
  assign y331 = ~1'b0 ;
  assign y332 = n838 ;
  assign y333 = ~1'b0 ;
  assign y334 = n840 ;
  assign y335 = ~1'b0 ;
  assign y336 = ~n841 ;
  assign y337 = n842 ;
  assign y338 = ~1'b0 ;
  assign y339 = n843 ;
  assign y340 = ~1'b0 ;
  assign y341 = n844 ;
  assign y342 = n847 ;
  assign y343 = n468 ;
  assign y344 = ~n852 ;
  assign y345 = n853 ;
  assign y346 = n857 ;
  assign y347 = ~n858 ;
  assign y348 = n719 ;
  assign y349 = n860 ;
  assign y350 = ~1'b0 ;
  assign y351 = ~n861 ;
  assign y352 = ~1'b0 ;
  assign y353 = n867 ;
  assign y354 = ~n871 ;
  assign y355 = ~n875 ;
  assign y356 = ~1'b0 ;
  assign y357 = ~1'b0 ;
  assign y358 = n876 ;
  assign y359 = n878 ;
  assign y360 = n882 ;
  assign y361 = ~1'b0 ;
  assign y362 = n884 ;
  assign y363 = n885 ;
  assign y364 = ~n890 ;
  assign y365 = ~1'b0 ;
  assign y366 = ~n892 ;
  assign y367 = ~n894 ;
  assign y368 = n897 ;
  assign y369 = ~n907 ;
  assign y370 = n911 ;
  assign y371 = ~1'b0 ;
  assign y372 = ~n913 ;
  assign y373 = ~n916 ;
  assign y374 = ~1'b0 ;
  assign y375 = ~1'b0 ;
  assign y376 = ~n922 ;
  assign y377 = n468 ;
  assign y378 = ~1'b0 ;
  assign y379 = ~n923 ;
  assign y380 = ~n926 ;
  assign y381 = 1'b0 ;
  assign y382 = ~1'b0 ;
  assign y383 = ~1'b0 ;
  assign y384 = n930 ;
  assign y385 = n323 ;
  assign y386 = ~n935 ;
  assign y387 = ~1'b0 ;
  assign y388 = n937 ;
  assign y389 = ~n939 ;
  assign y390 = ~n942 ;
  assign y391 = x83 ;
  assign y392 = ~n945 ;
  assign y393 = ~1'b0 ;
  assign y394 = ~n947 ;
  assign y395 = n951 ;
  assign y396 = ~1'b0 ;
  assign y397 = ~n952 ;
  assign y398 = ~n962 ;
  assign y399 = ~n964 ;
  assign y400 = n965 ;
  assign y401 = ~n973 ;
  assign y402 = n975 ;
  assign y403 = n982 ;
  assign y404 = n983 ;
  assign y405 = n986 ;
  assign y406 = ~n995 ;
  assign y407 = n997 ;
  assign y408 = ~n998 ;
  assign y409 = ~1'b0 ;
  assign y410 = ~n999 ;
  assign y411 = ~1'b0 ;
  assign y412 = n1003 ;
  assign y413 = ~n1011 ;
  assign y414 = ~n1013 ;
  assign y415 = ~n1019 ;
  assign y416 = ~n1024 ;
  assign y417 = n1026 ;
  assign y418 = n1031 ;
  assign y419 = ~n1038 ;
  assign y420 = ~n1039 ;
  assign y421 = ~n1040 ;
  assign y422 = ~n1042 ;
  assign y423 = n1045 ;
  assign y424 = ~1'b0 ;
  assign y425 = n1046 ;
  assign y426 = n1047 ;
  assign y427 = ~1'b0 ;
  assign y428 = ~n1053 ;
  assign y429 = n1054 ;
  assign y430 = ~n1057 ;
  assign y431 = ~1'b0 ;
  assign y432 = n1058 ;
  assign y433 = n1062 ;
  assign y434 = ~1'b0 ;
  assign y435 = ~n1064 ;
  assign y436 = ~n1065 ;
  assign y437 = n1067 ;
  assign y438 = n1068 ;
  assign y439 = ~1'b0 ;
  assign y440 = n709 ;
  assign y441 = ~1'b0 ;
  assign y442 = ~n1070 ;
  assign y443 = ~1'b0 ;
  assign y444 = n1071 ;
  assign y445 = ~1'b0 ;
  assign y446 = ~1'b0 ;
  assign y447 = ~1'b0 ;
  assign y448 = ~n1081 ;
  assign y449 = n1088 ;
  assign y450 = n1096 ;
  assign y451 = ~n1105 ;
  assign y452 = ~1'b0 ;
  assign y453 = 1'b0 ;
  assign y454 = ~1'b0 ;
  assign y455 = ~n1109 ;
  assign y456 = ~1'b0 ;
  assign y457 = ~n1111 ;
  assign y458 = ~n1117 ;
  assign y459 = ~1'b0 ;
  assign y460 = n1118 ;
  assign y461 = n1120 ;
  assign y462 = ~x75 ;
  assign y463 = ~n1129 ;
  assign y464 = n1132 ;
  assign y465 = ~1'b0 ;
  assign y466 = ~1'b0 ;
  assign y467 = n1135 ;
  assign y468 = n1137 ;
  assign y469 = ~1'b0 ;
  assign y470 = ~n1138 ;
  assign y471 = ~n297 ;
  assign y472 = n430 ;
  assign y473 = n1140 ;
  assign y474 = n1145 ;
  assign y475 = ~n1150 ;
  assign y476 = ~1'b0 ;
  assign y477 = ~n1157 ;
  assign y478 = ~n1164 ;
  assign y479 = ~n1166 ;
  assign y480 = ~1'b0 ;
  assign y481 = ~1'b0 ;
  assign y482 = ~n1169 ;
  assign y483 = n1170 ;
  assign y484 = ~1'b0 ;
  assign y485 = n1172 ;
  assign y486 = n1175 ;
  assign y487 = ~n1179 ;
  assign y488 = n1180 ;
  assign y489 = n1182 ;
  assign y490 = ~1'b0 ;
  assign y491 = n1183 ;
  assign y492 = n1189 ;
  assign y493 = ~1'b0 ;
  assign y494 = n1190 ;
  assign y495 = x34 ;
  assign y496 = ~1'b0 ;
  assign y497 = n1193 ;
  assign y498 = n1195 ;
  assign y499 = ~1'b0 ;
  assign y500 = ~1'b0 ;
  assign y501 = ~n1199 ;
  assign y502 = n1206 ;
  assign y503 = ~1'b0 ;
  assign y504 = ~n1208 ;
  assign y505 = ~n1211 ;
  assign y506 = ~n1213 ;
  assign y507 = n1215 ;
  assign y508 = ~n1219 ;
  assign y509 = n1222 ;
  assign y510 = ~1'b0 ;
  assign y511 = n1223 ;
  assign y512 = ~n1224 ;
  assign y513 = ~n1231 ;
  assign y514 = n1233 ;
  assign y515 = n1235 ;
  assign y516 = ~n1237 ;
  assign y517 = ~1'b0 ;
  assign y518 = n1242 ;
  assign y519 = n1244 ;
  assign y520 = ~1'b0 ;
  assign y521 = ~n1247 ;
  assign y522 = ~n1254 ;
  assign y523 = ~n1258 ;
  assign y524 = ~1'b0 ;
  assign y525 = n1259 ;
  assign y526 = ~n1261 ;
  assign y527 = ~1'b0 ;
  assign y528 = ~1'b0 ;
  assign y529 = n1264 ;
  assign y530 = n1266 ;
  assign y531 = n1271 ;
  assign y532 = ~n1273 ;
  assign y533 = ~n1276 ;
  assign y534 = ~1'b0 ;
  assign y535 = ~1'b0 ;
  assign y536 = ~1'b0 ;
  assign y537 = ~n1295 ;
  assign y538 = ~n1296 ;
  assign y539 = ~1'b0 ;
  assign y540 = ~n1304 ;
  assign y541 = ~n440 ;
  assign y542 = ~1'b0 ;
  assign y543 = ~1'b0 ;
  assign y544 = ~n1306 ;
  assign y545 = n1311 ;
  assign y546 = ~n1315 ;
  assign y547 = ~n1321 ;
  assign y548 = ~n1329 ;
  assign y549 = ~1'b0 ;
  assign y550 = ~1'b0 ;
  assign y551 = n1330 ;
  assign y552 = ~1'b0 ;
  assign y553 = n1333 ;
  assign y554 = n1340 ;
  assign y555 = n1341 ;
  assign y556 = n1351 ;
  assign y557 = ~1'b0 ;
  assign y558 = ~1'b0 ;
  assign y559 = ~1'b0 ;
  assign y560 = n1359 ;
  assign y561 = n1363 ;
  assign y562 = n1365 ;
  assign y563 = ~1'b0 ;
  assign y564 = ~1'b0 ;
  assign y565 = ~1'b0 ;
  assign y566 = ~n1367 ;
  assign y567 = n1370 ;
  assign y568 = ~1'b0 ;
  assign y569 = ~n1374 ;
  assign y570 = n1377 ;
  assign y571 = n1378 ;
  assign y572 = ~n1380 ;
  assign y573 = ~1'b0 ;
  assign y574 = ~1'b0 ;
  assign y575 = n468 ;
  assign y576 = ~1'b0 ;
  assign y577 = ~n1386 ;
  assign y578 = n1391 ;
  assign y579 = ~n1353 ;
  assign y580 = ~n1392 ;
  assign y581 = ~n1393 ;
  assign y582 = ~1'b0 ;
  assign y583 = n1394 ;
  assign y584 = ~1'b0 ;
  assign y585 = ~1'b0 ;
  assign y586 = ~n1396 ;
  assign y587 = ~n1398 ;
  assign y588 = ~n1401 ;
  assign y589 = n1405 ;
  assign y590 = ~1'b0 ;
  assign y591 = n1411 ;
  assign y592 = ~n1412 ;
  assign y593 = ~n1416 ;
  assign y594 = ~n1421 ;
  assign y595 = n1431 ;
  assign y596 = n1432 ;
  assign y597 = n157 ;
  assign y598 = ~1'b0 ;
  assign y599 = ~n1435 ;
  assign y600 = n1437 ;
  assign y601 = 1'b0 ;
  assign y602 = ~n1440 ;
  assign y603 = ~n1452 ;
  assign y604 = ~n1455 ;
  assign y605 = ~n1465 ;
  assign y606 = ~n1469 ;
  assign y607 = n1470 ;
  assign y608 = ~n1471 ;
  assign y609 = ~n1476 ;
  assign y610 = n1487 ;
  assign y611 = n1491 ;
  assign y612 = ~1'b0 ;
  assign y613 = n1493 ;
  assign y614 = ~n1502 ;
  assign y615 = ~1'b0 ;
  assign y616 = n1503 ;
  assign y617 = ~1'b0 ;
  assign y618 = n1507 ;
  assign y619 = ~n1509 ;
  assign y620 = ~1'b0 ;
  assign y621 = n1511 ;
  assign y622 = ~1'b0 ;
  assign y623 = ~1'b0 ;
  assign y624 = ~1'b0 ;
  assign y625 = ~1'b0 ;
  assign y626 = ~n1514 ;
  assign y627 = ~1'b0 ;
  assign y628 = 1'b0 ;
  assign y629 = ~1'b0 ;
  assign y630 = ~n1515 ;
  assign y631 = ~n1166 ;
  assign y632 = ~1'b0 ;
  assign y633 = ~n1517 ;
  assign y634 = ~n1518 ;
  assign y635 = ~n1523 ;
  assign y636 = n1524 ;
  assign y637 = ~n1531 ;
  assign y638 = ~n1534 ;
  assign y639 = n1536 ;
  assign y640 = ~n1540 ;
  assign y641 = ~n1543 ;
  assign y642 = ~n1550 ;
  assign y643 = ~1'b0 ;
  assign y644 = ~1'b0 ;
  assign y645 = ~n1552 ;
  assign y646 = ~1'b0 ;
  assign y647 = 1'b0 ;
  assign y648 = ~1'b0 ;
  assign y649 = ~n1556 ;
  assign y650 = ~n1560 ;
  assign y651 = n1563 ;
  assign y652 = ~n1566 ;
  assign y653 = ~1'b0 ;
  assign y654 = n1569 ;
  assign y655 = n1572 ;
  assign y656 = ~1'b0 ;
  assign y657 = ~1'b0 ;
  assign y658 = ~n1583 ;
  assign y659 = n1590 ;
  assign y660 = ~1'b0 ;
  assign y661 = ~n1594 ;
  assign y662 = n1597 ;
  assign y663 = ~n442 ;
  assign y664 = n1599 ;
  assign y665 = ~n1588 ;
  assign y666 = n1600 ;
  assign y667 = ~n1602 ;
  assign y668 = ~1'b0 ;
  assign y669 = n1603 ;
  assign y670 = ~1'b0 ;
  assign y671 = n1608 ;
  assign y672 = ~n1612 ;
  assign y673 = ~1'b0 ;
  assign y674 = ~n1616 ;
  assign y675 = ~n1623 ;
  assign y676 = n1625 ;
  assign y677 = x24 ;
  assign y678 = ~n1629 ;
  assign y679 = ~n1632 ;
  assign y680 = ~n1633 ;
  assign y681 = 1'b0 ;
  assign y682 = ~1'b0 ;
  assign y683 = n1642 ;
  assign y684 = ~n1645 ;
  assign y685 = ~1'b0 ;
  assign y686 = ~1'b0 ;
  assign y687 = n1647 ;
  assign y688 = ~1'b0 ;
  assign y689 = ~1'b0 ;
  assign y690 = ~n1652 ;
  assign y691 = n1654 ;
  assign y692 = ~n1657 ;
  assign y693 = ~1'b0 ;
  assign y694 = ~n855 ;
  assign y695 = n1664 ;
  assign y696 = ~1'b0 ;
  assign y697 = ~n1666 ;
  assign y698 = ~n1235 ;
  assign y699 = ~1'b0 ;
  assign y700 = ~1'b0 ;
  assign y701 = ~n1668 ;
  assign y702 = ~1'b0 ;
  assign y703 = ~1'b0 ;
  assign y704 = ~1'b0 ;
  assign y705 = n1674 ;
  assign y706 = n1676 ;
  assign y707 = ~n1681 ;
  assign y708 = ~n1686 ;
  assign y709 = ~n1689 ;
  assign y710 = ~n1693 ;
  assign y711 = ~n1695 ;
  assign y712 = ~n1700 ;
  assign y713 = n902 ;
  assign y714 = ~n1711 ;
  assign y715 = n1716 ;
  assign y716 = n1719 ;
  assign y717 = n1720 ;
  assign y718 = ~n1722 ;
  assign y719 = n1723 ;
  assign y720 = ~n1725 ;
  assign y721 = ~1'b0 ;
  assign y722 = n1728 ;
  assign y723 = ~n1740 ;
  assign y724 = ~1'b0 ;
  assign y725 = ~1'b0 ;
  assign y726 = ~1'b0 ;
  assign y727 = n1741 ;
  assign y728 = ~1'b0 ;
  assign y729 = n1743 ;
  assign y730 = ~n1747 ;
  assign y731 = n1748 ;
  assign y732 = n1755 ;
  assign y733 = ~n1756 ;
  assign y734 = ~n1759 ;
  assign y735 = n1765 ;
  assign y736 = ~1'b0 ;
  assign y737 = ~1'b0 ;
  assign y738 = ~n1767 ;
  assign y739 = ~1'b0 ;
  assign y740 = n1772 ;
  assign y741 = ~n1780 ;
  assign y742 = ~n1784 ;
  assign y743 = n1790 ;
  assign y744 = ~n1794 ;
  assign y745 = ~n1799 ;
  assign y746 = ~1'b0 ;
  assign y747 = n1803 ;
  assign y748 = ~1'b0 ;
  assign y749 = ~n1804 ;
  assign y750 = ~n1805 ;
  assign y751 = ~n1807 ;
  assign y752 = ~n1810 ;
  assign y753 = ~n1812 ;
  assign y754 = n1813 ;
  assign y755 = ~1'b0 ;
  assign y756 = ~1'b0 ;
  assign y757 = ~1'b0 ;
  assign y758 = 1'b0 ;
  assign y759 = n1817 ;
  assign y760 = ~n1819 ;
  assign y761 = n1824 ;
  assign y762 = ~1'b0 ;
  assign y763 = ~1'b0 ;
  assign y764 = ~1'b0 ;
  assign y765 = ~1'b0 ;
  assign y766 = ~1'b0 ;
  assign y767 = ~n1828 ;
  assign y768 = ~n174 ;
  assign y769 = ~n1832 ;
  assign y770 = n1835 ;
  assign y771 = n1844 ;
  assign y772 = ~1'b0 ;
  assign y773 = ~1'b0 ;
  assign y774 = n1849 ;
  assign y775 = n1851 ;
  assign y776 = n1858 ;
  assign y777 = ~n1860 ;
  assign y778 = ~n1861 ;
  assign y779 = ~n1862 ;
  assign y780 = ~n1863 ;
  assign y781 = ~1'b0 ;
  assign y782 = ~n1865 ;
  assign y783 = x46 ;
  assign y784 = ~n1874 ;
  assign y785 = ~n1876 ;
  assign y786 = ~n1877 ;
  assign y787 = ~n1880 ;
  assign y788 = ~1'b0 ;
  assign y789 = n1882 ;
  assign y790 = n1886 ;
  assign y791 = ~1'b0 ;
  assign y792 = n1891 ;
  assign y793 = ~n1895 ;
  assign y794 = ~n1906 ;
  assign y795 = n1124 ;
  assign y796 = ~n1909 ;
  assign y797 = ~1'b0 ;
  assign y798 = n1911 ;
  assign y799 = ~1'b0 ;
  assign y800 = n1912 ;
  assign y801 = ~1'b0 ;
  assign y802 = ~n1913 ;
  assign y803 = ~n1916 ;
  assign y804 = n1917 ;
  assign y805 = n1920 ;
  assign y806 = n1922 ;
  assign y807 = n679 ;
  assign y808 = n1927 ;
  assign y809 = ~1'b0 ;
  assign y810 = ~n1935 ;
  assign y811 = ~n1936 ;
  assign y812 = ~1'b0 ;
  assign y813 = ~1'b0 ;
  assign y814 = n1937 ;
  assign y815 = ~1'b0 ;
  assign y816 = ~n1943 ;
  assign y817 = ~n1950 ;
  assign y818 = ~n1953 ;
  assign y819 = ~1'b0 ;
  assign y820 = ~1'b0 ;
  assign y821 = ~1'b0 ;
  assign y822 = ~n1955 ;
  assign y823 = ~n1965 ;
  assign y824 = n1966 ;
  assign y825 = n1967 ;
  assign y826 = ~1'b0 ;
  assign y827 = n1970 ;
  assign y828 = n1971 ;
  assign y829 = x17 ;
  assign y830 = n1972 ;
  assign y831 = ~n1978 ;
  assign y832 = ~n1982 ;
  assign y833 = ~1'b0 ;
  assign y834 = n1988 ;
  assign y835 = ~n1991 ;
  assign y836 = n1995 ;
  assign y837 = ~n1996 ;
  assign y838 = n1507 ;
  assign y839 = ~1'b0 ;
  assign y840 = ~n1999 ;
  assign y841 = ~1'b0 ;
  assign y842 = n2003 ;
  assign y843 = ~n2005 ;
  assign y844 = ~1'b0 ;
  assign y845 = n2009 ;
  assign y846 = ~n2012 ;
  assign y847 = ~n2016 ;
  assign y848 = ~n2021 ;
  assign y849 = n2022 ;
  assign y850 = n2027 ;
  assign y851 = ~1'b0 ;
  assign y852 = ~1'b0 ;
  assign y853 = ~n2029 ;
  assign y854 = ~n2030 ;
  assign y855 = ~1'b0 ;
  assign y856 = ~n2033 ;
  assign y857 = ~n2036 ;
  assign y858 = ~n2039 ;
  assign y859 = ~1'b0 ;
  assign y860 = ~n2044 ;
  assign y861 = n2046 ;
  assign y862 = n2051 ;
  assign y863 = ~n2054 ;
  assign y864 = n2060 ;
  assign y865 = ~1'b0 ;
  assign y866 = ~n2062 ;
  assign y867 = ~n2066 ;
  assign y868 = n2067 ;
  assign y869 = ~n2068 ;
  assign y870 = ~n2070 ;
  assign y871 = ~1'b0 ;
  assign y872 = ~1'b0 ;
  assign y873 = n459 ;
  assign y874 = ~n2073 ;
  assign y875 = ~n2085 ;
  assign y876 = n2086 ;
  assign y877 = ~n2088 ;
  assign y878 = ~n2093 ;
  assign y879 = n2095 ;
  assign y880 = ~1'b0 ;
  assign y881 = ~n2096 ;
  assign y882 = n2098 ;
  assign y883 = ~n2105 ;
  assign y884 = n2107 ;
  assign y885 = ~1'b0 ;
  assign y886 = n1529 ;
  assign y887 = ~n2108 ;
  assign y888 = ~1'b0 ;
  assign y889 = n2111 ;
  assign y890 = ~1'b0 ;
  assign y891 = n2116 ;
  assign y892 = n2119 ;
  assign y893 = ~1'b0 ;
  assign y894 = 1'b0 ;
  assign y895 = ~n2120 ;
  assign y896 = n2128 ;
  assign y897 = ~n1761 ;
  assign y898 = ~n2134 ;
  assign y899 = ~1'b0 ;
  assign y900 = ~n2135 ;
  assign y901 = ~n2144 ;
  assign y902 = n2146 ;
  assign y903 = n2150 ;
  assign y904 = n2153 ;
  assign y905 = ~n358 ;
  assign y906 = ~n506 ;
  assign y907 = ~n2160 ;
  assign y908 = ~1'b0 ;
  assign y909 = ~n2167 ;
  assign y910 = n2179 ;
  assign y911 = 1'b0 ;
  assign y912 = n2180 ;
  assign y913 = ~1'b0 ;
  assign y914 = n2182 ;
  assign y915 = ~n2183 ;
  assign y916 = ~1'b0 ;
  assign y917 = ~1'b0 ;
  assign y918 = ~n2185 ;
  assign y919 = ~1'b0 ;
  assign y920 = ~n2189 ;
  assign y921 = ~1'b0 ;
  assign y922 = n2192 ;
  assign y923 = ~1'b0 ;
  assign y924 = ~1'b0 ;
  assign y925 = n2195 ;
  assign y926 = n2197 ;
  assign y927 = ~n2201 ;
  assign y928 = ~n2206 ;
  assign y929 = ~n2213 ;
  assign y930 = n368 ;
  assign y931 = ~1'b0 ;
  assign y932 = ~n2215 ;
  assign y933 = ~1'b0 ;
  assign y934 = ~n2218 ;
  assign y935 = ~n2221 ;
  assign y936 = ~n2231 ;
  assign y937 = n2232 ;
  assign y938 = n2234 ;
  assign y939 = ~1'b0 ;
  assign y940 = n2237 ;
  assign y941 = ~1'b0 ;
  assign y942 = ~n2240 ;
  assign y943 = n2249 ;
  assign y944 = n2255 ;
  assign y945 = ~n2257 ;
  assign y946 = n2259 ;
  assign y947 = ~1'b0 ;
  assign y948 = ~n2266 ;
  assign y949 = ~1'b0 ;
  assign y950 = ~n2267 ;
  assign y951 = ~n2274 ;
  assign y952 = ~n2275 ;
  assign y953 = ~1'b0 ;
  assign y954 = ~n2285 ;
  assign y955 = ~1'b0 ;
  assign y956 = n2287 ;
  assign y957 = n2288 ;
  assign y958 = ~n2289 ;
  assign y959 = ~n2293 ;
  assign y960 = ~n2300 ;
  assign y961 = ~1'b0 ;
  assign y962 = n2302 ;
  assign y963 = ~n2303 ;
  assign y964 = ~n2306 ;
  assign y965 = ~1'b0 ;
  assign y966 = ~n2308 ;
  assign y967 = ~n2310 ;
  assign y968 = ~1'b0 ;
  assign y969 = ~n2315 ;
  assign y970 = ~1'b0 ;
  assign y971 = ~n2318 ;
  assign y972 = ~n2323 ;
  assign y973 = ~1'b0 ;
  assign y974 = ~n2327 ;
  assign y975 = n2331 ;
  assign y976 = ~1'b0 ;
  assign y977 = ~n2332 ;
  assign y978 = n2334 ;
  assign y979 = ~1'b0 ;
  assign y980 = ~n2337 ;
  assign y981 = ~1'b0 ;
  assign y982 = ~1'b0 ;
  assign y983 = n2338 ;
  assign y984 = ~1'b0 ;
  assign y985 = ~n2339 ;
  assign y986 = ~n2344 ;
  assign y987 = ~1'b0 ;
  assign y988 = n2348 ;
  assign y989 = ~n2353 ;
  assign y990 = ~n1089 ;
  assign y991 = n2356 ;
  assign y992 = ~1'b0 ;
  assign y993 = ~n2357 ;
  assign y994 = ~1'b0 ;
  assign y995 = n2359 ;
  assign y996 = n2362 ;
  assign y997 = n2363 ;
  assign y998 = n1805 ;
  assign y999 = ~1'b0 ;
  assign y1000 = n2364 ;
  assign y1001 = ~n2371 ;
  assign y1002 = 1'b0 ;
  assign y1003 = ~n2372 ;
  assign y1004 = n2373 ;
  assign y1005 = ~n2374 ;
  assign y1006 = n2380 ;
  assign y1007 = ~1'b0 ;
  assign y1008 = n2381 ;
  assign y1009 = 1'b0 ;
  assign y1010 = ~1'b0 ;
  assign y1011 = 1'b0 ;
  assign y1012 = n2382 ;
  assign y1013 = n1147 ;
  assign y1014 = ~1'b0 ;
  assign y1015 = ~1'b0 ;
  assign y1016 = ~n2387 ;
  assign y1017 = ~1'b0 ;
  assign y1018 = n2388 ;
  assign y1019 = ~n2389 ;
  assign y1020 = n2391 ;
  assign y1021 = ~n2392 ;
  assign y1022 = ~n2395 ;
  assign y1023 = ~n2397 ;
  assign y1024 = ~1'b0 ;
  assign y1025 = ~n2398 ;
  assign y1026 = ~n2399 ;
  assign y1027 = ~n2412 ;
  assign y1028 = n2413 ;
  assign y1029 = 1'b0 ;
  assign y1030 = ~n2414 ;
  assign y1031 = ~n2424 ;
  assign y1032 = n2425 ;
  assign y1033 = ~n2427 ;
  assign y1034 = ~n2428 ;
  assign y1035 = ~n2429 ;
  assign y1036 = ~1'b0 ;
  assign y1037 = n556 ;
  assign y1038 = ~1'b0 ;
  assign y1039 = ~n2431 ;
  assign y1040 = n2436 ;
  assign y1041 = n2438 ;
  assign y1042 = ~1'b0 ;
  assign y1043 = n2441 ;
  assign y1044 = ~n2448 ;
  assign y1045 = n2449 ;
  assign y1046 = ~n2450 ;
  assign y1047 = n2451 ;
  assign y1048 = n2452 ;
  assign y1049 = ~n2456 ;
  assign y1050 = n2462 ;
  assign y1051 = n2464 ;
  assign y1052 = n2468 ;
  assign y1053 = ~n2476 ;
  assign y1054 = n2477 ;
  assign y1055 = ~n2479 ;
  assign y1056 = n2481 ;
  assign y1057 = ~n2482 ;
  assign y1058 = n2483 ;
  assign y1059 = ~n2487 ;
  assign y1060 = n2494 ;
  assign y1061 = ~n2412 ;
  assign y1062 = n2496 ;
  assign y1063 = n2504 ;
  assign y1064 = ~1'b0 ;
  assign y1065 = n2510 ;
  assign y1066 = n2512 ;
  assign y1067 = n2515 ;
  assign y1068 = n2516 ;
  assign y1069 = n2517 ;
  assign y1070 = ~n2520 ;
  assign y1071 = n2521 ;
  assign y1072 = ~n2525 ;
  assign y1073 = n2530 ;
  assign y1074 = n2537 ;
  assign y1075 = n2540 ;
  assign y1076 = n2553 ;
  assign y1077 = n2554 ;
  assign y1078 = ~n2557 ;
  assign y1079 = n533 ;
  assign y1080 = ~n2559 ;
  assign y1081 = n2560 ;
  assign y1082 = ~1'b0 ;
  assign y1083 = n2561 ;
  assign y1084 = ~n2563 ;
  assign y1085 = ~n2564 ;
  assign y1086 = ~n2569 ;
  assign y1087 = ~n2571 ;
  assign y1088 = ~n2577 ;
  assign y1089 = n2581 ;
  assign y1090 = ~1'b0 ;
  assign y1091 = n2582 ;
  assign y1092 = ~1'b0 ;
  assign y1093 = ~x81 ;
  assign y1094 = ~n2587 ;
  assign y1095 = ~n2593 ;
  assign y1096 = ~1'b0 ;
  assign y1097 = ~n708 ;
  assign y1098 = ~n2596 ;
  assign y1099 = ~1'b0 ;
  assign y1100 = n588 ;
  assign y1101 = n2597 ;
  assign y1102 = ~1'b0 ;
  assign y1103 = n2601 ;
  assign y1104 = ~n2602 ;
  assign y1105 = ~n1562 ;
  assign y1106 = n2603 ;
  assign y1107 = ~n2604 ;
  assign y1108 = ~n2607 ;
  assign y1109 = ~x6 ;
  assign y1110 = ~1'b0 ;
  assign y1111 = 1'b0 ;
  assign y1112 = n2610 ;
  assign y1113 = ~n2612 ;
  assign y1114 = ~n2621 ;
  assign y1115 = ~n2622 ;
  assign y1116 = ~1'b0 ;
  assign y1117 = n2624 ;
  assign y1118 = n2626 ;
  assign y1119 = ~1'b0 ;
  assign y1120 = ~n2627 ;
  assign y1121 = ~n2633 ;
  assign y1122 = ~1'b0 ;
  assign y1123 = n2221 ;
  assign y1124 = ~1'b0 ;
  assign y1125 = ~n2634 ;
  assign y1126 = n2636 ;
  assign y1127 = n2412 ;
  assign y1128 = ~1'b0 ;
  assign y1129 = ~1'b0 ;
  assign y1130 = ~n2638 ;
  assign y1131 = ~n2640 ;
  assign y1132 = ~n2647 ;
  assign y1133 = ~n2652 ;
  assign y1134 = ~1'b0 ;
  assign y1135 = n2654 ;
  assign y1136 = ~1'b0 ;
  assign y1137 = ~n2655 ;
  assign y1138 = ~1'b0 ;
  assign y1139 = ~n2665 ;
  assign y1140 = ~n2671 ;
  assign y1141 = n2676 ;
  assign y1142 = ~1'b0 ;
  assign y1143 = ~n2678 ;
  assign y1144 = n2680 ;
  assign y1145 = n2681 ;
  assign y1146 = n2686 ;
  assign y1147 = ~n2687 ;
  assign y1148 = ~1'b0 ;
  assign y1149 = ~n2689 ;
  assign y1150 = n677 ;
  assign y1151 = n2691 ;
  assign y1152 = n2692 ;
  assign y1153 = n2696 ;
  assign y1154 = n2712 ;
  assign y1155 = ~1'b0 ;
  assign y1156 = n2715 ;
  assign y1157 = ~1'b0 ;
  assign y1158 = ~1'b0 ;
  assign y1159 = n2717 ;
  assign y1160 = n2327 ;
  assign y1161 = n2722 ;
  assign y1162 = n2724 ;
  assign y1163 = ~1'b0 ;
  assign y1164 = n2726 ;
  assign y1165 = ~n2728 ;
  assign y1166 = n2730 ;
  assign y1167 = ~1'b0 ;
  assign y1168 = n2735 ;
  assign y1169 = ~n2737 ;
  assign y1170 = ~1'b0 ;
  assign y1171 = n2738 ;
  assign y1172 = n2742 ;
  assign y1173 = ~n2743 ;
  assign y1174 = 1'b0 ;
  assign y1175 = n2745 ;
  assign y1176 = n2750 ;
  assign y1177 = ~n2752 ;
  assign y1178 = ~1'b0 ;
  assign y1179 = ~n2763 ;
  assign y1180 = ~n2769 ;
  assign y1181 = n2776 ;
  assign y1182 = ~n2777 ;
  assign y1183 = n2780 ;
  assign y1184 = ~n2785 ;
  assign y1185 = ~n1572 ;
  assign y1186 = n2790 ;
  assign y1187 = ~1'b0 ;
  assign y1188 = ~1'b0 ;
  assign y1189 = ~n2792 ;
  assign y1190 = n2794 ;
  assign y1191 = ~n2797 ;
  assign y1192 = ~1'b0 ;
  assign y1193 = ~n2800 ;
  assign y1194 = ~n2804 ;
  assign y1195 = n2805 ;
  assign y1196 = n2806 ;
  assign y1197 = n2807 ;
  assign y1198 = ~n2812 ;
  assign y1199 = ~1'b0 ;
  assign y1200 = ~n2813 ;
  assign y1201 = ~n2814 ;
  assign y1202 = n2822 ;
  assign y1203 = ~n1588 ;
  assign y1204 = ~n2823 ;
  assign y1205 = n2824 ;
  assign y1206 = ~1'b0 ;
  assign y1207 = n2834 ;
  assign y1208 = ~n2838 ;
  assign y1209 = ~n2840 ;
  assign y1210 = n2846 ;
  assign y1211 = n2847 ;
  assign y1212 = n2849 ;
  assign y1213 = ~1'b0 ;
  assign y1214 = n2854 ;
  assign y1215 = n2855 ;
  assign y1216 = ~1'b0 ;
  assign y1217 = ~n2859 ;
  assign y1218 = ~1'b0 ;
  assign y1219 = n2862 ;
  assign y1220 = ~n2863 ;
  assign y1221 = ~1'b0 ;
  assign y1222 = ~n709 ;
  assign y1223 = ~n2866 ;
  assign y1224 = ~n2868 ;
  assign y1225 = ~1'b0 ;
  assign y1226 = ~1'b0 ;
  assign y1227 = n2869 ;
  assign y1228 = ~1'b0 ;
  assign y1229 = 1'b0 ;
  assign y1230 = ~n2872 ;
  assign y1231 = n2874 ;
  assign y1232 = ~1'b0 ;
  assign y1233 = n2875 ;
  assign y1234 = ~n2876 ;
  assign y1235 = ~1'b0 ;
  assign y1236 = ~n2878 ;
  assign y1237 = n2882 ;
  assign y1238 = ~1'b0 ;
  assign y1239 = n2883 ;
  assign y1240 = n2885 ;
  assign y1241 = ~1'b0 ;
  assign y1242 = ~n2886 ;
  assign y1243 = n2890 ;
  assign y1244 = n2898 ;
  assign y1245 = n2906 ;
  assign y1246 = ~1'b0 ;
  assign y1247 = ~1'b0 ;
  assign y1248 = ~n2912 ;
  assign y1249 = ~n2914 ;
  assign y1250 = n2915 ;
  assign y1251 = ~1'b0 ;
  assign y1252 = n2916 ;
  assign y1253 = n2920 ;
  assign y1254 = ~n2925 ;
  assign y1255 = ~n2928 ;
  assign y1256 = n2932 ;
  assign y1257 = n1629 ;
  assign y1258 = ~n2462 ;
  assign y1259 = ~n2936 ;
  assign y1260 = ~n2942 ;
  assign y1261 = ~1'b0 ;
  assign y1262 = ~n2945 ;
  assign y1263 = ~1'b0 ;
  assign y1264 = ~1'b0 ;
  assign y1265 = n2946 ;
  assign y1266 = ~n2947 ;
  assign y1267 = ~1'b0 ;
  assign y1268 = ~n1534 ;
  assign y1269 = ~n2948 ;
  assign y1270 = n2952 ;
  assign y1271 = ~1'b0 ;
  assign y1272 = n2955 ;
  assign y1273 = ~1'b0 ;
  assign y1274 = ~1'b0 ;
  assign y1275 = n2956 ;
  assign y1276 = n2957 ;
  assign y1277 = ~n2958 ;
  assign y1278 = n2959 ;
  assign y1279 = ~n2960 ;
  assign y1280 = n2970 ;
  assign y1281 = n2973 ;
  assign y1282 = ~1'b0 ;
  assign y1283 = ~n2974 ;
  assign y1284 = ~n2976 ;
  assign y1285 = n2979 ;
  assign y1286 = n2984 ;
  assign y1287 = n2985 ;
  assign y1288 = ~1'b0 ;
  assign y1289 = n2990 ;
  assign y1290 = 1'b0 ;
  assign y1291 = ~1'b0 ;
  assign y1292 = n2994 ;
  assign y1293 = ~1'b0 ;
  assign y1294 = ~1'b0 ;
  assign y1295 = 1'b0 ;
  assign y1296 = ~1'b0 ;
  assign y1297 = n3001 ;
  assign y1298 = n3003 ;
  assign y1299 = n3004 ;
  assign y1300 = n3008 ;
  assign y1301 = ~1'b0 ;
  assign y1302 = ~1'b0 ;
  assign y1303 = ~n3009 ;
  assign y1304 = n3013 ;
  assign y1305 = ~n3017 ;
  assign y1306 = ~n3020 ;
  assign y1307 = n3021 ;
  assign y1308 = n3022 ;
  assign y1309 = ~1'b0 ;
  assign y1310 = ~n3023 ;
  assign y1311 = ~1'b0 ;
  assign y1312 = ~n3029 ;
  assign y1313 = ~n143 ;
  assign y1314 = ~n3033 ;
  assign y1315 = ~1'b0 ;
  assign y1316 = ~n3041 ;
  assign y1317 = ~n3045 ;
  assign y1318 = ~n3046 ;
  assign y1319 = ~1'b0 ;
  assign y1320 = ~1'b0 ;
  assign y1321 = ~n3047 ;
  assign y1322 = ~n3051 ;
  assign y1323 = n3055 ;
  assign y1324 = n3058 ;
  assign y1325 = ~1'b0 ;
  assign y1326 = ~n3061 ;
  assign y1327 = 1'b0 ;
  assign y1328 = ~1'b0 ;
  assign y1329 = n3062 ;
  assign y1330 = ~1'b0 ;
  assign y1331 = ~n3065 ;
  assign y1332 = 1'b0 ;
  assign y1333 = n3066 ;
  assign y1334 = ~1'b0 ;
  assign y1335 = ~1'b0 ;
  assign y1336 = ~n3067 ;
  assign y1337 = ~1'b0 ;
  assign y1338 = ~1'b0 ;
  assign y1339 = n3068 ;
  assign y1340 = 1'b0 ;
  assign y1341 = ~1'b0 ;
  assign y1342 = 1'b0 ;
  assign y1343 = n3069 ;
  assign y1344 = ~1'b0 ;
  assign y1345 = ~n3071 ;
  assign y1346 = n3073 ;
  assign y1347 = n3075 ;
  assign y1348 = n3076 ;
  assign y1349 = n3080 ;
  assign y1350 = n3081 ;
  assign y1351 = ~1'b0 ;
  assign y1352 = ~n3084 ;
  assign y1353 = ~n3086 ;
  assign y1354 = 1'b0 ;
  assign y1355 = ~1'b0 ;
  assign y1356 = ~1'b0 ;
  assign y1357 = ~1'b0 ;
  assign y1358 = ~n3089 ;
  assign y1359 = n3091 ;
  assign y1360 = n3092 ;
  assign y1361 = ~n3095 ;
  assign y1362 = n3099 ;
  assign y1363 = ~1'b0 ;
  assign y1364 = ~n3100 ;
  assign y1365 = ~n3102 ;
  assign y1366 = 1'b0 ;
  assign y1367 = ~n2639 ;
  assign y1368 = ~n3105 ;
  assign y1369 = ~n3106 ;
  assign y1370 = ~n3109 ;
  assign y1371 = n3115 ;
  assign y1372 = ~n3116 ;
  assign y1373 = ~n3121 ;
  assign y1374 = n3122 ;
  assign y1375 = n3124 ;
  assign y1376 = n3133 ;
  assign y1377 = ~1'b0 ;
  assign y1378 = n3135 ;
  assign y1379 = 1'b0 ;
  assign y1380 = ~n3139 ;
  assign y1381 = n3140 ;
  assign y1382 = ~n3143 ;
  assign y1383 = n3153 ;
  assign y1384 = ~n3154 ;
  assign y1385 = ~1'b0 ;
  assign y1386 = ~1'b0 ;
  assign y1387 = ~n3156 ;
  assign y1388 = ~1'b0 ;
  assign y1389 = ~1'b0 ;
  assign y1390 = ~n3162 ;
  assign y1391 = n3164 ;
  assign y1392 = ~n928 ;
  assign y1393 = ~n3165 ;
  assign y1394 = n3169 ;
  assign y1395 = ~1'b0 ;
  assign y1396 = ~n3175 ;
  assign y1397 = ~1'b0 ;
  assign y1398 = ~n3177 ;
  assign y1399 = ~1'b0 ;
  assign y1400 = ~1'b0 ;
  assign y1401 = ~n3183 ;
  assign y1402 = ~n3185 ;
  assign y1403 = ~n3186 ;
  assign y1404 = ~1'b0 ;
  assign y1405 = ~n3188 ;
  assign y1406 = n3193 ;
  assign y1407 = ~1'b0 ;
  assign y1408 = ~1'b0 ;
  assign y1409 = n3195 ;
  assign y1410 = ~1'b0 ;
  assign y1411 = ~n3200 ;
  assign y1412 = ~n3203 ;
  assign y1413 = n3205 ;
  assign y1414 = n3207 ;
  assign y1415 = ~n3214 ;
  assign y1416 = ~n3215 ;
  assign y1417 = n3224 ;
  assign y1418 = n3227 ;
  assign y1419 = ~1'b0 ;
  assign y1420 = ~n3230 ;
  assign y1421 = ~1'b0 ;
  assign y1422 = n3231 ;
  assign y1423 = ~n3234 ;
  assign y1424 = ~n3236 ;
  assign y1425 = ~1'b0 ;
  assign y1426 = n496 ;
  assign y1427 = n3240 ;
  assign y1428 = ~n3243 ;
  assign y1429 = n3249 ;
  assign y1430 = n3262 ;
  assign y1431 = ~n3264 ;
  assign y1432 = ~n3273 ;
  assign y1433 = n3274 ;
  assign y1434 = ~1'b0 ;
  assign y1435 = n3279 ;
  assign y1436 = n3282 ;
  assign y1437 = ~n3286 ;
  assign y1438 = ~1'b0 ;
  assign y1439 = ~1'b0 ;
  assign y1440 = n3288 ;
  assign y1441 = ~1'b0 ;
  assign y1442 = n3292 ;
  assign y1443 = ~n3295 ;
  assign y1444 = ~n3298 ;
  assign y1445 = ~n3300 ;
  assign y1446 = ~n3302 ;
  assign y1447 = n3303 ;
  assign y1448 = n3310 ;
  assign y1449 = n3311 ;
  assign y1450 = ~n163 ;
  assign y1451 = ~n3314 ;
  assign y1452 = n3318 ;
  assign y1453 = ~1'b0 ;
  assign y1454 = ~1'b0 ;
  assign y1455 = n3319 ;
  assign y1456 = n3324 ;
  assign y1457 = n3326 ;
  assign y1458 = n3328 ;
  assign y1459 = n3331 ;
  assign y1460 = n3334 ;
  assign y1461 = ~1'b0 ;
  assign y1462 = ~n3335 ;
  assign y1463 = n3339 ;
  assign y1464 = ~1'b0 ;
  assign y1465 = n3340 ;
  assign y1466 = ~1'b0 ;
  assign y1467 = n3342 ;
  assign y1468 = n1578 ;
  assign y1469 = ~n3350 ;
  assign y1470 = ~1'b0 ;
  assign y1471 = ~1'b0 ;
  assign y1472 = ~1'b0 ;
  assign y1473 = ~n1714 ;
  assign y1474 = ~n3357 ;
  assign y1475 = ~1'b0 ;
  assign y1476 = ~1'b0 ;
  assign y1477 = n3359 ;
  assign y1478 = ~n3361 ;
  assign y1479 = 1'b0 ;
  assign y1480 = ~n3362 ;
  assign y1481 = ~1'b0 ;
  assign y1482 = ~n3366 ;
  assign y1483 = n3368 ;
  assign y1484 = n3369 ;
  assign y1485 = ~n3370 ;
  assign y1486 = ~1'b0 ;
  assign y1487 = n3372 ;
  assign y1488 = ~n3374 ;
  assign y1489 = n3376 ;
  assign y1490 = ~n3378 ;
  assign y1491 = ~1'b0 ;
  assign y1492 = ~n3381 ;
  assign y1493 = ~n3388 ;
  assign y1494 = n3389 ;
  assign y1495 = ~1'b0 ;
  assign y1496 = ~1'b0 ;
  assign y1497 = ~n3391 ;
  assign y1498 = ~1'b0 ;
  assign y1499 = ~1'b0 ;
  assign y1500 = n1338 ;
  assign y1501 = n3395 ;
  assign y1502 = n3401 ;
  assign y1503 = n3402 ;
  assign y1504 = ~n1722 ;
  assign y1505 = n3414 ;
  assign y1506 = n3417 ;
  assign y1507 = ~1'b0 ;
  assign y1508 = ~n3419 ;
  assign y1509 = n3420 ;
  assign y1510 = ~1'b0 ;
  assign y1511 = ~1'b0 ;
  assign y1512 = ~n3422 ;
  assign y1513 = n3424 ;
  assign y1514 = ~n3426 ;
  assign y1515 = n3429 ;
  assign y1516 = ~1'b0 ;
  assign y1517 = ~n3430 ;
  assign y1518 = n3434 ;
  assign y1519 = ~n3437 ;
  assign y1520 = n3438 ;
  assign y1521 = ~1'b0 ;
  assign y1522 = ~n3439 ;
  assign y1523 = ~n3444 ;
  assign y1524 = ~n3448 ;
  assign y1525 = ~1'b0 ;
  assign y1526 = n157 ;
  assign y1527 = n3449 ;
  assign y1528 = n3450 ;
  assign y1529 = ~n3453 ;
  assign y1530 = ~n3458 ;
  assign y1531 = n3463 ;
  assign y1532 = ~n3465 ;
  assign y1533 = ~1'b0 ;
  assign y1534 = ~n3468 ;
  assign y1535 = ~1'b0 ;
  assign y1536 = ~1'b0 ;
  assign y1537 = ~n3469 ;
  assign y1538 = ~1'b0 ;
  assign y1539 = n3474 ;
  assign y1540 = n3476 ;
  assign y1541 = n3477 ;
  assign y1542 = ~n3479 ;
  assign y1543 = ~1'b0 ;
  assign y1544 = ~1'b0 ;
  assign y1545 = ~1'b0 ;
  assign y1546 = ~1'b0 ;
  assign y1547 = n3485 ;
  assign y1548 = ~n257 ;
  assign y1549 = n3486 ;
  assign y1550 = ~1'b0 ;
  assign y1551 = n3487 ;
  assign y1552 = ~1'b0 ;
  assign y1553 = ~n3488 ;
  assign y1554 = n3491 ;
  assign y1555 = n3493 ;
  assign y1556 = n3494 ;
  assign y1557 = ~n3495 ;
  assign y1558 = ~1'b0 ;
  assign y1559 = ~n3497 ;
  assign y1560 = ~n3499 ;
  assign y1561 = ~1'b0 ;
  assign y1562 = n3501 ;
  assign y1563 = n2151 ;
  assign y1564 = ~n3502 ;
  assign y1565 = ~n3504 ;
  assign y1566 = ~n3505 ;
  assign y1567 = ~n3507 ;
  assign y1568 = ~1'b0 ;
  assign y1569 = ~n3508 ;
  assign y1570 = ~n3193 ;
  assign y1571 = ~1'b0 ;
  assign y1572 = 1'b0 ;
  assign y1573 = ~1'b0 ;
  assign y1574 = ~n3518 ;
  assign y1575 = ~n3526 ;
  assign y1576 = n1642 ;
  assign y1577 = ~n3528 ;
  assign y1578 = ~1'b0 ;
  assign y1579 = n3529 ;
  assign y1580 = ~n3530 ;
  assign y1581 = n3532 ;
  assign y1582 = ~1'b0 ;
  assign y1583 = n3536 ;
  assign y1584 = n3537 ;
  assign y1585 = n3539 ;
  assign y1586 = n3540 ;
  assign y1587 = ~1'b0 ;
  assign y1588 = ~n3542 ;
  assign y1589 = ~n3543 ;
  assign y1590 = n3058 ;
  assign y1591 = n3546 ;
  assign y1592 = n3547 ;
  assign y1593 = n3548 ;
  assign y1594 = n2969 ;
  assign y1595 = ~n3551 ;
  assign y1596 = ~n3557 ;
  assign y1597 = ~n3559 ;
  assign y1598 = ~1'b0 ;
  assign y1599 = ~n3561 ;
  assign y1600 = ~n3564 ;
  assign y1601 = n3567 ;
  assign y1602 = n3569 ;
  assign y1603 = ~n3571 ;
  assign y1604 = ~n3573 ;
  assign y1605 = ~n3577 ;
  assign y1606 = ~n3580 ;
  assign y1607 = ~1'b0 ;
  assign y1608 = n3583 ;
  assign y1609 = n3589 ;
  assign y1610 = n3595 ;
  assign y1611 = ~1'b0 ;
  assign y1612 = ~n3599 ;
  assign y1613 = ~1'b0 ;
  assign y1614 = ~n3601 ;
  assign y1615 = ~n3602 ;
  assign y1616 = ~n3605 ;
  assign y1617 = n3608 ;
  assign y1618 = ~n1329 ;
  assign y1619 = ~1'b0 ;
  assign y1620 = ~1'b0 ;
  assign y1621 = n3611 ;
  assign y1622 = n3615 ;
  assign y1623 = ~1'b0 ;
  assign y1624 = ~n3620 ;
  assign y1625 = ~n3635 ;
  assign y1626 = ~n3639 ;
  assign y1627 = n3642 ;
  assign y1628 = ~1'b0 ;
  assign y1629 = ~1'b0 ;
  assign y1630 = n2026 ;
  assign y1631 = ~n2904 ;
  assign y1632 = n3644 ;
  assign y1633 = ~1'b0 ;
  assign y1634 = ~n3511 ;
  assign y1635 = ~n3646 ;
  assign y1636 = n3648 ;
  assign y1637 = n3659 ;
  assign y1638 = ~1'b0 ;
  assign y1639 = n3664 ;
  assign y1640 = ~1'b0 ;
  assign y1641 = ~n3671 ;
  assign y1642 = n3673 ;
  assign y1643 = n3676 ;
  assign y1644 = n3677 ;
  assign y1645 = n3678 ;
  assign y1646 = n3690 ;
  assign y1647 = ~1'b0 ;
  assign y1648 = ~1'b0 ;
  assign y1649 = n3693 ;
  assign y1650 = n3694 ;
  assign y1651 = n3697 ;
  assign y1652 = ~1'b0 ;
  assign y1653 = n3700 ;
  assign y1654 = n3701 ;
  assign y1655 = ~n3702 ;
  assign y1656 = ~n3713 ;
  assign y1657 = ~1'b0 ;
  assign y1658 = ~1'b0 ;
  assign y1659 = n1511 ;
  assign y1660 = ~n3720 ;
  assign y1661 = ~n3724 ;
  assign y1662 = n1804 ;
  assign y1663 = n3726 ;
  assign y1664 = ~1'b0 ;
  assign y1665 = n3727 ;
  assign y1666 = n3734 ;
  assign y1667 = ~1'b0 ;
  assign y1668 = n3736 ;
  assign y1669 = ~n3119 ;
  assign y1670 = ~n3737 ;
  assign y1671 = ~n3741 ;
  assign y1672 = ~n3746 ;
  assign y1673 = ~n3752 ;
  assign y1674 = ~n3760 ;
  assign y1675 = ~1'b0 ;
  assign y1676 = ~n3404 ;
  assign y1677 = ~1'b0 ;
  assign y1678 = ~1'b0 ;
  assign y1679 = ~n3761 ;
  assign y1680 = ~n3762 ;
  assign y1681 = ~1'b0 ;
  assign y1682 = ~n3766 ;
  assign y1683 = ~1'b0 ;
  assign y1684 = n1481 ;
  assign y1685 = n3770 ;
  assign y1686 = n3775 ;
  assign y1687 = n3776 ;
  assign y1688 = ~1'b0 ;
  assign y1689 = ~n3780 ;
  assign y1690 = n2413 ;
  assign y1691 = n3781 ;
  assign y1692 = ~n3786 ;
  assign y1693 = n3788 ;
  assign y1694 = ~n3789 ;
  assign y1695 = ~1'b0 ;
  assign y1696 = ~1'b0 ;
  assign y1697 = n3790 ;
  assign y1698 = n3799 ;
  assign y1699 = ~1'b0 ;
  assign y1700 = ~n3804 ;
  assign y1701 = n3809 ;
  assign y1702 = ~n3811 ;
  assign y1703 = ~1'b0 ;
  assign y1704 = ~1'b0 ;
  assign y1705 = ~1'b0 ;
  assign y1706 = n3818 ;
  assign y1707 = ~n3823 ;
  assign y1708 = n3825 ;
  assign y1709 = ~n3834 ;
  assign y1710 = ~1'b0 ;
  assign y1711 = n3837 ;
  assign y1712 = ~1'b0 ;
  assign y1713 = n3854 ;
  assign y1714 = ~1'b0 ;
  assign y1715 = n2802 ;
  assign y1716 = ~1'b0 ;
  assign y1717 = ~n3857 ;
  assign y1718 = ~n3859 ;
  assign y1719 = ~n3865 ;
  assign y1720 = ~1'b0 ;
  assign y1721 = ~n3870 ;
  assign y1722 = n3873 ;
  assign y1723 = ~1'b0 ;
  assign y1724 = ~n3877 ;
  assign y1725 = ~n3879 ;
  assign y1726 = ~1'b0 ;
  assign y1727 = ~1'b0 ;
  assign y1728 = n3880 ;
  assign y1729 = ~1'b0 ;
  assign y1730 = 1'b0 ;
  assign y1731 = ~1'b0 ;
  assign y1732 = ~n3901 ;
  assign y1733 = n3908 ;
  assign y1734 = ~1'b0 ;
  assign y1735 = ~n3912 ;
  assign y1736 = ~n3922 ;
  assign y1737 = ~n3925 ;
  assign y1738 = n3927 ;
  assign y1739 = n3930 ;
  assign y1740 = ~1'b0 ;
  assign y1741 = n3931 ;
  assign y1742 = ~1'b0 ;
  assign y1743 = n3933 ;
  assign y1744 = ~1'b0 ;
  assign y1745 = ~1'b0 ;
  assign y1746 = ~1'b0 ;
  assign y1747 = n3935 ;
  assign y1748 = n3936 ;
  assign y1749 = n1331 ;
  assign y1750 = n3937 ;
  assign y1751 = ~n3940 ;
  assign y1752 = n3943 ;
  assign y1753 = n3944 ;
  assign y1754 = n2151 ;
  assign y1755 = ~1'b0 ;
  assign y1756 = n3945 ;
  assign y1757 = ~1'b0 ;
  assign y1758 = n3947 ;
  assign y1759 = n3949 ;
  assign y1760 = ~n1939 ;
  assign y1761 = n3950 ;
  assign y1762 = n3951 ;
  assign y1763 = ~1'b0 ;
  assign y1764 = ~n3958 ;
  assign y1765 = ~1'b0 ;
  assign y1766 = ~n3961 ;
  assign y1767 = ~1'b0 ;
  assign y1768 = ~n3962 ;
  assign y1769 = n3964 ;
  assign y1770 = n3966 ;
  assign y1771 = ~1'b0 ;
  assign y1772 = n3970 ;
  assign y1773 = n3974 ;
  assign y1774 = ~1'b0 ;
  assign y1775 = ~1'b0 ;
  assign y1776 = n3975 ;
  assign y1777 = ~n3981 ;
  assign y1778 = ~n3987 ;
  assign y1779 = n3992 ;
  assign y1780 = ~n3993 ;
  assign y1781 = ~n3995 ;
  assign y1782 = ~n3997 ;
  assign y1783 = n4002 ;
  assign y1784 = ~n4009 ;
  assign y1785 = n4010 ;
  assign y1786 = n4013 ;
  assign y1787 = ~n4015 ;
  assign y1788 = ~n4019 ;
  assign y1789 = n4020 ;
  assign y1790 = ~n4024 ;
  assign y1791 = n4028 ;
  assign y1792 = ~n4030 ;
  assign y1793 = n4050 ;
  assign y1794 = ~1'b0 ;
  assign y1795 = ~n1761 ;
  assign y1796 = n4051 ;
  assign y1797 = ~n4052 ;
  assign y1798 = ~n4058 ;
  assign y1799 = n4061 ;
  assign y1800 = ~1'b0 ;
  assign y1801 = n4064 ;
  assign y1802 = n4069 ;
  assign y1803 = n4070 ;
  assign y1804 = n4073 ;
  assign y1805 = ~1'b0 ;
  assign y1806 = ~1'b0 ;
  assign y1807 = ~n4077 ;
  assign y1808 = ~n4083 ;
  assign y1809 = ~n4089 ;
  assign y1810 = ~1'b0 ;
  assign y1811 = n4090 ;
  assign y1812 = n4091 ;
  assign y1813 = n4093 ;
  assign y1814 = ~n4094 ;
  assign y1815 = n4099 ;
  assign y1816 = n2479 ;
  assign y1817 = n4101 ;
  assign y1818 = ~n4102 ;
  assign y1819 = ~1'b0 ;
  assign y1820 = ~1'b0 ;
  assign y1821 = n4105 ;
  assign y1822 = n4107 ;
  assign y1823 = ~n4109 ;
  assign y1824 = ~n4117 ;
  assign y1825 = ~n4119 ;
  assign y1826 = ~1'b0 ;
  assign y1827 = ~1'b0 ;
  assign y1828 = ~1'b0 ;
  assign y1829 = ~1'b0 ;
  assign y1830 = ~n4120 ;
  assign y1831 = n3550 ;
  assign y1832 = ~n4134 ;
  assign y1833 = ~n4135 ;
  assign y1834 = n4137 ;
  assign y1835 = ~1'b0 ;
  assign y1836 = ~1'b0 ;
  assign y1837 = n4141 ;
  assign y1838 = ~1'b0 ;
  assign y1839 = n4149 ;
  assign y1840 = ~n4150 ;
  assign y1841 = ~n4151 ;
  assign y1842 = n4155 ;
  assign y1843 = ~1'b0 ;
  assign y1844 = ~n4156 ;
  assign y1845 = ~1'b0 ;
  assign y1846 = ~n4157 ;
  assign y1847 = ~1'b0 ;
  assign y1848 = n4161 ;
  assign y1849 = n4169 ;
  assign y1850 = n4174 ;
  assign y1851 = ~1'b0 ;
  assign y1852 = ~n4177 ;
  assign y1853 = ~1'b0 ;
  assign y1854 = ~n4183 ;
  assign y1855 = n4184 ;
  assign y1856 = n4187 ;
  assign y1857 = ~1'b0 ;
  assign y1858 = n4191 ;
  assign y1859 = ~n4192 ;
  assign y1860 = n4194 ;
  assign y1861 = n4195 ;
  assign y1862 = ~n4197 ;
  assign y1863 = ~n3636 ;
  assign y1864 = n4199 ;
  assign y1865 = ~1'b0 ;
  assign y1866 = n4200 ;
  assign y1867 = ~1'b0 ;
  assign y1868 = ~n3404 ;
  assign y1869 = ~n4201 ;
  assign y1870 = n4204 ;
  assign y1871 = ~1'b0 ;
  assign y1872 = n821 ;
  assign y1873 = ~n4205 ;
  assign y1874 = n4207 ;
  assign y1875 = ~n4208 ;
  assign y1876 = ~n4221 ;
  assign y1877 = ~1'b0 ;
  assign y1878 = n4222 ;
  assign y1879 = ~n4225 ;
  assign y1880 = 1'b0 ;
  assign y1881 = ~n4227 ;
  assign y1882 = n4230 ;
  assign y1883 = ~n4233 ;
  assign y1884 = ~n4235 ;
  assign y1885 = n4240 ;
  assign y1886 = n4242 ;
  assign y1887 = ~n4243 ;
  assign y1888 = ~1'b0 ;
  assign y1889 = ~1'b0 ;
  assign y1890 = n4244 ;
  assign y1891 = ~1'b0 ;
  assign y1892 = ~n4247 ;
  assign y1893 = ~1'b0 ;
  assign y1894 = n4251 ;
  assign y1895 = n4253 ;
  assign y1896 = n4255 ;
  assign y1897 = ~n2956 ;
  assign y1898 = ~1'b0 ;
  assign y1899 = ~1'b0 ;
  assign y1900 = ~n4259 ;
  assign y1901 = ~n4260 ;
  assign y1902 = ~n4261 ;
  assign y1903 = ~1'b0 ;
  assign y1904 = ~1'b0 ;
  assign y1905 = ~n4263 ;
  assign y1906 = n4265 ;
  assign y1907 = n4266 ;
  assign y1908 = ~n3733 ;
  assign y1909 = ~n4268 ;
  assign y1910 = ~n4280 ;
  assign y1911 = ~n4283 ;
  assign y1912 = ~n4287 ;
  assign y1913 = ~n4292 ;
  assign y1914 = ~n4293 ;
  assign y1915 = ~1'b0 ;
  assign y1916 = ~1'b0 ;
  assign y1917 = n4295 ;
  assign y1918 = n4296 ;
  assign y1919 = ~1'b0 ;
  assign y1920 = x112 ;
  assign y1921 = ~1'b0 ;
  assign y1922 = ~n4297 ;
  assign y1923 = n4299 ;
  assign y1924 = 1'b0 ;
  assign y1925 = ~1'b0 ;
  assign y1926 = ~n4300 ;
  assign y1927 = n4302 ;
  assign y1928 = ~1'b0 ;
  assign y1929 = ~n4303 ;
  assign y1930 = n4304 ;
  assign y1931 = ~n3988 ;
  assign y1932 = ~n519 ;
  assign y1933 = n3730 ;
  assign y1934 = ~n4308 ;
  assign y1935 = ~n4310 ;
  assign y1936 = ~n2014 ;
  assign y1937 = ~1'b0 ;
  assign y1938 = ~n4313 ;
  assign y1939 = ~n4314 ;
  assign y1940 = ~n4318 ;
  assign y1941 = ~1'b0 ;
  assign y1942 = ~n1481 ;
  assign y1943 = n2340 ;
  assign y1944 = 1'b0 ;
  assign y1945 = ~n4320 ;
  assign y1946 = ~n4325 ;
  assign y1947 = ~1'b0 ;
  assign y1948 = ~1'b0 ;
  assign y1949 = ~n4327 ;
  assign y1950 = n4330 ;
  assign y1951 = n4331 ;
  assign y1952 = ~1'b0 ;
  assign y1953 = n4333 ;
  assign y1954 = n747 ;
  assign y1955 = n4334 ;
  assign y1956 = 1'b0 ;
  assign y1957 = n4337 ;
  assign y1958 = n4338 ;
  assign y1959 = ~1'b0 ;
  assign y1960 = ~1'b0 ;
  assign y1961 = ~n4345 ;
  assign y1962 = ~1'b0 ;
  assign y1963 = n4348 ;
  assign y1964 = n4353 ;
  assign y1965 = ~n4354 ;
  assign y1966 = n4355 ;
  assign y1967 = ~n4360 ;
  assign y1968 = ~1'b0 ;
  assign y1969 = ~1'b0 ;
  assign y1970 = ~1'b0 ;
  assign y1971 = n4362 ;
  assign y1972 = ~n4365 ;
  assign y1973 = ~1'b0 ;
  assign y1974 = ~1'b0 ;
  assign y1975 = ~n1150 ;
  assign y1976 = ~n4366 ;
  assign y1977 = ~1'b0 ;
  assign y1978 = ~n4369 ;
  assign y1979 = ~1'b0 ;
  assign y1980 = 1'b0 ;
  assign y1981 = n4375 ;
  assign y1982 = ~n1231 ;
  assign y1983 = ~n1219 ;
  assign y1984 = ~1'b0 ;
  assign y1985 = ~1'b0 ;
  assign y1986 = n4382 ;
  assign y1987 = n4387 ;
  assign y1988 = ~1'b0 ;
  assign y1989 = n4388 ;
  assign y1990 = ~1'b0 ;
  assign y1991 = n4391 ;
  assign y1992 = n4393 ;
  assign y1993 = ~n4394 ;
  assign y1994 = ~1'b0 ;
  assign y1995 = ~1'b0 ;
  assign y1996 = n732 ;
  assign y1997 = n4396 ;
  assign y1998 = ~1'b0 ;
  assign y1999 = ~n4402 ;
  assign y2000 = ~1'b0 ;
  assign y2001 = n4407 ;
  assign y2002 = ~1'b0 ;
  assign y2003 = n4409 ;
  assign y2004 = n4412 ;
  assign y2005 = ~n2211 ;
  assign y2006 = ~n4415 ;
  assign y2007 = ~1'b0 ;
  assign y2008 = ~1'b0 ;
  assign y2009 = ~n4424 ;
  assign y2010 = n4427 ;
  assign y2011 = n4428 ;
  assign y2012 = ~n4434 ;
  assign y2013 = ~1'b0 ;
  assign y2014 = ~n4436 ;
  assign y2015 = ~n4438 ;
  assign y2016 = ~1'b0 ;
  assign y2017 = n4441 ;
  assign y2018 = n4443 ;
  assign y2019 = ~1'b0 ;
  assign y2020 = ~n4445 ;
  assign y2021 = n4451 ;
  assign y2022 = n4452 ;
  assign y2023 = n4454 ;
  assign y2024 = n4456 ;
  assign y2025 = n4458 ;
  assign y2026 = ~n4459 ;
  assign y2027 = ~n4465 ;
  assign y2028 = n4470 ;
  assign y2029 = n4471 ;
  assign y2030 = n4472 ;
  assign y2031 = ~1'b0 ;
  assign y2032 = ~1'b0 ;
  assign y2033 = n3887 ;
  assign y2034 = n4474 ;
  assign y2035 = n4476 ;
  assign y2036 = n4477 ;
  assign y2037 = n4478 ;
  assign y2038 = ~n4480 ;
  assign y2039 = ~1'b0 ;
  assign y2040 = ~1'b0 ;
  assign y2041 = ~1'b0 ;
  assign y2042 = ~n4481 ;
  assign y2043 = 1'b0 ;
  assign y2044 = ~n4486 ;
  assign y2045 = ~1'b0 ;
  assign y2046 = ~1'b0 ;
  assign y2047 = ~n4491 ;
  assign y2048 = ~n4493 ;
  assign y2049 = ~n4498 ;
  assign y2050 = ~1'b0 ;
  assign y2051 = ~1'b0 ;
  assign y2052 = ~1'b0 ;
  assign y2053 = n4510 ;
  assign y2054 = n4511 ;
  assign y2055 = ~1'b0 ;
  assign y2056 = ~n4512 ;
  assign y2057 = n4521 ;
  assign y2058 = n4523 ;
  assign y2059 = ~n4526 ;
  assign y2060 = ~1'b0 ;
  assign y2061 = ~n2246 ;
  assign y2062 = n4534 ;
  assign y2063 = ~1'b0 ;
  assign y2064 = ~n4540 ;
  assign y2065 = ~n630 ;
  assign y2066 = ~1'b0 ;
  assign y2067 = ~n4541 ;
  assign y2068 = n4542 ;
  assign y2069 = ~1'b0 ;
  assign y2070 = ~1'b0 ;
  assign y2071 = ~1'b0 ;
  assign y2072 = ~n152 ;
  assign y2073 = ~1'b0 ;
  assign y2074 = n4543 ;
  assign y2075 = ~n4547 ;
  assign y2076 = ~1'b0 ;
  assign y2077 = n4548 ;
  assign y2078 = ~n4549 ;
  assign y2079 = ~n4554 ;
  assign y2080 = n4562 ;
  assign y2081 = ~n4568 ;
  assign y2082 = ~n4569 ;
  assign y2083 = n4572 ;
  assign y2084 = n4576 ;
  assign y2085 = n4578 ;
  assign y2086 = n4581 ;
  assign y2087 = ~n569 ;
  assign y2088 = n1790 ;
  assign y2089 = ~n4585 ;
  assign y2090 = ~n4588 ;
  assign y2091 = ~1'b0 ;
  assign y2092 = ~1'b0 ;
  assign y2093 = n4593 ;
  assign y2094 = ~1'b0 ;
  assign y2095 = ~1'b0 ;
  assign y2096 = ~n4598 ;
  assign y2097 = ~1'b0 ;
  assign y2098 = n477 ;
  assign y2099 = ~n4602 ;
  assign y2100 = n4603 ;
  assign y2101 = ~n4605 ;
  assign y2102 = ~1'b0 ;
  assign y2103 = ~1'b0 ;
  assign y2104 = ~n4608 ;
  assign y2105 = n4610 ;
  assign y2106 = n4612 ;
  assign y2107 = ~1'b0 ;
  assign y2108 = ~n4613 ;
  assign y2109 = ~n4616 ;
  assign y2110 = ~n4618 ;
  assign y2111 = ~n4621 ;
  assign y2112 = n4624 ;
  assign y2113 = ~1'b0 ;
  assign y2114 = ~1'b0 ;
  assign y2115 = ~1'b0 ;
  assign y2116 = n851 ;
  assign y2117 = ~n4631 ;
  assign y2118 = ~n4635 ;
  assign y2119 = n4380 ;
  assign y2120 = ~n4638 ;
  assign y2121 = ~1'b0 ;
  assign y2122 = ~1'b0 ;
  assign y2123 = ~n4640 ;
  assign y2124 = ~n4647 ;
  assign y2125 = ~n4648 ;
  assign y2126 = ~1'b0 ;
  assign y2127 = ~1'b0 ;
  assign y2128 = ~n4649 ;
  assign y2129 = ~n4650 ;
  assign y2130 = n4655 ;
  assign y2131 = ~n4664 ;
  assign y2132 = n4665 ;
  assign y2133 = n4666 ;
  assign y2134 = ~1'b0 ;
  assign y2135 = n4669 ;
  assign y2136 = ~n4675 ;
  assign y2137 = n4676 ;
  assign y2138 = ~1'b0 ;
  assign y2139 = n4686 ;
  assign y2140 = ~1'b0 ;
  assign y2141 = n538 ;
  assign y2142 = ~1'b0 ;
  assign y2143 = n4690 ;
  assign y2144 = ~1'b0 ;
  assign y2145 = n4693 ;
  assign y2146 = ~1'b0 ;
  assign y2147 = n4694 ;
  assign y2148 = n4696 ;
  assign y2149 = n4697 ;
  assign y2150 = x94 ;
  assign y2151 = n4698 ;
  assign y2152 = n4707 ;
  assign y2153 = ~1'b0 ;
  assign y2154 = n4708 ;
  assign y2155 = ~n4712 ;
  assign y2156 = ~1'b0 ;
  assign y2157 = ~n4714 ;
  assign y2158 = ~n4716 ;
  assign y2159 = ~n4719 ;
  assign y2160 = ~1'b0 ;
  assign y2161 = ~1'b0 ;
  assign y2162 = ~1'b0 ;
  assign y2163 = ~n4724 ;
  assign y2164 = ~1'b0 ;
  assign y2165 = ~n4729 ;
  assign y2166 = ~1'b0 ;
  assign y2167 = ~n4730 ;
  assign y2168 = n4731 ;
  assign y2169 = n4734 ;
  assign y2170 = n4739 ;
  assign y2171 = ~n4740 ;
  assign y2172 = ~n4747 ;
  assign y2173 = n4748 ;
  assign y2174 = n4750 ;
  assign y2175 = ~1'b0 ;
  assign y2176 = ~n4753 ;
  assign y2177 = n3961 ;
  assign y2178 = n4761 ;
  assign y2179 = ~n4763 ;
  assign y2180 = ~n4767 ;
  assign y2181 = n4773 ;
  assign y2182 = n4774 ;
  assign y2183 = ~n4777 ;
  assign y2184 = n4778 ;
  assign y2185 = ~1'b0 ;
  assign y2186 = ~1'b0 ;
  assign y2187 = ~1'b0 ;
  assign y2188 = ~n4782 ;
  assign y2189 = ~1'b0 ;
  assign y2190 = ~n4783 ;
  assign y2191 = n4784 ;
  assign y2192 = ~1'b0 ;
  assign y2193 = n4786 ;
  assign y2194 = ~n4788 ;
  assign y2195 = ~n4790 ;
  assign y2196 = n4791 ;
  assign y2197 = ~n4792 ;
  assign y2198 = ~n4793 ;
  assign y2199 = ~1'b0 ;
  assign y2200 = ~1'b0 ;
  assign y2201 = ~n4797 ;
  assign y2202 = n4802 ;
  assign y2203 = ~n4808 ;
  assign y2204 = x54 ;
  assign y2205 = n4809 ;
  assign y2206 = ~n4811 ;
  assign y2207 = ~n4815 ;
  assign y2208 = n2103 ;
  assign y2209 = n4820 ;
  assign y2210 = ~1'b0 ;
  assign y2211 = ~1'b0 ;
  assign y2212 = n4821 ;
  assign y2213 = ~1'b0 ;
  assign y2214 = n4292 ;
  assign y2215 = ~n4822 ;
  assign y2216 = n4823 ;
  assign y2217 = ~1'b0 ;
  assign y2218 = ~n4826 ;
  assign y2219 = ~n4829 ;
  assign y2220 = ~1'b0 ;
  assign y2221 = ~n4832 ;
  assign y2222 = 1'b0 ;
  assign y2223 = ~1'b0 ;
  assign y2224 = n4834 ;
  assign y2225 = n4837 ;
  assign y2226 = n4840 ;
  assign y2227 = n4843 ;
  assign y2228 = n4266 ;
  assign y2229 = n4849 ;
  assign y2230 = ~1'b0 ;
  assign y2231 = n3482 ;
  assign y2232 = ~n4853 ;
  assign y2233 = n4859 ;
  assign y2234 = ~1'b0 ;
  assign y2235 = n4861 ;
  assign y2236 = ~n4872 ;
  assign y2237 = ~1'b0 ;
  assign y2238 = ~1'b0 ;
  assign y2239 = n4879 ;
  assign y2240 = n4880 ;
  assign y2241 = ~1'b0 ;
  assign y2242 = 1'b0 ;
  assign y2243 = ~n4883 ;
  assign y2244 = n4884 ;
  assign y2245 = n4886 ;
  assign y2246 = ~n4887 ;
  assign y2247 = n3365 ;
  assign y2248 = ~1'b0 ;
  assign y2249 = n4892 ;
  assign y2250 = ~1'b0 ;
  assign y2251 = ~1'b0 ;
  assign y2252 = ~1'b0 ;
  assign y2253 = ~1'b0 ;
  assign y2254 = ~1'b0 ;
  assign y2255 = ~n4893 ;
  assign y2256 = ~n4898 ;
  assign y2257 = ~n4901 ;
  assign y2258 = n4902 ;
  assign y2259 = ~1'b0 ;
  assign y2260 = ~1'b0 ;
  assign y2261 = ~1'b0 ;
  assign y2262 = ~n4905 ;
  assign y2263 = n4906 ;
  assign y2264 = ~n4910 ;
  assign y2265 = n4912 ;
  assign y2266 = n4917 ;
  assign y2267 = n4918 ;
  assign y2268 = ~n4924 ;
  assign y2269 = 1'b0 ;
  assign y2270 = n4925 ;
  assign y2271 = n4929 ;
  assign y2272 = ~n4933 ;
  assign y2273 = n4935 ;
  assign y2274 = ~1'b0 ;
  assign y2275 = ~n4938 ;
  assign y2276 = n4940 ;
  assign y2277 = ~n4941 ;
  assign y2278 = ~n4942 ;
  assign y2279 = ~n4944 ;
  assign y2280 = ~n4945 ;
  assign y2281 = ~n4955 ;
  assign y2282 = n4965 ;
  assign y2283 = n4966 ;
  assign y2284 = ~n4969 ;
  assign y2285 = ~1'b0 ;
  assign y2286 = ~1'b0 ;
  assign y2287 = ~n4970 ;
  assign y2288 = ~n4973 ;
  assign y2289 = n496 ;
  assign y2290 = ~n4978 ;
  assign y2291 = n4979 ;
  assign y2292 = ~1'b0 ;
  assign y2293 = n4985 ;
  assign y2294 = n4989 ;
  assign y2295 = ~n4990 ;
  assign y2296 = n4992 ;
  assign y2297 = ~1'b0 ;
  assign y2298 = n4995 ;
  assign y2299 = ~1'b0 ;
  assign y2300 = n4997 ;
  assign y2301 = ~n4999 ;
  assign y2302 = ~n5002 ;
  assign y2303 = ~1'b0 ;
  assign y2304 = ~n4516 ;
  assign y2305 = n5004 ;
  assign y2306 = ~1'b0 ;
  assign y2307 = ~1'b0 ;
  assign y2308 = ~n5005 ;
  assign y2309 = n5007 ;
  assign y2310 = ~n5009 ;
  assign y2311 = ~n5011 ;
  assign y2312 = ~1'b0 ;
  assign y2313 = ~1'b0 ;
  assign y2314 = n5012 ;
  assign y2315 = ~1'b0 ;
  assign y2316 = ~1'b0 ;
  assign y2317 = ~1'b0 ;
  assign y2318 = n5016 ;
  assign y2319 = ~n5020 ;
  assign y2320 = ~n5023 ;
  assign y2321 = ~1'b0 ;
  assign y2322 = n5031 ;
  assign y2323 = ~1'b0 ;
  assign y2324 = ~1'b0 ;
  assign y2325 = ~1'b0 ;
  assign y2326 = n5038 ;
  assign y2327 = n5040 ;
  assign y2328 = n5046 ;
  assign y2329 = ~n5049 ;
  assign y2330 = n5052 ;
  assign y2331 = ~1'b0 ;
  assign y2332 = ~1'b0 ;
  assign y2333 = n5053 ;
  assign y2334 = ~n3354 ;
  assign y2335 = n5054 ;
  assign y2336 = ~n5059 ;
  assign y2337 = ~1'b0 ;
  assign y2338 = ~1'b0 ;
  assign y2339 = n5062 ;
  assign y2340 = n5063 ;
  assign y2341 = ~n5067 ;
  assign y2342 = ~1'b0 ;
  assign y2343 = ~1'b0 ;
  assign y2344 = n5071 ;
  assign y2345 = n5074 ;
  assign y2346 = ~1'b0 ;
  assign y2347 = ~1'b0 ;
  assign y2348 = n5079 ;
  assign y2349 = ~1'b0 ;
  assign y2350 = n5080 ;
  assign y2351 = ~1'b0 ;
  assign y2352 = ~1'b0 ;
  assign y2353 = ~n5082 ;
  assign y2354 = ~n5083 ;
  assign y2355 = n5084 ;
  assign y2356 = ~1'b0 ;
  assign y2357 = ~1'b0 ;
  assign y2358 = n5091 ;
  assign y2359 = ~1'b0 ;
  assign y2360 = ~n5092 ;
  assign y2361 = n5098 ;
  assign y2362 = n5100 ;
  assign y2363 = ~1'b0 ;
  assign y2364 = ~n5102 ;
  assign y2365 = n5107 ;
  assign y2366 = ~1'b0 ;
  assign y2367 = ~1'b0 ;
  assign y2368 = ~n5111 ;
  assign y2369 = ~n5115 ;
  assign y2370 = ~n5117 ;
  assign y2371 = n5122 ;
  assign y2372 = n5132 ;
  assign y2373 = ~1'b0 ;
  assign y2374 = ~n5133 ;
  assign y2375 = ~n5134 ;
  assign y2376 = ~n5135 ;
  assign y2377 = n5137 ;
  assign y2378 = n5138 ;
  assign y2379 = ~1'b0 ;
  assign y2380 = ~n5140 ;
  assign y2381 = ~n5142 ;
  assign y2382 = n5143 ;
  assign y2383 = ~n5145 ;
  assign y2384 = ~n5146 ;
  assign y2385 = ~n5148 ;
  assign y2386 = ~1'b0 ;
  assign y2387 = ~1'b0 ;
  assign y2388 = ~1'b0 ;
  assign y2389 = ~n5152 ;
  assign y2390 = ~1'b0 ;
  assign y2391 = ~n5156 ;
  assign y2392 = 1'b0 ;
  assign y2393 = ~n5163 ;
  assign y2394 = n5165 ;
  assign y2395 = ~1'b0 ;
  assign y2396 = ~1'b0 ;
  assign y2397 = n5166 ;
  assign y2398 = ~1'b0 ;
  assign y2399 = ~1'b0 ;
  assign y2400 = n5167 ;
  assign y2401 = n5170 ;
  assign y2402 = n5171 ;
  assign y2403 = ~1'b0 ;
  assign y2404 = ~n5172 ;
  assign y2405 = n5177 ;
  assign y2406 = ~n5179 ;
  assign y2407 = ~n5187 ;
  assign y2408 = n5202 ;
  assign y2409 = ~1'b0 ;
  assign y2410 = n5203 ;
  assign y2411 = n5207 ;
  assign y2412 = ~n901 ;
  assign y2413 = ~1'b0 ;
  assign y2414 = n5215 ;
  assign y2415 = ~1'b0 ;
  assign y2416 = 1'b0 ;
  assign y2417 = ~1'b0 ;
  assign y2418 = n5219 ;
  assign y2419 = ~n5222 ;
  assign y2420 = ~1'b0 ;
  assign y2421 = ~1'b0 ;
  assign y2422 = n5224 ;
  assign y2423 = ~n5230 ;
  assign y2424 = ~n5231 ;
  assign y2425 = n5232 ;
  assign y2426 = ~1'b0 ;
  assign y2427 = ~n5235 ;
  assign y2428 = n5241 ;
  assign y2429 = ~n5242 ;
  assign y2430 = ~1'b0 ;
  assign y2431 = n5246 ;
  assign y2432 = ~1'b0 ;
  assign y2433 = ~1'b0 ;
  assign y2434 = n5261 ;
  assign y2435 = ~n5273 ;
  assign y2436 = ~1'b0 ;
  assign y2437 = ~1'b0 ;
  assign y2438 = n5274 ;
  assign y2439 = n4007 ;
  assign y2440 = ~n5276 ;
  assign y2441 = ~n5277 ;
  assign y2442 = n4204 ;
  assign y2443 = ~n5279 ;
  assign y2444 = ~1'b0 ;
  assign y2445 = n5283 ;
  assign y2446 = ~n5284 ;
  assign y2447 = 1'b0 ;
  assign y2448 = n5289 ;
  assign y2449 = ~1'b0 ;
  assign y2450 = ~n5294 ;
  assign y2451 = n5298 ;
  assign y2452 = n5302 ;
  assign y2453 = ~n5304 ;
  assign y2454 = ~n5305 ;
  assign y2455 = ~n5310 ;
  assign y2456 = ~1'b0 ;
  assign y2457 = ~n5311 ;
  assign y2458 = ~n476 ;
  assign y2459 = ~n5315 ;
  assign y2460 = ~n5317 ;
  assign y2461 = ~n5318 ;
  assign y2462 = n5323 ;
  assign y2463 = ~n5326 ;
  assign y2464 = n5327 ;
  assign y2465 = n5331 ;
  assign y2466 = ~n5340 ;
  assign y2467 = ~n5344 ;
  assign y2468 = ~1'b0 ;
  assign y2469 = ~1'b0 ;
  assign y2470 = ~1'b0 ;
  assign y2471 = ~n5347 ;
  assign y2472 = ~1'b0 ;
  assign y2473 = ~1'b0 ;
  assign y2474 = ~1'b0 ;
  assign y2475 = ~1'b0 ;
  assign y2476 = ~n5348 ;
  assign y2477 = ~n5349 ;
  assign y2478 = ~n5351 ;
  assign y2479 = n5354 ;
  assign y2480 = n5355 ;
  assign y2481 = ~1'b0 ;
  assign y2482 = n5360 ;
  assign y2483 = ~n5364 ;
  assign y2484 = ~n5368 ;
  assign y2485 = n5370 ;
  assign y2486 = ~1'b0 ;
  assign y2487 = ~1'b0 ;
  assign y2488 = ~1'b0 ;
  assign y2489 = ~n5375 ;
  assign y2490 = n2204 ;
  assign y2491 = ~n5376 ;
  assign y2492 = ~n5381 ;
  assign y2493 = n5387 ;
  assign y2494 = n583 ;
  assign y2495 = ~n5389 ;
  assign y2496 = n2409 ;
  assign y2497 = n5394 ;
  assign y2498 = n5400 ;
  assign y2499 = n5402 ;
  assign y2500 = ~n5404 ;
  assign y2501 = n5408 ;
  assign y2502 = n5410 ;
  assign y2503 = n5413 ;
  assign y2504 = n5419 ;
  assign y2505 = n5423 ;
  assign y2506 = ~1'b0 ;
  assign y2507 = ~1'b0 ;
  assign y2508 = n5427 ;
  assign y2509 = n5430 ;
  assign y2510 = n5431 ;
  assign y2511 = n5432 ;
  assign y2512 = ~1'b0 ;
  assign y2513 = n5435 ;
  assign y2514 = ~n5437 ;
  assign y2515 = 1'b0 ;
  assign y2516 = ~1'b0 ;
  assign y2517 = n5442 ;
  assign y2518 = n5446 ;
  assign y2519 = ~n5450 ;
  assign y2520 = ~1'b0 ;
  assign y2521 = ~n5451 ;
  assign y2522 = ~1'b0 ;
  assign y2523 = ~n5453 ;
  assign y2524 = ~n5461 ;
  assign y2525 = n5462 ;
  assign y2526 = ~1'b0 ;
  assign y2527 = ~1'b0 ;
  assign y2528 = ~1'b0 ;
  assign y2529 = ~n5466 ;
  assign y2530 = ~1'b0 ;
  assign y2531 = ~1'b0 ;
  assign y2532 = ~n5467 ;
  assign y2533 = n3124 ;
  assign y2534 = ~n5468 ;
  assign y2535 = ~n5471 ;
  assign y2536 = ~n5473 ;
  assign y2537 = ~1'b0 ;
  assign y2538 = n5479 ;
  assign y2539 = ~n5481 ;
  assign y2540 = ~n5484 ;
  assign y2541 = ~1'b0 ;
  assign y2542 = ~1'b0 ;
  assign y2543 = ~n5485 ;
  assign y2544 = n5487 ;
  assign y2545 = ~n5495 ;
  assign y2546 = ~n5497 ;
  assign y2547 = ~n5499 ;
  assign y2548 = ~n5503 ;
  assign y2549 = ~n5504 ;
  assign y2550 = n5506 ;
  assign y2551 = ~n5507 ;
  assign y2552 = ~n5508 ;
  assign y2553 = ~n5510 ;
  assign y2554 = n5516 ;
  assign y2555 = ~n5519 ;
  assign y2556 = ~n5523 ;
  assign y2557 = ~1'b0 ;
  assign y2558 = ~n5524 ;
  assign y2559 = ~1'b0 ;
  assign y2560 = ~n5529 ;
  assign y2561 = ~n5535 ;
  assign y2562 = ~1'b0 ;
  assign y2563 = ~n5537 ;
  assign y2564 = n5538 ;
  assign y2565 = ~1'b0 ;
  assign y2566 = n5542 ;
  assign y2567 = n5544 ;
  assign y2568 = ~1'b0 ;
  assign y2569 = ~1'b0 ;
  assign y2570 = ~n5554 ;
  assign y2571 = ~n5561 ;
  assign y2572 = n5568 ;
  assign y2573 = ~n1247 ;
  assign y2574 = ~1'b0 ;
  assign y2575 = ~1'b0 ;
  assign y2576 = ~n5569 ;
  assign y2577 = ~1'b0 ;
  assign y2578 = 1'b0 ;
  assign y2579 = n5573 ;
  assign y2580 = ~n5574 ;
  assign y2581 = ~1'b0 ;
  assign y2582 = n5575 ;
  assign y2583 = ~1'b0 ;
  assign y2584 = n5577 ;
  assign y2585 = ~n5578 ;
  assign y2586 = ~1'b0 ;
  assign y2587 = ~n5582 ;
  assign y2588 = n5588 ;
  assign y2589 = n5592 ;
  assign y2590 = ~n5595 ;
  assign y2591 = ~n5597 ;
  assign y2592 = ~n5598 ;
  assign y2593 = ~n4547 ;
  assign y2594 = ~n5599 ;
  assign y2595 = ~1'b0 ;
  assign y2596 = ~1'b0 ;
  assign y2597 = 1'b0 ;
  assign y2598 = n5600 ;
  assign y2599 = n152 ;
  assign y2600 = ~n5603 ;
  assign y2601 = ~n5605 ;
  assign y2602 = ~1'b0 ;
  assign y2603 = ~n5606 ;
  assign y2604 = n5608 ;
  assign y2605 = 1'b0 ;
  assign y2606 = n5611 ;
  assign y2607 = n5620 ;
  assign y2608 = ~n5622 ;
  assign y2609 = ~n5623 ;
  assign y2610 = ~1'b0 ;
  assign y2611 = ~n5630 ;
  assign y2612 = ~1'b0 ;
  assign y2613 = ~n5642 ;
  assign y2614 = n5643 ;
  assign y2615 = n5644 ;
  assign y2616 = ~1'b0 ;
  assign y2617 = ~1'b0 ;
  assign y2618 = ~n3681 ;
  assign y2619 = ~1'b0 ;
  assign y2620 = ~1'b0 ;
  assign y2621 = ~n4107 ;
  assign y2622 = ~n5646 ;
  assign y2623 = ~1'b0 ;
  assign y2624 = ~1'b0 ;
  assign y2625 = n5647 ;
  assign y2626 = ~n5648 ;
  assign y2627 = ~1'b0 ;
  assign y2628 = ~n5651 ;
  assign y2629 = n5657 ;
  assign y2630 = n5661 ;
  assign y2631 = ~1'b0 ;
  assign y2632 = n5666 ;
  assign y2633 = n5669 ;
  assign y2634 = ~n5670 ;
  assign y2635 = ~n5671 ;
  assign y2636 = ~1'b0 ;
  assign y2637 = ~n5674 ;
  assign y2638 = ~n5677 ;
  assign y2639 = n5680 ;
  assign y2640 = ~n5683 ;
  assign y2641 = ~n5687 ;
  assign y2642 = n5692 ;
  assign y2643 = ~n5694 ;
  assign y2644 = ~n5696 ;
  assign y2645 = ~n5698 ;
  assign y2646 = ~n5699 ;
  assign y2647 = ~n5707 ;
  assign y2648 = ~1'b0 ;
  assign y2649 = ~n5709 ;
  assign y2650 = n5716 ;
  assign y2651 = ~n5718 ;
  assign y2652 = ~n5720 ;
  assign y2653 = n5721 ;
  assign y2654 = ~n5722 ;
  assign y2655 = ~1'b0 ;
  assign y2656 = ~n5726 ;
  assign y2657 = ~n5728 ;
  assign y2658 = ~n5730 ;
  assign y2659 = ~n5731 ;
  assign y2660 = ~1'b0 ;
  assign y2661 = ~1'b0 ;
  assign y2662 = ~n5735 ;
  assign y2663 = ~n391 ;
  assign y2664 = ~1'b0 ;
  assign y2665 = ~n5738 ;
  assign y2666 = ~n5739 ;
  assign y2667 = ~n5740 ;
  assign y2668 = ~n5741 ;
  assign y2669 = n5742 ;
  assign y2670 = ~1'b0 ;
  assign y2671 = n5745 ;
  assign y2672 = ~1'b0 ;
  assign y2673 = ~n5747 ;
  assign y2674 = ~1'b0 ;
  assign y2675 = ~n5752 ;
  assign y2676 = ~n5759 ;
  assign y2677 = ~1'b0 ;
  assign y2678 = ~n5760 ;
  assign y2679 = ~n5762 ;
  assign y2680 = n5763 ;
  assign y2681 = n5768 ;
  assign y2682 = ~1'b0 ;
  assign y2683 = n5772 ;
  assign y2684 = ~n5784 ;
  assign y2685 = ~1'b0 ;
  assign y2686 = ~n5790 ;
  assign y2687 = ~n5792 ;
  assign y2688 = ~n5794 ;
  assign y2689 = ~n5798 ;
  assign y2690 = ~1'b0 ;
  assign y2691 = ~n5802 ;
  assign y2692 = ~1'b0 ;
  assign y2693 = ~n5805 ;
  assign y2694 = ~n5809 ;
  assign y2695 = n5814 ;
  assign y2696 = ~n5816 ;
  assign y2697 = n5819 ;
  assign y2698 = n5820 ;
  assign y2699 = ~n5825 ;
  assign y2700 = ~1'b0 ;
  assign y2701 = n5827 ;
  assign y2702 = ~1'b0 ;
  assign y2703 = n5828 ;
  assign y2704 = n5834 ;
  assign y2705 = n5836 ;
  assign y2706 = ~n5841 ;
  assign y2707 = n5842 ;
  assign y2708 = ~n5845 ;
  assign y2709 = 1'b0 ;
  assign y2710 = n5848 ;
  assign y2711 = n5849 ;
  assign y2712 = ~n5850 ;
  assign y2713 = n5854 ;
  assign y2714 = n5858 ;
  assign y2715 = ~1'b0 ;
  assign y2716 = ~1'b0 ;
  assign y2717 = n5859 ;
  assign y2718 = n978 ;
  assign y2719 = n5862 ;
  assign y2720 = 1'b0 ;
  assign y2721 = ~1'b0 ;
  assign y2722 = ~1'b0 ;
  assign y2723 = ~1'b0 ;
  assign y2724 = ~n5865 ;
  assign y2725 = ~n5867 ;
  assign y2726 = ~n5870 ;
  assign y2727 = n5872 ;
  assign y2728 = ~n5876 ;
  assign y2729 = n5879 ;
  assign y2730 = ~n5886 ;
  assign y2731 = ~n5891 ;
  assign y2732 = ~1'b0 ;
  assign y2733 = ~n5899 ;
  assign y2734 = ~n5904 ;
  assign y2735 = n5905 ;
  assign y2736 = ~1'b0 ;
  assign y2737 = ~n5906 ;
  assign y2738 = n1439 ;
  assign y2739 = ~n4324 ;
  assign y2740 = n5909 ;
  assign y2741 = ~n5911 ;
  assign y2742 = ~1'b0 ;
  assign y2743 = ~n5920 ;
  assign y2744 = n5921 ;
  assign y2745 = ~n5925 ;
  assign y2746 = ~1'b0 ;
  assign y2747 = ~n5928 ;
  assign y2748 = ~1'b0 ;
  assign y2749 = ~1'b0 ;
  assign y2750 = ~n2204 ;
  assign y2751 = ~1'b0 ;
  assign y2752 = ~n5930 ;
  assign y2753 = n5931 ;
  assign y2754 = ~n5933 ;
  assign y2755 = ~1'b0 ;
  assign y2756 = ~n177 ;
  assign y2757 = ~1'b0 ;
  assign y2758 = n5934 ;
  assign y2759 = ~1'b0 ;
  assign y2760 = ~1'b0 ;
  assign y2761 = n5937 ;
  assign y2762 = ~n5941 ;
  assign y2763 = n5942 ;
  assign y2764 = ~1'b0 ;
  assign y2765 = n5945 ;
  assign y2766 = ~1'b0 ;
  assign y2767 = ~1'b0 ;
  assign y2768 = n5950 ;
  assign y2769 = n5951 ;
  assign y2770 = ~n5952 ;
  assign y2771 = n5954 ;
  assign y2772 = n5959 ;
  assign y2773 = n5961 ;
  assign y2774 = 1'b0 ;
  assign y2775 = n5963 ;
  assign y2776 = n5966 ;
  assign y2777 = ~1'b0 ;
  assign y2778 = ~1'b0 ;
  assign y2779 = n5967 ;
  assign y2780 = 1'b0 ;
  assign y2781 = n5969 ;
  assign y2782 = ~1'b0 ;
  assign y2783 = n5972 ;
  assign y2784 = ~1'b0 ;
  assign y2785 = ~n5977 ;
  assign y2786 = ~n5983 ;
  assign y2787 = ~n468 ;
  assign y2788 = n5985 ;
  assign y2789 = n5989 ;
  assign y2790 = ~n5992 ;
  assign y2791 = n5993 ;
  assign y2792 = n5997 ;
  assign y2793 = ~n6002 ;
  assign y2794 = ~1'b0 ;
  assign y2795 = ~1'b0 ;
  assign y2796 = ~n458 ;
  assign y2797 = n6003 ;
  assign y2798 = ~1'b0 ;
  assign y2799 = n6006 ;
  assign y2800 = ~n6017 ;
  assign y2801 = n6019 ;
  assign y2802 = n6020 ;
  assign y2803 = ~1'b0 ;
  assign y2804 = ~n6023 ;
  assign y2805 = ~n6025 ;
  assign y2806 = n6029 ;
  assign y2807 = ~n6034 ;
  assign y2808 = ~n6036 ;
  assign y2809 = n6038 ;
  assign y2810 = ~n6043 ;
  assign y2811 = n6044 ;
  assign y2812 = ~n6045 ;
  assign y2813 = ~1'b0 ;
  assign y2814 = ~1'b0 ;
  assign y2815 = n6047 ;
  assign y2816 = ~n2899 ;
  assign y2817 = ~1'b0 ;
  assign y2818 = ~n6052 ;
  assign y2819 = ~n6053 ;
  assign y2820 = ~1'b0 ;
  assign y2821 = ~n6055 ;
  assign y2822 = n6056 ;
  assign y2823 = n6059 ;
  assign y2824 = n6060 ;
  assign y2825 = n6062 ;
  assign y2826 = ~n6066 ;
  assign y2827 = n6072 ;
  assign y2828 = n6078 ;
  assign y2829 = ~n6086 ;
  assign y2830 = ~1'b0 ;
  assign y2831 = n6088 ;
  assign y2832 = ~n6092 ;
  assign y2833 = ~n6094 ;
  assign y2834 = n6097 ;
  assign y2835 = ~n6099 ;
  assign y2836 = n6104 ;
  assign y2837 = ~1'b0 ;
  assign y2838 = n6107 ;
  assign y2839 = ~1'b0 ;
  assign y2840 = ~1'b0 ;
  assign y2841 = n6110 ;
  assign y2842 = ~n6111 ;
  assign y2843 = ~1'b0 ;
  assign y2844 = ~1'b0 ;
  assign y2845 = ~1'b0 ;
  assign y2846 = n6115 ;
  assign y2847 = ~1'b0 ;
  assign y2848 = n6118 ;
  assign y2849 = ~n6122 ;
  assign y2850 = ~n6126 ;
  assign y2851 = ~n6129 ;
  assign y2852 = ~n6136 ;
  assign y2853 = n6138 ;
  assign y2854 = n6140 ;
  assign y2855 = ~n6156 ;
  assign y2856 = n6161 ;
  assign y2857 = ~1'b0 ;
  assign y2858 = n6166 ;
  assign y2859 = n6171 ;
  assign y2860 = ~n6177 ;
  assign y2861 = ~n6179 ;
  assign y2862 = n6182 ;
  assign y2863 = ~1'b0 ;
  assign y2864 = ~n6185 ;
  assign y2865 = n6190 ;
  assign y2866 = ~1'b0 ;
  assign y2867 = ~1'b0 ;
  assign y2868 = ~n6193 ;
  assign y2869 = ~n6201 ;
  assign y2870 = ~n6202 ;
  assign y2871 = ~n1597 ;
  assign y2872 = ~1'b0 ;
  assign y2873 = ~1'b0 ;
  assign y2874 = n6204 ;
  assign y2875 = n6205 ;
  assign y2876 = ~n6206 ;
  assign y2877 = n6213 ;
  assign y2878 = ~n6220 ;
  assign y2879 = n6224 ;
  assign y2880 = ~1'b0 ;
  assign y2881 = ~n6229 ;
  assign y2882 = n6233 ;
  assign y2883 = n6236 ;
  assign y2884 = n6238 ;
  assign y2885 = n6245 ;
  assign y2886 = 1'b0 ;
  assign y2887 = ~1'b0 ;
  assign y2888 = n6247 ;
  assign y2889 = n6249 ;
  assign y2890 = ~1'b0 ;
  assign y2891 = ~n6251 ;
  assign y2892 = 1'b0 ;
  assign y2893 = ~n5850 ;
  assign y2894 = ~n6254 ;
  assign y2895 = ~n6258 ;
  assign y2896 = ~1'b0 ;
  assign y2897 = ~n2433 ;
  assign y2898 = n6263 ;
  assign y2899 = ~1'b0 ;
  assign y2900 = ~n6269 ;
  assign y2901 = 1'b0 ;
  assign y2902 = ~n6275 ;
  assign y2903 = ~n6277 ;
  assign y2904 = ~n6286 ;
  assign y2905 = n6288 ;
  assign y2906 = ~n6289 ;
  assign y2907 = ~n6293 ;
  assign y2908 = ~n6299 ;
  assign y2909 = ~n6305 ;
  assign y2910 = n6307 ;
  assign y2911 = n6309 ;
  assign y2912 = ~n6311 ;
  assign y2913 = ~n6317 ;
  assign y2914 = ~n6319 ;
  assign y2915 = n6323 ;
  assign y2916 = ~1'b0 ;
  assign y2917 = n6324 ;
  assign y2918 = n6326 ;
  assign y2919 = ~n6331 ;
  assign y2920 = ~n6333 ;
  assign y2921 = ~n6336 ;
  assign y2922 = n6340 ;
  assign y2923 = ~n6342 ;
  assign y2924 = ~1'b0 ;
  assign y2925 = n6343 ;
  assign y2926 = n6347 ;
  assign y2927 = ~n6348 ;
  assign y2928 = ~1'b0 ;
  assign y2929 = 1'b0 ;
  assign y2930 = n6350 ;
  assign y2931 = n6359 ;
  assign y2932 = ~1'b0 ;
  assign y2933 = ~1'b0 ;
  assign y2934 = ~n6366 ;
  assign y2935 = ~1'b0 ;
  assign y2936 = ~n6367 ;
  assign y2937 = ~n6372 ;
  assign y2938 = n6376 ;
  assign y2939 = ~n6389 ;
  assign y2940 = n6392 ;
  assign y2941 = n6396 ;
  assign y2942 = n6397 ;
  assign y2943 = n6403 ;
  assign y2944 = n6409 ;
  assign y2945 = ~n6415 ;
  assign y2946 = n6419 ;
  assign y2947 = n6421 ;
  assign y2948 = ~1'b0 ;
  assign y2949 = 1'b0 ;
  assign y2950 = n6424 ;
  assign y2951 = n6428 ;
  assign y2952 = n6436 ;
  assign y2953 = ~n6438 ;
  assign y2954 = ~1'b0 ;
  assign y2955 = n6444 ;
  assign y2956 = ~1'b0 ;
  assign y2957 = 1'b0 ;
  assign y2958 = ~1'b0 ;
  assign y2959 = ~n6445 ;
  assign y2960 = n6449 ;
  assign y2961 = ~1'b0 ;
  assign y2962 = ~1'b0 ;
  assign y2963 = ~n6450 ;
  assign y2964 = n6452 ;
  assign y2965 = ~1'b0 ;
  assign y2966 = n586 ;
  assign y2967 = ~1'b0 ;
  assign y2968 = ~n6459 ;
  assign y2969 = n6463 ;
  assign y2970 = ~1'b0 ;
  assign y2971 = ~n6464 ;
  assign y2972 = ~n6468 ;
  assign y2973 = ~n6470 ;
  assign y2974 = ~n6473 ;
  assign y2975 = n6478 ;
  assign y2976 = ~1'b0 ;
  assign y2977 = ~n6275 ;
  assign y2978 = ~n6481 ;
  assign y2979 = ~n6484 ;
  assign y2980 = n6486 ;
  assign y2981 = 1'b0 ;
  assign y2982 = ~1'b0 ;
  assign y2983 = ~1'b0 ;
  assign y2984 = n6487 ;
  assign y2985 = ~1'b0 ;
  assign y2986 = n6491 ;
  assign y2987 = ~n6494 ;
  assign y2988 = ~1'b0 ;
  assign y2989 = n6495 ;
  assign y2990 = n6500 ;
  assign y2991 = n6504 ;
  assign y2992 = n6509 ;
  assign y2993 = ~1'b0 ;
  assign y2994 = n5492 ;
  assign y2995 = 1'b0 ;
  assign y2996 = ~n6515 ;
  assign y2997 = n377 ;
  assign y2998 = n6518 ;
  assign y2999 = ~n6520 ;
  assign y3000 = ~n6525 ;
  assign y3001 = n672 ;
  assign y3002 = ~n6526 ;
  assign y3003 = ~1'b0 ;
  assign y3004 = ~1'b0 ;
  assign y3005 = ~1'b0 ;
  assign y3006 = ~n6527 ;
  assign y3007 = ~n6535 ;
  assign y3008 = ~1'b0 ;
  assign y3009 = n6540 ;
  assign y3010 = ~1'b0 ;
  assign y3011 = ~1'b0 ;
  assign y3012 = ~n6544 ;
  assign y3013 = ~1'b0 ;
  assign y3014 = ~n4666 ;
  assign y3015 = n6547 ;
  assign y3016 = ~1'b0 ;
  assign y3017 = n1157 ;
  assign y3018 = ~n6549 ;
  assign y3019 = n6550 ;
  assign y3020 = n6563 ;
  assign y3021 = n6566 ;
  assign y3022 = n6580 ;
  assign y3023 = ~n6582 ;
  assign y3024 = ~1'b0 ;
  assign y3025 = ~1'b0 ;
  assign y3026 = n6585 ;
  assign y3027 = n6586 ;
  assign y3028 = ~n6588 ;
  assign y3029 = ~n6590 ;
  assign y3030 = ~n6592 ;
  assign y3031 = ~1'b0 ;
  assign y3032 = ~n3602 ;
  assign y3033 = ~n6597 ;
  assign y3034 = ~n6603 ;
  assign y3035 = ~1'b0 ;
  assign y3036 = n6604 ;
  assign y3037 = ~1'b0 ;
  assign y3038 = ~1'b0 ;
  assign y3039 = n6605 ;
  assign y3040 = ~n6606 ;
  assign y3041 = n6608 ;
  assign y3042 = ~1'b0 ;
  assign y3043 = ~1'b0 ;
  assign y3044 = n6609 ;
  assign y3045 = ~n6611 ;
  assign y3046 = ~1'b0 ;
  assign y3047 = ~n6612 ;
  assign y3048 = n4578 ;
  assign y3049 = ~n6614 ;
  assign y3050 = n6615 ;
  assign y3051 = n6616 ;
  assign y3052 = ~n6618 ;
  assign y3053 = n1880 ;
  assign y3054 = ~n6620 ;
  assign y3055 = n6621 ;
  assign y3056 = n6625 ;
  assign y3057 = ~1'b0 ;
  assign y3058 = n6626 ;
  assign y3059 = ~n6630 ;
  assign y3060 = ~n5736 ;
  assign y3061 = n6634 ;
  assign y3062 = n1406 ;
  assign y3063 = ~1'b0 ;
  assign y3064 = n6646 ;
  assign y3065 = ~1'b0 ;
  assign y3066 = ~n6648 ;
  assign y3067 = n6650 ;
  assign y3068 = ~1'b0 ;
  assign y3069 = 1'b0 ;
  assign y3070 = ~1'b0 ;
  assign y3071 = ~1'b0 ;
  assign y3072 = ~n6655 ;
  assign y3073 = ~1'b0 ;
  assign y3074 = n6658 ;
  assign y3075 = ~n6659 ;
  assign y3076 = n6663 ;
  assign y3077 = ~n6667 ;
  assign y3078 = ~1'b0 ;
  assign y3079 = ~1'b0 ;
  assign y3080 = n5635 ;
  assign y3081 = ~n6671 ;
  assign y3082 = ~n6672 ;
  assign y3083 = ~n6674 ;
  assign y3084 = ~n6676 ;
  assign y3085 = ~1'b0 ;
  assign y3086 = n6677 ;
  assign y3087 = ~n6684 ;
  assign y3088 = n6688 ;
  assign y3089 = ~1'b0 ;
  assign y3090 = ~1'b0 ;
  assign y3091 = ~1'b0 ;
  assign y3092 = n6689 ;
  assign y3093 = n6690 ;
  assign y3094 = n2635 ;
  assign y3095 = ~1'b0 ;
  assign y3096 = ~n6693 ;
  assign y3097 = ~1'b0 ;
  assign y3098 = n6695 ;
  assign y3099 = ~n6698 ;
  assign y3100 = n6702 ;
  assign y3101 = n6714 ;
  assign y3102 = ~1'b0 ;
  assign y3103 = n6719 ;
  assign y3104 = ~n6721 ;
  assign y3105 = ~1'b0 ;
  assign y3106 = ~1'b0 ;
  assign y3107 = n6725 ;
  assign y3108 = ~1'b0 ;
  assign y3109 = ~1'b0 ;
  assign y3110 = ~1'b0 ;
  assign y3111 = ~1'b0 ;
  assign y3112 = ~n6727 ;
  assign y3113 = ~1'b0 ;
  assign y3114 = ~1'b0 ;
  assign y3115 = ~n6728 ;
  assign y3116 = ~n2494 ;
  assign y3117 = n6729 ;
  assign y3118 = ~1'b0 ;
  assign y3119 = n6735 ;
  assign y3120 = n6737 ;
  assign y3121 = ~1'b0 ;
  assign y3122 = ~n6739 ;
  assign y3123 = ~n6744 ;
  assign y3124 = ~n6746 ;
  assign y3125 = ~n6747 ;
  assign y3126 = ~1'b0 ;
  assign y3127 = ~1'b0 ;
  assign y3128 = n6748 ;
  assign y3129 = n6755 ;
  assign y3130 = n6757 ;
  assign y3131 = ~1'b0 ;
  assign y3132 = ~1'b0 ;
  assign y3133 = n6758 ;
  assign y3134 = ~n6760 ;
  assign y3135 = n6771 ;
  assign y3136 = ~n6776 ;
  assign y3137 = n2479 ;
  assign y3138 = ~1'b0 ;
  assign y3139 = ~n6784 ;
  assign y3140 = ~1'b0 ;
  assign y3141 = ~n6787 ;
  assign y3142 = n5737 ;
  assign y3143 = ~n6789 ;
  assign y3144 = ~1'b0 ;
  assign y3145 = ~n6791 ;
  assign y3146 = n6793 ;
  assign y3147 = ~n6794 ;
  assign y3148 = n6796 ;
  assign y3149 = ~n6797 ;
  assign y3150 = n6800 ;
  assign y3151 = ~n6801 ;
  assign y3152 = ~n6802 ;
  assign y3153 = ~1'b0 ;
  assign y3154 = ~1'b0 ;
  assign y3155 = ~1'b0 ;
  assign y3156 = ~n6804 ;
  assign y3157 = 1'b0 ;
  assign y3158 = n6805 ;
  assign y3159 = n6809 ;
  assign y3160 = n6813 ;
  assign y3161 = n6815 ;
  assign y3162 = ~n6818 ;
  assign y3163 = ~n6823 ;
  assign y3164 = n6827 ;
  assign y3165 = ~n6828 ;
  assign y3166 = ~n6833 ;
  assign y3167 = ~n6834 ;
  assign y3168 = n6835 ;
  assign y3169 = ~n5647 ;
  assign y3170 = ~n6836 ;
  assign y3171 = ~n6839 ;
  assign y3172 = ~n3276 ;
  assign y3173 = n6840 ;
  assign y3174 = ~1'b0 ;
  assign y3175 = n6848 ;
  assign y3176 = n6854 ;
  assign y3177 = ~n6857 ;
  assign y3178 = ~n6860 ;
  assign y3179 = ~1'b0 ;
  assign y3180 = n6861 ;
  assign y3181 = n6867 ;
  assign y3182 = n6869 ;
  assign y3183 = ~1'b0 ;
  assign y3184 = n2337 ;
  assign y3185 = ~1'b0 ;
  assign y3186 = ~1'b0 ;
  assign y3187 = ~1'b0 ;
  assign y3188 = n6871 ;
  assign y3189 = n6872 ;
  assign y3190 = ~1'b0 ;
  assign y3191 = ~1'b0 ;
  assign y3192 = ~n6873 ;
  assign y3193 = n6876 ;
  assign y3194 = n6883 ;
  assign y3195 = n6886 ;
  assign y3196 = ~1'b0 ;
  assign y3197 = n6888 ;
  assign y3198 = ~1'b0 ;
  assign y3199 = ~n6896 ;
  assign y3200 = n6898 ;
  assign y3201 = ~1'b0 ;
  assign y3202 = 1'b0 ;
  assign y3203 = n6899 ;
  assign y3204 = ~1'b0 ;
  assign y3205 = ~1'b0 ;
  assign y3206 = ~1'b0 ;
  assign y3207 = ~1'b0 ;
  assign y3208 = n6900 ;
  assign y3209 = ~1'b0 ;
  assign y3210 = ~1'b0 ;
  assign y3211 = ~n6905 ;
  assign y3212 = ~1'b0 ;
  assign y3213 = n3757 ;
  assign y3214 = ~n6909 ;
  assign y3215 = n6913 ;
  assign y3216 = ~n2303 ;
  assign y3217 = n6914 ;
  assign y3218 = ~n6916 ;
  assign y3219 = ~1'b0 ;
  assign y3220 = ~n6921 ;
  assign y3221 = n6922 ;
  assign y3222 = ~n6923 ;
  assign y3223 = ~1'b0 ;
  assign y3224 = n6924 ;
  assign y3225 = ~1'b0 ;
  assign y3226 = ~n1295 ;
  assign y3227 = ~1'b0 ;
  assign y3228 = ~n6926 ;
  assign y3229 = 1'b0 ;
  assign y3230 = ~1'b0 ;
  assign y3231 = ~n6928 ;
  assign y3232 = n6933 ;
  assign y3233 = n6934 ;
  assign y3234 = n6936 ;
  assign y3235 = ~1'b0 ;
  assign y3236 = ~1'b0 ;
  assign y3237 = ~n6938 ;
  assign y3238 = ~n6940 ;
  assign y3239 = n6941 ;
  assign y3240 = ~n6944 ;
  assign y3241 = n6949 ;
  assign y3242 = ~1'b0 ;
  assign y3243 = ~n6951 ;
  assign y3244 = n6954 ;
  assign y3245 = ~1'b0 ;
  assign y3246 = n6956 ;
  assign y3247 = n2123 ;
  assign y3248 = ~n6961 ;
  assign y3249 = ~n6963 ;
  assign y3250 = ~n6964 ;
  assign y3251 = n6965 ;
  assign y3252 = n6966 ;
  assign y3253 = n6969 ;
  assign y3254 = ~n3824 ;
  assign y3255 = ~n6970 ;
  assign y3256 = ~1'b0 ;
  assign y3257 = ~1'b0 ;
  assign y3258 = n3606 ;
  assign y3259 = ~1'b0 ;
  assign y3260 = n6971 ;
  assign y3261 = ~n6972 ;
  assign y3262 = ~n2093 ;
  assign y3263 = ~n6973 ;
  assign y3264 = n6974 ;
  assign y3265 = ~n6975 ;
  assign y3266 = ~n6977 ;
  assign y3267 = ~1'b0 ;
  assign y3268 = 1'b0 ;
  assign y3269 = ~n713 ;
  assign y3270 = n6979 ;
  assign y3271 = n6984 ;
  assign y3272 = n6985 ;
  assign y3273 = ~1'b0 ;
  assign y3274 = n2484 ;
  assign y3275 = ~n6988 ;
  assign y3276 = n6989 ;
  assign y3277 = n6994 ;
  assign y3278 = 1'b0 ;
  assign y3279 = ~1'b0 ;
  assign y3280 = ~n6995 ;
  assign y3281 = n6996 ;
  assign y3282 = ~1'b0 ;
  assign y3283 = ~1'b0 ;
  assign y3284 = n6997 ;
  assign y3285 = ~n6998 ;
  assign y3286 = ~n7000 ;
  assign y3287 = ~n7001 ;
  assign y3288 = ~1'b0 ;
  assign y3289 = n7002 ;
  assign y3290 = ~n7006 ;
  assign y3291 = n7007 ;
  assign y3292 = ~1'b0 ;
  assign y3293 = ~n7008 ;
  assign y3294 = n7010 ;
  assign y3295 = n7011 ;
  assign y3296 = ~n7016 ;
  assign y3297 = ~n7024 ;
  assign y3298 = n7028 ;
  assign y3299 = ~1'b0 ;
  assign y3300 = ~n7030 ;
  assign y3301 = n7031 ;
  assign y3302 = ~n7037 ;
  assign y3303 = n7038 ;
  assign y3304 = ~1'b0 ;
  assign y3305 = ~n7039 ;
  assign y3306 = n7040 ;
  assign y3307 = ~1'b0 ;
  assign y3308 = ~1'b0 ;
  assign y3309 = ~n7041 ;
  assign y3310 = n7029 ;
  assign y3311 = ~n7047 ;
  assign y3312 = ~1'b0 ;
  assign y3313 = n7048 ;
  assign y3314 = ~n7050 ;
  assign y3315 = ~n7051 ;
  assign y3316 = n900 ;
  assign y3317 = n7054 ;
  assign y3318 = n7057 ;
  assign y3319 = ~n7066 ;
  assign y3320 = ~1'b0 ;
  assign y3321 = ~n7068 ;
  assign y3322 = ~1'b0 ;
  assign y3323 = n7071 ;
  assign y3324 = n7080 ;
  assign y3325 = ~1'b0 ;
  assign y3326 = ~n7086 ;
  assign y3327 = n7093 ;
  assign y3328 = n7096 ;
  assign y3329 = n7099 ;
  assign y3330 = ~n7100 ;
  assign y3331 = ~n7101 ;
  assign y3332 = ~1'b0 ;
  assign y3333 = ~1'b0 ;
  assign y3334 = ~n7102 ;
  assign y3335 = n7105 ;
  assign y3336 = ~1'b0 ;
  assign y3337 = ~n7108 ;
  assign y3338 = ~1'b0 ;
  assign y3339 = ~1'b0 ;
  assign y3340 = ~n7112 ;
  assign y3341 = 1'b0 ;
  assign y3342 = ~n7114 ;
  assign y3343 = n7116 ;
  assign y3344 = ~n7118 ;
  assign y3345 = ~n7119 ;
  assign y3346 = n7120 ;
  assign y3347 = ~1'b0 ;
  assign y3348 = ~1'b0 ;
  assign y3349 = ~1'b0 ;
  assign y3350 = ~1'b0 ;
  assign y3351 = ~n225 ;
  assign y3352 = ~n7121 ;
  assign y3353 = 1'b0 ;
  assign y3354 = ~1'b0 ;
  assign y3355 = n7131 ;
  assign y3356 = ~n7134 ;
  assign y3357 = n7143 ;
  assign y3358 = ~n7148 ;
  assign y3359 = n7150 ;
  assign y3360 = n7156 ;
  assign y3361 = n7158 ;
  assign y3362 = ~n7161 ;
  assign y3363 = ~n7167 ;
  assign y3364 = n7171 ;
  assign y3365 = ~n7177 ;
  assign y3366 = ~1'b0 ;
  assign y3367 = ~n7178 ;
  assign y3368 = n7185 ;
  assign y3369 = ~1'b0 ;
  assign y3370 = ~1'b0 ;
  assign y3371 = n5667 ;
  assign y3372 = n7189 ;
  assign y3373 = n7190 ;
  assign y3374 = n7191 ;
  assign y3375 = ~1'b0 ;
  assign y3376 = ~1'b0 ;
  assign y3377 = n2924 ;
  assign y3378 = n7192 ;
  assign y3379 = ~1'b0 ;
  assign y3380 = n7194 ;
  assign y3381 = ~n7195 ;
  assign y3382 = n7196 ;
  assign y3383 = ~n7157 ;
  assign y3384 = ~1'b0 ;
  assign y3385 = n7198 ;
  assign y3386 = ~1'b0 ;
  assign y3387 = ~1'b0 ;
  assign y3388 = ~1'b0 ;
  assign y3389 = n7204 ;
  assign y3390 = n7205 ;
  assign y3391 = ~n7206 ;
  assign y3392 = ~1'b0 ;
  assign y3393 = ~1'b0 ;
  assign y3394 = ~n7207 ;
  assign y3395 = ~n7216 ;
  assign y3396 = ~n7218 ;
  assign y3397 = ~n7220 ;
  assign y3398 = ~n7226 ;
  assign y3399 = ~n7229 ;
  assign y3400 = n7230 ;
  assign y3401 = n7233 ;
  assign y3402 = ~n7235 ;
  assign y3403 = n7236 ;
  assign y3404 = ~1'b0 ;
  assign y3405 = n7239 ;
  assign y3406 = ~1'b0 ;
  assign y3407 = ~1'b0 ;
  assign y3408 = ~n7242 ;
  assign y3409 = 1'b0 ;
  assign y3410 = ~n7243 ;
  assign y3411 = ~1'b0 ;
  assign y3412 = n7244 ;
  assign y3413 = ~n7245 ;
  assign y3414 = ~n7247 ;
  assign y3415 = ~n7248 ;
  assign y3416 = ~1'b0 ;
  assign y3417 = ~1'b0 ;
  assign y3418 = ~1'b0 ;
  assign y3419 = ~n7253 ;
  assign y3420 = ~1'b0 ;
  assign y3421 = 1'b0 ;
  assign y3422 = ~n7255 ;
  assign y3423 = ~n7260 ;
  assign y3424 = n7263 ;
  assign y3425 = n7273 ;
  assign y3426 = ~n7275 ;
  assign y3427 = ~1'b0 ;
  assign y3428 = ~1'b0 ;
  assign y3429 = ~1'b0 ;
  assign y3430 = ~1'b0 ;
  assign y3431 = n412 ;
  assign y3432 = ~n7282 ;
  assign y3433 = n643 ;
  assign y3434 = n7284 ;
  assign y3435 = ~1'b0 ;
  assign y3436 = n6049 ;
  assign y3437 = n7285 ;
  assign y3438 = n7295 ;
  assign y3439 = n7297 ;
  assign y3440 = ~1'b0 ;
  assign y3441 = ~1'b0 ;
  assign y3442 = ~1'b0 ;
  assign y3443 = 1'b0 ;
  assign y3444 = n7298 ;
  assign y3445 = ~n7299 ;
  assign y3446 = ~1'b0 ;
  assign y3447 = ~1'b0 ;
  assign y3448 = n7307 ;
  assign y3449 = ~n5203 ;
  assign y3450 = ~1'b0 ;
  assign y3451 = n7313 ;
  assign y3452 = n7315 ;
  assign y3453 = 1'b0 ;
  assign y3454 = n7316 ;
  assign y3455 = ~n7320 ;
  assign y3456 = ~1'b0 ;
  assign y3457 = ~n7322 ;
  assign y3458 = ~1'b0 ;
  assign y3459 = ~n7325 ;
  assign y3460 = ~n5996 ;
  assign y3461 = ~n7326 ;
  assign y3462 = n7328 ;
  assign y3463 = n7330 ;
  assign y3464 = ~n7331 ;
  assign y3465 = ~n7333 ;
  assign y3466 = n7338 ;
  assign y3467 = ~1'b0 ;
  assign y3468 = n7339 ;
  assign y3469 = ~1'b0 ;
  assign y3470 = n7341 ;
  assign y3471 = ~1'b0 ;
  assign y3472 = n709 ;
  assign y3473 = n7344 ;
  assign y3474 = 1'b0 ;
  assign y3475 = ~n7346 ;
  assign y3476 = ~1'b0 ;
  assign y3477 = ~n7351 ;
  assign y3478 = n7354 ;
  assign y3479 = n7359 ;
  assign y3480 = ~n7362 ;
  assign y3481 = ~n7364 ;
  assign y3482 = ~1'b0 ;
  assign y3483 = 1'b0 ;
  assign y3484 = ~1'b0 ;
  assign y3485 = ~n7366 ;
  assign y3486 = ~1'b0 ;
  assign y3487 = ~n7367 ;
  assign y3488 = n7368 ;
  assign y3489 = ~1'b0 ;
  assign y3490 = n7373 ;
  assign y3491 = ~n7376 ;
  assign y3492 = n7378 ;
  assign y3493 = ~1'b0 ;
  assign y3494 = ~n7381 ;
  assign y3495 = ~n7382 ;
  assign y3496 = ~1'b0 ;
  assign y3497 = ~n7394 ;
  assign y3498 = ~n795 ;
  assign y3499 = ~n7396 ;
  assign y3500 = n7401 ;
  assign y3501 = ~1'b0 ;
  assign y3502 = ~n5915 ;
  assign y3503 = n7403 ;
  assign y3504 = ~1'b0 ;
  assign y3505 = ~n7406 ;
  assign y3506 = ~1'b0 ;
  assign y3507 = ~n4727 ;
  assign y3508 = n7410 ;
  assign y3509 = ~n7412 ;
  assign y3510 = ~n7415 ;
  assign y3511 = n7423 ;
  assign y3512 = ~1'b0 ;
  assign y3513 = n7424 ;
  assign y3514 = ~1'b0 ;
  assign y3515 = ~n7430 ;
  assign y3516 = 1'b0 ;
  assign y3517 = ~n7431 ;
  assign y3518 = ~n7434 ;
  assign y3519 = n1157 ;
  assign y3520 = ~1'b0 ;
  assign y3521 = ~1'b0 ;
  assign y3522 = ~n7439 ;
  assign y3523 = ~1'b0 ;
  assign y3524 = ~1'b0 ;
  assign y3525 = ~n3680 ;
  assign y3526 = ~1'b0 ;
  assign y3527 = n7441 ;
  assign y3528 = ~1'b0 ;
  assign y3529 = ~n7444 ;
  assign y3530 = n7446 ;
  assign y3531 = n7447 ;
  assign y3532 = n7450 ;
  assign y3533 = n7451 ;
  assign y3534 = ~n7455 ;
  assign y3535 = n7459 ;
  assign y3536 = ~1'b0 ;
  assign y3537 = ~n7461 ;
  assign y3538 = ~1'b0 ;
  assign y3539 = n7468 ;
  assign y3540 = n7469 ;
  assign y3541 = ~n7473 ;
  assign y3542 = ~n7476 ;
  assign y3543 = ~1'b0 ;
  assign y3544 = n7478 ;
  assign y3545 = n2603 ;
  assign y3546 = ~n7479 ;
  assign y3547 = ~n7485 ;
  assign y3548 = ~n7486 ;
  assign y3549 = n7492 ;
  assign y3550 = ~1'b0 ;
  assign y3551 = n7495 ;
  assign y3552 = n7496 ;
  assign y3553 = n7498 ;
  assign y3554 = ~1'b0 ;
  assign y3555 = n7500 ;
  assign y3556 = ~1'b0 ;
  assign y3557 = ~n3193 ;
  assign y3558 = n7501 ;
  assign y3559 = ~n7505 ;
  assign y3560 = n7511 ;
  assign y3561 = ~1'b0 ;
  assign y3562 = ~1'b0 ;
  assign y3563 = n7513 ;
  assign y3564 = ~n7516 ;
  assign y3565 = ~n7526 ;
  assign y3566 = 1'b0 ;
  assign y3567 = ~n7528 ;
  assign y3568 = 1'b0 ;
  assign y3569 = n1295 ;
  assign y3570 = ~1'b0 ;
  assign y3571 = ~1'b0 ;
  assign y3572 = ~1'b0 ;
  assign y3573 = ~1'b0 ;
  assign y3574 = n7529 ;
  assign y3575 = n7535 ;
  assign y3576 = ~1'b0 ;
  assign y3577 = ~1'b0 ;
  assign y3578 = n7540 ;
  assign y3579 = n901 ;
  assign y3580 = ~n7543 ;
  assign y3581 = n7546 ;
  assign y3582 = n7548 ;
  assign y3583 = n7549 ;
  assign y3584 = 1'b0 ;
  assign y3585 = ~n7554 ;
  assign y3586 = n7557 ;
  assign y3587 = ~1'b0 ;
  assign y3588 = n7143 ;
  assign y3589 = ~n7559 ;
  assign y3590 = n7566 ;
  assign y3591 = ~1'b0 ;
  assign y3592 = n7569 ;
  assign y3593 = ~n7570 ;
  assign y3594 = n7574 ;
  assign y3595 = ~n7582 ;
  assign y3596 = n7585 ;
  assign y3597 = ~n7586 ;
  assign y3598 = 1'b0 ;
  assign y3599 = ~n3015 ;
  assign y3600 = n7587 ;
  assign y3601 = n7592 ;
  assign y3602 = ~n7594 ;
  assign y3603 = n7603 ;
  assign y3604 = ~n7604 ;
  assign y3605 = ~1'b0 ;
  assign y3606 = n7610 ;
  assign y3607 = ~1'b0 ;
  assign y3608 = n7612 ;
  assign y3609 = ~1'b0 ;
  assign y3610 = ~n7614 ;
  assign y3611 = ~1'b0 ;
  assign y3612 = ~n7615 ;
  assign y3613 = ~1'b0 ;
  assign y3614 = ~1'b0 ;
  assign y3615 = ~n7617 ;
  assign y3616 = n7622 ;
  assign y3617 = n7623 ;
  assign y3618 = ~1'b0 ;
  assign y3619 = ~1'b0 ;
  assign y3620 = ~n7624 ;
  assign y3621 = n7625 ;
  assign y3622 = ~n2130 ;
  assign y3623 = n7627 ;
  assign y3624 = ~n7639 ;
  assign y3625 = n7641 ;
  assign y3626 = ~1'b0 ;
  assign y3627 = n7643 ;
  assign y3628 = ~n7645 ;
  assign y3629 = ~1'b0 ;
  assign y3630 = ~n7649 ;
  assign y3631 = ~1'b0 ;
  assign y3632 = ~n7650 ;
  assign y3633 = ~1'b0 ;
  assign y3634 = n141 ;
  assign y3635 = ~n7653 ;
  assign y3636 = n7655 ;
  assign y3637 = ~1'b0 ;
  assign y3638 = ~n7656 ;
  assign y3639 = ~1'b0 ;
  assign y3640 = ~1'b0 ;
  assign y3641 = ~n7658 ;
  assign y3642 = ~n7661 ;
  assign y3643 = ~n7664 ;
  assign y3644 = ~n7665 ;
  assign y3645 = ~1'b0 ;
  assign y3646 = ~1'b0 ;
  assign y3647 = n7671 ;
  assign y3648 = n7677 ;
  assign y3649 = ~n7680 ;
  assign y3650 = n7682 ;
  assign y3651 = ~n7684 ;
  assign y3652 = ~1'b0 ;
  assign y3653 = ~n7685 ;
  assign y3654 = ~n7693 ;
  assign y3655 = ~1'b0 ;
  assign y3656 = ~1'b0 ;
  assign y3657 = ~1'b0 ;
  assign y3658 = ~1'b0 ;
  assign y3659 = ~n7698 ;
  assign y3660 = n479 ;
  assign y3661 = ~n7699 ;
  assign y3662 = n7703 ;
  assign y3663 = ~n7705 ;
  assign y3664 = ~n583 ;
  assign y3665 = ~1'b0 ;
  assign y3666 = ~1'b0 ;
  assign y3667 = n7706 ;
  assign y3668 = ~1'b0 ;
  assign y3669 = n3109 ;
  assign y3670 = ~1'b0 ;
  assign y3671 = ~n7707 ;
  assign y3672 = ~1'b0 ;
  assign y3673 = ~1'b0 ;
  assign y3674 = ~1'b0 ;
  assign y3675 = n7708 ;
  assign y3676 = ~1'b0 ;
  assign y3677 = n3641 ;
  assign y3678 = n7712 ;
  assign y3679 = ~n7715 ;
  assign y3680 = ~n297 ;
  assign y3681 = ~n7716 ;
  assign y3682 = ~n7718 ;
  assign y3683 = ~n7719 ;
  assign y3684 = ~n7720 ;
  assign y3685 = ~n7723 ;
  assign y3686 = n7727 ;
  assign y3687 = ~n7731 ;
  assign y3688 = ~n7732 ;
  assign y3689 = ~1'b0 ;
  assign y3690 = n7737 ;
  assign y3691 = ~1'b0 ;
  assign y3692 = n7738 ;
  assign y3693 = ~n7742 ;
  assign y3694 = n7749 ;
  assign y3695 = ~n7757 ;
  assign y3696 = n7761 ;
  assign y3697 = 1'b0 ;
  assign y3698 = ~1'b0 ;
  assign y3699 = ~1'b0 ;
  assign y3700 = ~n7762 ;
  assign y3701 = n7766 ;
  assign y3702 = n7773 ;
  assign y3703 = n7774 ;
  assign y3704 = ~1'b0 ;
  assign y3705 = n7777 ;
  assign y3706 = ~1'b0 ;
  assign y3707 = n3365 ;
  assign y3708 = ~n7778 ;
  assign y3709 = ~n7779 ;
  assign y3710 = ~1'b0 ;
  assign y3711 = ~n7780 ;
  assign y3712 = ~n7783 ;
  assign y3713 = n7784 ;
  assign y3714 = ~1'b0 ;
  assign y3715 = ~1'b0 ;
  assign y3716 = ~n7787 ;
  assign y3717 = n7791 ;
  assign y3718 = n7799 ;
  assign y3719 = n7801 ;
  assign y3720 = 1'b0 ;
  assign y3721 = ~n7804 ;
  assign y3722 = ~1'b0 ;
  assign y3723 = ~n7811 ;
  assign y3724 = ~n7818 ;
  assign y3725 = ~n7821 ;
  assign y3726 = ~1'b0 ;
  assign y3727 = n3991 ;
  assign y3728 = 1'b0 ;
  assign y3729 = n7824 ;
  assign y3730 = 1'b0 ;
  assign y3731 = n7830 ;
  assign y3732 = ~n7831 ;
  assign y3733 = ~n7834 ;
  assign y3734 = ~1'b0 ;
  assign y3735 = ~1'b0 ;
  assign y3736 = n7837 ;
  assign y3737 = n7838 ;
  assign y3738 = n2559 ;
  assign y3739 = ~n7840 ;
  assign y3740 = ~1'b0 ;
  assign y3741 = ~1'b0 ;
  assign y3742 = n7842 ;
  assign y3743 = ~n3993 ;
  assign y3744 = n7847 ;
  assign y3745 = ~n7849 ;
  assign y3746 = ~1'b0 ;
  assign y3747 = ~n7851 ;
  assign y3748 = ~n7854 ;
  assign y3749 = n7855 ;
  assign y3750 = ~1'b0 ;
  assign y3751 = 1'b0 ;
  assign y3752 = n7857 ;
  assign y3753 = n7858 ;
  assign y3754 = ~n7860 ;
  assign y3755 = ~n7867 ;
  assign y3756 = n7869 ;
  assign y3757 = ~1'b0 ;
  assign y3758 = ~1'b0 ;
  assign y3759 = ~1'b0 ;
  assign y3760 = n2819 ;
  assign y3761 = ~1'b0 ;
  assign y3762 = n7874 ;
  assign y3763 = ~1'b0 ;
  assign y3764 = ~n7876 ;
  assign y3765 = ~1'b0 ;
  assign y3766 = ~1'b0 ;
  assign y3767 = ~n7879 ;
  assign y3768 = ~n7884 ;
  assign y3769 = ~n7888 ;
  assign y3770 = ~n7890 ;
  assign y3771 = n7891 ;
  assign y3772 = ~n7894 ;
  assign y3773 = n3015 ;
  assign y3774 = ~n7898 ;
  assign y3775 = ~n7900 ;
  assign y3776 = ~n7902 ;
  assign y3777 = n2412 ;
  assign y3778 = ~n7905 ;
  assign y3779 = n7906 ;
  assign y3780 = ~1'b0 ;
  assign y3781 = ~n7918 ;
  assign y3782 = ~1'b0 ;
  assign y3783 = ~n7923 ;
  assign y3784 = n7929 ;
  assign y3785 = ~n7931 ;
  assign y3786 = ~1'b0 ;
  assign y3787 = ~n7936 ;
  assign y3788 = ~1'b0 ;
  assign y3789 = ~n956 ;
  assign y3790 = ~n7939 ;
  assign y3791 = ~n7940 ;
  assign y3792 = n7948 ;
  assign y3793 = n7951 ;
  assign y3794 = n7954 ;
  assign y3795 = ~n7956 ;
  assign y3796 = 1'b0 ;
  assign y3797 = ~n7957 ;
  assign y3798 = n7958 ;
  assign y3799 = ~n7959 ;
  assign y3800 = n7961 ;
  assign y3801 = ~n7963 ;
  assign y3802 = ~1'b0 ;
  assign y3803 = ~n7964 ;
  assign y3804 = ~1'b0 ;
  assign y3805 = ~1'b0 ;
  assign y3806 = ~n7966 ;
  assign y3807 = ~1'b0 ;
  assign y3808 = n7967 ;
  assign y3809 = ~1'b0 ;
  assign y3810 = n7970 ;
  assign y3811 = ~1'b0 ;
  assign y3812 = ~n7972 ;
  assign y3813 = ~n7974 ;
  assign y3814 = n7982 ;
  assign y3815 = n7988 ;
  assign y3816 = ~1'b0 ;
  assign y3817 = ~1'b0 ;
  assign y3818 = ~n7995 ;
  assign y3819 = ~n7997 ;
  assign y3820 = n8003 ;
  assign y3821 = ~1'b0 ;
  assign y3822 = 1'b0 ;
  assign y3823 = ~n8006 ;
  assign y3824 = ~1'b0 ;
  assign y3825 = ~1'b0 ;
  assign y3826 = ~n8007 ;
  assign y3827 = n8009 ;
  assign y3828 = ~1'b0 ;
  assign y3829 = ~1'b0 ;
  assign y3830 = n8012 ;
  assign y3831 = n8013 ;
  assign y3832 = ~1'b0 ;
  assign y3833 = ~1'b0 ;
  assign y3834 = ~1'b0 ;
  assign y3835 = n8015 ;
  assign y3836 = ~n8021 ;
  assign y3837 = ~n8025 ;
  assign y3838 = ~n8026 ;
  assign y3839 = ~n8029 ;
  assign y3840 = ~1'b0 ;
  assign y3841 = n8030 ;
  assign y3842 = ~n8031 ;
  assign y3843 = ~n8035 ;
  assign y3844 = 1'b0 ;
  assign y3845 = n2654 ;
  assign y3846 = n8038 ;
  assign y3847 = n8040 ;
  assign y3848 = n8041 ;
  assign y3849 = ~1'b0 ;
  assign y3850 = n8053 ;
  assign y3851 = ~n8054 ;
  assign y3852 = ~1'b0 ;
  assign y3853 = ~1'b0 ;
  assign y3854 = n8056 ;
  assign y3855 = n8063 ;
  assign y3856 = ~1'b0 ;
  assign y3857 = ~1'b0 ;
  assign y3858 = n8065 ;
  assign y3859 = ~n8068 ;
  assign y3860 = n8070 ;
  assign y3861 = ~n8071 ;
  assign y3862 = n8075 ;
  assign y3863 = ~1'b0 ;
  assign y3864 = ~1'b0 ;
  assign y3865 = ~1'b0 ;
  assign y3866 = n8077 ;
  assign y3867 = ~1'b0 ;
  assign y3868 = ~1'b0 ;
  assign y3869 = n8078 ;
  assign y3870 = ~1'b0 ;
  assign y3871 = ~n8081 ;
  assign y3872 = ~1'b0 ;
  assign y3873 = n8083 ;
  assign y3874 = ~n8089 ;
  assign y3875 = ~1'b0 ;
  assign y3876 = ~n8090 ;
  assign y3877 = ~1'b0 ;
  assign y3878 = n8094 ;
  assign y3879 = n8098 ;
  assign y3880 = n8100 ;
  assign y3881 = n8101 ;
  assign y3882 = ~1'b0 ;
  assign y3883 = ~n8104 ;
  assign y3884 = n4036 ;
  assign y3885 = ~n8107 ;
  assign y3886 = n8111 ;
  assign y3887 = n8113 ;
  assign y3888 = ~n8114 ;
  assign y3889 = ~n8118 ;
  assign y3890 = ~n8119 ;
  assign y3891 = ~1'b0 ;
  assign y3892 = ~1'b0 ;
  assign y3893 = n8122 ;
  assign y3894 = ~n8123 ;
  assign y3895 = n8127 ;
  assign y3896 = ~n8128 ;
  assign y3897 = ~1'b0 ;
  assign y3898 = ~n8131 ;
  assign y3899 = ~1'b0 ;
  assign y3900 = ~n8134 ;
  assign y3901 = n8139 ;
  assign y3902 = n8140 ;
  assign y3903 = n8142 ;
  assign y3904 = ~1'b0 ;
  assign y3905 = ~n8147 ;
  assign y3906 = ~1'b0 ;
  assign y3907 = ~1'b0 ;
  assign y3908 = n8148 ;
  assign y3909 = n8149 ;
  assign y3910 = ~n8153 ;
  assign y3911 = ~1'b0 ;
  assign y3912 = n8156 ;
  assign y3913 = ~n8162 ;
  assign y3914 = ~1'b0 ;
  assign y3915 = ~1'b0 ;
  assign y3916 = ~n8167 ;
  assign y3917 = n8171 ;
  assign y3918 = ~n8174 ;
  assign y3919 = ~n8177 ;
  assign y3920 = ~n8181 ;
  assign y3921 = ~1'b0 ;
  assign y3922 = n8184 ;
  assign y3923 = n8187 ;
  assign y3924 = ~n8197 ;
  assign y3925 = n8198 ;
  assign y3926 = ~1'b0 ;
  assign y3927 = ~n8199 ;
  assign y3928 = ~1'b0 ;
  assign y3929 = ~1'b0 ;
  assign y3930 = ~n8201 ;
  assign y3931 = n8203 ;
  assign y3932 = ~n6385 ;
  assign y3933 = ~n8204 ;
  assign y3934 = ~n8206 ;
  assign y3935 = ~n8208 ;
  assign y3936 = n5297 ;
  assign y3937 = ~1'b0 ;
  assign y3938 = ~1'b0 ;
  assign y3939 = ~n8209 ;
  assign y3940 = n8215 ;
  assign y3941 = ~1'b0 ;
  assign y3942 = ~n8217 ;
  assign y3943 = n4782 ;
  assign y3944 = n8219 ;
  assign y3945 = n8220 ;
  assign y3946 = n4723 ;
  assign y3947 = ~n8221 ;
  assign y3948 = ~1'b0 ;
  assign y3949 = ~n8223 ;
  assign y3950 = n6201 ;
  assign y3951 = ~n8229 ;
  assign y3952 = ~1'b0 ;
  assign y3953 = n1687 ;
  assign y3954 = ~n8231 ;
  assign y3955 = n8235 ;
  assign y3956 = ~n8239 ;
  assign y3957 = ~1'b0 ;
  assign y3958 = ~1'b0 ;
  assign y3959 = n7096 ;
  assign y3960 = n8240 ;
  assign y3961 = ~n8243 ;
  assign y3962 = ~1'b0 ;
  assign y3963 = n8245 ;
  assign y3964 = ~1'b0 ;
  assign y3965 = ~1'b0 ;
  assign y3966 = ~n8246 ;
  assign y3967 = ~n8251 ;
  assign y3968 = ~n8255 ;
  assign y3969 = ~n8265 ;
  assign y3970 = n2998 ;
  assign y3971 = ~n8271 ;
  assign y3972 = ~1'b0 ;
  assign y3973 = n8273 ;
  assign y3974 = ~n8278 ;
  assign y3975 = n8285 ;
  assign y3976 = n8287 ;
  assign y3977 = ~n8290 ;
  assign y3978 = ~n8293 ;
  assign y3979 = n8294 ;
  assign y3980 = n8297 ;
  assign y3981 = ~1'b0 ;
  assign y3982 = ~1'b0 ;
  assign y3983 = 1'b0 ;
  assign y3984 = ~1'b0 ;
  assign y3985 = ~n8298 ;
  assign y3986 = ~n8301 ;
  assign y3987 = ~1'b0 ;
  assign y3988 = ~n3961 ;
  assign y3989 = ~n8303 ;
  assign y3990 = n8310 ;
  assign y3991 = n8312 ;
  assign y3992 = ~n8317 ;
  assign y3993 = n4063 ;
  assign y3994 = n2414 ;
  assign y3995 = ~n8319 ;
  assign y3996 = n8321 ;
  assign y3997 = ~n8323 ;
  assign y3998 = ~1'b0 ;
  assign y3999 = ~n8325 ;
  assign y4000 = ~1'b0 ;
  assign y4001 = n8327 ;
  assign y4002 = ~n7779 ;
  assign y4003 = n8328 ;
  assign y4004 = n8330 ;
  assign y4005 = ~n8331 ;
  assign y4006 = ~n6655 ;
  assign y4007 = n8333 ;
  assign y4008 = ~n8337 ;
  assign y4009 = ~1'b0 ;
  assign y4010 = ~n7521 ;
  assign y4011 = ~1'b0 ;
  assign y4012 = n8346 ;
  assign y4013 = ~n8351 ;
  assign y4014 = n6159 ;
  assign y4015 = n8352 ;
  assign y4016 = ~n8353 ;
  assign y4017 = ~n8355 ;
  assign y4018 = n8357 ;
  assign y4019 = n8358 ;
  assign y4020 = ~1'b0 ;
  assign y4021 = ~1'b0 ;
  assign y4022 = ~n6759 ;
  assign y4023 = ~1'b0 ;
  assign y4024 = ~n8362 ;
  assign y4025 = ~n8365 ;
  assign y4026 = ~n8376 ;
  assign y4027 = ~n8381 ;
  assign y4028 = ~n8384 ;
  assign y4029 = ~n8388 ;
  assign y4030 = n8397 ;
  assign y4031 = n666 ;
  assign y4032 = n8404 ;
  assign y4033 = ~n8265 ;
  assign y4034 = ~n8405 ;
  assign y4035 = ~1'b0 ;
  assign y4036 = n8407 ;
  assign y4037 = n8411 ;
  assign y4038 = n8412 ;
  assign y4039 = n8414 ;
  assign y4040 = ~n8416 ;
  assign y4041 = ~n1212 ;
  assign y4042 = ~1'b0 ;
  assign y4043 = ~n8418 ;
  assign y4044 = ~1'b0 ;
  assign y4045 = ~1'b0 ;
  assign y4046 = n8420 ;
  assign y4047 = ~1'b0 ;
  assign y4048 = ~n8424 ;
  assign y4049 = ~1'b0 ;
  assign y4050 = ~1'b0 ;
  assign y4051 = ~1'b0 ;
  assign y4052 = ~1'b0 ;
  assign y4053 = n8425 ;
  assign y4054 = n8427 ;
  assign y4055 = n8432 ;
  assign y4056 = ~1'b0 ;
  assign y4057 = ~1'b0 ;
  assign y4058 = n8435 ;
  assign y4059 = ~n8437 ;
  assign y4060 = ~1'b0 ;
  assign y4061 = n7185 ;
  assign y4062 = ~n8442 ;
  assign y4063 = ~n8445 ;
  assign y4064 = ~n8446 ;
  assign y4065 = ~1'b0 ;
  assign y4066 = ~1'b0 ;
  assign y4067 = ~n3159 ;
  assign y4068 = n8448 ;
  assign y4069 = ~1'b0 ;
  assign y4070 = ~1'b0 ;
  assign y4071 = ~1'b0 ;
  assign y4072 = 1'b0 ;
  assign y4073 = ~n8451 ;
  assign y4074 = ~n8456 ;
  assign y4075 = n8458 ;
  assign y4076 = ~n8466 ;
  assign y4077 = n8468 ;
  assign y4078 = 1'b0 ;
  assign y4079 = n8469 ;
  assign y4080 = n8471 ;
  assign y4081 = ~1'b0 ;
  assign y4082 = ~n8472 ;
  assign y4083 = n900 ;
  assign y4084 = ~1'b0 ;
  assign y4085 = ~n8481 ;
  assign y4086 = ~n8482 ;
  assign y4087 = ~1'b0 ;
  assign y4088 = ~1'b0 ;
  assign y4089 = n8483 ;
  assign y4090 = ~n8486 ;
  assign y4091 = ~n8487 ;
  assign y4092 = ~1'b0 ;
  assign y4093 = ~n8489 ;
  assign y4094 = ~n8490 ;
  assign y4095 = ~n8491 ;
  assign y4096 = ~1'b0 ;
  assign y4097 = ~n8495 ;
  assign y4098 = 1'b0 ;
  assign y4099 = n8498 ;
  assign y4100 = ~n7368 ;
  assign y4101 = ~n8499 ;
  assign y4102 = n8501 ;
  assign y4103 = ~n8503 ;
  assign y4104 = ~1'b0 ;
  assign y4105 = 1'b0 ;
  assign y4106 = ~n8506 ;
  assign y4107 = n8510 ;
  assign y4108 = ~1'b0 ;
  assign y4109 = ~n2235 ;
  assign y4110 = n8512 ;
  assign y4111 = n8513 ;
  assign y4112 = n8514 ;
  assign y4113 = ~n8518 ;
  assign y4114 = ~1'b0 ;
  assign y4115 = ~1'b0 ;
  assign y4116 = ~1'b0 ;
  assign y4117 = n8521 ;
  assign y4118 = n8522 ;
  assign y4119 = ~1'b0 ;
  assign y4120 = ~1'b0 ;
  assign y4121 = n8524 ;
  assign y4122 = n8525 ;
  assign y4123 = ~n8531 ;
  assign y4124 = ~1'b0 ;
  assign y4125 = ~n8537 ;
  assign y4126 = ~n8539 ;
  assign y4127 = ~1'b0 ;
  assign y4128 = ~n8548 ;
  assign y4129 = ~n8550 ;
  assign y4130 = n8552 ;
  assign y4131 = n8554 ;
  assign y4132 = ~1'b0 ;
  assign y4133 = ~n8556 ;
  assign y4134 = ~n8561 ;
  assign y4135 = ~1'b0 ;
  assign y4136 = ~1'b0 ;
  assign y4137 = n8562 ;
  assign y4138 = ~1'b0 ;
  assign y4139 = n8566 ;
  assign y4140 = ~1'b0 ;
  assign y4141 = ~n8567 ;
  assign y4142 = ~n8568 ;
  assign y4143 = ~n8571 ;
  assign y4144 = n8581 ;
  assign y4145 = n8582 ;
  assign y4146 = ~1'b0 ;
  assign y4147 = ~n8584 ;
  assign y4148 = n3738 ;
  assign y4149 = n8585 ;
  assign y4150 = ~n8587 ;
  assign y4151 = ~n8592 ;
  assign y4152 = n8593 ;
  assign y4153 = n8594 ;
  assign y4154 = n8598 ;
  assign y4155 = n742 ;
  assign y4156 = n8602 ;
  assign y4157 = ~n8605 ;
  assign y4158 = n8611 ;
  assign y4159 = ~1'b0 ;
  assign y4160 = ~n8615 ;
  assign y4161 = n8625 ;
  assign y4162 = ~n8627 ;
  assign y4163 = n8628 ;
  assign y4164 = ~1'b0 ;
  assign y4165 = n8632 ;
  assign y4166 = n8633 ;
  assign y4167 = 1'b0 ;
  assign y4168 = n8637 ;
  assign y4169 = n8638 ;
  assign y4170 = ~n4588 ;
  assign y4171 = n3003 ;
  assign y4172 = n8639 ;
  assign y4173 = ~1'b0 ;
  assign y4174 = ~1'b0 ;
  assign y4175 = ~1'b0 ;
  assign y4176 = ~1'b0 ;
  assign y4177 = ~1'b0 ;
  assign y4178 = ~n8644 ;
  assign y4179 = ~1'b0 ;
  assign y4180 = ~1'b0 ;
  assign y4181 = ~1'b0 ;
  assign y4182 = n8646 ;
  assign y4183 = ~n8648 ;
  assign y4184 = ~n8651 ;
  assign y4185 = n8657 ;
  assign y4186 = ~1'b0 ;
  assign y4187 = ~n8659 ;
  assign y4188 = ~1'b0 ;
  assign y4189 = n8664 ;
  assign y4190 = n8666 ;
  assign y4191 = ~n8668 ;
  assign y4192 = ~n8669 ;
  assign y4193 = n8674 ;
  assign y4194 = ~1'b0 ;
  assign y4195 = ~1'b0 ;
  assign y4196 = ~n8676 ;
  assign y4197 = ~n8680 ;
  assign y4198 = n8682 ;
  assign y4199 = n8686 ;
  assign y4200 = ~n8688 ;
  assign y4201 = n8697 ;
  assign y4202 = n8700 ;
  assign y4203 = n8702 ;
  assign y4204 = n8705 ;
  assign y4205 = ~n586 ;
  assign y4206 = n8709 ;
  assign y4207 = ~n8711 ;
  assign y4208 = n8716 ;
  assign y4209 = n8725 ;
  assign y4210 = n8726 ;
  assign y4211 = ~1'b0 ;
  assign y4212 = ~n8728 ;
  assign y4213 = ~1'b0 ;
  assign y4214 = ~n8735 ;
  assign y4215 = n8737 ;
  assign y4216 = n8739 ;
  assign y4217 = ~1'b0 ;
  assign y4218 = ~1'b0 ;
  assign y4219 = ~n8741 ;
  assign y4220 = ~n8742 ;
  assign y4221 = ~1'b0 ;
  assign y4222 = ~n8744 ;
  assign y4223 = n8747 ;
  assign y4224 = n8750 ;
  assign y4225 = ~1'b0 ;
  assign y4226 = n8753 ;
  assign y4227 = n8756 ;
  assign y4228 = n2222 ;
  assign y4229 = ~n8758 ;
  assign y4230 = ~1'b0 ;
  assign y4231 = n8766 ;
  assign y4232 = ~n8767 ;
  assign y4233 = ~1'b0 ;
  assign y4234 = ~1'b0 ;
  assign y4235 = ~1'b0 ;
  assign y4236 = ~n8773 ;
  assign y4237 = ~1'b0 ;
  assign y4238 = n8776 ;
  assign y4239 = ~n8781 ;
  assign y4240 = 1'b0 ;
  assign y4241 = ~n8787 ;
  assign y4242 = ~1'b0 ;
  assign y4243 = n8788 ;
  assign y4244 = ~1'b0 ;
  assign y4245 = n8789 ;
  assign y4246 = ~1'b0 ;
  assign y4247 = n8794 ;
  assign y4248 = ~1'b0 ;
  assign y4249 = n8795 ;
  assign y4250 = n8802 ;
  assign y4251 = ~1'b0 ;
  assign y4252 = ~1'b0 ;
  assign y4253 = ~n8803 ;
  assign y4254 = n8805 ;
  assign y4255 = n8807 ;
  assign y4256 = ~n8808 ;
  assign y4257 = 1'b0 ;
  assign y4258 = n339 ;
  assign y4259 = ~n8809 ;
  assign y4260 = ~n8812 ;
  assign y4261 = ~n8813 ;
  assign y4262 = n8814 ;
  assign y4263 = ~1'b0 ;
  assign y4264 = n8815 ;
  assign y4265 = ~n8820 ;
  assign y4266 = ~1'b0 ;
  assign y4267 = ~n8821 ;
  assign y4268 = ~n8824 ;
  assign y4269 = ~1'b0 ;
  assign y4270 = ~1'b0 ;
  assign y4271 = n8828 ;
  assign y4272 = n8832 ;
  assign y4273 = ~1'b0 ;
  assign y4274 = ~1'b0 ;
  assign y4275 = ~1'b0 ;
  assign y4276 = ~1'b0 ;
  assign y4277 = ~1'b0 ;
  assign y4278 = ~n8835 ;
  assign y4279 = n8836 ;
  assign y4280 = ~n5662 ;
  assign y4281 = n8837 ;
  assign y4282 = ~1'b0 ;
  assign y4283 = n8842 ;
  assign y4284 = n8843 ;
  assign y4285 = n8848 ;
  assign y4286 = n8849 ;
  assign y4287 = n4817 ;
  assign y4288 = ~n8852 ;
  assign y4289 = ~n8856 ;
  assign y4290 = ~n8859 ;
  assign y4291 = ~1'b0 ;
  assign y4292 = n7649 ;
  assign y4293 = n8860 ;
  assign y4294 = n8865 ;
  assign y4295 = ~1'b0 ;
  assign y4296 = ~n8866 ;
  assign y4297 = n8867 ;
  assign y4298 = n8874 ;
  assign y4299 = ~n8876 ;
  assign y4300 = n8877 ;
  assign y4301 = n8883 ;
  assign y4302 = ~1'b0 ;
  assign y4303 = n8885 ;
  assign y4304 = n1511 ;
  assign y4305 = ~n8886 ;
  assign y4306 = ~n8887 ;
  assign y4307 = n8888 ;
  assign y4308 = n8889 ;
  assign y4309 = n8890 ;
  assign y4310 = ~1'b0 ;
  assign y4311 = n8893 ;
  assign y4312 = ~1'b0 ;
  assign y4313 = n8895 ;
  assign y4314 = ~n8897 ;
  assign y4315 = ~1'b0 ;
  assign y4316 = ~n8898 ;
  assign y4317 = n8902 ;
  assign y4318 = ~1'b0 ;
  assign y4319 = ~n8906 ;
  assign y4320 = ~1'b0 ;
  assign y4321 = 1'b0 ;
  assign y4322 = ~1'b0 ;
  assign y4323 = ~n8909 ;
  assign y4324 = ~1'b0 ;
  assign y4325 = ~1'b0 ;
  assign y4326 = n3761 ;
  assign y4327 = ~n8915 ;
  assign y4328 = n8916 ;
  assign y4329 = n8919 ;
  assign y4330 = n8926 ;
  assign y4331 = ~n8928 ;
  assign y4332 = ~n8929 ;
  assign y4333 = ~n8931 ;
  assign y4334 = n8932 ;
  assign y4335 = ~n8934 ;
  assign y4336 = n5038 ;
  assign y4337 = ~n8938 ;
  assign y4338 = ~n8940 ;
  assign y4339 = ~1'b0 ;
  assign y4340 = ~n8945 ;
  assign y4341 = ~n1383 ;
  assign y4342 = ~n8950 ;
  assign y4343 = ~n8951 ;
  assign y4344 = ~n8952 ;
  assign y4345 = ~n6932 ;
  assign y4346 = ~1'b0 ;
  assign y4347 = ~n8956 ;
  assign y4348 = ~n8958 ;
  assign y4349 = ~n8960 ;
  assign y4350 = ~1'b0 ;
  assign y4351 = n6561 ;
  assign y4352 = ~n8964 ;
  assign y4353 = n903 ;
  assign y4354 = ~1'b0 ;
  assign y4355 = n8968 ;
  assign y4356 = n8969 ;
  assign y4357 = ~1'b0 ;
  assign y4358 = n8970 ;
  assign y4359 = ~n1588 ;
  assign y4360 = ~n8971 ;
  assign y4361 = ~n7043 ;
  assign y4362 = ~1'b0 ;
  assign y4363 = ~1'b0 ;
  assign y4364 = ~n8978 ;
  assign y4365 = ~n8979 ;
  assign y4366 = ~1'b0 ;
  assign y4367 = ~1'b0 ;
  assign y4368 = n8984 ;
  assign y4369 = ~n8985 ;
  assign y4370 = n7854 ;
  assign y4371 = ~1'b0 ;
  assign y4372 = n8988 ;
  assign y4373 = ~1'b0 ;
  assign y4374 = n8991 ;
  assign y4375 = ~n8992 ;
  assign y4376 = ~1'b0 ;
  assign y4377 = ~n5102 ;
  assign y4378 = ~n1992 ;
  assign y4379 = n8995 ;
  assign y4380 = n9001 ;
  assign y4381 = n9004 ;
  assign y4382 = ~1'b0 ;
  assign y4383 = ~n9005 ;
  assign y4384 = n9006 ;
  assign y4385 = n9012 ;
  assign y4386 = n9016 ;
  assign y4387 = ~1'b0 ;
  assign y4388 = n9017 ;
  assign y4389 = ~n9019 ;
  assign y4390 = ~1'b0 ;
  assign y4391 = n9021 ;
  assign y4392 = ~n9026 ;
  assign y4393 = n9030 ;
  assign y4394 = n9032 ;
  assign y4395 = ~n9034 ;
  assign y4396 = ~n9036 ;
  assign y4397 = ~1'b0 ;
  assign y4398 = ~1'b0 ;
  assign y4399 = ~n9039 ;
  assign y4400 = ~1'b0 ;
  assign y4401 = ~n9040 ;
  assign y4402 = n9043 ;
  assign y4403 = ~1'b0 ;
  assign y4404 = n9046 ;
  assign y4405 = ~n6523 ;
  assign y4406 = ~n1396 ;
  assign y4407 = ~n9049 ;
  assign y4408 = ~n9051 ;
  assign y4409 = ~n9057 ;
  assign y4410 = n9058 ;
  assign y4411 = n9060 ;
  assign y4412 = ~1'b0 ;
  assign y4413 = ~n9061 ;
  assign y4414 = ~n9065 ;
  assign y4415 = ~n9067 ;
  assign y4416 = n9068 ;
  assign y4417 = n9070 ;
  assign y4418 = ~1'b0 ;
  assign y4419 = ~n9072 ;
  assign y4420 = ~n9073 ;
  assign y4421 = ~n9075 ;
  assign y4422 = n9077 ;
  assign y4423 = ~n9079 ;
  assign y4424 = ~1'b0 ;
  assign y4425 = ~n9082 ;
  assign y4426 = ~n9086 ;
  assign y4427 = n9087 ;
  assign y4428 = n9091 ;
  assign y4429 = ~n9092 ;
  assign y4430 = n9098 ;
  assign y4431 = ~1'b0 ;
  assign y4432 = ~1'b0 ;
  assign y4433 = ~n9099 ;
  assign y4434 = ~1'b0 ;
  assign y4435 = ~n9100 ;
  assign y4436 = n9105 ;
  assign y4437 = 1'b0 ;
  assign y4438 = n2596 ;
  assign y4439 = ~1'b0 ;
  assign y4440 = ~n9106 ;
  assign y4441 = ~n9109 ;
  assign y4442 = n9112 ;
  assign y4443 = ~1'b0 ;
  assign y4444 = ~n9114 ;
  assign y4445 = ~n9116 ;
  assign y4446 = n9119 ;
  assign y4447 = ~n9123 ;
  assign y4448 = n9124 ;
  assign y4449 = ~n9125 ;
  assign y4450 = n9128 ;
  assign y4451 = ~n9129 ;
  assign y4452 = ~n9131 ;
  assign y4453 = ~n9134 ;
  assign y4454 = ~n9136 ;
  assign y4455 = n9139 ;
  assign y4456 = ~1'b0 ;
  assign y4457 = ~1'b0 ;
  assign y4458 = n805 ;
  assign y4459 = n9143 ;
  assign y4460 = ~n9144 ;
  assign y4461 = n9147 ;
  assign y4462 = ~1'b0 ;
  assign y4463 = n8416 ;
  assign y4464 = ~1'b0 ;
  assign y4465 = ~n9148 ;
  assign y4466 = n9151 ;
  assign y4467 = n9158 ;
  assign y4468 = n9161 ;
  assign y4469 = n9162 ;
  assign y4470 = n9165 ;
  assign y4471 = ~1'b0 ;
  assign y4472 = n9170 ;
  assign y4473 = ~1'b0 ;
  assign y4474 = ~n9171 ;
  assign y4475 = n9180 ;
  assign y4476 = ~1'b0 ;
  assign y4477 = n9187 ;
  assign y4478 = ~1'b0 ;
  assign y4479 = n9191 ;
  assign y4480 = ~n7575 ;
  assign y4481 = ~n9196 ;
  assign y4482 = ~1'b0 ;
  assign y4483 = ~n9197 ;
  assign y4484 = ~1'b0 ;
  assign y4485 = n9200 ;
  assign y4486 = ~n9202 ;
  assign y4487 = ~n9203 ;
  assign y4488 = ~n9209 ;
  assign y4489 = n9213 ;
  assign y4490 = ~1'b0 ;
  assign y4491 = 1'b0 ;
  assign y4492 = n9000 ;
  assign y4493 = n9215 ;
  assign y4494 = n9216 ;
  assign y4495 = ~n9217 ;
  assign y4496 = ~1'b0 ;
  assign y4497 = n9223 ;
  assign y4498 = ~n9227 ;
  assign y4499 = ~n9229 ;
  assign y4500 = ~1'b0 ;
  assign y4501 = ~1'b0 ;
  assign y4502 = n3097 ;
  assign y4503 = n9240 ;
  assign y4504 = ~n7045 ;
  assign y4505 = ~n9248 ;
  assign y4506 = n9249 ;
  assign y4507 = ~n9253 ;
  assign y4508 = ~n9255 ;
  assign y4509 = n9259 ;
  assign y4510 = ~n9261 ;
  assign y4511 = ~1'b0 ;
  assign y4512 = ~1'b0 ;
  assign y4513 = ~n9262 ;
  assign y4514 = n6412 ;
  assign y4515 = ~1'b0 ;
  assign y4516 = 1'b0 ;
  assign y4517 = ~n9267 ;
  assign y4518 = n9276 ;
  assign y4519 = 1'b0 ;
  assign y4520 = ~n9277 ;
  assign y4521 = ~1'b0 ;
  assign y4522 = n9278 ;
  assign y4523 = n9279 ;
  assign y4524 = ~n2330 ;
  assign y4525 = ~n9283 ;
  assign y4526 = ~n9286 ;
  assign y4527 = n9287 ;
  assign y4528 = ~1'b0 ;
  assign y4529 = ~n9288 ;
  assign y4530 = ~n9290 ;
  assign y4531 = ~n9293 ;
  assign y4532 = ~1'b0 ;
  assign y4533 = n4985 ;
  assign y4534 = ~1'b0 ;
  assign y4535 = ~1'b0 ;
  assign y4536 = n9297 ;
  assign y4537 = ~n9298 ;
  assign y4538 = ~1'b0 ;
  assign y4539 = ~1'b0 ;
  assign y4540 = ~1'b0 ;
  assign y4541 = n9299 ;
  assign y4542 = n9302 ;
  assign y4543 = ~1'b0 ;
  assign y4544 = ~n9304 ;
  assign y4545 = ~n1422 ;
  assign y4546 = ~n9305 ;
  assign y4547 = ~1'b0 ;
  assign y4548 = ~n9307 ;
  assign y4549 = ~1'b0 ;
  assign y4550 = n9312 ;
  assign y4551 = ~1'b0 ;
  assign y4552 = ~n9313 ;
  assign y4553 = ~n9315 ;
  assign y4554 = ~n9317 ;
  assign y4555 = n9322 ;
  assign y4556 = n9325 ;
  assign y4557 = ~n9330 ;
  assign y4558 = n9338 ;
  assign y4559 = 1'b0 ;
  assign y4560 = ~n8299 ;
  assign y4561 = n2228 ;
  assign y4562 = ~n9344 ;
  assign y4563 = ~n9349 ;
  assign y4564 = ~1'b0 ;
  assign y4565 = n6148 ;
  assign y4566 = n9353 ;
  assign y4567 = n9356 ;
  assign y4568 = n9358 ;
  assign y4569 = ~n607 ;
  assign y4570 = ~n9360 ;
  assign y4571 = ~n9362 ;
  assign y4572 = ~n9366 ;
  assign y4573 = n4159 ;
  assign y4574 = n9368 ;
  assign y4575 = ~n3762 ;
  assign y4576 = n9370 ;
  assign y4577 = ~n9372 ;
  assign y4578 = n9373 ;
  assign y4579 = ~1'b0 ;
  assign y4580 = n9375 ;
  assign y4581 = ~1'b0 ;
  assign y4582 = n9377 ;
  assign y4583 = ~1'b0 ;
  assign y4584 = n9379 ;
  assign y4585 = n9381 ;
  assign y4586 = n9390 ;
  assign y4587 = ~1'b0 ;
  assign y4588 = ~1'b0 ;
  assign y4589 = n9391 ;
  assign y4590 = n9397 ;
  assign y4591 = n9399 ;
  assign y4592 = ~1'b0 ;
  assign y4593 = ~n2005 ;
  assign y4594 = n9400 ;
  assign y4595 = n9409 ;
  assign y4596 = ~n9412 ;
  assign y4597 = ~n9417 ;
  assign y4598 = ~1'b0 ;
  assign y4599 = ~1'b0 ;
  assign y4600 = ~1'b0 ;
  assign y4601 = n4613 ;
  assign y4602 = n9418 ;
  assign y4603 = ~n9423 ;
  assign y4604 = n9425 ;
  assign y4605 = ~n9427 ;
  assign y4606 = ~n9428 ;
  assign y4607 = ~1'b0 ;
  assign y4608 = ~1'b0 ;
  assign y4609 = n9429 ;
  assign y4610 = n9436 ;
  assign y4611 = n3758 ;
  assign y4612 = ~n9439 ;
  assign y4613 = ~1'b0 ;
  assign y4614 = n9441 ;
  assign y4615 = ~1'b0 ;
  assign y4616 = ~n9442 ;
  assign y4617 = ~1'b0 ;
  assign y4618 = n9445 ;
  assign y4619 = n9446 ;
  assign y4620 = ~n9450 ;
  assign y4621 = ~n9451 ;
  assign y4622 = ~1'b0 ;
  assign y4623 = ~n9453 ;
  assign y4624 = ~1'b0 ;
  assign y4625 = ~n9455 ;
  assign y4626 = n9456 ;
  assign y4627 = ~1'b0 ;
  assign y4628 = n9458 ;
  assign y4629 = ~n9460 ;
  assign y4630 = ~n9463 ;
  assign y4631 = n9465 ;
  assign y4632 = ~n9469 ;
  assign y4633 = ~n9471 ;
  assign y4634 = ~1'b0 ;
  assign y4635 = ~1'b0 ;
  assign y4636 = ~n900 ;
  assign y4637 = ~1'b0 ;
  assign y4638 = ~1'b0 ;
  assign y4639 = ~n9472 ;
  assign y4640 = ~1'b0 ;
  assign y4641 = ~n9473 ;
  assign y4642 = ~n9479 ;
  assign y4643 = ~n9484 ;
  assign y4644 = ~n9486 ;
  assign y4645 = ~1'b0 ;
  assign y4646 = n9490 ;
  assign y4647 = n9495 ;
  assign y4648 = ~1'b0 ;
  assign y4649 = n1033 ;
  assign y4650 = n9497 ;
  assign y4651 = n9498 ;
  assign y4652 = ~1'b0 ;
  assign y4653 = n9508 ;
  assign y4654 = ~n9510 ;
  assign y4655 = n9512 ;
  assign y4656 = n9513 ;
  assign y4657 = ~n9515 ;
  assign y4658 = n9518 ;
  assign y4659 = ~n9520 ;
  assign y4660 = ~1'b0 ;
  assign y4661 = n9522 ;
  assign y4662 = n9523 ;
  assign y4663 = ~n9527 ;
  assign y4664 = n9538 ;
  assign y4665 = ~n9540 ;
  assign y4666 = 1'b0 ;
  assign y4667 = ~1'b0 ;
  assign y4668 = n9542 ;
  assign y4669 = ~n9546 ;
  assign y4670 = n9550 ;
  assign y4671 = ~n9551 ;
  assign y4672 = ~1'b0 ;
  assign y4673 = ~1'b0 ;
  assign y4674 = n9552 ;
  assign y4675 = n9555 ;
  assign y4676 = ~n9556 ;
  assign y4677 = ~n9557 ;
  assign y4678 = ~1'b0 ;
  assign y4679 = ~n2156 ;
  assign y4680 = ~n9559 ;
  assign y4681 = n9566 ;
  assign y4682 = ~n9568 ;
  assign y4683 = ~n9573 ;
  assign y4684 = ~1'b0 ;
  assign y4685 = n9577 ;
  assign y4686 = ~1'b0 ;
  assign y4687 = n9578 ;
  assign y4688 = ~1'b0 ;
  assign y4689 = ~1'b0 ;
  assign y4690 = ~n1664 ;
  assign y4691 = ~1'b0 ;
  assign y4692 = ~1'b0 ;
  assign y4693 = n9581 ;
  assign y4694 = n9584 ;
  assign y4695 = ~n9594 ;
  assign y4696 = ~1'b0 ;
  assign y4697 = n9596 ;
  assign y4698 = n9598 ;
  assign y4699 = n9601 ;
  assign y4700 = ~n9604 ;
  assign y4701 = ~n9607 ;
  assign y4702 = ~1'b0 ;
  assign y4703 = ~1'b0 ;
  assign y4704 = 1'b0 ;
  assign y4705 = ~1'b0 ;
  assign y4706 = ~n9613 ;
  assign y4707 = n9615 ;
  assign y4708 = ~n9618 ;
  assign y4709 = ~n9627 ;
  assign y4710 = ~1'b0 ;
  assign y4711 = ~1'b0 ;
  assign y4712 = n9632 ;
  assign y4713 = n9635 ;
  assign y4714 = ~1'b0 ;
  assign y4715 = ~1'b0 ;
  assign y4716 = ~n9637 ;
  assign y4717 = ~n9642 ;
  assign y4718 = n9644 ;
  assign y4719 = ~n9646 ;
  assign y4720 = ~1'b0 ;
  assign y4721 = n9647 ;
  assign y4722 = ~1'b0 ;
  assign y4723 = ~n9650 ;
  assign y4724 = n9652 ;
  assign y4725 = n1143 ;
  assign y4726 = ~1'b0 ;
  assign y4727 = ~n9657 ;
  assign y4728 = ~1'b0 ;
  assign y4729 = ~n9660 ;
  assign y4730 = ~n9661 ;
  assign y4731 = ~n9662 ;
  assign y4732 = n9664 ;
  assign y4733 = n9665 ;
  assign y4734 = ~n9670 ;
  assign y4735 = ~1'b0 ;
  assign y4736 = n9671 ;
  assign y4737 = ~1'b0 ;
  assign y4738 = 1'b0 ;
  assign y4739 = ~n9672 ;
  assign y4740 = ~n9675 ;
  assign y4741 = n9677 ;
  assign y4742 = ~n9678 ;
  assign y4743 = ~1'b0 ;
  assign y4744 = ~n9680 ;
  assign y4745 = n9686 ;
  assign y4746 = 1'b0 ;
  assign y4747 = ~n9689 ;
  assign y4748 = ~1'b0 ;
  assign y4749 = n9690 ;
  assign y4750 = ~n9694 ;
  assign y4751 = ~1'b0 ;
  assign y4752 = ~n9695 ;
  assign y4753 = ~1'b0 ;
  assign y4754 = ~n5203 ;
  assign y4755 = n9696 ;
  assign y4756 = n9698 ;
  assign y4757 = ~1'b0 ;
  assign y4758 = ~n9701 ;
  assign y4759 = ~1'b0 ;
  assign y4760 = ~n9703 ;
  assign y4761 = n9706 ;
  assign y4762 = ~1'b0 ;
  assign y4763 = ~n9708 ;
  assign y4764 = ~1'b0 ;
  assign y4765 = ~1'b0 ;
  assign y4766 = ~n9710 ;
  assign y4767 = n9714 ;
  assign y4768 = ~n9716 ;
  assign y4769 = ~1'b0 ;
  assign y4770 = n9717 ;
  assign y4771 = ~n9718 ;
  assign y4772 = ~1'b0 ;
  assign y4773 = 1'b0 ;
  assign y4774 = ~n9720 ;
  assign y4775 = ~1'b0 ;
  assign y4776 = ~1'b0 ;
  assign y4777 = n3973 ;
  assign y4778 = n9727 ;
  assign y4779 = x64 ;
  assign y4780 = n9733 ;
  assign y4781 = ~n9734 ;
  assign y4782 = ~n9752 ;
  assign y4783 = ~n9755 ;
  assign y4784 = ~n9759 ;
  assign y4785 = ~n2321 ;
  assign y4786 = ~n9763 ;
  assign y4787 = n9765 ;
  assign y4788 = ~n9766 ;
  assign y4789 = ~1'b0 ;
  assign y4790 = 1'b0 ;
  assign y4791 = ~n9771 ;
  assign y4792 = ~1'b0 ;
  assign y4793 = ~n9773 ;
  assign y4794 = n9774 ;
  assign y4795 = ~1'b0 ;
  assign y4796 = n9775 ;
  assign y4797 = n9776 ;
  assign y4798 = ~n9779 ;
  assign y4799 = n9780 ;
  assign y4800 = ~1'b0 ;
  assign y4801 = ~1'b0 ;
  assign y4802 = ~n9783 ;
  assign y4803 = ~1'b0 ;
  assign y4804 = n9786 ;
  assign y4805 = ~1'b0 ;
  assign y4806 = ~n7902 ;
  assign y4807 = ~n9789 ;
  assign y4808 = n9793 ;
  assign y4809 = ~n9795 ;
  assign y4810 = n6523 ;
  assign y4811 = ~1'b0 ;
  assign y4812 = n9797 ;
  assign y4813 = ~1'b0 ;
  assign y4814 = n9801 ;
  assign y4815 = n9802 ;
  assign y4816 = n9807 ;
  assign y4817 = ~n9808 ;
  assign y4818 = ~n9811 ;
  assign y4819 = ~n9812 ;
  assign y4820 = n9815 ;
  assign y4821 = ~n9819 ;
  assign y4822 = 1'b0 ;
  assign y4823 = ~n9820 ;
  assign y4824 = ~n9821 ;
  assign y4825 = ~n9824 ;
  assign y4826 = n9829 ;
  assign y4827 = n9832 ;
  assign y4828 = ~1'b0 ;
  assign y4829 = ~n9834 ;
  assign y4830 = ~1'b0 ;
  assign y4831 = ~n9842 ;
  assign y4832 = ~1'b0 ;
  assign y4833 = n9843 ;
  assign y4834 = ~n9848 ;
  assign y4835 = n9851 ;
  assign y4836 = ~n9855 ;
  assign y4837 = ~n9861 ;
  assign y4838 = ~1'b0 ;
  assign y4839 = ~1'b0 ;
  assign y4840 = ~1'b0 ;
  assign y4841 = ~n9864 ;
  assign y4842 = ~1'b0 ;
  assign y4843 = ~n9867 ;
  assign y4844 = n9868 ;
  assign y4845 = n9873 ;
  assign y4846 = n9874 ;
  assign y4847 = ~n9878 ;
  assign y4848 = n9879 ;
  assign y4849 = ~n9882 ;
  assign y4850 = ~n9884 ;
  assign y4851 = n9886 ;
  assign y4852 = ~n9891 ;
  assign y4853 = n9892 ;
  assign y4854 = ~n4923 ;
  assign y4855 = 1'b0 ;
  assign y4856 = n9895 ;
  assign y4857 = n9901 ;
  assign y4858 = n9902 ;
  assign y4859 = ~1'b0 ;
  assign y4860 = ~n9906 ;
  assign y4861 = ~n9908 ;
  assign y4862 = n9909 ;
  assign y4863 = ~n9913 ;
  assign y4864 = ~n9917 ;
  assign y4865 = n9919 ;
  assign y4866 = ~1'b0 ;
  assign y4867 = n9920 ;
  assign y4868 = ~n9927 ;
  assign y4869 = ~n9937 ;
  assign y4870 = ~1'b0 ;
  assign y4871 = ~n5665 ;
  assign y4872 = ~1'b0 ;
  assign y4873 = ~1'b0 ;
  assign y4874 = n9941 ;
  assign y4875 = ~1'b0 ;
  assign y4876 = ~n9942 ;
  assign y4877 = ~n9944 ;
  assign y4878 = ~1'b0 ;
  assign y4879 = n9946 ;
  assign y4880 = ~1'b0 ;
  assign y4881 = n9947 ;
  assign y4882 = 1'b0 ;
  assign y4883 = n9961 ;
  assign y4884 = ~n9966 ;
  assign y4885 = ~n9967 ;
  assign y4886 = n9969 ;
  assign y4887 = ~1'b0 ;
  assign y4888 = ~n9972 ;
  assign y4889 = ~1'b0 ;
  assign y4890 = n5911 ;
  assign y4891 = ~n9973 ;
  assign y4892 = ~1'b0 ;
  assign y4893 = ~n9977 ;
  assign y4894 = ~1'b0 ;
  assign y4895 = ~1'b0 ;
  assign y4896 = ~n9978 ;
  assign y4897 = n9980 ;
  assign y4898 = ~n9986 ;
  assign y4899 = ~n4973 ;
  assign y4900 = ~1'b0 ;
  assign y4901 = ~n3646 ;
  assign y4902 = ~1'b0 ;
  assign y4903 = ~1'b0 ;
  assign y4904 = ~n9992 ;
  assign y4905 = ~1'b0 ;
  assign y4906 = ~1'b0 ;
  assign y4907 = ~n9995 ;
  assign y4908 = ~1'b0 ;
  assign y4909 = ~n9997 ;
  assign y4910 = ~n9999 ;
  assign y4911 = ~n10003 ;
  assign y4912 = n4778 ;
  assign y4913 = ~n10007 ;
  assign y4914 = ~1'b0 ;
  assign y4915 = ~n10010 ;
  assign y4916 = ~n10013 ;
  assign y4917 = n10022 ;
  assign y4918 = n8092 ;
  assign y4919 = ~1'b0 ;
  assign y4920 = ~1'b0 ;
  assign y4921 = ~n10027 ;
  assign y4922 = n10029 ;
  assign y4923 = ~n10033 ;
  assign y4924 = ~1'b0 ;
  assign y4925 = ~n10035 ;
  assign y4926 = ~n10036 ;
  assign y4927 = ~n10040 ;
  assign y4928 = ~1'b0 ;
  assign y4929 = n9160 ;
  assign y4930 = 1'b0 ;
  assign y4931 = n10041 ;
  assign y4932 = n10043 ;
  assign y4933 = n10046 ;
  assign y4934 = n10047 ;
  assign y4935 = ~n10049 ;
  assign y4936 = ~n10051 ;
  assign y4937 = n10055 ;
  assign y4938 = ~n10057 ;
  assign y4939 = n10066 ;
  assign y4940 = ~n10069 ;
  assign y4941 = ~1'b0 ;
  assign y4942 = ~n10070 ;
  assign y4943 = ~1'b0 ;
  assign y4944 = ~n10073 ;
  assign y4945 = ~n10075 ;
  assign y4946 = ~n10077 ;
  assign y4947 = n10079 ;
  assign y4948 = n10084 ;
  assign y4949 = ~1'b0 ;
  assign y4950 = ~n10087 ;
  assign y4951 = n10089 ;
  assign y4952 = ~1'b0 ;
  assign y4953 = ~n10090 ;
  assign y4954 = ~n10096 ;
  assign y4955 = ~n10098 ;
  assign y4956 = n10101 ;
  assign y4957 = ~1'b0 ;
  assign y4958 = ~n10108 ;
  assign y4959 = n10110 ;
  assign y4960 = ~n10112 ;
  assign y4961 = ~n10115 ;
  assign y4962 = ~n10116 ;
  assign y4963 = 1'b0 ;
  assign y4964 = ~1'b0 ;
  assign y4965 = n10118 ;
  assign y4966 = ~n10120 ;
  assign y4967 = ~1'b0 ;
  assign y4968 = ~n10124 ;
  assign y4969 = ~1'b0 ;
  assign y4970 = ~n10125 ;
  assign y4971 = n10129 ;
  assign y4972 = ~1'b0 ;
  assign y4973 = ~n10131 ;
  assign y4974 = n275 ;
  assign y4975 = ~n10132 ;
  assign y4976 = n10133 ;
  assign y4977 = n10134 ;
  assign y4978 = ~x50 ;
  assign y4979 = ~n9240 ;
  assign y4980 = n10138 ;
  assign y4981 = n6437 ;
  assign y4982 = ~n10146 ;
  assign y4983 = ~n10150 ;
  assign y4984 = ~n10157 ;
  assign y4985 = ~n10159 ;
  assign y4986 = ~n10162 ;
  assign y4987 = ~n10165 ;
  assign y4988 = ~1'b0 ;
  assign y4989 = ~n10166 ;
  assign y4990 = ~n10169 ;
  assign y4991 = ~n10174 ;
  assign y4992 = ~n10178 ;
  assign y4993 = ~1'b0 ;
  assign y4994 = ~1'b0 ;
  assign y4995 = ~1'b0 ;
  assign y4996 = ~n10179 ;
  assign y4997 = n10180 ;
  assign y4998 = ~n10182 ;
  assign y4999 = ~n10185 ;
  assign y5000 = n10187 ;
  assign y5001 = ~n10192 ;
  assign y5002 = ~n10196 ;
  assign y5003 = n3139 ;
  assign y5004 = ~1'b0 ;
  assign y5005 = ~n10199 ;
  assign y5006 = n10200 ;
  assign y5007 = n10201 ;
  assign y5008 = ~n10202 ;
  assign y5009 = ~n10203 ;
  assign y5010 = ~n10207 ;
  assign y5011 = ~1'b0 ;
  assign y5012 = ~n10208 ;
  assign y5013 = n10211 ;
  assign y5014 = n10213 ;
  assign y5015 = n10219 ;
  assign y5016 = n10220 ;
  assign y5017 = ~n10224 ;
  assign y5018 = ~n10226 ;
  assign y5019 = ~1'b0 ;
  assign y5020 = 1'b0 ;
  assign y5021 = n10229 ;
  assign y5022 = n10233 ;
  assign y5023 = ~1'b0 ;
  assign y5024 = ~n10235 ;
  assign y5025 = ~n10237 ;
  assign y5026 = ~n10241 ;
  assign y5027 = ~1'b0 ;
  assign y5028 = ~n10244 ;
  assign y5029 = n10250 ;
  assign y5030 = ~1'b0 ;
  assign y5031 = ~n10251 ;
  assign y5032 = n10252 ;
  assign y5033 = n10254 ;
  assign y5034 = ~1'b0 ;
  assign y5035 = n10257 ;
  assign y5036 = ~1'b0 ;
  assign y5037 = ~n10259 ;
  assign y5038 = ~n10260 ;
  assign y5039 = ~1'b0 ;
  assign y5040 = ~1'b0 ;
  assign y5041 = ~1'b0 ;
  assign y5042 = ~1'b0 ;
  assign y5043 = ~1'b0 ;
  assign y5044 = n10262 ;
  assign y5045 = ~n10268 ;
  assign y5046 = ~n10269 ;
  assign y5047 = n7621 ;
  assign y5048 = ~1'b0 ;
  assign y5049 = n10270 ;
  assign y5050 = ~n10271 ;
  assign y5051 = ~n10275 ;
  assign y5052 = ~1'b0 ;
  assign y5053 = ~n10280 ;
  assign y5054 = ~n10287 ;
  assign y5055 = n10288 ;
  assign y5056 = ~1'b0 ;
  assign y5057 = n10290 ;
  assign y5058 = ~n10293 ;
  assign y5059 = ~1'b0 ;
  assign y5060 = ~1'b0 ;
  assign y5061 = ~1'b0 ;
  assign y5062 = n10296 ;
  assign y5063 = ~n10299 ;
  assign y5064 = n10300 ;
  assign y5065 = ~n4013 ;
  assign y5066 = ~n10307 ;
  assign y5067 = n10317 ;
  assign y5068 = ~n10322 ;
  assign y5069 = n10323 ;
  assign y5070 = n3868 ;
  assign y5071 = n10327 ;
  assign y5072 = ~1'b0 ;
  assign y5073 = ~1'b0 ;
  assign y5074 = ~1'b0 ;
  assign y5075 = ~1'b0 ;
  assign y5076 = ~n6953 ;
  assign y5077 = n10328 ;
  assign y5078 = ~n10332 ;
  assign y5079 = ~1'b0 ;
  assign y5080 = n10336 ;
  assign y5081 = n10340 ;
  assign y5082 = ~n10346 ;
  assign y5083 = ~n10348 ;
  assign y5084 = ~n10351 ;
  assign y5085 = ~n10355 ;
  assign y5086 = n10363 ;
  assign y5087 = ~n10365 ;
  assign y5088 = n8229 ;
  assign y5089 = n10366 ;
  assign y5090 = n10370 ;
  assign y5091 = ~n10371 ;
  assign y5092 = n10372 ;
  assign y5093 = n10373 ;
  assign y5094 = ~n4596 ;
  assign y5095 = ~1'b0 ;
  assign y5096 = n10375 ;
  assign y5097 = ~1'b0 ;
  assign y5098 = 1'b0 ;
  assign y5099 = ~1'b0 ;
  assign y5100 = ~n10381 ;
  assign y5101 = ~1'b0 ;
  assign y5102 = ~n10386 ;
  assign y5103 = ~1'b0 ;
  assign y5104 = ~1'b0 ;
  assign y5105 = n676 ;
  assign y5106 = ~1'b0 ;
  assign y5107 = ~n10387 ;
  assign y5108 = ~n1189 ;
  assign y5109 = n417 ;
  assign y5110 = ~n10388 ;
  assign y5111 = ~1'b0 ;
  assign y5112 = n10392 ;
  assign y5113 = ~1'b0 ;
  assign y5114 = ~1'b0 ;
  assign y5115 = n10394 ;
  assign y5116 = ~n10395 ;
  assign y5117 = n10398 ;
  assign y5118 = n10401 ;
  assign y5119 = 1'b0 ;
  assign y5120 = ~n10402 ;
  assign y5121 = n10407 ;
  assign y5122 = n8705 ;
  assign y5123 = n10411 ;
  assign y5124 = n10413 ;
  assign y5125 = ~n10414 ;
  assign y5126 = ~n10415 ;
  assign y5127 = n10420 ;
  assign y5128 = ~n10422 ;
  assign y5129 = ~n10424 ;
  assign y5130 = ~1'b0 ;
  assign y5131 = n10425 ;
  assign y5132 = ~n10427 ;
  assign y5133 = ~n10431 ;
  assign y5134 = n10433 ;
  assign y5135 = n10435 ;
  assign y5136 = n10441 ;
  assign y5137 = ~n10443 ;
  assign y5138 = ~n10444 ;
  assign y5139 = n10447 ;
  assign y5140 = ~1'b0 ;
  assign y5141 = ~n2737 ;
  assign y5142 = ~n10448 ;
  assign y5143 = ~1'b0 ;
  assign y5144 = ~n10452 ;
  assign y5145 = n10453 ;
  assign y5146 = ~1'b0 ;
  assign y5147 = ~1'b0 ;
  assign y5148 = n10457 ;
  assign y5149 = ~n10459 ;
  assign y5150 = ~n8599 ;
  assign y5151 = ~1'b0 ;
  assign y5152 = ~n10460 ;
  assign y5153 = n10462 ;
  assign y5154 = ~n10466 ;
  assign y5155 = ~1'b0 ;
  assign y5156 = ~n10471 ;
  assign y5157 = ~1'b0 ;
  assign y5158 = n10476 ;
  assign y5159 = ~1'b0 ;
  assign y5160 = ~n10477 ;
  assign y5161 = ~n10478 ;
  assign y5162 = ~n10481 ;
  assign y5163 = n10491 ;
  assign y5164 = n10492 ;
  assign y5165 = ~n10494 ;
  assign y5166 = ~n10496 ;
  assign y5167 = ~1'b0 ;
  assign y5168 = n10497 ;
  assign y5169 = ~n2278 ;
  assign y5170 = n3240 ;
  assign y5171 = ~n10503 ;
  assign y5172 = n10504 ;
  assign y5173 = n10509 ;
  assign y5174 = n10515 ;
  assign y5175 = ~n10517 ;
  assign y5176 = ~n10519 ;
  assign y5177 = ~1'b0 ;
  assign y5178 = ~n10520 ;
  assign y5179 = n10523 ;
  assign y5180 = n10525 ;
  assign y5181 = ~n10529 ;
  assign y5182 = ~1'b0 ;
  assign y5183 = ~1'b0 ;
  assign y5184 = ~1'b0 ;
  assign y5185 = ~n10532 ;
  assign y5186 = n5624 ;
  assign y5187 = ~n10535 ;
  assign y5188 = n10536 ;
  assign y5189 = n10538 ;
  assign y5190 = n10541 ;
  assign y5191 = ~1'b0 ;
  assign y5192 = n10542 ;
  assign y5193 = ~n10544 ;
  assign y5194 = n10547 ;
  assign y5195 = n10554 ;
  assign y5196 = ~x87 ;
  assign y5197 = n10555 ;
  assign y5198 = ~n2489 ;
  assign y5199 = ~n10557 ;
  assign y5200 = ~1'b0 ;
  assign y5201 = ~1'b0 ;
  assign y5202 = ~n10562 ;
  assign y5203 = ~n2168 ;
  assign y5204 = ~n10566 ;
  assign y5205 = n10568 ;
  assign y5206 = ~n8393 ;
  assign y5207 = ~1'b0 ;
  assign y5208 = ~n10571 ;
  assign y5209 = ~n10575 ;
  assign y5210 = n10580 ;
  assign y5211 = n10581 ;
  assign y5212 = ~n10582 ;
  assign y5213 = n10583 ;
  assign y5214 = n10586 ;
  assign y5215 = n10589 ;
  assign y5216 = ~n10592 ;
  assign y5217 = ~n10596 ;
  assign y5218 = n10598 ;
  assign y5219 = ~n10600 ;
  assign y5220 = ~1'b0 ;
  assign y5221 = ~1'b0 ;
  assign y5222 = n10602 ;
  assign y5223 = 1'b0 ;
  assign y5224 = ~1'b0 ;
  assign y5225 = n10603 ;
  assign y5226 = n10609 ;
  assign y5227 = ~1'b0 ;
  assign y5228 = ~n10610 ;
  assign y5229 = ~1'b0 ;
  assign y5230 = ~n10614 ;
  assign y5231 = n10616 ;
  assign y5232 = 1'b0 ;
  assign y5233 = ~n10619 ;
  assign y5234 = ~n10627 ;
  assign y5235 = ~n10628 ;
  assign y5236 = n10630 ;
  assign y5237 = n10632 ;
  assign y5238 = ~1'b0 ;
  assign y5239 = n10634 ;
  assign y5240 = ~n10635 ;
  assign y5241 = ~n7527 ;
  assign y5242 = n10637 ;
  assign y5243 = n2723 ;
  assign y5244 = ~1'b0 ;
  assign y5245 = ~n10638 ;
  assign y5246 = ~n10644 ;
  assign y5247 = ~n3253 ;
  assign y5248 = ~n10645 ;
  assign y5249 = ~1'b0 ;
  assign y5250 = n10647 ;
  assign y5251 = ~n10650 ;
  assign y5252 = n10659 ;
  assign y5253 = n10660 ;
  assign y5254 = n10665 ;
  assign y5255 = ~n10669 ;
  assign y5256 = n10671 ;
  assign y5257 = ~n10674 ;
  assign y5258 = ~1'b0 ;
  assign y5259 = ~n10675 ;
  assign y5260 = n10677 ;
  assign y5261 = n10678 ;
  assign y5262 = ~n10679 ;
  assign y5263 = ~n10681 ;
  assign y5264 = n10685 ;
  assign y5265 = ~n10686 ;
  assign y5266 = n10690 ;
  assign y5267 = n10691 ;
  assign y5268 = n2412 ;
  assign y5269 = n10700 ;
  assign y5270 = n4474 ;
  assign y5271 = n10702 ;
  assign y5272 = ~n10703 ;
  assign y5273 = n10704 ;
  assign y5274 = 1'b0 ;
  assign y5275 = ~1'b0 ;
  assign y5276 = ~n10705 ;
  assign y5277 = ~n5457 ;
  assign y5278 = n10709 ;
  assign y5279 = ~n10710 ;
  assign y5280 = n7463 ;
  assign y5281 = ~1'b0 ;
  assign y5282 = ~1'b0 ;
  assign y5283 = ~n10714 ;
  assign y5284 = n4973 ;
  assign y5285 = ~1'b0 ;
  assign y5286 = n10716 ;
  assign y5287 = ~1'b0 ;
  assign y5288 = ~n3130 ;
  assign y5289 = ~n10721 ;
  assign y5290 = 1'b0 ;
  assign y5291 = n10722 ;
  assign y5292 = ~n10725 ;
  assign y5293 = ~n10726 ;
  assign y5294 = ~1'b0 ;
  assign y5295 = ~1'b0 ;
  assign y5296 = n10727 ;
  assign y5297 = ~1'b0 ;
  assign y5298 = ~n10732 ;
  assign y5299 = n2170 ;
  assign y5300 = n10736 ;
  assign y5301 = ~n10737 ;
  assign y5302 = ~1'b0 ;
  assign y5303 = ~n10739 ;
  assign y5304 = n10744 ;
  assign y5305 = ~1'b0 ;
  assign y5306 = ~n10750 ;
  assign y5307 = ~1'b0 ;
  assign y5308 = n6569 ;
  assign y5309 = ~n10751 ;
  assign y5310 = n10754 ;
  assign y5311 = ~1'b0 ;
  assign y5312 = ~1'b0 ;
  assign y5313 = ~n10755 ;
  assign y5314 = ~n10757 ;
  assign y5315 = n10765 ;
  assign y5316 = n10773 ;
  assign y5317 = n10774 ;
  assign y5318 = n10777 ;
  assign y5319 = ~n10780 ;
  assign y5320 = ~n10783 ;
  assign y5321 = ~1'b0 ;
  assign y5322 = ~1'b0 ;
  assign y5323 = n10793 ;
  assign y5324 = ~n10801 ;
  assign y5325 = ~n10803 ;
  assign y5326 = n4759 ;
  assign y5327 = ~n3389 ;
  assign y5328 = n10805 ;
  assign y5329 = ~1'b0 ;
  assign y5330 = ~1'b0 ;
  assign y5331 = ~n10812 ;
  assign y5332 = ~1'b0 ;
  assign y5333 = ~1'b0 ;
  assign y5334 = ~1'b0 ;
  assign y5335 = n10816 ;
  assign y5336 = ~1'b0 ;
  assign y5337 = ~n10817 ;
  assign y5338 = ~1'b0 ;
  assign y5339 = n10818 ;
  assign y5340 = n10819 ;
  assign y5341 = ~n10826 ;
  assign y5342 = n10828 ;
  assign y5343 = n10829 ;
  assign y5344 = ~1'b0 ;
  assign y5345 = ~n10833 ;
  assign y5346 = ~n10835 ;
  assign y5347 = ~1'b0 ;
  assign y5348 = n10836 ;
  assign y5349 = ~1'b0 ;
  assign y5350 = ~1'b0 ;
  assign y5351 = n10839 ;
  assign y5352 = ~n10844 ;
  assign y5353 = n10845 ;
  assign y5354 = ~n10847 ;
  assign y5355 = ~1'b0 ;
  assign y5356 = ~n10848 ;
  assign y5357 = n10849 ;
  assign y5358 = ~n10852 ;
  assign y5359 = ~1'b0 ;
  assign y5360 = ~n10854 ;
  assign y5361 = ~1'b0 ;
  assign y5362 = ~n10858 ;
  assign y5363 = n10859 ;
  assign y5364 = 1'b0 ;
  assign y5365 = ~n10861 ;
  assign y5366 = ~n10864 ;
  assign y5367 = ~1'b0 ;
  assign y5368 = ~n10866 ;
  assign y5369 = n10867 ;
  assign y5370 = n10868 ;
  assign y5371 = ~n10871 ;
  assign y5372 = n272 ;
  assign y5373 = ~1'b0 ;
  assign y5374 = ~n10872 ;
  assign y5375 = ~n10875 ;
  assign y5376 = ~n10877 ;
  assign y5377 = ~n10884 ;
  assign y5378 = ~n10889 ;
  assign y5379 = ~n10892 ;
  assign y5380 = ~n10894 ;
  assign y5381 = n10895 ;
  assign y5382 = n10896 ;
  assign y5383 = ~n10899 ;
  assign y5384 = ~1'b0 ;
  assign y5385 = n10901 ;
  assign y5386 = n10903 ;
  assign y5387 = n10906 ;
  assign y5388 = n10913 ;
  assign y5389 = n3080 ;
  assign y5390 = ~n10916 ;
  assign y5391 = ~n10918 ;
  assign y5392 = n10920 ;
  assign y5393 = ~1'b0 ;
  assign y5394 = ~n2489 ;
  assign y5395 = n10921 ;
  assign y5396 = ~n10924 ;
  assign y5397 = ~1'b0 ;
  assign y5398 = ~1'b0 ;
  assign y5399 = ~n10925 ;
  assign y5400 = ~n10928 ;
  assign y5401 = ~1'b0 ;
  assign y5402 = n10929 ;
  assign y5403 = n2183 ;
  assign y5404 = n10931 ;
  assign y5405 = ~n5451 ;
  assign y5406 = ~1'b0 ;
  assign y5407 = n10932 ;
  assign y5408 = ~1'b0 ;
  assign y5409 = ~1'b0 ;
  assign y5410 = n10935 ;
  assign y5411 = n10936 ;
  assign y5412 = ~1'b0 ;
  assign y5413 = n10939 ;
  assign y5414 = ~n10940 ;
  assign y5415 = ~1'b0 ;
  assign y5416 = ~n10944 ;
  assign y5417 = 1'b0 ;
  assign y5418 = n10948 ;
  assign y5419 = ~n10952 ;
  assign y5420 = n5063 ;
  assign y5421 = ~1'b0 ;
  assign y5422 = n10957 ;
  assign y5423 = n10958 ;
  assign y5424 = 1'b0 ;
  assign y5425 = ~n4664 ;
  assign y5426 = ~n10960 ;
  assign y5427 = n6904 ;
  assign y5428 = ~n10966 ;
  assign y5429 = n9911 ;
  assign y5430 = ~n10967 ;
  assign y5431 = n10969 ;
  assign y5432 = ~1'b0 ;
  assign y5433 = n10970 ;
  assign y5434 = ~n10973 ;
  assign y5435 = n10974 ;
  assign y5436 = ~n10979 ;
  assign y5437 = n7012 ;
  assign y5438 = n10980 ;
  assign y5439 = ~1'b0 ;
  assign y5440 = n10984 ;
  assign y5441 = ~1'b0 ;
  assign y5442 = ~1'b0 ;
  assign y5443 = ~n10989 ;
  assign y5444 = n10990 ;
  assign y5445 = ~n10991 ;
  assign y5446 = ~1'b0 ;
  assign y5447 = n10993 ;
  assign y5448 = ~1'b0 ;
  assign y5449 = ~1'b0 ;
  assign y5450 = ~n10514 ;
  assign y5451 = ~n10994 ;
  assign y5452 = ~1'b0 ;
  assign y5453 = n10997 ;
  assign y5454 = n10999 ;
  assign y5455 = n11000 ;
  assign y5456 = ~n11001 ;
  assign y5457 = ~n11003 ;
  assign y5458 = ~n11006 ;
  assign y5459 = ~n11013 ;
  assign y5460 = ~n11015 ;
  assign y5461 = ~1'b0 ;
  assign y5462 = ~1'b0 ;
  assign y5463 = n11019 ;
  assign y5464 = ~n11021 ;
  assign y5465 = ~n11023 ;
  assign y5466 = ~n11025 ;
  assign y5467 = n11027 ;
  assign y5468 = ~n11029 ;
  assign y5469 = n11033 ;
  assign y5470 = n1512 ;
  assign y5471 = n11040 ;
  assign y5472 = ~1'b0 ;
  assign y5473 = ~n11043 ;
  assign y5474 = n11044 ;
  assign y5475 = 1'b0 ;
  assign y5476 = n3888 ;
  assign y5477 = ~1'b0 ;
  assign y5478 = ~n11046 ;
  assign y5479 = ~1'b0 ;
  assign y5480 = ~n11054 ;
  assign y5481 = n11056 ;
  assign y5482 = 1'b0 ;
  assign y5483 = ~n11061 ;
  assign y5484 = ~1'b0 ;
  assign y5485 = ~1'b0 ;
  assign y5486 = ~n4853 ;
  assign y5487 = ~1'b0 ;
  assign y5488 = n11064 ;
  assign y5489 = n5830 ;
  assign y5490 = n11065 ;
  assign y5491 = ~1'b0 ;
  assign y5492 = n11066 ;
  assign y5493 = n11069 ;
  assign y5494 = ~1'b0 ;
  assign y5495 = ~n11074 ;
  assign y5496 = n11076 ;
  assign y5497 = ~n309 ;
  assign y5498 = n11079 ;
  assign y5499 = n11085 ;
  assign y5500 = ~n11089 ;
  assign y5501 = n11090 ;
  assign y5502 = ~n11094 ;
  assign y5503 = ~n11098 ;
  assign y5504 = n11100 ;
  assign y5505 = ~1'b0 ;
  assign y5506 = n11102 ;
  assign y5507 = n11103 ;
  assign y5508 = n7280 ;
  assign y5509 = n11106 ;
  assign y5510 = n11107 ;
  assign y5511 = 1'b0 ;
  assign y5512 = 1'b0 ;
  assign y5513 = ~n11110 ;
  assign y5514 = ~n11114 ;
  assign y5515 = n11115 ;
  assign y5516 = ~n11119 ;
  assign y5517 = 1'b0 ;
  assign y5518 = ~1'b0 ;
  assign y5519 = ~n11123 ;
  assign y5520 = ~n11126 ;
  assign y5521 = ~1'b0 ;
  assign y5522 = n3505 ;
  assign y5523 = ~n11128 ;
  assign y5524 = ~n8237 ;
  assign y5525 = ~1'b0 ;
  assign y5526 = ~n11131 ;
  assign y5527 = n11133 ;
  assign y5528 = ~n11142 ;
  assign y5529 = ~1'b0 ;
  assign y5530 = ~n4333 ;
  assign y5531 = ~n11144 ;
  assign y5532 = ~n11147 ;
  assign y5533 = ~n11149 ;
  assign y5534 = ~1'b0 ;
  assign y5535 = n11150 ;
  assign y5536 = ~1'b0 ;
  assign y5537 = n11158 ;
  assign y5538 = ~n11163 ;
  assign y5539 = ~n11165 ;
  assign y5540 = ~n11167 ;
  assign y5541 = ~1'b0 ;
  assign y5542 = n11174 ;
  assign y5543 = n11175 ;
  assign y5544 = ~n11180 ;
  assign y5545 = ~n11185 ;
  assign y5546 = ~1'b0 ;
  assign y5547 = ~n11187 ;
  assign y5548 = n11191 ;
  assign y5549 = n11192 ;
  assign y5550 = ~n11194 ;
  assign y5551 = ~1'b0 ;
  assign y5552 = ~n11197 ;
  assign y5553 = ~1'b0 ;
  assign y5554 = n11200 ;
  assign y5555 = ~n11204 ;
  assign y5556 = n11207 ;
  assign y5557 = n11211 ;
  assign y5558 = ~n9176 ;
  assign y5559 = ~1'b0 ;
  assign y5560 = ~1'b0 ;
  assign y5561 = n11213 ;
  assign y5562 = ~n11217 ;
  assign y5563 = ~n11219 ;
  assign y5564 = ~1'b0 ;
  assign y5565 = n11221 ;
  assign y5566 = ~1'b0 ;
  assign y5567 = ~1'b0 ;
  assign y5568 = ~1'b0 ;
  assign y5569 = ~n9345 ;
  assign y5570 = ~n11229 ;
  assign y5571 = ~1'b0 ;
  assign y5572 = ~n11239 ;
  assign y5573 = ~1'b0 ;
  assign y5574 = n11243 ;
  assign y5575 = ~n11248 ;
  assign y5576 = n11253 ;
  assign y5577 = n11254 ;
  assign y5578 = ~1'b0 ;
  assign y5579 = ~n11256 ;
  assign y5580 = n11258 ;
  assign y5581 = ~n11260 ;
  assign y5582 = n11262 ;
  assign y5583 = ~n11263 ;
  assign y5584 = ~1'b0 ;
  assign y5585 = ~n7783 ;
  assign y5586 = ~n11264 ;
  assign y5587 = ~1'b0 ;
  assign y5588 = ~n11265 ;
  assign y5589 = ~1'b0 ;
  assign y5590 = n11276 ;
  assign y5591 = ~1'b0 ;
  assign y5592 = n11278 ;
  assign y5593 = n11286 ;
  assign y5594 = ~n11289 ;
  assign y5595 = n11293 ;
  assign y5596 = ~n11294 ;
  assign y5597 = ~n11295 ;
  assign y5598 = ~1'b0 ;
  assign y5599 = ~n11297 ;
  assign y5600 = ~1'b0 ;
  assign y5601 = ~n11298 ;
  assign y5602 = ~n11302 ;
  assign y5603 = n11304 ;
  assign y5604 = ~1'b0 ;
  assign y5605 = ~n11310 ;
  assign y5606 = ~1'b0 ;
  assign y5607 = ~n11311 ;
  assign y5608 = ~n11313 ;
  assign y5609 = n11315 ;
  assign y5610 = ~1'b0 ;
  assign y5611 = ~1'b0 ;
  assign y5612 = ~1'b0 ;
  assign y5613 = ~n11316 ;
  assign y5614 = n11320 ;
  assign y5615 = ~n10905 ;
  assign y5616 = n11322 ;
  assign y5617 = ~n11330 ;
  assign y5618 = n11331 ;
  assign y5619 = n11340 ;
  assign y5620 = ~n11341 ;
  assign y5621 = ~1'b0 ;
  assign y5622 = ~n11348 ;
  assign y5623 = ~1'b0 ;
  assign y5624 = n11350 ;
  assign y5625 = ~1'b0 ;
  assign y5626 = ~n11353 ;
  assign y5627 = ~n11357 ;
  assign y5628 = n11358 ;
  assign y5629 = ~n11361 ;
  assign y5630 = ~1'b0 ;
  assign y5631 = n11364 ;
  assign y5632 = n11365 ;
  assign y5633 = ~n11368 ;
  assign y5634 = n11371 ;
  assign y5635 = ~1'b0 ;
  assign y5636 = ~1'b0 ;
  assign y5637 = ~n11375 ;
  assign y5638 = ~n11382 ;
  assign y5639 = ~n6614 ;
  assign y5640 = ~x54 ;
  assign y5641 = 1'b0 ;
  assign y5642 = ~1'b0 ;
  assign y5643 = n11384 ;
  assign y5644 = n11387 ;
  assign y5645 = n11393 ;
  assign y5646 = n11396 ;
  assign y5647 = ~1'b0 ;
  assign y5648 = ~1'b0 ;
  assign y5649 = n11399 ;
  assign y5650 = n11400 ;
  assign y5651 = ~n11404 ;
  assign y5652 = ~n11408 ;
  assign y5653 = ~n11410 ;
  assign y5654 = ~1'b0 ;
  assign y5655 = ~n5630 ;
  assign y5656 = n11411 ;
  assign y5657 = ~n11412 ;
  assign y5658 = ~1'b0 ;
  assign y5659 = ~1'b0 ;
  assign y5660 = ~1'b0 ;
  assign y5661 = n11415 ;
  assign y5662 = ~1'b0 ;
  assign y5663 = ~1'b0 ;
  assign y5664 = ~n11419 ;
  assign y5665 = n11422 ;
  assign y5666 = ~n11423 ;
  assign y5667 = ~n11424 ;
  assign y5668 = ~n11428 ;
  assign y5669 = n11429 ;
  assign y5670 = ~1'b0 ;
  assign y5671 = ~1'b0 ;
  assign y5672 = n11438 ;
  assign y5673 = ~n3618 ;
  assign y5674 = ~n11440 ;
  assign y5675 = ~n11442 ;
  assign y5676 = ~n8787 ;
  assign y5677 = ~n11444 ;
  assign y5678 = n11452 ;
  assign y5679 = ~n11453 ;
  assign y5680 = ~n1121 ;
  assign y5681 = ~1'b0 ;
  assign y5682 = ~1'b0 ;
  assign y5683 = ~n11457 ;
  assign y5684 = ~1'b0 ;
  assign y5685 = ~n11466 ;
  assign y5686 = ~1'b0 ;
  assign y5687 = ~1'b0 ;
  assign y5688 = n11472 ;
  assign y5689 = ~1'b0 ;
  assign y5690 = ~n11478 ;
  assign y5691 = ~n11479 ;
  assign y5692 = n11482 ;
  assign y5693 = ~n11483 ;
  assign y5694 = ~n11484 ;
  assign y5695 = n11485 ;
  assign y5696 = ~n11487 ;
  assign y5697 = n11488 ;
  assign y5698 = n11491 ;
  assign y5699 = n5726 ;
  assign y5700 = ~n11495 ;
  assign y5701 = ~n11496 ;
  assign y5702 = ~n11498 ;
  assign y5703 = ~1'b0 ;
  assign y5704 = ~n11500 ;
  assign y5705 = n11502 ;
  assign y5706 = ~1'b0 ;
  assign y5707 = n8431 ;
  assign y5708 = ~1'b0 ;
  assign y5709 = ~1'b0 ;
  assign y5710 = ~1'b0 ;
  assign y5711 = n11504 ;
  assign y5712 = n11505 ;
  assign y5713 = n11506 ;
  assign y5714 = ~n11510 ;
  assign y5715 = ~n11512 ;
  assign y5716 = n11514 ;
  assign y5717 = ~n11518 ;
  assign y5718 = ~n11526 ;
  assign y5719 = ~1'b0 ;
  assign y5720 = ~n11527 ;
  assign y5721 = n11528 ;
  assign y5722 = 1'b0 ;
  assign y5723 = n11532 ;
  assign y5724 = n11534 ;
  assign y5725 = ~n11539 ;
  assign y5726 = n2091 ;
  assign y5727 = n11541 ;
  assign y5728 = ~1'b0 ;
  assign y5729 = ~n11542 ;
  assign y5730 = 1'b0 ;
  assign y5731 = 1'b0 ;
  assign y5732 = ~n11544 ;
  assign y5733 = ~n11545 ;
  assign y5734 = n11548 ;
  assign y5735 = ~n11552 ;
  assign y5736 = ~1'b0 ;
  assign y5737 = ~1'b0 ;
  assign y5738 = n11561 ;
  assign y5739 = ~n11563 ;
  assign y5740 = n11566 ;
  assign y5741 = n11572 ;
  assign y5742 = ~1'b0 ;
  assign y5743 = n11577 ;
  assign y5744 = n10809 ;
  assign y5745 = ~n11580 ;
  assign y5746 = ~n11582 ;
  assign y5747 = ~n11584 ;
  assign y5748 = ~n11585 ;
  assign y5749 = ~1'b0 ;
  assign y5750 = ~1'b0 ;
  assign y5751 = n11586 ;
  assign y5752 = ~n11588 ;
  assign y5753 = n11589 ;
  assign y5754 = n11590 ;
  assign y5755 = n11591 ;
  assign y5756 = ~n11592 ;
  assign y5757 = ~n7248 ;
  assign y5758 = ~1'b0 ;
  assign y5759 = n11595 ;
  assign y5760 = n9184 ;
  assign y5761 = ~n11596 ;
  assign y5762 = ~1'b0 ;
  assign y5763 = n11601 ;
  assign y5764 = ~1'b0 ;
  assign y5765 = n11602 ;
  assign y5766 = ~n11605 ;
  assign y5767 = ~n11609 ;
  assign y5768 = ~1'b0 ;
  assign y5769 = ~1'b0 ;
  assign y5770 = ~n11610 ;
  assign y5771 = ~n11611 ;
  assign y5772 = ~n11613 ;
  assign y5773 = 1'b0 ;
  assign y5774 = n11618 ;
  assign y5775 = ~1'b0 ;
  assign y5776 = ~n11621 ;
  assign y5777 = n11622 ;
  assign y5778 = n11634 ;
  assign y5779 = n11640 ;
  assign y5780 = ~n11645 ;
  assign y5781 = n11652 ;
  assign y5782 = ~1'b0 ;
  assign y5783 = ~1'b0 ;
  assign y5784 = n11653 ;
  assign y5785 = ~n11655 ;
  assign y5786 = n11657 ;
  assign y5787 = n11659 ;
  assign y5788 = ~n11667 ;
  assign y5789 = ~1'b0 ;
  assign y5790 = ~1'b0 ;
  assign y5791 = n11668 ;
  assign y5792 = ~1'b0 ;
  assign y5793 = n11670 ;
  assign y5794 = n11672 ;
  assign y5795 = 1'b0 ;
  assign y5796 = ~1'b0 ;
  assign y5797 = 1'b0 ;
  assign y5798 = ~1'b0 ;
  assign y5799 = n11673 ;
  assign y5800 = ~n11675 ;
  assign y5801 = n11679 ;
  assign y5802 = n11681 ;
  assign y5803 = ~n11689 ;
  assign y5804 = 1'b0 ;
  assign y5805 = ~1'b0 ;
  assign y5806 = ~1'b0 ;
  assign y5807 = ~1'b0 ;
  assign y5808 = n11694 ;
  assign y5809 = n540 ;
  assign y5810 = ~n11698 ;
  assign y5811 = ~n11699 ;
  assign y5812 = ~1'b0 ;
  assign y5813 = ~n11703 ;
  assign y5814 = ~n5751 ;
  assign y5815 = ~n11704 ;
  assign y5816 = n11706 ;
  assign y5817 = n6907 ;
  assign y5818 = ~n11710 ;
  assign y5819 = ~n11713 ;
  assign y5820 = ~n11714 ;
  assign y5821 = n11719 ;
  assign y5822 = ~n11720 ;
  assign y5823 = n11725 ;
  assign y5824 = ~n11730 ;
  assign y5825 = ~n11738 ;
  assign y5826 = ~1'b0 ;
  assign y5827 = n11739 ;
  assign y5828 = n11740 ;
  assign y5829 = n11741 ;
  assign y5830 = ~n11745 ;
  assign y5831 = ~1'b0 ;
  assign y5832 = ~n3741 ;
  assign y5833 = n11747 ;
  assign y5834 = n11750 ;
  assign y5835 = n11751 ;
  assign y5836 = ~1'b0 ;
  assign y5837 = n11755 ;
  assign y5838 = ~n11756 ;
  assign y5839 = ~1'b0 ;
  assign y5840 = ~n11758 ;
  assign y5841 = ~1'b0 ;
  assign y5842 = ~n11764 ;
  assign y5843 = ~1'b0 ;
  assign y5844 = ~n11766 ;
  assign y5845 = ~n11770 ;
  assign y5846 = ~n11772 ;
  assign y5847 = n11773 ;
  assign y5848 = ~1'b0 ;
  assign y5849 = ~n11774 ;
  assign y5850 = ~n11783 ;
  assign y5851 = n11784 ;
  assign y5852 = ~1'b0 ;
  assign y5853 = n11786 ;
  assign y5854 = ~n11787 ;
  assign y5855 = n11790 ;
  assign y5856 = n11793 ;
  assign y5857 = ~1'b0 ;
  assign y5858 = ~n11796 ;
  assign y5859 = n11800 ;
  assign y5860 = ~n11801 ;
  assign y5861 = ~n11803 ;
  assign y5862 = ~1'b0 ;
  assign y5863 = ~n11805 ;
  assign y5864 = n11807 ;
  assign y5865 = ~1'b0 ;
  assign y5866 = ~n11808 ;
  assign y5867 = ~1'b0 ;
  assign y5868 = n11809 ;
  assign y5869 = ~1'b0 ;
  assign y5870 = ~1'b0 ;
  assign y5871 = ~1'b0 ;
  assign y5872 = ~n11815 ;
  assign y5873 = ~n11818 ;
  assign y5874 = ~n11820 ;
  assign y5875 = ~1'b0 ;
  assign y5876 = n11822 ;
  assign y5877 = n1102 ;
  assign y5878 = ~1'b0 ;
  assign y5879 = ~n11824 ;
  assign y5880 = ~1'b0 ;
  assign y5881 = ~1'b0 ;
  assign y5882 = n10602 ;
  assign y5883 = ~1'b0 ;
  assign y5884 = ~n11829 ;
  assign y5885 = n1609 ;
  assign y5886 = ~1'b0 ;
  assign y5887 = n11835 ;
  assign y5888 = n11840 ;
  assign y5889 = n11842 ;
  assign y5890 = ~1'b0 ;
  assign y5891 = 1'b0 ;
  assign y5892 = ~1'b0 ;
  assign y5893 = ~n1470 ;
  assign y5894 = ~n11844 ;
  assign y5895 = ~n11848 ;
  assign y5896 = n11849 ;
  assign y5897 = ~n11851 ;
  assign y5898 = ~n11853 ;
  assign y5899 = ~n11855 ;
  assign y5900 = n1627 ;
  assign y5901 = n11857 ;
  assign y5902 = n7705 ;
  assign y5903 = ~1'b0 ;
  assign y5904 = n11866 ;
  assign y5905 = ~n11872 ;
  assign y5906 = n11873 ;
  assign y5907 = n11875 ;
  assign y5908 = ~n11884 ;
  assign y5909 = ~1'b0 ;
  assign y5910 = ~1'b0 ;
  assign y5911 = ~n9878 ;
  assign y5912 = n11885 ;
  assign y5913 = ~n11889 ;
  assign y5914 = ~n11893 ;
  assign y5915 = ~1'b0 ;
  assign y5916 = n11904 ;
  assign y5917 = ~n11906 ;
  assign y5918 = ~n11915 ;
  assign y5919 = ~1'b0 ;
  assign y5920 = n9790 ;
  assign y5921 = n11916 ;
  assign y5922 = ~1'b0 ;
  assign y5923 = ~1'b0 ;
  assign y5924 = ~1'b0 ;
  assign y5925 = 1'b0 ;
  assign y5926 = ~1'b0 ;
  assign y5927 = ~1'b0 ;
  assign y5928 = ~n11919 ;
  assign y5929 = ~n11924 ;
  assign y5930 = n10580 ;
  assign y5931 = ~n11925 ;
  assign y5932 = n11927 ;
  assign y5933 = ~1'b0 ;
  assign y5934 = ~1'b0 ;
  assign y5935 = ~n11928 ;
  assign y5936 = 1'b0 ;
  assign y5937 = n2912 ;
  assign y5938 = ~1'b0 ;
  assign y5939 = ~n11932 ;
  assign y5940 = ~n11935 ;
  assign y5941 = ~n11936 ;
  assign y5942 = 1'b0 ;
  assign y5943 = ~1'b0 ;
  assign y5944 = ~n11937 ;
  assign y5945 = ~1'b0 ;
  assign y5946 = ~n11941 ;
  assign y5947 = ~n11944 ;
  assign y5948 = n11945 ;
  assign y5949 = ~n11947 ;
  assign y5950 = n11951 ;
  assign y5951 = ~n11953 ;
  assign y5952 = n11955 ;
  assign y5953 = ~1'b0 ;
  assign y5954 = ~1'b0 ;
  assign y5955 = ~n11958 ;
  assign y5956 = ~1'b0 ;
  assign y5957 = n11959 ;
  assign y5958 = ~n11961 ;
  assign y5959 = ~1'b0 ;
  assign y5960 = ~1'b0 ;
  assign y5961 = ~1'b0 ;
  assign y5962 = ~1'b0 ;
  assign y5963 = ~1'b0 ;
  assign y5964 = ~n7600 ;
  assign y5965 = n11962 ;
  assign y5966 = ~1'b0 ;
  assign y5967 = ~1'b0 ;
  assign y5968 = ~n11963 ;
  assign y5969 = ~n11964 ;
  assign y5970 = n11968 ;
  assign y5971 = ~n11969 ;
  assign y5972 = n11970 ;
  assign y5973 = n11972 ;
  assign y5974 = n11973 ;
  assign y5975 = ~n11974 ;
  assign y5976 = ~n11977 ;
  assign y5977 = ~1'b0 ;
  assign y5978 = ~1'b0 ;
  assign y5979 = n11983 ;
  assign y5980 = n11993 ;
  assign y5981 = ~n11994 ;
  assign y5982 = n8235 ;
  assign y5983 = ~n11996 ;
  assign y5984 = ~1'b0 ;
  assign y5985 = ~n11998 ;
  assign y5986 = n12000 ;
  assign y5987 = n12006 ;
  assign y5988 = ~n12009 ;
  assign y5989 = n12016 ;
  assign y5990 = ~1'b0 ;
  assign y5991 = ~1'b0 ;
  assign y5992 = n12018 ;
  assign y5993 = ~n12021 ;
  assign y5994 = ~1'b0 ;
  assign y5995 = ~n12028 ;
  assign y5996 = ~n12032 ;
  assign y5997 = ~n12035 ;
  assign y5998 = 1'b0 ;
  assign y5999 = n12038 ;
  assign y6000 = n12041 ;
  assign y6001 = n12043 ;
  assign y6002 = n12047 ;
  assign y6003 = ~n12054 ;
  assign y6004 = ~1'b0 ;
  assign y6005 = ~n12059 ;
  assign y6006 = n12061 ;
  assign y6007 = n12062 ;
  assign y6008 = 1'b0 ;
  assign y6009 = ~n12063 ;
  assign y6010 = n9696 ;
  assign y6011 = n12064 ;
  assign y6012 = n12066 ;
  assign y6013 = n12067 ;
  assign y6014 = ~n12072 ;
  assign y6015 = ~n12074 ;
  assign y6016 = ~n12076 ;
  assign y6017 = ~1'b0 ;
  assign y6018 = ~1'b0 ;
  assign y6019 = ~n12077 ;
  assign y6020 = 1'b0 ;
  assign y6021 = n12079 ;
  assign y6022 = ~n12080 ;
  assign y6023 = ~n12081 ;
  assign y6024 = n12083 ;
  assign y6025 = ~1'b0 ;
  assign y6026 = 1'b0 ;
  assign y6027 = n7415 ;
  assign y6028 = ~n12084 ;
  assign y6029 = ~1'b0 ;
  assign y6030 = ~1'b0 ;
  assign y6031 = ~1'b0 ;
  assign y6032 = ~n12087 ;
  assign y6033 = n12091 ;
  assign y6034 = ~1'b0 ;
  assign y6035 = n12092 ;
  assign y6036 = ~n12094 ;
  assign y6037 = ~1'b0 ;
  assign y6038 = n12097 ;
  assign y6039 = ~n12098 ;
  assign y6040 = ~n10699 ;
  assign y6041 = ~n12100 ;
  assign y6042 = n12102 ;
  assign y6043 = ~1'b0 ;
  assign y6044 = ~n12123 ;
  assign y6045 = ~n12128 ;
  assign y6046 = ~n12129 ;
  assign y6047 = ~n12131 ;
  assign y6048 = ~n12132 ;
  assign y6049 = ~1'b0 ;
  assign y6050 = n12134 ;
  assign y6051 = ~n12135 ;
  assign y6052 = ~1'b0 ;
  assign y6053 = n12142 ;
  assign y6054 = n12143 ;
  assign y6055 = n12148 ;
  assign y6056 = ~1'b0 ;
  assign y6057 = n12149 ;
  assign y6058 = ~1'b0 ;
  assign y6059 = ~1'b0 ;
  assign y6060 = n12150 ;
  assign y6061 = n12154 ;
  assign y6062 = n12156 ;
  assign y6063 = ~n12157 ;
  assign y6064 = ~n5586 ;
  assign y6065 = ~1'b0 ;
  assign y6066 = ~n12160 ;
  assign y6067 = n12165 ;
  assign y6068 = n12167 ;
  assign y6069 = n12168 ;
  assign y6070 = n12172 ;
  assign y6071 = ~n12175 ;
  assign y6072 = ~n12181 ;
  assign y6073 = n12183 ;
  assign y6074 = ~1'b0 ;
  assign y6075 = n12186 ;
  assign y6076 = n12188 ;
  assign y6077 = ~n12199 ;
  assign y6078 = n12200 ;
  assign y6079 = ~1'b0 ;
  assign y6080 = ~1'b0 ;
  assign y6081 = ~n12203 ;
  assign y6082 = ~n12206 ;
  assign y6083 = ~n12210 ;
  assign y6084 = ~n2144 ;
  assign y6085 = ~1'b0 ;
  assign y6086 = ~1'b0 ;
  assign y6087 = n12216 ;
  assign y6088 = ~1'b0 ;
  assign y6089 = ~n12217 ;
  assign y6090 = n12220 ;
  assign y6091 = ~n6534 ;
  assign y6092 = n12224 ;
  assign y6093 = n12229 ;
  assign y6094 = ~n12231 ;
  assign y6095 = ~n3388 ;
  assign y6096 = ~n12232 ;
  assign y6097 = ~1'b0 ;
  assign y6098 = ~n12233 ;
  assign y6099 = ~n12238 ;
  assign y6100 = n12239 ;
  assign y6101 = n12242 ;
  assign y6102 = ~1'b0 ;
  assign y6103 = ~1'b0 ;
  assign y6104 = ~1'b0 ;
  assign y6105 = n12243 ;
  assign y6106 = n12246 ;
  assign y6107 = ~1'b0 ;
  assign y6108 = ~1'b0 ;
  assign y6109 = ~1'b0 ;
  assign y6110 = ~n11410 ;
  assign y6111 = ~1'b0 ;
  assign y6112 = n12251 ;
  assign y6113 = n12256 ;
  assign y6114 = n12257 ;
  assign y6115 = ~1'b0 ;
  assign y6116 = ~1'b0 ;
  assign y6117 = ~1'b0 ;
  assign y6118 = ~1'b0 ;
  assign y6119 = n12263 ;
  assign y6120 = ~n12264 ;
  assign y6121 = 1'b0 ;
  assign y6122 = n12266 ;
  assign y6123 = ~n12268 ;
  assign y6124 = ~n12269 ;
  assign y6125 = ~n208 ;
  assign y6126 = ~n12271 ;
  assign y6127 = ~n600 ;
  assign y6128 = ~1'b0 ;
  assign y6129 = ~1'b0 ;
  assign y6130 = n2630 ;
  assign y6131 = 1'b0 ;
  assign y6132 = ~1'b0 ;
  assign y6133 = ~n12272 ;
  assign y6134 = ~1'b0 ;
  assign y6135 = ~1'b0 ;
  assign y6136 = ~1'b0 ;
  assign y6137 = ~1'b0 ;
  assign y6138 = ~1'b0 ;
  assign y6139 = ~1'b0 ;
  assign y6140 = 1'b0 ;
  assign y6141 = n12273 ;
  assign y6142 = n12274 ;
  assign y6143 = ~n12276 ;
  assign y6144 = ~n12281 ;
  assign y6145 = ~n12283 ;
  assign y6146 = n12284 ;
  assign y6147 = ~1'b0 ;
  assign y6148 = n12289 ;
  assign y6149 = ~n12291 ;
  assign y6150 = ~1'b0 ;
  assign y6151 = n8910 ;
  assign y6152 = ~n12292 ;
  assign y6153 = ~1'b0 ;
  assign y6154 = n12297 ;
  assign y6155 = ~1'b0 ;
  assign y6156 = ~n12299 ;
  assign y6157 = ~n2414 ;
  assign y6158 = ~1'b0 ;
  assign y6159 = n12304 ;
  assign y6160 = ~1'b0 ;
  assign y6161 = ~n8126 ;
  assign y6162 = n12306 ;
  assign y6163 = ~1'b0 ;
  assign y6164 = n12307 ;
  assign y6165 = ~1'b0 ;
  assign y6166 = n12308 ;
  assign y6167 = ~1'b0 ;
  assign y6168 = ~n12310 ;
  assign y6169 = ~1'b0 ;
  assign y6170 = ~n12317 ;
  assign y6171 = n12337 ;
  assign y6172 = ~1'b0 ;
  assign y6173 = ~n12338 ;
  assign y6174 = n12339 ;
  assign y6175 = ~n12340 ;
  assign y6176 = ~n12344 ;
  assign y6177 = n12353 ;
  assign y6178 = ~n12357 ;
  assign y6179 = n12361 ;
  assign y6180 = ~1'b0 ;
  assign y6181 = n12362 ;
  assign y6182 = ~n12363 ;
  assign y6183 = ~n12365 ;
  assign y6184 = n12367 ;
  assign y6185 = n12369 ;
  assign y6186 = n12372 ;
  assign y6187 = ~n12377 ;
  assign y6188 = n12380 ;
  assign y6189 = ~1'b0 ;
  assign y6190 = ~1'b0 ;
  assign y6191 = n12383 ;
  assign y6192 = ~n12386 ;
  assign y6193 = n12387 ;
  assign y6194 = ~n12390 ;
  assign y6195 = ~1'b0 ;
  assign y6196 = ~n11990 ;
  assign y6197 = n12391 ;
  assign y6198 = n12395 ;
  assign y6199 = n12396 ;
  assign y6200 = n12397 ;
  assign y6201 = ~n12399 ;
  assign y6202 = n12402 ;
  assign y6203 = ~1'b0 ;
  assign y6204 = ~n12404 ;
  assign y6205 = n12405 ;
  assign y6206 = ~n12406 ;
  assign y6207 = ~1'b0 ;
  assign y6208 = ~n12408 ;
  assign y6209 = ~1'b0 ;
  assign y6210 = ~1'b0 ;
  assign y6211 = n3532 ;
  assign y6212 = ~n12414 ;
  assign y6213 = n12416 ;
  assign y6214 = ~1'b0 ;
  assign y6215 = n12417 ;
  assign y6216 = ~1'b0 ;
  assign y6217 = n12421 ;
  assign y6218 = n12423 ;
  assign y6219 = ~n12424 ;
  assign y6220 = ~1'b0 ;
  assign y6221 = ~n12427 ;
  assign y6222 = ~n12428 ;
  assign y6223 = ~1'b0 ;
  assign y6224 = n12432 ;
  assign y6225 = ~1'b0 ;
  assign y6226 = ~1'b0 ;
  assign y6227 = ~1'b0 ;
  assign y6228 = n12434 ;
  assign y6229 = ~n12438 ;
  assign y6230 = ~1'b0 ;
  assign y6231 = ~n12439 ;
  assign y6232 = ~n10782 ;
  assign y6233 = ~1'b0 ;
  assign y6234 = ~n12440 ;
  assign y6235 = ~1'b0 ;
  assign y6236 = n12442 ;
  assign y6237 = n12444 ;
  assign y6238 = n12446 ;
  assign y6239 = n12452 ;
  assign y6240 = ~n12457 ;
  assign y6241 = ~n12458 ;
  assign y6242 = ~n12465 ;
  assign y6243 = n12468 ;
  assign y6244 = ~1'b0 ;
  assign y6245 = ~1'b0 ;
  assign y6246 = n12470 ;
  assign y6247 = ~1'b0 ;
  assign y6248 = n12479 ;
  assign y6249 = ~1'b0 ;
  assign y6250 = ~n12483 ;
  assign y6251 = n12485 ;
  assign y6252 = ~n12486 ;
  assign y6253 = ~1'b0 ;
  assign y6254 = ~n12487 ;
  assign y6255 = n12491 ;
  assign y6256 = n12500 ;
  assign y6257 = ~n12501 ;
  assign y6258 = ~n12503 ;
  assign y6259 = ~n12504 ;
  assign y6260 = ~1'b0 ;
  assign y6261 = ~n12507 ;
  assign y6262 = n12511 ;
  assign y6263 = ~n12513 ;
  assign y6264 = ~1'b0 ;
  assign y6265 = ~1'b0 ;
  assign y6266 = n12518 ;
  assign y6267 = ~1'b0 ;
  assign y6268 = ~1'b0 ;
  assign y6269 = ~n12522 ;
  assign y6270 = 1'b0 ;
  assign y6271 = ~n12524 ;
  assign y6272 = 1'b0 ;
  assign y6273 = ~n12525 ;
  assign y6274 = n12527 ;
  assign y6275 = ~1'b0 ;
  assign y6276 = n12530 ;
  assign y6277 = n12532 ;
  assign y6278 = ~n12534 ;
  assign y6279 = n12535 ;
  assign y6280 = ~n12538 ;
  assign y6281 = ~n12539 ;
  assign y6282 = ~1'b0 ;
  assign y6283 = 1'b0 ;
  assign y6284 = ~1'b0 ;
  assign y6285 = n12543 ;
  assign y6286 = n9214 ;
  assign y6287 = ~n12545 ;
  assign y6288 = 1'b0 ;
  assign y6289 = n12546 ;
  assign y6290 = ~n12548 ;
  assign y6291 = n12551 ;
  assign y6292 = ~1'b0 ;
  assign y6293 = ~n12554 ;
  assign y6294 = ~1'b0 ;
  assign y6295 = n12556 ;
  assign y6296 = ~n12558 ;
  assign y6297 = ~n12559 ;
  assign y6298 = ~n12565 ;
  assign y6299 = n12566 ;
  assign y6300 = ~n12567 ;
  assign y6301 = ~n12571 ;
  assign y6302 = n7055 ;
  assign y6303 = ~n12573 ;
  assign y6304 = n12582 ;
  assign y6305 = n12587 ;
  assign y6306 = n12589 ;
  assign y6307 = ~n12590 ;
  assign y6308 = ~n12591 ;
  assign y6309 = n12593 ;
  assign y6310 = ~1'b0 ;
  assign y6311 = n12594 ;
  assign y6312 = ~1'b0 ;
  assign y6313 = n12595 ;
  assign y6314 = ~n10275 ;
  assign y6315 = n12599 ;
  assign y6316 = ~n12602 ;
  assign y6317 = ~n12604 ;
  assign y6318 = n12605 ;
  assign y6319 = ~1'b0 ;
  assign y6320 = n12606 ;
  assign y6321 = n12609 ;
  assign y6322 = ~n12610 ;
  assign y6323 = ~1'b0 ;
  assign y6324 = n7968 ;
  assign y6325 = ~1'b0 ;
  assign y6326 = ~n12612 ;
  assign y6327 = n12613 ;
  assign y6328 = ~n12616 ;
  assign y6329 = n12618 ;
  assign y6330 = ~1'b0 ;
  assign y6331 = ~n12620 ;
  assign y6332 = ~n12621 ;
  assign y6333 = ~n12624 ;
  assign y6334 = ~n12625 ;
  assign y6335 = 1'b0 ;
  assign y6336 = n12627 ;
  assign y6337 = ~n12630 ;
  assign y6338 = n12635 ;
  assign y6339 = ~n12637 ;
  assign y6340 = ~n12641 ;
  assign y6341 = ~n12645 ;
  assign y6342 = ~n12647 ;
  assign y6343 = ~n12649 ;
  assign y6344 = 1'b0 ;
  assign y6345 = ~n12653 ;
  assign y6346 = ~n1296 ;
  assign y6347 = ~1'b0 ;
  assign y6348 = n12654 ;
  assign y6349 = ~n12656 ;
  assign y6350 = ~n12658 ;
  assign y6351 = n12667 ;
  assign y6352 = n12668 ;
  assign y6353 = n12669 ;
  assign y6354 = n12670 ;
  assign y6355 = ~n12674 ;
  assign y6356 = n12676 ;
  assign y6357 = ~n12677 ;
  assign y6358 = ~n12678 ;
  assign y6359 = ~n12679 ;
  assign y6360 = ~1'b0 ;
  assign y6361 = ~n12680 ;
  assign y6362 = ~1'b0 ;
  assign y6363 = n12681 ;
  assign y6364 = ~n12682 ;
  assign y6365 = n12684 ;
  assign y6366 = ~n12688 ;
  assign y6367 = ~n12690 ;
  assign y6368 = ~1'b0 ;
  assign y6369 = n12695 ;
  assign y6370 = n12709 ;
  assign y6371 = n12710 ;
  assign y6372 = ~n12716 ;
  assign y6373 = n12719 ;
  assign y6374 = n12723 ;
  assign y6375 = ~1'b0 ;
  assign y6376 = ~n12725 ;
  assign y6377 = n12727 ;
  assign y6378 = ~n12733 ;
  assign y6379 = ~1'b0 ;
  assign y6380 = ~n12740 ;
  assign y6381 = ~n12742 ;
  assign y6382 = ~n12743 ;
  assign y6383 = n12750 ;
  assign y6384 = ~1'b0 ;
  assign y6385 = ~n12754 ;
  assign y6386 = ~n12755 ;
  assign y6387 = ~n12756 ;
  assign y6388 = n12763 ;
  assign y6389 = ~1'b0 ;
  assign y6390 = ~1'b0 ;
  assign y6391 = ~n12764 ;
  assign y6392 = n12767 ;
  assign y6393 = n12768 ;
  assign y6394 = n12770 ;
  assign y6395 = ~n12776 ;
  assign y6396 = ~n12777 ;
  assign y6397 = ~1'b0 ;
  assign y6398 = n12779 ;
  assign y6399 = ~n12785 ;
  assign y6400 = ~n12788 ;
  assign y6401 = n12789 ;
  assign y6402 = ~1'b0 ;
  assign y6403 = ~1'b0 ;
  assign y6404 = ~1'b0 ;
  assign y6405 = ~1'b0 ;
  assign y6406 = ~1'b0 ;
  assign y6407 = ~n12795 ;
  assign y6408 = n5962 ;
  assign y6409 = ~n12800 ;
  assign y6410 = ~1'b0 ;
  assign y6411 = ~1'b0 ;
  assign y6412 = n12803 ;
  assign y6413 = ~n12805 ;
  assign y6414 = ~n12810 ;
  assign y6415 = n6794 ;
  assign y6416 = ~n12822 ;
  assign y6417 = n12833 ;
  assign y6418 = ~n12836 ;
  assign y6419 = ~n12838 ;
  assign y6420 = ~n12840 ;
  assign y6421 = n829 ;
  assign y6422 = ~n12842 ;
  assign y6423 = 1'b0 ;
  assign y6424 = n12843 ;
  assign y6425 = n12844 ;
  assign y6426 = n12845 ;
  assign y6427 = ~n12850 ;
  assign y6428 = n12853 ;
  assign y6429 = ~1'b0 ;
  assign y6430 = n12854 ;
  assign y6431 = ~1'b0 ;
  assign y6432 = ~1'b0 ;
  assign y6433 = ~n12858 ;
  assign y6434 = ~n12862 ;
  assign y6435 = n12863 ;
  assign y6436 = n12864 ;
  assign y6437 = n12867 ;
  assign y6438 = ~n6043 ;
  assign y6439 = ~n12869 ;
  assign y6440 = ~1'b0 ;
  assign y6441 = n12873 ;
  assign y6442 = ~1'b0 ;
  assign y6443 = ~n12876 ;
  assign y6444 = ~1'b0 ;
  assign y6445 = ~n12878 ;
  assign y6446 = ~1'b0 ;
  assign y6447 = n12879 ;
  assign y6448 = n11188 ;
  assign y6449 = ~1'b0 ;
  assign y6450 = ~n11307 ;
  assign y6451 = ~n12885 ;
  assign y6452 = ~1'b0 ;
  assign y6453 = n12893 ;
  assign y6454 = ~1'b0 ;
  assign y6455 = ~1'b0 ;
  assign y6456 = ~n12895 ;
  assign y6457 = ~1'b0 ;
  assign y6458 = ~1'b0 ;
  assign y6459 = n12896 ;
  assign y6460 = ~1'b0 ;
  assign y6461 = n12898 ;
  assign y6462 = ~n12899 ;
  assign y6463 = ~n12902 ;
  assign y6464 = ~n6716 ;
  assign y6465 = ~n12908 ;
  assign y6466 = n12909 ;
  assign y6467 = ~n12910 ;
  assign y6468 = ~n12911 ;
  assign y6469 = ~n12915 ;
  assign y6470 = ~1'b0 ;
  assign y6471 = n12922 ;
  assign y6472 = n12923 ;
  assign y6473 = ~n12924 ;
  assign y6474 = n12925 ;
  assign y6475 = ~n12931 ;
  assign y6476 = ~1'b0 ;
  assign y6477 = ~n12933 ;
  assign y6478 = ~n12937 ;
  assign y6479 = ~1'b0 ;
  assign y6480 = n12938 ;
  assign y6481 = n12939 ;
  assign y6482 = n12941 ;
  assign y6483 = n12947 ;
  assign y6484 = ~1'b0 ;
  assign y6485 = ~n12948 ;
  assign y6486 = n12950 ;
  assign y6487 = ~1'b0 ;
  assign y6488 = n12951 ;
  assign y6489 = ~n12952 ;
  assign y6490 = ~1'b0 ;
  assign y6491 = ~n12955 ;
  assign y6492 = n12958 ;
  assign y6493 = ~n12959 ;
  assign y6494 = ~n12961 ;
  assign y6495 = ~n12963 ;
  assign y6496 = n12964 ;
  assign y6497 = ~n12965 ;
  assign y6498 = ~1'b0 ;
  assign y6499 = n12967 ;
  assign y6500 = ~1'b0 ;
  assign y6501 = ~1'b0 ;
  assign y6502 = ~n12972 ;
  assign y6503 = ~1'b0 ;
  assign y6504 = n12974 ;
  assign y6505 = n12977 ;
  assign y6506 = ~1'b0 ;
  assign y6507 = n12978 ;
  assign y6508 = n8602 ;
  assign y6509 = ~n12982 ;
  assign y6510 = n12983 ;
  assign y6511 = ~n12984 ;
  assign y6512 = ~n12986 ;
  assign y6513 = ~n12987 ;
  assign y6514 = ~n12989 ;
  assign y6515 = ~n12990 ;
  assign y6516 = n12992 ;
  assign y6517 = n12994 ;
  assign y6518 = n12996 ;
  assign y6519 = ~n12997 ;
  assign y6520 = n13001 ;
  assign y6521 = ~n13004 ;
  assign y6522 = n8845 ;
  assign y6523 = ~n13009 ;
  assign y6524 = n13012 ;
  assign y6525 = ~n1119 ;
  assign y6526 = n13014 ;
  assign y6527 = n13015 ;
  assign y6528 = n13021 ;
  assign y6529 = ~n13022 ;
  assign y6530 = ~1'b0 ;
  assign y6531 = n3298 ;
  assign y6532 = n8068 ;
  assign y6533 = ~1'b0 ;
  assign y6534 = ~1'b0 ;
  assign y6535 = ~n13024 ;
  assign y6536 = ~1'b0 ;
  assign y6537 = ~1'b0 ;
  assign y6538 = ~n13030 ;
  assign y6539 = n13035 ;
  assign y6540 = ~n13038 ;
  assign y6541 = ~n13040 ;
  assign y6542 = ~n13043 ;
  assign y6543 = n13044 ;
  assign y6544 = ~1'b0 ;
  assign y6545 = n13052 ;
  assign y6546 = ~n13056 ;
  assign y6547 = n13057 ;
  assign y6548 = ~n13058 ;
  assign y6549 = ~n13060 ;
  assign y6550 = ~n11378 ;
  assign y6551 = n13062 ;
  assign y6552 = ~1'b0 ;
  assign y6553 = ~n13069 ;
  assign y6554 = ~1'b0 ;
  assign y6555 = ~n13072 ;
  assign y6556 = n13075 ;
  assign y6557 = ~n13078 ;
  assign y6558 = ~n13085 ;
  assign y6559 = ~1'b0 ;
  assign y6560 = ~1'b0 ;
  assign y6561 = n13088 ;
  assign y6562 = n13095 ;
  assign y6563 = ~1'b0 ;
  assign y6564 = ~n13102 ;
  assign y6565 = ~n13104 ;
  assign y6566 = ~n13106 ;
  assign y6567 = ~n4463 ;
  assign y6568 = ~1'b0 ;
  assign y6569 = n13107 ;
  assign y6570 = n13111 ;
  assign y6571 = ~n13113 ;
  assign y6572 = ~n2622 ;
  assign y6573 = ~1'b0 ;
  assign y6574 = ~n13118 ;
  assign y6575 = ~n13120 ;
  assign y6576 = n13125 ;
  assign y6577 = ~n13126 ;
  assign y6578 = ~1'b0 ;
  assign y6579 = n13129 ;
  assign y6580 = n13130 ;
  assign y6581 = n13131 ;
  assign y6582 = n13132 ;
  assign y6583 = ~n13133 ;
  assign y6584 = ~n13138 ;
  assign y6585 = 1'b0 ;
  assign y6586 = ~n13140 ;
  assign y6587 = 1'b0 ;
  assign y6588 = ~1'b0 ;
  assign y6589 = ~n13141 ;
  assign y6590 = ~n13146 ;
  assign y6591 = ~n13149 ;
  assign y6592 = ~n13150 ;
  assign y6593 = n13152 ;
  assign y6594 = ~1'b0 ;
  assign y6595 = ~1'b0 ;
  assign y6596 = ~1'b0 ;
  assign y6597 = n13153 ;
  assign y6598 = n13156 ;
  assign y6599 = ~1'b0 ;
  assign y6600 = ~n13159 ;
  assign y6601 = ~n13163 ;
  assign y6602 = ~n13164 ;
  assign y6603 = ~1'b0 ;
  assign y6604 = ~n13167 ;
  assign y6605 = ~n13168 ;
  assign y6606 = n3758 ;
  assign y6607 = ~n13170 ;
  assign y6608 = n13172 ;
  assign y6609 = ~1'b0 ;
  assign y6610 = ~n13174 ;
  assign y6611 = ~1'b0 ;
  assign y6612 = ~n6661 ;
  assign y6613 = ~1'b0 ;
  assign y6614 = ~1'b0 ;
  assign y6615 = ~n496 ;
  assign y6616 = ~n13177 ;
  assign y6617 = ~1'b0 ;
  assign y6618 = n13179 ;
  assign y6619 = ~n13181 ;
  assign y6620 = n13184 ;
  assign y6621 = 1'b0 ;
  assign y6622 = ~n13191 ;
  assign y6623 = n7308 ;
  assign y6624 = ~1'b0 ;
  assign y6625 = ~n13192 ;
  assign y6626 = n13193 ;
  assign y6627 = ~1'b0 ;
  assign y6628 = n13196 ;
  assign y6629 = ~n13197 ;
  assign y6630 = ~n13198 ;
  assign y6631 = ~n13200 ;
  assign y6632 = n13202 ;
  assign y6633 = n13206 ;
  assign y6634 = ~1'b0 ;
  assign y6635 = ~n13213 ;
  assign y6636 = ~1'b0 ;
  assign y6637 = n13214 ;
  assign y6638 = ~1'b0 ;
  assign y6639 = ~n13217 ;
  assign y6640 = n13218 ;
  assign y6641 = ~n13219 ;
  assign y6642 = n13220 ;
  assign y6643 = n13238 ;
  assign y6644 = ~1'b0 ;
  assign y6645 = n13241 ;
  assign y6646 = n13242 ;
  assign y6647 = ~n13244 ;
  assign y6648 = 1'b0 ;
  assign y6649 = ~n13248 ;
  assign y6650 = ~1'b0 ;
  assign y6651 = ~n13250 ;
  assign y6652 = ~1'b0 ;
  assign y6653 = n13254 ;
  assign y6654 = ~1'b0 ;
  assign y6655 = ~n13259 ;
  assign y6656 = ~1'b0 ;
  assign y6657 = ~n13260 ;
  assign y6658 = ~1'b0 ;
  assign y6659 = ~1'b0 ;
  assign y6660 = n13261 ;
  assign y6661 = ~n13266 ;
  assign y6662 = n13270 ;
  assign y6663 = ~1'b0 ;
  assign y6664 = n13275 ;
  assign y6665 = ~1'b0 ;
  assign y6666 = ~n13276 ;
  assign y6667 = n13277 ;
  assign y6668 = n13280 ;
  assign y6669 = ~n13281 ;
  assign y6670 = ~1'b0 ;
  assign y6671 = ~1'b0 ;
  assign y6672 = n4053 ;
  assign y6673 = ~1'b0 ;
  assign y6674 = n13282 ;
  assign y6675 = ~n13287 ;
  assign y6676 = ~n13289 ;
  assign y6677 = ~n13290 ;
  assign y6678 = n560 ;
  assign y6679 = ~1'b0 ;
  assign y6680 = n13293 ;
  assign y6681 = n13294 ;
  assign y6682 = ~1'b0 ;
  assign y6683 = ~1'b0 ;
  assign y6684 = n13303 ;
  assign y6685 = ~n13304 ;
  assign y6686 = n13306 ;
  assign y6687 = 1'b0 ;
  assign y6688 = ~1'b0 ;
  assign y6689 = n13307 ;
  assign y6690 = ~n13312 ;
  assign y6691 = ~1'b0 ;
  assign y6692 = ~1'b0 ;
  assign y6693 = ~n13313 ;
  assign y6694 = n13314 ;
  assign y6695 = n13317 ;
  assign y6696 = n2670 ;
  assign y6697 = ~n13319 ;
  assign y6698 = n13327 ;
  assign y6699 = ~n13332 ;
  assign y6700 = ~1'b0 ;
  assign y6701 = ~n13334 ;
  assign y6702 = ~1'b0 ;
  assign y6703 = ~1'b0 ;
  assign y6704 = ~n13337 ;
  assign y6705 = n13338 ;
  assign y6706 = n13342 ;
  assign y6707 = n13350 ;
  assign y6708 = n6347 ;
  assign y6709 = ~n13351 ;
  assign y6710 = n13352 ;
  assign y6711 = 1'b0 ;
  assign y6712 = ~1'b0 ;
  assign y6713 = ~n13354 ;
  assign y6714 = ~1'b0 ;
  assign y6715 = n13355 ;
  assign y6716 = n13356 ;
  assign y6717 = ~n13359 ;
  assign y6718 = n13362 ;
  assign y6719 = ~1'b0 ;
  assign y6720 = ~1'b0 ;
  assign y6721 = ~n13363 ;
  assign y6722 = ~1'b0 ;
  assign y6723 = n13365 ;
  assign y6724 = ~1'b0 ;
  assign y6725 = ~1'b0 ;
  assign y6726 = ~1'b0 ;
  assign y6727 = ~1'b0 ;
  assign y6728 = n13366 ;
  assign y6729 = n13372 ;
  assign y6730 = n13374 ;
  assign y6731 = n13375 ;
  assign y6732 = n13377 ;
  assign y6733 = ~n13379 ;
  assign y6734 = ~1'b0 ;
  assign y6735 = ~1'b0 ;
  assign y6736 = n12690 ;
  assign y6737 = n13380 ;
  assign y6738 = n13383 ;
  assign y6739 = n13385 ;
  assign y6740 = 1'b0 ;
  assign y6741 = n13388 ;
  assign y6742 = ~n13390 ;
  assign y6743 = n13394 ;
  assign y6744 = ~n13395 ;
  assign y6745 = ~n13398 ;
  assign y6746 = ~n13399 ;
  assign y6747 = ~n13401 ;
  assign y6748 = n13404 ;
  assign y6749 = ~n13406 ;
  assign y6750 = ~1'b0 ;
  assign y6751 = n13410 ;
  assign y6752 = ~1'b0 ;
  assign y6753 = n3269 ;
  assign y6754 = n13415 ;
  assign y6755 = n13421 ;
  assign y6756 = ~n13434 ;
  assign y6757 = n3641 ;
  assign y6758 = ~1'b0 ;
  assign y6759 = ~1'b0 ;
  assign y6760 = n13435 ;
  assign y6761 = ~n6598 ;
  assign y6762 = ~n13436 ;
  assign y6763 = n13441 ;
  assign y6764 = ~n13445 ;
  assign y6765 = ~1'b0 ;
  assign y6766 = ~n13446 ;
  assign y6767 = n13451 ;
  assign y6768 = ~n13452 ;
  assign y6769 = n13454 ;
  assign y6770 = n13455 ;
  assign y6771 = n13457 ;
  assign y6772 = n13459 ;
  assign y6773 = n13461 ;
  assign y6774 = ~n13462 ;
  assign y6775 = n13467 ;
  assign y6776 = ~n13468 ;
  assign y6777 = ~1'b0 ;
  assign y6778 = n13473 ;
  assign y6779 = ~1'b0 ;
  assign y6780 = ~1'b0 ;
  assign y6781 = ~1'b0 ;
  assign y6782 = ~1'b0 ;
  assign y6783 = n13475 ;
  assign y6784 = ~1'b0 ;
  assign y6785 = ~1'b0 ;
  assign y6786 = n13484 ;
  assign y6787 = ~n13486 ;
  assign y6788 = ~1'b0 ;
  assign y6789 = ~n13490 ;
  assign y6790 = n13495 ;
  assign y6791 = ~n13500 ;
  assign y6792 = n13503 ;
  assign y6793 = n13506 ;
  assign y6794 = ~1'b0 ;
  assign y6795 = n13507 ;
  assign y6796 = ~n13508 ;
  assign y6797 = n13509 ;
  assign y6798 = ~n13513 ;
  assign y6799 = n13514 ;
  assign y6800 = 1'b0 ;
  assign y6801 = ~n13519 ;
  assign y6802 = ~1'b0 ;
  assign y6803 = ~1'b0 ;
  assign y6804 = ~n13522 ;
  assign y6805 = ~n13527 ;
  assign y6806 = n13528 ;
  assign y6807 = ~1'b0 ;
  assign y6808 = 1'b0 ;
  assign y6809 = ~n13530 ;
  assign y6810 = ~n13532 ;
  assign y6811 = ~1'b0 ;
  assign y6812 = ~1'b0 ;
  assign y6813 = n13535 ;
  assign y6814 = n13536 ;
  assign y6815 = ~n13538 ;
  assign y6816 = ~1'b0 ;
  assign y6817 = ~n6036 ;
  assign y6818 = n13541 ;
  assign y6819 = ~1'b0 ;
  assign y6820 = n13543 ;
  assign y6821 = ~n13544 ;
  assign y6822 = ~1'b0 ;
  assign y6823 = ~n13545 ;
  assign y6824 = ~1'b0 ;
  assign y6825 = n13554 ;
  assign y6826 = ~n13555 ;
  assign y6827 = ~n1541 ;
  assign y6828 = n6830 ;
  assign y6829 = ~1'b0 ;
  assign y6830 = n13557 ;
  assign y6831 = ~1'b0 ;
  assign y6832 = n13560 ;
  assign y6833 = ~n13563 ;
  assign y6834 = n13566 ;
  assign y6835 = ~n13572 ;
  assign y6836 = ~1'b0 ;
  assign y6837 = ~1'b0 ;
  assign y6838 = ~n13574 ;
  assign y6839 = ~n13576 ;
  assign y6840 = ~n13579 ;
  assign y6841 = n1204 ;
  assign y6842 = n10352 ;
  assign y6843 = n13580 ;
  assign y6844 = ~1'b0 ;
  assign y6845 = n13582 ;
  assign y6846 = ~n13585 ;
  assign y6847 = ~n13586 ;
  assign y6848 = ~1'b0 ;
  assign y6849 = n3820 ;
  assign y6850 = n13588 ;
  assign y6851 = ~1'b0 ;
  assign y6852 = ~1'b0 ;
  assign y6853 = ~1'b0 ;
  assign y6854 = ~1'b0 ;
  assign y6855 = ~n13589 ;
  assign y6856 = ~n13590 ;
  assign y6857 = ~n13591 ;
  assign y6858 = ~n13598 ;
  assign y6859 = ~1'b0 ;
  assign y6860 = ~1'b0 ;
  assign y6861 = ~n13600 ;
  assign y6862 = ~1'b0 ;
  assign y6863 = n13608 ;
  assign y6864 = n13609 ;
  assign y6865 = ~1'b0 ;
  assign y6866 = n13610 ;
  assign y6867 = ~n13611 ;
  assign y6868 = n9847 ;
  assign y6869 = ~x113 ;
  assign y6870 = ~1'b0 ;
  assign y6871 = 1'b0 ;
  assign y6872 = n10782 ;
  assign y6873 = ~n13623 ;
  assign y6874 = ~1'b0 ;
  assign y6875 = n13629 ;
  assign y6876 = ~1'b0 ;
  assign y6877 = ~n13630 ;
  assign y6878 = ~1'b0 ;
  assign y6879 = ~1'b0 ;
  assign y6880 = ~1'b0 ;
  assign y6881 = ~1'b0 ;
  assign y6882 = ~n13631 ;
  assign y6883 = ~1'b0 ;
  assign y6884 = n3694 ;
  assign y6885 = ~1'b0 ;
  assign y6886 = ~n13632 ;
  assign y6887 = ~n13633 ;
  assign y6888 = ~n13634 ;
  assign y6889 = n13639 ;
  assign y6890 = n13640 ;
  assign y6891 = n13642 ;
  assign y6892 = n13645 ;
  assign y6893 = ~1'b0 ;
  assign y6894 = ~1'b0 ;
  assign y6895 = n13647 ;
  assign y6896 = ~n13650 ;
  assign y6897 = ~1'b0 ;
  assign y6898 = n13652 ;
  assign y6899 = ~n13653 ;
  assign y6900 = ~1'b0 ;
  assign y6901 = n10592 ;
  assign y6902 = ~1'b0 ;
  assign y6903 = n13654 ;
  assign y6904 = n13660 ;
  assign y6905 = n4763 ;
  assign y6906 = 1'b0 ;
  assign y6907 = ~n13661 ;
  assign y6908 = ~1'b0 ;
  assign y6909 = n13662 ;
  assign y6910 = ~n13664 ;
  assign y6911 = ~1'b0 ;
  assign y6912 = n13666 ;
  assign y6913 = ~1'b0 ;
  assign y6914 = ~n13667 ;
  assign y6915 = ~1'b0 ;
  assign y6916 = ~1'b0 ;
  assign y6917 = ~n13668 ;
  assign y6918 = ~n13672 ;
  assign y6919 = n13677 ;
  assign y6920 = ~n13678 ;
  assign y6921 = n13688 ;
  assign y6922 = ~1'b0 ;
  assign y6923 = ~n13689 ;
  assign y6924 = n13691 ;
  assign y6925 = n13693 ;
  assign y6926 = ~n13698 ;
  assign y6927 = ~n13702 ;
  assign y6928 = ~1'b0 ;
  assign y6929 = ~n7145 ;
  assign y6930 = ~n5850 ;
  assign y6931 = ~n13703 ;
  assign y6932 = ~n13706 ;
  assign y6933 = n777 ;
  assign y6934 = n13714 ;
  assign y6935 = ~n13716 ;
  assign y6936 = ~1'b0 ;
  assign y6937 = 1'b0 ;
  assign y6938 = n13719 ;
  assign y6939 = n13721 ;
  assign y6940 = n13727 ;
  assign y6941 = n2126 ;
  assign y6942 = ~n13728 ;
  assign y6943 = 1'b0 ;
  assign y6944 = n13731 ;
  assign y6945 = ~n13735 ;
  assign y6946 = ~n13736 ;
  assign y6947 = n13739 ;
  assign y6948 = ~n13743 ;
  assign y6949 = ~n13745 ;
  assign y6950 = ~1'b0 ;
  assign y6951 = n13748 ;
  assign y6952 = ~n13752 ;
  assign y6953 = ~1'b0 ;
  assign y6954 = ~n13756 ;
  assign y6955 = n13761 ;
  assign y6956 = ~n13763 ;
  assign y6957 = ~n9506 ;
  assign y6958 = n351 ;
  assign y6959 = ~n13764 ;
  assign y6960 = n10339 ;
  assign y6961 = ~1'b0 ;
  assign y6962 = ~1'b0 ;
  assign y6963 = ~1'b0 ;
  assign y6964 = n13765 ;
  assign y6965 = ~1'b0 ;
  assign y6966 = ~1'b0 ;
  assign y6967 = ~n12753 ;
  assign y6968 = ~1'b0 ;
  assign y6969 = n13768 ;
  assign y6970 = n13769 ;
  assign y6971 = n13772 ;
  assign y6972 = ~1'b0 ;
  assign y6973 = ~n12774 ;
  assign y6974 = ~n13774 ;
  assign y6975 = n13780 ;
  assign y6976 = ~n8720 ;
  assign y6977 = ~n13781 ;
  assign y6978 = n13782 ;
  assign y6979 = n13783 ;
  assign y6980 = ~n5092 ;
  assign y6981 = ~1'b0 ;
  assign y6982 = ~1'b0 ;
  assign y6983 = ~n13785 ;
  assign y6984 = ~1'b0 ;
  assign y6985 = ~1'b0 ;
  assign y6986 = ~n13786 ;
  assign y6987 = ~1'b0 ;
  assign y6988 = n13792 ;
  assign y6989 = ~n13795 ;
  assign y6990 = n13796 ;
  assign y6991 = ~1'b0 ;
  assign y6992 = ~n13800 ;
  assign y6993 = ~n13804 ;
  assign y6994 = 1'b0 ;
  assign y6995 = ~n13805 ;
  assign y6996 = ~1'b0 ;
  assign y6997 = ~n13808 ;
  assign y6998 = ~1'b0 ;
  assign y6999 = n13809 ;
  assign y7000 = ~n13810 ;
  assign y7001 = n13815 ;
  assign y7002 = ~n13816 ;
  assign y7003 = n13817 ;
  assign y7004 = n13827 ;
  assign y7005 = ~1'b0 ;
  assign y7006 = ~n13830 ;
  assign y7007 = ~n13833 ;
  assign y7008 = n13834 ;
  assign y7009 = n13839 ;
  assign y7010 = n487 ;
  assign y7011 = n450 ;
  assign y7012 = n13840 ;
  assign y7013 = ~1'b0 ;
  assign y7014 = ~1'b0 ;
  assign y7015 = ~n13841 ;
  assign y7016 = n13844 ;
  assign y7017 = ~n13849 ;
  assign y7018 = ~n11744 ;
  assign y7019 = n13851 ;
  assign y7020 = ~1'b0 ;
  assign y7021 = n13853 ;
  assign y7022 = n13855 ;
  assign y7023 = n13859 ;
  assign y7024 = n13861 ;
  assign y7025 = ~n13863 ;
  assign y7026 = ~n13870 ;
  assign y7027 = n13874 ;
  assign y7028 = n11488 ;
  assign y7029 = ~n13876 ;
  assign y7030 = n13880 ;
  assign y7031 = ~n13884 ;
  assign y7032 = ~n13885 ;
  assign y7033 = ~1'b0 ;
  assign y7034 = ~n13888 ;
  assign y7035 = n13890 ;
  assign y7036 = n13892 ;
  assign y7037 = ~n13894 ;
  assign y7038 = ~n13896 ;
  assign y7039 = ~1'b0 ;
  assign y7040 = ~1'b0 ;
  assign y7041 = ~1'b0 ;
  assign y7042 = ~1'b0 ;
  assign y7043 = ~n13898 ;
  assign y7044 = n13899 ;
  assign y7045 = n13900 ;
  assign y7046 = n13902 ;
  assign y7047 = ~1'b0 ;
  assign y7048 = 1'b0 ;
  assign y7049 = n13905 ;
  assign y7050 = ~1'b0 ;
  assign y7051 = ~1'b0 ;
  assign y7052 = n10291 ;
  assign y7053 = n13908 ;
  assign y7054 = ~1'b0 ;
  assign y7055 = n13909 ;
  assign y7056 = n13910 ;
  assign y7057 = ~n13911 ;
  assign y7058 = n13912 ;
  assign y7059 = ~n13914 ;
  assign y7060 = ~n13916 ;
  assign y7061 = ~n13917 ;
  assign y7062 = n3690 ;
  assign y7063 = n13922 ;
  assign y7064 = ~n13924 ;
  assign y7065 = n13926 ;
  assign y7066 = ~1'b0 ;
  assign y7067 = ~n13929 ;
  assign y7068 = ~n13930 ;
  assign y7069 = n13931 ;
  assign y7070 = ~n13932 ;
  assign y7071 = ~1'b0 ;
  assign y7072 = ~n13934 ;
  assign y7073 = n13936 ;
  assign y7074 = n13941 ;
  assign y7075 = ~1'b0 ;
  assign y7076 = ~1'b0 ;
  assign y7077 = ~1'b0 ;
  assign y7078 = n13942 ;
  assign y7079 = ~1'b0 ;
  assign y7080 = ~n9073 ;
  assign y7081 = n13943 ;
  assign y7082 = n13947 ;
  assign y7083 = ~n13949 ;
  assign y7084 = n13950 ;
  assign y7085 = n1200 ;
  assign y7086 = n12626 ;
  assign y7087 = n13955 ;
  assign y7088 = ~n13957 ;
  assign y7089 = n13959 ;
  assign y7090 = 1'b0 ;
  assign y7091 = ~n13960 ;
  assign y7092 = ~n13699 ;
  assign y7093 = ~n13961 ;
  assign y7094 = ~n13962 ;
  assign y7095 = n13963 ;
  assign y7096 = n13964 ;
  assign y7097 = n13966 ;
  assign y7098 = ~n13971 ;
  assign y7099 = n13973 ;
  assign y7100 = ~n13975 ;
  assign y7101 = ~n2268 ;
  assign y7102 = n13976 ;
  assign y7103 = n13979 ;
  assign y7104 = n13984 ;
  assign y7105 = n13986 ;
  assign y7106 = n13987 ;
  assign y7107 = n9288 ;
  assign y7108 = n13988 ;
  assign y7109 = n11067 ;
  assign y7110 = n13997 ;
  assign y7111 = ~n14004 ;
  assign y7112 = ~n14006 ;
  assign y7113 = n14011 ;
  assign y7114 = n3474 ;
  assign y7115 = ~1'b0 ;
  assign y7116 = ~1'b0 ;
  assign y7117 = n14012 ;
  assign y7118 = 1'b0 ;
  assign y7119 = ~1'b0 ;
  assign y7120 = ~1'b0 ;
  assign y7121 = ~n6759 ;
  assign y7122 = ~n14020 ;
  assign y7123 = ~n14023 ;
  assign y7124 = ~n14024 ;
  assign y7125 = ~1'b0 ;
  assign y7126 = ~1'b0 ;
  assign y7127 = ~n14029 ;
  assign y7128 = ~n14031 ;
  assign y7129 = ~1'b0 ;
  assign y7130 = ~1'b0 ;
  assign y7131 = ~1'b0 ;
  assign y7132 = ~n14033 ;
  assign y7133 = n14034 ;
  assign y7134 = n14038 ;
  assign y7135 = ~n14039 ;
  assign y7136 = ~n14041 ;
  assign y7137 = ~1'b0 ;
  assign y7138 = n14046 ;
  assign y7139 = ~n14054 ;
  assign y7140 = ~n11762 ;
  assign y7141 = ~n10747 ;
  assign y7142 = ~1'b0 ;
  assign y7143 = n14055 ;
  assign y7144 = ~n7902 ;
  assign y7145 = ~n14057 ;
  assign y7146 = ~n14059 ;
  assign y7147 = ~1'b0 ;
  assign y7148 = ~n14063 ;
  assign y7149 = n14068 ;
  assign y7150 = ~n14072 ;
  assign y7151 = n14082 ;
  assign y7152 = ~n14084 ;
  assign y7153 = ~n14086 ;
  assign y7154 = n14088 ;
  assign y7155 = ~n14089 ;
  assign y7156 = ~n12030 ;
  assign y7157 = ~n14092 ;
  assign y7158 = ~1'b0 ;
  assign y7159 = ~1'b0 ;
  assign y7160 = ~n14096 ;
  assign y7161 = n14097 ;
  assign y7162 = n14102 ;
  assign y7163 = ~n14104 ;
  assign y7164 = n14107 ;
  assign y7165 = ~n14109 ;
  assign y7166 = ~n14110 ;
  assign y7167 = n14113 ;
  assign y7168 = n3367 ;
  assign y7169 = ~1'b0 ;
  assign y7170 = n14115 ;
  assign y7171 = ~n14116 ;
  assign y7172 = ~n14117 ;
  assign y7173 = ~n14121 ;
  assign y7174 = ~n14130 ;
  assign y7175 = n14134 ;
  assign y7176 = n2956 ;
  assign y7177 = n14135 ;
  assign y7178 = ~1'b0 ;
  assign y7179 = ~n14142 ;
  assign y7180 = n14144 ;
  assign y7181 = ~1'b0 ;
  assign y7182 = n14152 ;
  assign y7183 = ~1'b0 ;
  assign y7184 = n14153 ;
  assign y7185 = ~1'b0 ;
  assign y7186 = n14160 ;
  assign y7187 = ~n14162 ;
  assign y7188 = n14164 ;
  assign y7189 = n14169 ;
  assign y7190 = n10460 ;
  assign y7191 = n9899 ;
  assign y7192 = ~n14170 ;
  assign y7193 = ~n14171 ;
  assign y7194 = ~n14175 ;
  assign y7195 = ~n14177 ;
  assign y7196 = n14179 ;
  assign y7197 = n5638 ;
  assign y7198 = n14182 ;
  assign y7199 = n14184 ;
  assign y7200 = ~1'b0 ;
  assign y7201 = ~1'b0 ;
  assign y7202 = ~n14190 ;
  assign y7203 = ~n14192 ;
  assign y7204 = n4428 ;
  assign y7205 = ~1'b0 ;
  assign y7206 = ~n14195 ;
  assign y7207 = ~n14202 ;
  assign y7208 = n14204 ;
  assign y7209 = n14205 ;
  assign y7210 = n14206 ;
  assign y7211 = ~1'b0 ;
  assign y7212 = ~n14207 ;
  assign y7213 = n14209 ;
  assign y7214 = ~n14212 ;
  assign y7215 = ~n14215 ;
  assign y7216 = ~1'b0 ;
  assign y7217 = ~1'b0 ;
  assign y7218 = n14220 ;
  assign y7219 = ~n14221 ;
  assign y7220 = 1'b0 ;
  assign y7221 = ~1'b0 ;
  assign y7222 = ~1'b0 ;
  assign y7223 = ~1'b0 ;
  assign y7224 = ~n14225 ;
  assign y7225 = ~n14226 ;
  assign y7226 = ~n14227 ;
  assign y7227 = ~n14230 ;
  assign y7228 = ~n14239 ;
  assign y7229 = ~n14242 ;
  assign y7230 = ~n14248 ;
  assign y7231 = ~1'b0 ;
  assign y7232 = ~n14249 ;
  assign y7233 = ~n14251 ;
  assign y7234 = n14252 ;
  assign y7235 = ~n14253 ;
  assign y7236 = ~n14258 ;
  assign y7237 = ~n14264 ;
  assign y7238 = n14266 ;
  assign y7239 = ~1'b0 ;
  assign y7240 = n14277 ;
  assign y7241 = n14282 ;
  assign y7242 = ~n14284 ;
  assign y7243 = ~1'b0 ;
  assign y7244 = ~n14287 ;
  assign y7245 = ~1'b0 ;
  assign y7246 = n14289 ;
  assign y7247 = ~n14291 ;
  assign y7248 = ~1'b0 ;
  assign y7249 = n14293 ;
  assign y7250 = ~n14295 ;
  assign y7251 = ~n14297 ;
  assign y7252 = ~1'b0 ;
  assign y7253 = n5958 ;
  assign y7254 = ~1'b0 ;
  assign y7255 = ~n14298 ;
  assign y7256 = ~1'b0 ;
  assign y7257 = n14301 ;
  assign y7258 = ~n14303 ;
  assign y7259 = ~n7906 ;
  assign y7260 = n4426 ;
  assign y7261 = ~n14305 ;
  assign y7262 = ~n14308 ;
  assign y7263 = n14311 ;
  assign y7264 = ~n14313 ;
  assign y7265 = ~1'b0 ;
  assign y7266 = ~1'b0 ;
  assign y7267 = ~n14314 ;
  assign y7268 = ~1'b0 ;
  assign y7269 = n14317 ;
  assign y7270 = ~n14318 ;
  assign y7271 = n14321 ;
  assign y7272 = ~n14322 ;
  assign y7273 = ~n14324 ;
  assign y7274 = ~1'b0 ;
  assign y7275 = ~1'b0 ;
  assign y7276 = ~n14326 ;
  assign y7277 = ~n2969 ;
  assign y7278 = n14327 ;
  assign y7279 = n14329 ;
  assign y7280 = ~1'b0 ;
  assign y7281 = n14338 ;
  assign y7282 = n14341 ;
  assign y7283 = n14344 ;
  assign y7284 = n14345 ;
  assign y7285 = ~1'b0 ;
  assign y7286 = ~n14348 ;
  assign y7287 = ~1'b0 ;
  assign y7288 = ~1'b0 ;
  assign y7289 = ~n3229 ;
  assign y7290 = ~1'b0 ;
  assign y7291 = ~1'b0 ;
  assign y7292 = n14349 ;
  assign y7293 = n14354 ;
  assign y7294 = ~n14355 ;
  assign y7295 = n14358 ;
  assign y7296 = ~1'b0 ;
  assign y7297 = ~n14361 ;
  assign y7298 = ~n14366 ;
  assign y7299 = n1343 ;
  assign y7300 = ~n14370 ;
  assign y7301 = ~1'b0 ;
  assign y7302 = ~n14377 ;
  assign y7303 = ~n14379 ;
  assign y7304 = n14385 ;
  assign y7305 = n14392 ;
  assign y7306 = 1'b0 ;
  assign y7307 = ~n14398 ;
  assign y7308 = ~1'b0 ;
  assign y7309 = ~n14399 ;
  assign y7310 = n14401 ;
  assign y7311 = ~1'b0 ;
  assign y7312 = ~1'b0 ;
  assign y7313 = ~n14402 ;
  assign y7314 = ~1'b0 ;
  assign y7315 = n14406 ;
  assign y7316 = ~n8366 ;
  assign y7317 = n14408 ;
  assign y7318 = ~n14410 ;
  assign y7319 = ~n7963 ;
  assign y7320 = ~n14416 ;
  assign y7321 = ~1'b0 ;
  assign y7322 = ~n14421 ;
  assign y7323 = n14425 ;
  assign y7324 = ~n14429 ;
  assign y7325 = n14430 ;
  assign y7326 = ~1'b0 ;
  assign y7327 = ~n14432 ;
  assign y7328 = ~n6034 ;
  assign y7329 = ~1'b0 ;
  assign y7330 = ~n9438 ;
  assign y7331 = n14436 ;
  assign y7332 = ~1'b0 ;
  assign y7333 = ~n14438 ;
  assign y7334 = ~n14443 ;
  assign y7335 = ~n14452 ;
  assign y7336 = ~1'b0 ;
  assign y7337 = 1'b0 ;
  assign y7338 = ~1'b0 ;
  assign y7339 = n14453 ;
  assign y7340 = n14454 ;
  assign y7341 = n14461 ;
  assign y7342 = n14463 ;
  assign y7343 = n14465 ;
  assign y7344 = ~n14467 ;
  assign y7345 = ~1'b0 ;
  assign y7346 = ~1'b0 ;
  assign y7347 = ~n14468 ;
  assign y7348 = ~n14470 ;
  assign y7349 = n14471 ;
  assign y7350 = ~1'b0 ;
  assign y7351 = ~1'b0 ;
  assign y7352 = n14472 ;
  assign y7353 = ~1'b0 ;
  assign y7354 = ~1'b0 ;
  assign y7355 = ~n14473 ;
  assign y7356 = ~n10485 ;
  assign y7357 = n5345 ;
  assign y7358 = ~n14477 ;
  assign y7359 = ~1'b0 ;
  assign y7360 = n14481 ;
  assign y7361 = n14482 ;
  assign y7362 = ~1'b0 ;
  assign y7363 = 1'b0 ;
  assign y7364 = n14483 ;
  assign y7365 = n14485 ;
  assign y7366 = ~n13882 ;
  assign y7367 = ~n1353 ;
  assign y7368 = ~1'b0 ;
  assign y7369 = ~n14486 ;
  assign y7370 = n14487 ;
  assign y7371 = ~1'b0 ;
  assign y7372 = ~1'b0 ;
  assign y7373 = ~n14492 ;
  assign y7374 = ~1'b0 ;
  assign y7375 = ~n461 ;
  assign y7376 = n14499 ;
  assign y7377 = ~1'b0 ;
  assign y7378 = n14504 ;
  assign y7379 = ~n14508 ;
  assign y7380 = ~n14511 ;
  assign y7381 = n14513 ;
  assign y7382 = ~1'b0 ;
  assign y7383 = ~1'b0 ;
  assign y7384 = n8097 ;
  assign y7385 = ~n14516 ;
  assign y7386 = ~n14517 ;
  assign y7387 = ~n3824 ;
  assign y7388 = ~n14522 ;
  assign y7389 = ~1'b0 ;
  assign y7390 = ~1'b0 ;
  assign y7391 = n14523 ;
  assign y7392 = n14524 ;
  assign y7393 = ~n13942 ;
  assign y7394 = ~n14527 ;
  assign y7395 = ~n14533 ;
  assign y7396 = ~n14536 ;
  assign y7397 = ~1'b0 ;
  assign y7398 = ~n14541 ;
  assign y7399 = ~1'b0 ;
  assign y7400 = n14543 ;
  assign y7401 = ~1'b0 ;
  assign y7402 = ~n456 ;
  assign y7403 = ~n14547 ;
  assign y7404 = ~n14550 ;
  assign y7405 = ~n14553 ;
  assign y7406 = ~1'b0 ;
  assign y7407 = n14554 ;
  assign y7408 = ~1'b0 ;
  assign y7409 = ~1'b0 ;
  assign y7410 = n8896 ;
  assign y7411 = ~1'b0 ;
  assign y7412 = ~1'b0 ;
  assign y7413 = n14556 ;
  assign y7414 = ~1'b0 ;
  assign y7415 = n14559 ;
  assign y7416 = ~n14560 ;
  assign y7417 = n4610 ;
  assign y7418 = ~1'b0 ;
  assign y7419 = ~n3674 ;
  assign y7420 = ~1'b0 ;
  assign y7421 = n8021 ;
  assign y7422 = ~n14567 ;
  assign y7423 = ~n14568 ;
  assign y7424 = ~n14570 ;
  assign y7425 = ~1'b0 ;
  assign y7426 = 1'b0 ;
  assign y7427 = ~n14572 ;
  assign y7428 = n14579 ;
  assign y7429 = 1'b0 ;
  assign y7430 = ~n14580 ;
  assign y7431 = ~1'b0 ;
  assign y7432 = ~n14582 ;
  assign y7433 = ~n3789 ;
  assign y7434 = ~n14588 ;
  assign y7435 = ~n14594 ;
  assign y7436 = ~1'b0 ;
  assign y7437 = n14600 ;
  assign y7438 = ~1'b0 ;
  assign y7439 = ~n14601 ;
  assign y7440 = ~1'b0 ;
  assign y7441 = ~1'b0 ;
  assign y7442 = 1'b0 ;
  assign y7443 = ~n14609 ;
  assign y7444 = n14615 ;
  assign y7445 = n14617 ;
  assign y7446 = n14623 ;
  assign y7447 = n14627 ;
  assign y7448 = n12812 ;
  assign y7449 = ~1'b0 ;
  assign y7450 = ~n14629 ;
  assign y7451 = 1'b0 ;
  assign y7452 = ~1'b0 ;
  assign y7453 = ~n12941 ;
  assign y7454 = n14630 ;
  assign y7455 = ~n14632 ;
  assign y7456 = n14633 ;
  assign y7457 = ~n14636 ;
  assign y7458 = ~n14637 ;
  assign y7459 = n4809 ;
  assign y7460 = ~n14639 ;
  assign y7461 = ~n14642 ;
  assign y7462 = ~n14645 ;
  assign y7463 = n14647 ;
  assign y7464 = ~n14649 ;
  assign y7465 = ~1'b0 ;
  assign y7466 = n14650 ;
  assign y7467 = ~n14658 ;
  assign y7468 = ~1'b0 ;
  assign y7469 = ~1'b0 ;
  assign y7470 = ~1'b0 ;
  assign y7471 = n14662 ;
  assign y7472 = ~n14665 ;
  assign y7473 = ~n14667 ;
  assign y7474 = ~n14669 ;
  assign y7475 = ~n14670 ;
  assign y7476 = ~n14672 ;
  assign y7477 = ~n14677 ;
  assign y7478 = n14678 ;
  assign y7479 = n14679 ;
  assign y7480 = ~1'b0 ;
  assign y7481 = ~n14682 ;
  assign y7482 = ~n14683 ;
  assign y7483 = ~1'b0 ;
  assign y7484 = ~n10152 ;
  assign y7485 = n14687 ;
  assign y7486 = n9894 ;
  assign y7487 = ~n14691 ;
  assign y7488 = n14692 ;
  assign y7489 = ~n14695 ;
  assign y7490 = ~n8850 ;
  assign y7491 = ~n14698 ;
  assign y7492 = ~n14699 ;
  assign y7493 = ~n14701 ;
  assign y7494 = ~1'b0 ;
  assign y7495 = n14702 ;
  assign y7496 = n14704 ;
  assign y7497 = ~n14706 ;
  assign y7498 = n14711 ;
  assign y7499 = ~n484 ;
  assign y7500 = n14714 ;
  assign y7501 = ~n14716 ;
  assign y7502 = ~n14717 ;
  assign y7503 = ~1'b0 ;
  assign y7504 = ~1'b0 ;
  assign y7505 = ~n14719 ;
  assign y7506 = n14720 ;
  assign y7507 = ~1'b0 ;
  assign y7508 = n14722 ;
  assign y7509 = ~n14724 ;
  assign y7510 = n14729 ;
  assign y7511 = ~1'b0 ;
  assign y7512 = ~n14731 ;
  assign y7513 = n14734 ;
  assign y7514 = ~n14739 ;
  assign y7515 = n10506 ;
  assign y7516 = ~n14741 ;
  assign y7517 = ~n14758 ;
  assign y7518 = ~n14760 ;
  assign y7519 = n14761 ;
  assign y7520 = ~n14762 ;
  assign y7521 = ~n14764 ;
  assign y7522 = ~n14768 ;
  assign y7523 = n14772 ;
  assign y7524 = ~n14774 ;
  assign y7525 = n14776 ;
  assign y7526 = ~n14780 ;
  assign y7527 = n14782 ;
  assign y7528 = n14786 ;
  assign y7529 = n14787 ;
  assign y7530 = n14789 ;
  assign y7531 = ~n14792 ;
  assign y7532 = n14799 ;
  assign y7533 = ~1'b0 ;
  assign y7534 = ~1'b0 ;
  assign y7535 = n14800 ;
  assign y7536 = ~1'b0 ;
  assign y7537 = ~1'b0 ;
  assign y7538 = n14805 ;
  assign y7539 = n14814 ;
  assign y7540 = n6653 ;
  assign y7541 = ~1'b0 ;
  assign y7542 = ~n14816 ;
  assign y7543 = ~n14818 ;
  assign y7544 = ~1'b0 ;
  assign y7545 = n14821 ;
  assign y7546 = ~n14823 ;
  assign y7547 = ~n4345 ;
  assign y7548 = ~n14828 ;
  assign y7549 = n14829 ;
  assign y7550 = ~1'b0 ;
  assign y7551 = ~1'b0 ;
  assign y7552 = n14837 ;
  assign y7553 = ~n14843 ;
  assign y7554 = 1'b0 ;
  assign y7555 = ~1'b0 ;
  assign y7556 = n14848 ;
  assign y7557 = ~n4650 ;
  assign y7558 = n14852 ;
  assign y7559 = ~n14853 ;
  assign y7560 = n14858 ;
  assign y7561 = n14859 ;
  assign y7562 = n14863 ;
  assign y7563 = ~n14875 ;
  assign y7564 = n14879 ;
  assign y7565 = ~n14880 ;
  assign y7566 = n14882 ;
  assign y7567 = ~n14886 ;
  assign y7568 = ~1'b0 ;
  assign y7569 = n14887 ;
  assign y7570 = ~n14889 ;
  assign y7571 = n14891 ;
  assign y7572 = n14894 ;
  assign y7573 = n14895 ;
  assign y7574 = n14896 ;
  assign y7575 = n14898 ;
  assign y7576 = n14902 ;
  assign y7577 = n14905 ;
  assign y7578 = ~1'b0 ;
  assign y7579 = ~n14910 ;
  assign y7580 = ~1'b0 ;
  assign y7581 = ~n14916 ;
  assign y7582 = ~1'b0 ;
  assign y7583 = ~1'b0 ;
  assign y7584 = n14918 ;
  assign y7585 = n14922 ;
  assign y7586 = ~n6000 ;
  assign y7587 = n14924 ;
  assign y7588 = ~1'b0 ;
  assign y7589 = n4578 ;
  assign y7590 = n14927 ;
  assign y7591 = ~1'b0 ;
  assign y7592 = ~n14929 ;
  assign y7593 = n14932 ;
  assign y7594 = n14935 ;
  assign y7595 = ~1'b0 ;
  assign y7596 = ~n14936 ;
  assign y7597 = ~n14942 ;
  assign y7598 = ~1'b0 ;
  assign y7599 = ~n14945 ;
  assign y7600 = n14946 ;
  assign y7601 = ~n14948 ;
  assign y7602 = n14950 ;
  assign y7603 = ~1'b0 ;
  assign y7604 = n14953 ;
  assign y7605 = n14954 ;
  assign y7606 = ~1'b0 ;
  assign y7607 = ~1'b0 ;
  assign y7608 = ~n14959 ;
  assign y7609 = ~n14961 ;
  assign y7610 = ~n14963 ;
  assign y7611 = n14965 ;
  assign y7612 = ~n14966 ;
  assign y7613 = n14967 ;
  assign y7614 = ~n14971 ;
  assign y7615 = ~1'b0 ;
  assign y7616 = n14973 ;
  assign y7617 = ~n14975 ;
  assign y7618 = ~n14977 ;
  assign y7619 = ~n14978 ;
  assign y7620 = n14981 ;
  assign y7621 = ~1'b0 ;
  assign y7622 = ~1'b0 ;
  assign y7623 = ~n8595 ;
  assign y7624 = ~1'b0 ;
  assign y7625 = n14982 ;
  assign y7626 = ~n14988 ;
  assign y7627 = ~1'b0 ;
  assign y7628 = n14990 ;
  assign y7629 = ~1'b0 ;
  assign y7630 = ~n14992 ;
  assign y7631 = ~n14993 ;
  assign y7632 = ~n14996 ;
  assign y7633 = ~n14997 ;
  assign y7634 = ~n14999 ;
  assign y7635 = ~n15001 ;
  assign y7636 = ~n15003 ;
  assign y7637 = ~1'b0 ;
  assign y7638 = ~n15010 ;
  assign y7639 = ~1'b0 ;
  assign y7640 = n15011 ;
  assign y7641 = n15014 ;
  assign y7642 = ~n15017 ;
  assign y7643 = n15021 ;
  assign y7644 = ~n15024 ;
  assign y7645 = ~1'b0 ;
  assign y7646 = n15026 ;
  assign y7647 = n15032 ;
  assign y7648 = n15035 ;
  assign y7649 = n15039 ;
  assign y7650 = n15045 ;
  assign y7651 = ~1'b0 ;
  assign y7652 = ~n15048 ;
  assign y7653 = ~n15050 ;
  assign y7654 = n15054 ;
  assign y7655 = n15055 ;
  assign y7656 = ~n15056 ;
  assign y7657 = n15062 ;
  assign y7658 = ~1'b0 ;
  assign y7659 = ~1'b0 ;
  assign y7660 = ~n15064 ;
  assign y7661 = n15070 ;
  assign y7662 = ~1'b0 ;
  assign y7663 = ~n15071 ;
  assign y7664 = n15072 ;
  assign y7665 = ~n6118 ;
  assign y7666 = ~n15075 ;
  assign y7667 = ~n15077 ;
  assign y7668 = ~n15081 ;
  assign y7669 = n15082 ;
  assign y7670 = n15083 ;
  assign y7671 = ~1'b0 ;
  assign y7672 = ~1'b0 ;
  assign y7673 = ~n15087 ;
  assign y7674 = n15088 ;
  assign y7675 = ~1'b0 ;
  assign y7676 = ~1'b0 ;
  assign y7677 = n15091 ;
  assign y7678 = n15092 ;
  assign y7679 = ~n15094 ;
  assign y7680 = ~1'b0 ;
  assign y7681 = ~n15095 ;
  assign y7682 = n15100 ;
  assign y7683 = ~n15101 ;
  assign y7684 = ~1'b0 ;
  assign y7685 = ~n15104 ;
  assign y7686 = ~1'b0 ;
  assign y7687 = ~n15113 ;
  assign y7688 = n15114 ;
  assign y7689 = ~n15118 ;
  assign y7690 = n15119 ;
  assign y7691 = ~n15120 ;
  assign y7692 = ~1'b0 ;
  assign y7693 = n15121 ;
  assign y7694 = ~n15122 ;
  assign y7695 = n15124 ;
  assign y7696 = ~n15127 ;
  assign y7697 = ~n15128 ;
  assign y7698 = n15130 ;
  assign y7699 = n15131 ;
  assign y7700 = n7370 ;
  assign y7701 = ~n15132 ;
  assign y7702 = n15133 ;
  assign y7703 = ~1'b0 ;
  assign y7704 = ~n15139 ;
  assign y7705 = n15141 ;
  assign y7706 = ~n15143 ;
  assign y7707 = ~n15144 ;
  assign y7708 = ~1'b0 ;
  assign y7709 = ~1'b0 ;
  assign y7710 = ~n15148 ;
  assign y7711 = n15151 ;
  assign y7712 = ~1'b0 ;
  assign y7713 = ~n15154 ;
  assign y7714 = n15160 ;
  assign y7715 = ~1'b0 ;
  assign y7716 = n15161 ;
  assign y7717 = ~1'b0 ;
  assign y7718 = ~n15166 ;
  assign y7719 = n15168 ;
  assign y7720 = n15170 ;
  assign y7721 = ~1'b0 ;
  assign y7722 = ~1'b0 ;
  assign y7723 = ~n2810 ;
  assign y7724 = 1'b0 ;
  assign y7725 = ~n15172 ;
  assign y7726 = ~n15177 ;
  assign y7727 = ~1'b0 ;
  assign y7728 = ~n15182 ;
  assign y7729 = ~1'b0 ;
  assign y7730 = ~n15184 ;
  assign y7731 = n15188 ;
  assign y7732 = ~n7548 ;
  assign y7733 = n15189 ;
  assign y7734 = ~n15197 ;
  assign y7735 = n13724 ;
  assign y7736 = n13698 ;
  assign y7737 = ~n15198 ;
  assign y7738 = n15200 ;
  assign y7739 = ~1'b0 ;
  assign y7740 = n15205 ;
  assign y7741 = ~1'b0 ;
  assign y7742 = ~1'b0 ;
  assign y7743 = n15207 ;
  assign y7744 = n15208 ;
  assign y7745 = ~n15212 ;
  assign y7746 = ~n15213 ;
  assign y7747 = ~1'b0 ;
  assign y7748 = 1'b0 ;
  assign y7749 = ~1'b0 ;
  assign y7750 = n15214 ;
  assign y7751 = ~n15215 ;
  assign y7752 = n409 ;
  assign y7753 = n15216 ;
  assign y7754 = ~n15217 ;
  assign y7755 = n15218 ;
  assign y7756 = ~1'b0 ;
  assign y7757 = n15220 ;
  assign y7758 = n15225 ;
  assign y7759 = ~n15226 ;
  assign y7760 = n15228 ;
  assign y7761 = ~n15231 ;
  assign y7762 = n15232 ;
  assign y7763 = ~1'b0 ;
  assign y7764 = n15234 ;
  assign y7765 = n15235 ;
  assign y7766 = n6545 ;
  assign y7767 = 1'b0 ;
  assign y7768 = n15236 ;
  assign y7769 = ~1'b0 ;
  assign y7770 = ~n4526 ;
  assign y7771 = ~n9370 ;
  assign y7772 = ~n15237 ;
  assign y7773 = ~n15241 ;
  assign y7774 = ~1'b0 ;
  assign y7775 = ~1'b0 ;
  assign y7776 = n15243 ;
  assign y7777 = n15245 ;
  assign y7778 = ~n15249 ;
  assign y7779 = ~n15251 ;
  assign y7780 = n15255 ;
  assign y7781 = n15256 ;
  assign y7782 = n15257 ;
  assign y7783 = ~1'b0 ;
  assign y7784 = ~1'b0 ;
  assign y7785 = ~n15259 ;
  assign y7786 = n15264 ;
  assign y7787 = ~n15265 ;
  assign y7788 = ~1'b0 ;
  assign y7789 = ~1'b0 ;
  assign y7790 = n9037 ;
  assign y7791 = ~1'b0 ;
  assign y7792 = ~n15268 ;
  assign y7793 = n15269 ;
  assign y7794 = ~1'b0 ;
  assign y7795 = n15271 ;
  assign y7796 = n15273 ;
  assign y7797 = n15277 ;
  assign y7798 = n15278 ;
  assign y7799 = n15285 ;
  assign y7800 = n15287 ;
  assign y7801 = n15288 ;
  assign y7802 = n15289 ;
  assign y7803 = n5603 ;
  assign y7804 = ~n15292 ;
  assign y7805 = n15295 ;
  assign y7806 = n15299 ;
  assign y7807 = ~n15304 ;
  assign y7808 = ~n15305 ;
  assign y7809 = ~1'b0 ;
  assign y7810 = ~n2409 ;
  assign y7811 = ~1'b0 ;
  assign y7812 = n15307 ;
  assign y7813 = ~n15312 ;
  assign y7814 = n15313 ;
  assign y7815 = ~1'b0 ;
  assign y7816 = ~n15317 ;
  assign y7817 = ~n15319 ;
  assign y7818 = ~n15321 ;
  assign y7819 = ~1'b0 ;
  assign y7820 = ~n15323 ;
  assign y7821 = n15325 ;
  assign y7822 = ~n7420 ;
  assign y7823 = ~n15327 ;
  assign y7824 = ~1'b0 ;
  assign y7825 = n15332 ;
  assign y7826 = n15333 ;
  assign y7827 = ~n15337 ;
  assign y7828 = ~1'b0 ;
  assign y7829 = ~1'b0 ;
  assign y7830 = ~1'b0 ;
  assign y7831 = n15346 ;
  assign y7832 = ~n15348 ;
  assign y7833 = n15350 ;
  assign y7834 = ~1'b0 ;
  assign y7835 = ~n15354 ;
  assign y7836 = n15361 ;
  assign y7837 = ~n15365 ;
  assign y7838 = n15366 ;
  assign y7839 = n4700 ;
  assign y7840 = n15367 ;
  assign y7841 = n15368 ;
  assign y7842 = n15370 ;
  assign y7843 = n15373 ;
  assign y7844 = n15374 ;
  assign y7845 = ~n15377 ;
  assign y7846 = 1'b0 ;
  assign y7847 = ~n15379 ;
  assign y7848 = ~n15380 ;
  assign y7849 = ~1'b0 ;
  assign y7850 = ~n15381 ;
  assign y7851 = ~n15384 ;
  assign y7852 = 1'b0 ;
  assign y7853 = n15386 ;
  assign y7854 = n15387 ;
  assign y7855 = ~n15388 ;
  assign y7856 = ~n15389 ;
  assign y7857 = ~n15391 ;
  assign y7858 = n15396 ;
  assign y7859 = ~1'b0 ;
  assign y7860 = ~1'b0 ;
  assign y7861 = ~n15397 ;
  assign y7862 = ~n2020 ;
  assign y7863 = ~n1819 ;
  assign y7864 = n11348 ;
  assign y7865 = n15400 ;
  assign y7866 = ~1'b0 ;
  assign y7867 = ~1'b0 ;
  assign y7868 = n15402 ;
  assign y7869 = ~n15405 ;
  assign y7870 = ~1'b0 ;
  assign y7871 = n2103 ;
  assign y7872 = ~1'b0 ;
  assign y7873 = ~1'b0 ;
  assign y7874 = n15412 ;
  assign y7875 = 1'b0 ;
  assign y7876 = ~n15417 ;
  assign y7877 = n15421 ;
  assign y7878 = ~n15425 ;
  assign y7879 = n15426 ;
  assign y7880 = ~n1487 ;
  assign y7881 = ~1'b0 ;
  assign y7882 = ~1'b0 ;
  assign y7883 = ~n15428 ;
  assign y7884 = n15432 ;
  assign y7885 = ~n9935 ;
  assign y7886 = ~n15435 ;
  assign y7887 = n5537 ;
  assign y7888 = n15437 ;
  assign y7889 = ~n5050 ;
  assign y7890 = n10216 ;
  assign y7891 = n15440 ;
  assign y7892 = ~n15442 ;
  assign y7893 = ~1'b0 ;
  assign y7894 = n15443 ;
  assign y7895 = n15444 ;
  assign y7896 = ~1'b0 ;
  assign y7897 = ~1'b0 ;
  assign y7898 = n15446 ;
  assign y7899 = n15448 ;
  assign y7900 = n13307 ;
  assign y7901 = ~1'b0 ;
  assign y7902 = n15450 ;
  assign y7903 = n15456 ;
  assign y7904 = ~n15457 ;
  assign y7905 = ~n15459 ;
  assign y7906 = ~n15460 ;
  assign y7907 = ~n15462 ;
  assign y7908 = n511 ;
  assign y7909 = ~1'b0 ;
  assign y7910 = n15463 ;
  assign y7911 = n15464 ;
  assign y7912 = n15469 ;
  assign y7913 = ~1'b0 ;
  assign y7914 = ~1'b0 ;
  assign y7915 = n15471 ;
  assign y7916 = ~n15477 ;
  assign y7917 = ~1'b0 ;
  assign y7918 = ~n15481 ;
  assign y7919 = ~1'b0 ;
  assign y7920 = ~n15482 ;
  assign y7921 = ~1'b0 ;
  assign y7922 = n15484 ;
  assign y7923 = ~n15489 ;
  assign y7924 = ~1'b0 ;
  assign y7925 = n15490 ;
  assign y7926 = ~n15495 ;
  assign y7927 = ~n15502 ;
  assign y7928 = ~1'b0 ;
  assign y7929 = n15506 ;
  assign y7930 = ~1'b0 ;
  assign y7931 = ~n15507 ;
  assign y7932 = ~n9320 ;
  assign y7933 = ~1'b0 ;
  assign y7934 = ~1'b0 ;
  assign y7935 = ~n14159 ;
  assign y7936 = n15510 ;
  assign y7937 = n15514 ;
  assign y7938 = n15515 ;
  assign y7939 = ~n15516 ;
  assign y7940 = ~n15517 ;
  assign y7941 = ~1'b0 ;
  assign y7942 = ~1'b0 ;
  assign y7943 = ~1'b0 ;
  assign y7944 = ~1'b0 ;
  assign y7945 = n15520 ;
  assign y7946 = n15521 ;
  assign y7947 = n3311 ;
  assign y7948 = n15522 ;
  assign y7949 = ~1'b0 ;
  assign y7950 = ~n15525 ;
  assign y7951 = ~n1102 ;
  assign y7952 = ~n15527 ;
  assign y7953 = ~n15528 ;
  assign y7954 = n15534 ;
  assign y7955 = n15536 ;
  assign y7956 = ~n15537 ;
  assign y7957 = ~1'b0 ;
  assign y7958 = ~1'b0 ;
  assign y7959 = ~n15538 ;
  assign y7960 = n15539 ;
  assign y7961 = ~n15540 ;
  assign y7962 = ~1'b0 ;
  assign y7963 = n15542 ;
  assign y7964 = n15549 ;
  assign y7965 = n15550 ;
  assign y7966 = 1'b0 ;
  assign y7967 = ~n15552 ;
  assign y7968 = ~n15554 ;
  assign y7969 = ~n15556 ;
  assign y7970 = 1'b0 ;
  assign y7971 = n15558 ;
  assign y7972 = ~n15560 ;
  assign y7973 = ~n7221 ;
  assign y7974 = n15564 ;
  assign y7975 = ~1'b0 ;
  assign y7976 = ~1'b0 ;
  assign y7977 = n15568 ;
  assign y7978 = n15570 ;
  assign y7979 = ~n15571 ;
  assign y7980 = ~n15572 ;
  assign y7981 = ~n15579 ;
  assign y7982 = ~1'b0 ;
  assign y7983 = ~n15583 ;
  assign y7984 = ~1'b0 ;
  assign y7985 = ~n15587 ;
  assign y7986 = ~1'b0 ;
  assign y7987 = ~n15592 ;
  assign y7988 = n15593 ;
  assign y7989 = ~n15594 ;
  assign y7990 = ~1'b0 ;
  assign y7991 = ~1'b0 ;
  assign y7992 = n15595 ;
  assign y7993 = ~1'b0 ;
  assign y7994 = n15600 ;
  assign y7995 = n15608 ;
  assign y7996 = ~n15612 ;
  assign y7997 = n15614 ;
  assign y7998 = ~1'b0 ;
  assign y7999 = ~n15615 ;
  assign y8000 = ~n15617 ;
  assign y8001 = ~1'b0 ;
  assign y8002 = ~1'b0 ;
  assign y8003 = ~n15619 ;
  assign y8004 = ~n15622 ;
  assign y8005 = n15627 ;
  assign y8006 = ~n15631 ;
  assign y8007 = ~n15636 ;
  assign y8008 = n15639 ;
  assign y8009 = ~1'b0 ;
  assign y8010 = ~n15643 ;
  assign y8011 = ~n15645 ;
  assign y8012 = n15648 ;
  assign y8013 = n5431 ;
  assign y8014 = ~n15651 ;
  assign y8015 = ~n15653 ;
  assign y8016 = ~1'b0 ;
  assign y8017 = n15658 ;
  assign y8018 = n15660 ;
  assign y8019 = ~n15661 ;
  assign y8020 = ~1'b0 ;
  assign y8021 = n15665 ;
  assign y8022 = ~1'b0 ;
  assign y8023 = n15668 ;
  assign y8024 = n15671 ;
  assign y8025 = ~n5189 ;
  assign y8026 = ~1'b0 ;
  assign y8027 = ~n15673 ;
  assign y8028 = ~1'b0 ;
  assign y8029 = ~1'b0 ;
  assign y8030 = ~n15675 ;
  assign y8031 = n15679 ;
  assign y8032 = n15682 ;
  assign y8033 = ~1'b0 ;
  assign y8034 = ~n15689 ;
  assign y8035 = ~1'b0 ;
  assign y8036 = n15691 ;
  assign y8037 = ~n15692 ;
  assign y8038 = n15694 ;
  assign y8039 = ~1'b0 ;
  assign y8040 = ~1'b0 ;
  assign y8041 = ~1'b0 ;
  assign y8042 = ~n15696 ;
  assign y8043 = ~1'b0 ;
  assign y8044 = n15699 ;
  assign y8045 = n15701 ;
  assign y8046 = n15702 ;
  assign y8047 = ~1'b0 ;
  assign y8048 = ~n15714 ;
  assign y8049 = ~n15716 ;
  assign y8050 = n15722 ;
  assign y8051 = ~n15724 ;
  assign y8052 = ~1'b0 ;
  assign y8053 = ~n15725 ;
  assign y8054 = ~1'b0 ;
  assign y8055 = ~1'b0 ;
  assign y8056 = ~1'b0 ;
  assign y8057 = n15726 ;
  assign y8058 = ~1'b0 ;
  assign y8059 = ~n5135 ;
  assign y8060 = ~1'b0 ;
  assign y8061 = n9348 ;
  assign y8062 = n15732 ;
  assign y8063 = n15733 ;
  assign y8064 = ~n15734 ;
  assign y8065 = ~n15739 ;
  assign y8066 = ~1'b0 ;
  assign y8067 = ~1'b0 ;
  assign y8068 = n15741 ;
  assign y8069 = ~n15743 ;
  assign y8070 = n15749 ;
  assign y8071 = ~n15753 ;
  assign y8072 = ~1'b0 ;
  assign y8073 = ~1'b0 ;
  assign y8074 = n7419 ;
  assign y8075 = ~1'b0 ;
  assign y8076 = ~n15757 ;
  assign y8077 = ~n15759 ;
  assign y8078 = ~1'b0 ;
  assign y8079 = n3741 ;
  assign y8080 = ~n15763 ;
  assign y8081 = ~n15764 ;
  assign y8082 = ~1'b0 ;
  assign y8083 = ~1'b0 ;
  assign y8084 = 1'b0 ;
  assign y8085 = ~n15765 ;
  assign y8086 = n15766 ;
  assign y8087 = ~1'b0 ;
  assign y8088 = ~n15767 ;
  assign y8089 = ~n15771 ;
  assign y8090 = ~1'b0 ;
  assign y8091 = ~1'b0 ;
  assign y8092 = n15772 ;
  assign y8093 = ~n15773 ;
  assign y8094 = ~1'b0 ;
  assign y8095 = ~n15774 ;
  assign y8096 = n15776 ;
  assign y8097 = ~1'b0 ;
  assign y8098 = ~n6017 ;
  assign y8099 = ~1'b0 ;
  assign y8100 = ~n15777 ;
  assign y8101 = ~1'b0 ;
  assign y8102 = ~n15778 ;
  assign y8103 = ~1'b0 ;
  assign y8104 = ~1'b0 ;
  assign y8105 = n15779 ;
  assign y8106 = n15784 ;
  assign y8107 = n15788 ;
  assign y8108 = n15791 ;
  assign y8109 = ~n15797 ;
  assign y8110 = ~n15806 ;
  assign y8111 = n15813 ;
  assign y8112 = ~n15814 ;
  assign y8113 = ~n15817 ;
  assign y8114 = n15820 ;
  assign y8115 = ~n15821 ;
  assign y8116 = ~n15822 ;
  assign y8117 = n15825 ;
  assign y8118 = n15828 ;
  assign y8119 = ~n15831 ;
  assign y8120 = ~n15833 ;
  assign y8121 = ~n15839 ;
  assign y8122 = ~n15841 ;
  assign y8123 = ~1'b0 ;
  assign y8124 = n7897 ;
  assign y8125 = n15845 ;
  assign y8126 = n15847 ;
  assign y8127 = ~1'b0 ;
  assign y8128 = ~n15853 ;
  assign y8129 = ~n15858 ;
  assign y8130 = ~n15862 ;
  assign y8131 = ~n3314 ;
  assign y8132 = n15864 ;
  assign y8133 = n15865 ;
  assign y8134 = n15869 ;
  assign y8135 = ~n5500 ;
  assign y8136 = ~n15870 ;
  assign y8137 = ~n15873 ;
  assign y8138 = ~1'b0 ;
  assign y8139 = n15876 ;
  assign y8140 = ~1'b0 ;
  assign y8141 = ~1'b0 ;
  assign y8142 = n15880 ;
  assign y8143 = n15881 ;
  assign y8144 = n15884 ;
  assign y8145 = n15885 ;
  assign y8146 = ~n15887 ;
  assign y8147 = ~n15888 ;
  assign y8148 = n15889 ;
  assign y8149 = ~n15890 ;
  assign y8150 = n15891 ;
  assign y8151 = n15900 ;
  assign y8152 = n15907 ;
  assign y8153 = ~n15908 ;
  assign y8154 = ~n15910 ;
  assign y8155 = ~n15915 ;
  assign y8156 = n5834 ;
  assign y8157 = ~n15916 ;
  assign y8158 = n15919 ;
  assign y8159 = ~n15922 ;
  assign y8160 = ~1'b0 ;
  assign y8161 = ~1'b0 ;
  assign y8162 = ~1'b0 ;
  assign y8163 = ~1'b0 ;
  assign y8164 = ~n15924 ;
  assign y8165 = ~1'b0 ;
  assign y8166 = ~n15927 ;
  assign y8167 = ~n15928 ;
  assign y8168 = ~n15930 ;
  assign y8169 = n15931 ;
  assign y8170 = ~1'b0 ;
  assign y8171 = n15934 ;
  assign y8172 = ~n15938 ;
  assign y8173 = ~n15940 ;
  assign y8174 = ~1'b0 ;
  assign y8175 = ~1'b0 ;
  assign y8176 = n15944 ;
  assign y8177 = ~1'b0 ;
  assign y8178 = ~n15947 ;
  assign y8179 = ~1'b0 ;
  assign y8180 = n15948 ;
  assign y8181 = n15950 ;
  assign y8182 = ~1'b0 ;
  assign y8183 = ~1'b0 ;
  assign y8184 = ~1'b0 ;
  assign y8185 = ~1'b0 ;
  assign y8186 = ~n8149 ;
  assign y8187 = ~n15951 ;
  assign y8188 = n10901 ;
  assign y8189 = ~n15953 ;
  assign y8190 = ~n15954 ;
  assign y8191 = n9794 ;
  assign y8192 = n15955 ;
  assign y8193 = ~1'b0 ;
  assign y8194 = ~n15957 ;
  assign y8195 = n15958 ;
  assign y8196 = n15959 ;
  assign y8197 = n15971 ;
  assign y8198 = ~1'b0 ;
  assign y8199 = ~1'b0 ;
  assign y8200 = ~1'b0 ;
  assign y8201 = ~n15972 ;
  assign y8202 = ~n15976 ;
  assign y8203 = ~n15979 ;
  assign y8204 = ~n15981 ;
  assign y8205 = ~1'b0 ;
  assign y8206 = ~1'b0 ;
  assign y8207 = ~1'b0 ;
  assign y8208 = ~n15982 ;
  assign y8209 = ~1'b0 ;
  assign y8210 = ~1'b0 ;
  assign y8211 = ~n15983 ;
  assign y8212 = ~1'b0 ;
  assign y8213 = ~n15984 ;
  assign y8214 = n15986 ;
  assign y8215 = ~n15991 ;
  assign y8216 = ~n15994 ;
  assign y8217 = ~n15998 ;
  assign y8218 = ~n15999 ;
  assign y8219 = n4024 ;
  assign y8220 = n1237 ;
  assign y8221 = ~1'b0 ;
  assign y8222 = n16003 ;
  assign y8223 = ~n16004 ;
  assign y8224 = ~1'b0 ;
  assign y8225 = n10388 ;
  assign y8226 = n16006 ;
  assign y8227 = ~n16007 ;
  assign y8228 = ~n16012 ;
  assign y8229 = ~n16018 ;
  assign y8230 = n16022 ;
  assign y8231 = ~n16023 ;
  assign y8232 = n16026 ;
  assign y8233 = ~n16039 ;
  assign y8234 = ~1'b0 ;
  assign y8235 = ~n16040 ;
  assign y8236 = ~n16044 ;
  assign y8237 = ~n16046 ;
  assign y8238 = ~1'b0 ;
  assign y8239 = ~1'b0 ;
  assign y8240 = ~1'b0 ;
  assign y8241 = ~n10163 ;
  assign y8242 = ~n16053 ;
  assign y8243 = ~1'b0 ;
  assign y8244 = ~n16054 ;
  assign y8245 = n16057 ;
  assign y8246 = ~1'b0 ;
  assign y8247 = ~1'b0 ;
  assign y8248 = ~1'b0 ;
  assign y8249 = n16059 ;
  assign y8250 = n2295 ;
  assign y8251 = ~1'b0 ;
  assign y8252 = ~1'b0 ;
  assign y8253 = n16065 ;
  assign y8254 = ~n16069 ;
  assign y8255 = n16071 ;
  assign y8256 = n16072 ;
  assign y8257 = ~n16074 ;
  assign y8258 = ~n16076 ;
  assign y8259 = ~n16077 ;
  assign y8260 = n16078 ;
  assign y8261 = ~n16082 ;
  assign y8262 = ~n16083 ;
  assign y8263 = ~n16084 ;
  assign y8264 = ~1'b0 ;
  assign y8265 = ~1'b0 ;
  assign y8266 = ~n14596 ;
  assign y8267 = ~n16087 ;
  assign y8268 = ~1'b0 ;
  assign y8269 = n16092 ;
  assign y8270 = ~n9681 ;
  assign y8271 = ~1'b0 ;
  assign y8272 = ~n16093 ;
  assign y8273 = n11706 ;
  assign y8274 = n16099 ;
  assign y8275 = ~1'b0 ;
  assign y8276 = n16102 ;
  assign y8277 = ~n16104 ;
  assign y8278 = n16106 ;
  assign y8279 = ~1'b0 ;
  assign y8280 = n16107 ;
  assign y8281 = ~n16112 ;
  assign y8282 = n16113 ;
  assign y8283 = n16115 ;
  assign y8284 = ~1'b0 ;
  assign y8285 = n16116 ;
  assign y8286 = n16118 ;
  assign y8287 = n16123 ;
  assign y8288 = ~1'b0 ;
  assign y8289 = n16125 ;
  assign y8290 = ~1'b0 ;
  assign y8291 = n16129 ;
  assign y8292 = ~n1448 ;
  assign y8293 = ~1'b0 ;
  assign y8294 = n16130 ;
  assign y8295 = n16132 ;
  assign y8296 = ~1'b0 ;
  assign y8297 = ~n16135 ;
  assign y8298 = ~1'b0 ;
  assign y8299 = ~n16140 ;
  assign y8300 = n16142 ;
  assign y8301 = ~1'b0 ;
  assign y8302 = ~n16146 ;
  assign y8303 = ~1'b0 ;
  assign y8304 = ~1'b0 ;
  assign y8305 = n16147 ;
  assign y8306 = ~n16153 ;
  assign y8307 = ~1'b0 ;
  assign y8308 = ~1'b0 ;
  assign y8309 = n16154 ;
  assign y8310 = ~1'b0 ;
  assign y8311 = n16156 ;
  assign y8312 = n16157 ;
  assign y8313 = n16158 ;
  assign y8314 = n16160 ;
  assign y8315 = ~n16162 ;
  assign y8316 = ~1'b0 ;
  assign y8317 = ~n9578 ;
  assign y8318 = n16164 ;
  assign y8319 = ~n16168 ;
  assign y8320 = ~1'b0 ;
  assign y8321 = n16170 ;
  assign y8322 = ~1'b0 ;
  assign y8323 = ~n16171 ;
  assign y8324 = ~n16174 ;
  assign y8325 = ~n16176 ;
  assign y8326 = ~n16177 ;
  assign y8327 = ~1'b0 ;
  assign y8328 = ~1'b0 ;
  assign y8329 = ~n16184 ;
  assign y8330 = n16187 ;
  assign y8331 = ~1'b0 ;
  assign y8332 = ~n16194 ;
  assign y8333 = ~n16197 ;
  assign y8334 = ~n16198 ;
  assign y8335 = ~1'b0 ;
  assign y8336 = ~1'b0 ;
  assign y8337 = n16199 ;
  assign y8338 = 1'b0 ;
  assign y8339 = ~n16200 ;
  assign y8340 = ~1'b0 ;
  assign y8341 = n16201 ;
  assign y8342 = n16204 ;
  assign y8343 = ~1'b0 ;
  assign y8344 = n16208 ;
  assign y8345 = n16210 ;
  assign y8346 = n16211 ;
  assign y8347 = ~1'b0 ;
  assign y8348 = ~1'b0 ;
  assign y8349 = n16212 ;
  assign y8350 = 1'b0 ;
  assign y8351 = n16213 ;
  assign y8352 = n16215 ;
  assign y8353 = n16218 ;
  assign y8354 = ~1'b0 ;
  assign y8355 = n16219 ;
  assign y8356 = n16221 ;
  assign y8357 = ~n5805 ;
  assign y8358 = ~1'b0 ;
  assign y8359 = ~n16225 ;
  assign y8360 = ~1'b0 ;
  assign y8361 = ~1'b0 ;
  assign y8362 = n16227 ;
  assign y8363 = ~1'b0 ;
  assign y8364 = 1'b0 ;
  assign y8365 = n16228 ;
  assign y8366 = n16233 ;
  assign y8367 = ~n6158 ;
  assign y8368 = ~n16236 ;
  assign y8369 = ~1'b0 ;
  assign y8370 = n16237 ;
  assign y8371 = ~1'b0 ;
  assign y8372 = ~1'b0 ;
  assign y8373 = ~1'b0 ;
  assign y8374 = n16238 ;
  assign y8375 = ~1'b0 ;
  assign y8376 = ~n8027 ;
  assign y8377 = ~n16242 ;
  assign y8378 = ~n16243 ;
  assign y8379 = ~1'b0 ;
  assign y8380 = n16244 ;
  assign y8381 = ~1'b0 ;
  assign y8382 = n16245 ;
  assign y8383 = ~1'b0 ;
  assign y8384 = n16247 ;
  assign y8385 = ~n16251 ;
  assign y8386 = n16252 ;
  assign y8387 = n16255 ;
  assign y8388 = ~n16256 ;
  assign y8389 = n16258 ;
  assign y8390 = n16260 ;
  assign y8391 = n10080 ;
  assign y8392 = n16261 ;
  assign y8393 = ~n16265 ;
  assign y8394 = ~1'b0 ;
  assign y8395 = ~n16270 ;
  assign y8396 = n16272 ;
  assign y8397 = ~1'b0 ;
  assign y8398 = ~n16275 ;
  assign y8399 = ~n16278 ;
  assign y8400 = n15113 ;
  assign y8401 = ~1'b0 ;
  assign y8402 = n16280 ;
  assign y8403 = n16282 ;
  assign y8404 = ~n16285 ;
  assign y8405 = n16289 ;
  assign y8406 = ~n16293 ;
  assign y8407 = ~n16294 ;
  assign y8408 = ~n16300 ;
  assign y8409 = n16301 ;
  assign y8410 = ~1'b0 ;
  assign y8411 = ~n16302 ;
  assign y8412 = ~n16306 ;
  assign y8413 = n16307 ;
  assign y8414 = ~1'b0 ;
  assign y8415 = ~n16309 ;
  assign y8416 = n16310 ;
  assign y8417 = n16311 ;
  assign y8418 = ~1'b0 ;
  assign y8419 = ~n16312 ;
  assign y8420 = ~1'b0 ;
  assign y8421 = ~n16318 ;
  assign y8422 = ~n16320 ;
  assign y8423 = ~1'b0 ;
  assign y8424 = ~1'b0 ;
  assign y8425 = ~1'b0 ;
  assign y8426 = n16322 ;
  assign y8427 = ~1'b0 ;
  assign y8428 = n16329 ;
  assign y8429 = n16335 ;
  assign y8430 = ~n16338 ;
  assign y8431 = ~n16346 ;
  assign y8432 = ~n16347 ;
  assign y8433 = n16349 ;
  assign y8434 = n16350 ;
  assign y8435 = ~1'b0 ;
  assign y8436 = ~1'b0 ;
  assign y8437 = ~n16352 ;
  assign y8438 = ~n16353 ;
  assign y8439 = n16356 ;
  assign y8440 = ~n16360 ;
  assign y8441 = ~n16361 ;
  assign y8442 = ~1'b0 ;
  assign y8443 = ~n16366 ;
  assign y8444 = 1'b0 ;
  assign y8445 = ~n16367 ;
  assign y8446 = ~1'b0 ;
  assign y8447 = n16368 ;
  assign y8448 = n16369 ;
  assign y8449 = n16370 ;
  assign y8450 = ~n16371 ;
  assign y8451 = ~n16372 ;
  assign y8452 = 1'b0 ;
  assign y8453 = ~1'b0 ;
  assign y8454 = ~1'b0 ;
  assign y8455 = ~1'b0 ;
  assign y8456 = ~1'b0 ;
  assign y8457 = ~n16373 ;
  assign y8458 = ~n16375 ;
  assign y8459 = n16378 ;
  assign y8460 = n9410 ;
  assign y8461 = n16379 ;
  assign y8462 = ~1'b0 ;
  assign y8463 = ~n16381 ;
  assign y8464 = n16382 ;
  assign y8465 = n16385 ;
  assign y8466 = n3190 ;
  assign y8467 = n16386 ;
  assign y8468 = ~1'b0 ;
  assign y8469 = ~n16388 ;
  assign y8470 = ~n16390 ;
  assign y8471 = n16391 ;
  assign y8472 = n16392 ;
  assign y8473 = n6263 ;
  assign y8474 = n16393 ;
  assign y8475 = ~1'b0 ;
  assign y8476 = ~1'b0 ;
  assign y8477 = ~n16394 ;
  assign y8478 = ~1'b0 ;
  assign y8479 = ~n16399 ;
  assign y8480 = ~n16400 ;
  assign y8481 = n16401 ;
  assign y8482 = ~n16402 ;
  assign y8483 = n16404 ;
  assign y8484 = ~n16410 ;
  assign y8485 = ~n16414 ;
  assign y8486 = n16417 ;
  assign y8487 = ~1'b0 ;
  assign y8488 = n16418 ;
  assign y8489 = ~n16419 ;
  assign y8490 = ~n16420 ;
  assign y8491 = ~1'b0 ;
  assign y8492 = n11178 ;
  assign y8493 = ~n16423 ;
  assign y8494 = n16425 ;
  assign y8495 = ~n16427 ;
  assign y8496 = ~n16428 ;
  assign y8497 = ~1'b0 ;
  assign y8498 = ~1'b0 ;
  assign y8499 = ~1'b0 ;
  assign y8500 = ~n16429 ;
  assign y8501 = ~n16430 ;
  assign y8502 = ~n16436 ;
  assign y8503 = ~n16437 ;
  assign y8504 = n16438 ;
  assign y8505 = n16440 ;
  assign y8506 = ~1'b0 ;
  assign y8507 = n16441 ;
  assign y8508 = n16442 ;
  assign y8509 = ~n16443 ;
  assign y8510 = ~1'b0 ;
  assign y8511 = n16451 ;
  assign y8512 = ~n16453 ;
  assign y8513 = ~1'b0 ;
  assign y8514 = ~1'b0 ;
  assign y8515 = ~1'b0 ;
  assign y8516 = ~1'b0 ;
  assign y8517 = n16455 ;
  assign y8518 = ~n16460 ;
  assign y8519 = ~1'b0 ;
  assign y8520 = n16464 ;
  assign y8521 = n16465 ;
  assign y8522 = ~1'b0 ;
  assign y8523 = ~n16472 ;
  assign y8524 = n16474 ;
  assign y8525 = ~1'b0 ;
  assign y8526 = ~n11414 ;
  assign y8527 = n16475 ;
  assign y8528 = n16480 ;
  assign y8529 = ~n16484 ;
  assign y8530 = n16487 ;
  assign y8531 = n16488 ;
  assign y8532 = n16489 ;
  assign y8533 = ~1'b0 ;
  assign y8534 = ~1'b0 ;
  assign y8535 = ~1'b0 ;
  assign y8536 = ~n16490 ;
  assign y8537 = ~1'b0 ;
  assign y8538 = ~n16491 ;
  assign y8539 = ~n16492 ;
  assign y8540 = ~1'b0 ;
  assign y8541 = n16498 ;
  assign y8542 = n16499 ;
  assign y8543 = ~n16501 ;
  assign y8544 = ~n16502 ;
  assign y8545 = n16506 ;
  assign y8546 = ~n16508 ;
  assign y8547 = ~n16509 ;
  assign y8548 = n16514 ;
  assign y8549 = ~1'b0 ;
  assign y8550 = ~n16515 ;
  assign y8551 = ~1'b0 ;
  assign y8552 = ~n16517 ;
  assign y8553 = ~n16519 ;
  assign y8554 = n16521 ;
  assign y8555 = ~1'b0 ;
  assign y8556 = ~1'b0 ;
  assign y8557 = n16523 ;
  assign y8558 = ~n16526 ;
  assign y8559 = ~n16527 ;
  assign y8560 = n16528 ;
  assign y8561 = ~n16530 ;
  assign y8562 = ~1'b0 ;
  assign y8563 = ~n16533 ;
  assign y8564 = ~1'b0 ;
  assign y8565 = ~n16537 ;
  assign y8566 = ~1'b0 ;
  assign y8567 = ~n16541 ;
  assign y8568 = ~1'b0 ;
  assign y8569 = n16542 ;
  assign y8570 = ~1'b0 ;
  assign y8571 = ~1'b0 ;
  assign y8572 = ~n16543 ;
  assign y8573 = ~n16545 ;
  assign y8574 = ~n13293 ;
  assign y8575 = n16547 ;
  assign y8576 = ~n16549 ;
  assign y8577 = ~1'b0 ;
  assign y8578 = ~1'b0 ;
  assign y8579 = n16550 ;
  assign y8580 = n16554 ;
  assign y8581 = ~n1444 ;
  assign y8582 = 1'b0 ;
  assign y8583 = ~1'b0 ;
  assign y8584 = ~1'b0 ;
  assign y8585 = ~1'b0 ;
  assign y8586 = ~1'b0 ;
  assign y8587 = n15035 ;
  assign y8588 = n16555 ;
  assign y8589 = ~n16557 ;
  assign y8590 = n16560 ;
  assign y8591 = ~n9068 ;
  assign y8592 = ~n16562 ;
  assign y8593 = n16563 ;
  assign y8594 = n16567 ;
  assign y8595 = 1'b0 ;
  assign y8596 = ~n16568 ;
  assign y8597 = ~1'b0 ;
  assign y8598 = ~n16569 ;
  assign y8599 = n16572 ;
  assign y8600 = ~1'b0 ;
  assign y8601 = ~1'b0 ;
  assign y8602 = n1330 ;
  assign y8603 = ~1'b0 ;
  assign y8604 = ~n16575 ;
  assign y8605 = ~n16578 ;
  assign y8606 = n16580 ;
  assign y8607 = ~1'b0 ;
  assign y8608 = ~n10842 ;
  assign y8609 = n16582 ;
  assign y8610 = n16583 ;
  assign y8611 = n16590 ;
  assign y8612 = ~n16592 ;
  assign y8613 = ~n16595 ;
  assign y8614 = ~1'b0 ;
  assign y8615 = n16596 ;
  assign y8616 = 1'b0 ;
  assign y8617 = n16598 ;
  assign y8618 = ~n16601 ;
  assign y8619 = ~n16602 ;
  assign y8620 = ~n16603 ;
  assign y8621 = ~n16605 ;
  assign y8622 = ~1'b0 ;
  assign y8623 = ~n16610 ;
  assign y8624 = ~1'b0 ;
  assign y8625 = ~1'b0 ;
  assign y8626 = n2289 ;
  assign y8627 = ~n16614 ;
  assign y8628 = n16615 ;
  assign y8629 = ~n16617 ;
  assign y8630 = ~1'b0 ;
  assign y8631 = n16620 ;
  assign y8632 = n16623 ;
  assign y8633 = ~1'b0 ;
  assign y8634 = ~n16624 ;
  assign y8635 = 1'b0 ;
  assign y8636 = ~1'b0 ;
  assign y8637 = ~1'b0 ;
  assign y8638 = ~1'b0 ;
  assign y8639 = ~n16626 ;
  assign y8640 = n16627 ;
  assign y8641 = n175 ;
  assign y8642 = ~n16633 ;
  assign y8643 = n16635 ;
  assign y8644 = 1'b0 ;
  assign y8645 = ~1'b0 ;
  assign y8646 = ~n16636 ;
  assign y8647 = n16638 ;
  assign y8648 = 1'b0 ;
  assign y8649 = ~1'b0 ;
  assign y8650 = n16641 ;
  assign y8651 = ~n16643 ;
  assign y8652 = ~1'b0 ;
  assign y8653 = n16644 ;
  assign y8654 = ~n16650 ;
  assign y8655 = ~n195 ;
  assign y8656 = n16652 ;
  assign y8657 = ~n16656 ;
  assign y8658 = ~1'b0 ;
  assign y8659 = ~1'b0 ;
  assign y8660 = ~n16660 ;
  assign y8661 = ~n16664 ;
  assign y8662 = n16665 ;
  assign y8663 = ~1'b0 ;
  assign y8664 = ~1'b0 ;
  assign y8665 = n8187 ;
  assign y8666 = n16669 ;
  assign y8667 = ~n16671 ;
  assign y8668 = n16682 ;
  assign y8669 = ~1'b0 ;
  assign y8670 = n16685 ;
  assign y8671 = ~n16687 ;
  assign y8672 = ~n6997 ;
  assign y8673 = ~n16693 ;
  assign y8674 = n16696 ;
  assign y8675 = ~1'b0 ;
  assign y8676 = ~1'b0 ;
  assign y8677 = n16703 ;
  assign y8678 = ~n16705 ;
  assign y8679 = n16707 ;
  assign y8680 = ~n16708 ;
  assign y8681 = n16709 ;
  assign y8682 = ~1'b0 ;
  assign y8683 = ~1'b0 ;
  assign y8684 = ~1'b0 ;
  assign y8685 = ~1'b0 ;
  assign y8686 = ~1'b0 ;
  assign y8687 = ~1'b0 ;
  assign y8688 = ~n16710 ;
  assign y8689 = ~n16711 ;
  assign y8690 = n16716 ;
  assign y8691 = n16727 ;
  assign y8692 = ~1'b0 ;
  assign y8693 = ~n16733 ;
  assign y8694 = n9242 ;
  assign y8695 = ~n16737 ;
  assign y8696 = ~1'b0 ;
  assign y8697 = ~1'b0 ;
  assign y8698 = n16739 ;
  assign y8699 = ~1'b0 ;
  assign y8700 = n16740 ;
  assign y8701 = ~n16751 ;
  assign y8702 = ~n16753 ;
  assign y8703 = n16757 ;
  assign y8704 = n16760 ;
  assign y8705 = n16762 ;
  assign y8706 = n16764 ;
  assign y8707 = ~n16765 ;
  assign y8708 = ~n16766 ;
  assign y8709 = ~1'b0 ;
  assign y8710 = ~1'b0 ;
  assign y8711 = ~1'b0 ;
  assign y8712 = n16767 ;
  assign y8713 = ~n16770 ;
  assign y8714 = ~1'b0 ;
  assign y8715 = ~1'b0 ;
  assign y8716 = ~1'b0 ;
  assign y8717 = ~n3257 ;
  assign y8718 = ~n16777 ;
  assign y8719 = ~1'b0 ;
  assign y8720 = ~1'b0 ;
  assign y8721 = ~n16782 ;
  assign y8722 = ~n16785 ;
  assign y8723 = n16786 ;
  assign y8724 = n16790 ;
  assign y8725 = ~n16791 ;
  assign y8726 = ~n16680 ;
  assign y8727 = n16795 ;
  assign y8728 = ~1'b0 ;
  assign y8729 = ~1'b0 ;
  assign y8730 = ~1'b0 ;
  assign y8731 = ~n16798 ;
  assign y8732 = n16801 ;
  assign y8733 = ~n16802 ;
  assign y8734 = ~1'b0 ;
  assign y8735 = ~n14684 ;
  assign y8736 = ~1'b0 ;
  assign y8737 = ~n16804 ;
  assign y8738 = n16808 ;
  assign y8739 = n16809 ;
  assign y8740 = ~n16811 ;
  assign y8741 = n16812 ;
  assign y8742 = ~n16815 ;
  assign y8743 = n16818 ;
  assign y8744 = ~n632 ;
  assign y8745 = ~n16821 ;
  assign y8746 = ~1'b0 ;
  assign y8747 = ~n16822 ;
  assign y8748 = n16823 ;
  assign y8749 = ~n16829 ;
  assign y8750 = n16840 ;
  assign y8751 = n16841 ;
  assign y8752 = ~n16843 ;
  assign y8753 = n16844 ;
  assign y8754 = n16847 ;
  assign y8755 = ~n16848 ;
  assign y8756 = ~n2774 ;
  assign y8757 = n9663 ;
  assign y8758 = n16849 ;
  assign y8759 = ~n16852 ;
  assign y8760 = n16854 ;
  assign y8761 = ~n12087 ;
  assign y8762 = ~n16855 ;
  assign y8763 = n16856 ;
  assign y8764 = ~1'b0 ;
  assign y8765 = ~n16857 ;
  assign y8766 = ~1'b0 ;
  assign y8767 = n16861 ;
  assign y8768 = ~n16862 ;
  assign y8769 = n16864 ;
  assign y8770 = n16866 ;
  assign y8771 = ~1'b0 ;
  assign y8772 = n16870 ;
  assign y8773 = n16873 ;
  assign y8774 = ~n16874 ;
  assign y8775 = ~1'b0 ;
  assign y8776 = n16875 ;
  assign y8777 = n16877 ;
  assign y8778 = n16882 ;
  assign y8779 = n16883 ;
  assign y8780 = n16891 ;
  assign y8781 = n16896 ;
  assign y8782 = ~n16898 ;
  assign y8783 = n16901 ;
  assign y8784 = ~n16911 ;
  assign y8785 = n16917 ;
  assign y8786 = ~n16920 ;
  assign y8787 = n16922 ;
  assign y8788 = ~1'b0 ;
  assign y8789 = ~n16924 ;
  assign y8790 = ~n16929 ;
  assign y8791 = ~n16930 ;
  assign y8792 = ~n16934 ;
  assign y8793 = ~1'b0 ;
  assign y8794 = ~n16936 ;
  assign y8795 = n16937 ;
  assign y8796 = ~n16366 ;
  assign y8797 = 1'b0 ;
  assign y8798 = ~n16938 ;
  assign y8799 = n2613 ;
  assign y8800 = ~1'b0 ;
  assign y8801 = n16940 ;
  assign y8802 = n16944 ;
  assign y8803 = n16946 ;
  assign y8804 = ~n16948 ;
  assign y8805 = ~1'b0 ;
  assign y8806 = ~1'b0 ;
  assign y8807 = ~n16950 ;
  assign y8808 = ~n16952 ;
  assign y8809 = ~n16953 ;
  assign y8810 = n16954 ;
  assign y8811 = ~n16958 ;
  assign y8812 = ~1'b0 ;
  assign y8813 = n16959 ;
  assign y8814 = n16960 ;
  assign y8815 = ~n16961 ;
  assign y8816 = ~n16966 ;
  assign y8817 = ~n16968 ;
  assign y8818 = ~1'b0 ;
  assign y8819 = n16972 ;
  assign y8820 = ~n16979 ;
  assign y8821 = n16983 ;
  assign y8822 = ~n16984 ;
  assign y8823 = ~1'b0 ;
  assign y8824 = n16985 ;
  assign y8825 = ~n16987 ;
  assign y8826 = ~n16988 ;
  assign y8827 = ~n16989 ;
  assign y8828 = ~n16991 ;
  assign y8829 = ~1'b0 ;
  assign y8830 = ~n16994 ;
  assign y8831 = n16995 ;
  assign y8832 = ~n16998 ;
  assign y8833 = ~n17000 ;
  assign y8834 = ~n17001 ;
  assign y8835 = ~1'b0 ;
  assign y8836 = ~n17004 ;
  assign y8837 = ~n17008 ;
  assign y8838 = ~1'b0 ;
  assign y8839 = ~n17010 ;
  assign y8840 = ~n17021 ;
  assign y8841 = ~n17026 ;
  assign y8842 = ~1'b0 ;
  assign y8843 = ~n17027 ;
  assign y8844 = n17032 ;
  assign y8845 = n17035 ;
  assign y8846 = ~1'b0 ;
  assign y8847 = n17037 ;
  assign y8848 = ~n17041 ;
  assign y8849 = n17043 ;
  assign y8850 = ~n17048 ;
  assign y8851 = ~1'b0 ;
  assign y8852 = ~n17054 ;
  assign y8853 = n17055 ;
  assign y8854 = 1'b0 ;
  assign y8855 = ~n17063 ;
  assign y8856 = n17068 ;
  assign y8857 = ~1'b0 ;
  assign y8858 = n17070 ;
  assign y8859 = ~n17078 ;
  assign y8860 = n17081 ;
  assign y8861 = n17084 ;
  assign y8862 = ~1'b0 ;
  assign y8863 = ~n17087 ;
  assign y8864 = ~1'b0 ;
  assign y8865 = ~1'b0 ;
  assign y8866 = ~n17090 ;
  assign y8867 = n17091 ;
  assign y8868 = 1'b0 ;
  assign y8869 = n17098 ;
  assign y8870 = ~n17102 ;
  assign y8871 = 1'b0 ;
  assign y8872 = ~n17104 ;
  assign y8873 = ~1'b0 ;
  assign y8874 = n17106 ;
  assign y8875 = ~n17110 ;
  assign y8876 = n17111 ;
  assign y8877 = ~n17117 ;
  assign y8878 = n7762 ;
  assign y8879 = ~1'b0 ;
  assign y8880 = n17118 ;
  assign y8881 = n17119 ;
  assign y8882 = n17123 ;
  assign y8883 = ~n17124 ;
  assign y8884 = ~n17125 ;
  assign y8885 = n17128 ;
  assign y8886 = n17129 ;
  assign y8887 = ~1'b0 ;
  assign y8888 = ~n17131 ;
  assign y8889 = n17138 ;
  assign y8890 = ~n17141 ;
  assign y8891 = n4562 ;
  assign y8892 = ~n17142 ;
  assign y8893 = ~1'b0 ;
  assign y8894 = ~n17144 ;
  assign y8895 = n17145 ;
  assign y8896 = ~n17148 ;
  assign y8897 = ~n17151 ;
  assign y8898 = n17152 ;
  assign y8899 = n17157 ;
  assign y8900 = n17158 ;
  assign y8901 = ~n17160 ;
  assign y8902 = ~n17161 ;
  assign y8903 = n17167 ;
  assign y8904 = ~1'b0 ;
  assign y8905 = n4884 ;
  assign y8906 = ~n17169 ;
  assign y8907 = ~1'b0 ;
  assign y8908 = n17171 ;
  assign y8909 = n8085 ;
  assign y8910 = n3540 ;
  assign y8911 = ~1'b0 ;
  assign y8912 = ~n17174 ;
  assign y8913 = ~1'b0 ;
  assign y8914 = n17178 ;
  assign y8915 = ~n17180 ;
  assign y8916 = ~1'b0 ;
  assign y8917 = ~n17182 ;
  assign y8918 = ~n13785 ;
  assign y8919 = ~n6368 ;
  assign y8920 = ~n17188 ;
  assign y8921 = ~n17189 ;
  assign y8922 = ~1'b0 ;
  assign y8923 = ~1'b0 ;
  assign y8924 = ~n17192 ;
  assign y8925 = ~1'b0 ;
  assign y8926 = ~n17194 ;
  assign y8927 = ~n5111 ;
  assign y8928 = n17196 ;
  assign y8929 = ~n17198 ;
  assign y8930 = ~n17202 ;
  assign y8931 = n17203 ;
  assign y8932 = ~n17204 ;
  assign y8933 = ~1'b0 ;
  assign y8934 = n17209 ;
  assign y8935 = ~n17210 ;
  assign y8936 = ~n17212 ;
  assign y8937 = ~n17216 ;
  assign y8938 = ~n17221 ;
  assign y8939 = ~n17223 ;
  assign y8940 = ~n17232 ;
  assign y8941 = ~n17234 ;
  assign y8942 = n17236 ;
  assign y8943 = ~1'b0 ;
  assign y8944 = ~n17238 ;
  assign y8945 = n17240 ;
  assign y8946 = ~n17246 ;
  assign y8947 = ~n17254 ;
  assign y8948 = ~n10235 ;
  assign y8949 = ~n17255 ;
  assign y8950 = ~1'b0 ;
  assign y8951 = ~n17256 ;
  assign y8952 = n17257 ;
  assign y8953 = ~n17262 ;
  assign y8954 = n17265 ;
  assign y8955 = ~n17269 ;
  assign y8956 = 1'b0 ;
  assign y8957 = n17272 ;
  assign y8958 = 1'b0 ;
  assign y8959 = n17273 ;
  assign y8960 = ~n17274 ;
  assign y8961 = ~n17277 ;
  assign y8962 = n17281 ;
  assign y8963 = ~n17285 ;
  assign y8964 = ~n17287 ;
  assign y8965 = ~1'b0 ;
  assign y8966 = ~1'b0 ;
  assign y8967 = ~n17289 ;
  assign y8968 = ~n17292 ;
  assign y8969 = ~n17294 ;
  assign y8970 = ~n17295 ;
  assign y8971 = 1'b0 ;
  assign y8972 = n17297 ;
  assign y8973 = ~1'b0 ;
  assign y8974 = n17302 ;
  assign y8975 = n17304 ;
  assign y8976 = ~n17306 ;
  assign y8977 = n17307 ;
  assign y8978 = ~1'b0 ;
  assign y8979 = ~1'b0 ;
  assign y8980 = ~1'b0 ;
  assign y8981 = n17308 ;
  assign y8982 = n17312 ;
  assign y8983 = ~1'b0 ;
  assign y8984 = ~1'b0 ;
  assign y8985 = ~n17316 ;
  assign y8986 = ~1'b0 ;
  assign y8987 = ~1'b0 ;
  assign y8988 = ~n17324 ;
  assign y8989 = ~1'b0 ;
  assign y8990 = ~n17329 ;
  assign y8991 = n17333 ;
  assign y8992 = ~n17335 ;
  assign y8993 = n17339 ;
  assign y8994 = n17341 ;
  assign y8995 = ~n17342 ;
  assign y8996 = ~n17344 ;
  assign y8997 = ~n17345 ;
  assign y8998 = ~n17346 ;
  assign y8999 = ~n17348 ;
  assign y9000 = n14801 ;
  assign y9001 = ~1'b0 ;
  assign y9002 = n17354 ;
  assign y9003 = ~n17360 ;
  assign y9004 = ~n17361 ;
  assign y9005 = n17363 ;
  assign y9006 = n17364 ;
  assign y9007 = n17370 ;
  assign y9008 = n17371 ;
  assign y9009 = n17372 ;
  assign y9010 = ~n17374 ;
  assign y9011 = ~1'b0 ;
  assign y9012 = ~1'b0 ;
  assign y9013 = ~n17375 ;
  assign y9014 = n17378 ;
  assign y9015 = n17379 ;
  assign y9016 = n17380 ;
  assign y9017 = ~n17382 ;
  assign y9018 = ~n17386 ;
  assign y9019 = ~n17388 ;
  assign y9020 = ~1'b0 ;
  assign y9021 = ~1'b0 ;
  assign y9022 = n11292 ;
  assign y9023 = n17391 ;
  assign y9024 = n17392 ;
  assign y9025 = ~1'b0 ;
  assign y9026 = ~n17394 ;
  assign y9027 = ~n17396 ;
  assign y9028 = ~n17398 ;
  assign y9029 = ~n17402 ;
  assign y9030 = ~n17409 ;
  assign y9031 = ~n17411 ;
  assign y9032 = ~n17414 ;
  assign y9033 = ~1'b0 ;
  assign y9034 = ~n17418 ;
  assign y9035 = ~n17419 ;
  assign y9036 = ~1'b0 ;
  assign y9037 = ~1'b0 ;
  assign y9038 = 1'b0 ;
  assign y9039 = n17424 ;
  assign y9040 = n17425 ;
  assign y9041 = ~1'b0 ;
  assign y9042 = ~1'b0 ;
  assign y9043 = ~1'b0 ;
  assign y9044 = ~1'b0 ;
  assign y9045 = ~1'b0 ;
  assign y9046 = ~1'b0 ;
  assign y9047 = n560 ;
  assign y9048 = ~1'b0 ;
  assign y9049 = ~1'b0 ;
  assign y9050 = ~n17427 ;
  assign y9051 = n17431 ;
  assign y9052 = ~1'b0 ;
  assign y9053 = ~n17434 ;
  assign y9054 = ~1'b0 ;
  assign y9055 = ~n17435 ;
  assign y9056 = n17436 ;
  assign y9057 = n17439 ;
  assign y9058 = n17441 ;
  assign y9059 = 1'b0 ;
  assign y9060 = n17446 ;
  assign y9061 = ~n17447 ;
  assign y9062 = ~1'b0 ;
  assign y9063 = n8496 ;
  assign y9064 = n17448 ;
  assign y9065 = n17450 ;
  assign y9066 = ~n17453 ;
  assign y9067 = ~1'b0 ;
  assign y9068 = n17460 ;
  assign y9069 = n17461 ;
  assign y9070 = n17462 ;
  assign y9071 = ~n17463 ;
  assign y9072 = ~n17467 ;
  assign y9073 = n17468 ;
  assign y9074 = n17473 ;
  assign y9075 = ~n17478 ;
  assign y9076 = 1'b0 ;
  assign y9077 = ~1'b0 ;
  assign y9078 = ~1'b0 ;
  assign y9079 = ~1'b0 ;
  assign y9080 = ~n17479 ;
  assign y9081 = ~n17480 ;
  assign y9082 = ~n17481 ;
  assign y9083 = 1'b0 ;
  assign y9084 = ~1'b0 ;
  assign y9085 = n17483 ;
  assign y9086 = ~1'b0 ;
  assign y9087 = ~n17485 ;
  assign y9088 = ~n17488 ;
  assign y9089 = n17491 ;
  assign y9090 = ~1'b0 ;
  assign y9091 = n17493 ;
  assign y9092 = ~1'b0 ;
  assign y9093 = n5300 ;
  assign y9094 = ~1'b0 ;
  assign y9095 = ~1'b0 ;
  assign y9096 = n17495 ;
  assign y9097 = ~n17496 ;
  assign y9098 = ~n17497 ;
  assign y9099 = ~n13202 ;
  assign y9100 = n17499 ;
  assign y9101 = ~n17500 ;
  assign y9102 = n1761 ;
  assign y9103 = ~n17506 ;
  assign y9104 = ~1'b0 ;
  assign y9105 = ~n17508 ;
  assign y9106 = ~1'b0 ;
  assign y9107 = ~n17511 ;
  assign y9108 = ~n17512 ;
  assign y9109 = n17513 ;
  assign y9110 = ~1'b0 ;
  assign y9111 = ~n17516 ;
  assign y9112 = n11243 ;
  assign y9113 = ~1'b0 ;
  assign y9114 = ~1'b0 ;
  assign y9115 = 1'b0 ;
  assign y9116 = 1'b0 ;
  assign y9117 = ~n17519 ;
  assign y9118 = n17520 ;
  assign y9119 = ~n611 ;
  assign y9120 = ~n17522 ;
  assign y9121 = ~1'b0 ;
  assign y9122 = n17523 ;
  assign y9123 = ~n17524 ;
  assign y9124 = ~n17525 ;
  assign y9125 = ~n17527 ;
  assign y9126 = n17528 ;
  assign y9127 = ~1'b0 ;
  assign y9128 = 1'b0 ;
  assign y9129 = ~n17529 ;
  assign y9130 = n17530 ;
  assign y9131 = ~n17536 ;
  assign y9132 = ~1'b0 ;
  assign y9133 = n17538 ;
  assign y9134 = n17539 ;
  assign y9135 = ~1'b0 ;
  assign y9136 = n17543 ;
  assign y9137 = ~1'b0 ;
  assign y9138 = ~1'b0 ;
  assign y9139 = ~1'b0 ;
  assign y9140 = ~1'b0 ;
  assign y9141 = ~n17544 ;
  assign y9142 = n17550 ;
  assign y9143 = n17555 ;
  assign y9144 = ~1'b0 ;
  assign y9145 = ~1'b0 ;
  assign y9146 = ~1'b0 ;
  assign y9147 = ~n17556 ;
  assign y9148 = n17558 ;
  assign y9149 = ~1'b0 ;
  assign y9150 = n17560 ;
  assign y9151 = n17562 ;
  assign y9152 = n853 ;
  assign y9153 = n17567 ;
  assign y9154 = n17568 ;
  assign y9155 = ~n17570 ;
  assign y9156 = ~n17572 ;
  assign y9157 = ~n17574 ;
  assign y9158 = ~n7535 ;
  assign y9159 = ~n6323 ;
  assign y9160 = ~n17576 ;
  assign y9161 = ~n17578 ;
  assign y9162 = n17581 ;
  assign y9163 = n17582 ;
  assign y9164 = ~n17583 ;
  assign y9165 = ~n17587 ;
  assign y9166 = ~1'b0 ;
  assign y9167 = ~n17589 ;
  assign y9168 = n17593 ;
  assign y9169 = ~n17594 ;
  assign y9170 = n17596 ;
  assign y9171 = ~1'b0 ;
  assign y9172 = ~n17598 ;
  assign y9173 = ~n17599 ;
  assign y9174 = ~n17601 ;
  assign y9175 = n17602 ;
  assign y9176 = n17603 ;
  assign y9177 = ~n17604 ;
  assign y9178 = n17607 ;
  assign y9179 = 1'b0 ;
  assign y9180 = ~n17612 ;
  assign y9181 = n17613 ;
  assign y9182 = ~n17614 ;
  assign y9183 = n17615 ;
  assign y9184 = ~1'b0 ;
  assign y9185 = n17617 ;
  assign y9186 = n17618 ;
  assign y9187 = ~n14321 ;
  assign y9188 = n4308 ;
  assign y9189 = n17619 ;
  assign y9190 = 1'b0 ;
  assign y9191 = ~1'b0 ;
  assign y9192 = ~n17623 ;
  assign y9193 = ~n17625 ;
  assign y9194 = ~n7568 ;
  assign y9195 = ~n17628 ;
  assign y9196 = n11474 ;
  assign y9197 = ~1'b0 ;
  assign y9198 = 1'b0 ;
  assign y9199 = ~1'b0 ;
  assign y9200 = ~n17630 ;
  assign y9201 = n17631 ;
  assign y9202 = n17632 ;
  assign y9203 = ~n17634 ;
  assign y9204 = n17643 ;
  assign y9205 = ~1'b0 ;
  assign y9206 = 1'b0 ;
  assign y9207 = ~n17644 ;
  assign y9208 = n17646 ;
  assign y9209 = ~n17647 ;
  assign y9210 = ~n17648 ;
  assign y9211 = ~n17654 ;
  assign y9212 = ~n17656 ;
  assign y9213 = ~n17660 ;
  assign y9214 = ~1'b0 ;
  assign y9215 = ~n17661 ;
  assign y9216 = n17662 ;
  assign y9217 = ~1'b0 ;
  assign y9218 = ~1'b0 ;
  assign y9219 = n17664 ;
  assign y9220 = n5080 ;
  assign y9221 = ~1'b0 ;
  assign y9222 = ~1'b0 ;
  assign y9223 = n17667 ;
  assign y9224 = ~n17670 ;
  assign y9225 = n17673 ;
  assign y9226 = ~1'b0 ;
  assign y9227 = ~1'b0 ;
  assign y9228 = n17683 ;
  assign y9229 = n17685 ;
  assign y9230 = ~n17687 ;
  assign y9231 = ~1'b0 ;
  assign y9232 = n17688 ;
  assign y9233 = ~1'b0 ;
  assign y9234 = ~1'b0 ;
  assign y9235 = n17690 ;
  assign y9236 = n709 ;
  assign y9237 = ~n17692 ;
  assign y9238 = ~n17702 ;
  assign y9239 = n17706 ;
  assign y9240 = ~n1853 ;
  assign y9241 = n17711 ;
  assign y9242 = ~n17715 ;
  assign y9243 = n17717 ;
  assign y9244 = n17718 ;
  assign y9245 = ~n17719 ;
  assign y9246 = n17720 ;
  assign y9247 = n17722 ;
  assign y9248 = ~n17726 ;
  assign y9249 = ~n17727 ;
  assign y9250 = n17728 ;
  assign y9251 = n17733 ;
  assign y9252 = ~n17736 ;
  assign y9253 = ~1'b0 ;
  assign y9254 = n17741 ;
  assign y9255 = ~1'b0 ;
  assign y9256 = n17747 ;
  assign y9257 = ~n17748 ;
  assign y9258 = ~1'b0 ;
  assign y9259 = n17749 ;
  assign y9260 = ~1'b0 ;
  assign y9261 = ~1'b0 ;
  assign y9262 = ~n17753 ;
  assign y9263 = n17757 ;
  assign y9264 = n17759 ;
  assign y9265 = n17761 ;
  assign y9266 = ~n17763 ;
  assign y9267 = ~1'b0 ;
  assign y9268 = ~1'b0 ;
  assign y9269 = 1'b0 ;
  assign y9270 = ~1'b0 ;
  assign y9271 = ~n17765 ;
  assign y9272 = n17766 ;
  assign y9273 = ~n17773 ;
  assign y9274 = ~n17776 ;
  assign y9275 = ~n17777 ;
  assign y9276 = ~1'b0 ;
  assign y9277 = n17780 ;
  assign y9278 = ~n17783 ;
  assign y9279 = n17784 ;
  assign y9280 = ~n17785 ;
  assign y9281 = ~1'b0 ;
  assign y9282 = ~1'b0 ;
  assign y9283 = n17789 ;
  assign y9284 = ~1'b0 ;
  assign y9285 = ~1'b0 ;
  assign y9286 = n17020 ;
  assign y9287 = ~n17791 ;
  assign y9288 = n17794 ;
  assign y9289 = n17797 ;
  assign y9290 = ~1'b0 ;
  assign y9291 = ~1'b0 ;
  assign y9292 = ~n17799 ;
  assign y9293 = ~n17800 ;
  assign y9294 = ~n17802 ;
  assign y9295 = n17803 ;
  assign y9296 = n17804 ;
  assign y9297 = n17811 ;
  assign y9298 = ~n17813 ;
  assign y9299 = ~n17817 ;
  assign y9300 = ~n17819 ;
  assign y9301 = ~1'b0 ;
  assign y9302 = n17821 ;
  assign y9303 = n17825 ;
  assign y9304 = n17827 ;
  assign y9305 = ~1'b0 ;
  assign y9306 = n17829 ;
  assign y9307 = ~n17830 ;
  assign y9308 = n17832 ;
  assign y9309 = ~n17837 ;
  assign y9310 = ~1'b0 ;
  assign y9311 = ~1'b0 ;
  assign y9312 = ~1'b0 ;
  assign y9313 = n17840 ;
  assign y9314 = ~1'b0 ;
  assign y9315 = ~n17841 ;
  assign y9316 = n17843 ;
  assign y9317 = ~1'b0 ;
  assign y9318 = ~1'b0 ;
  assign y9319 = n17847 ;
  assign y9320 = n17848 ;
  assign y9321 = n17858 ;
  assign y9322 = n17860 ;
  assign y9323 = ~n17863 ;
  assign y9324 = ~n17865 ;
  assign y9325 = ~n17866 ;
  assign y9326 = ~n6817 ;
  assign y9327 = ~1'b0 ;
  assign y9328 = n17867 ;
  assign y9329 = n17872 ;
  assign y9330 = n17873 ;
  assign y9331 = ~n17874 ;
  assign y9332 = ~n17878 ;
  assign y9333 = n17881 ;
  assign y9334 = ~n17882 ;
  assign y9335 = n3389 ;
  assign y9336 = ~1'b0 ;
  assign y9337 = n17885 ;
  assign y9338 = ~n17887 ;
  assign y9339 = ~n17891 ;
  assign y9340 = n17893 ;
  assign y9341 = ~n17897 ;
  assign y9342 = ~1'b0 ;
  assign y9343 = n17898 ;
  assign y9344 = ~1'b0 ;
  assign y9345 = n17901 ;
  assign y9346 = n17906 ;
  assign y9347 = ~1'b0 ;
  assign y9348 = n17907 ;
  assign y9349 = ~n17908 ;
  assign y9350 = ~1'b0 ;
  assign y9351 = ~n17910 ;
  assign y9352 = ~n2958 ;
  assign y9353 = ~n17912 ;
  assign y9354 = ~1'b0 ;
  assign y9355 = ~n17913 ;
  assign y9356 = ~n5276 ;
  assign y9357 = ~n17917 ;
  assign y9358 = n17918 ;
  assign y9359 = n17920 ;
  assign y9360 = ~1'b0 ;
  assign y9361 = n17923 ;
  assign y9362 = n8038 ;
  assign y9363 = ~n17935 ;
  assign y9364 = n17936 ;
  assign y9365 = ~1'b0 ;
  assign y9366 = n17938 ;
  assign y9367 = ~1'b0 ;
  assign y9368 = n17764 ;
  assign y9369 = ~n17940 ;
  assign y9370 = ~n17943 ;
  assign y9371 = ~1'b0 ;
  assign y9372 = ~n17948 ;
  assign y9373 = ~1'b0 ;
  assign y9374 = n17952 ;
  assign y9375 = ~n17957 ;
  assign y9376 = n17958 ;
  assign y9377 = ~n17965 ;
  assign y9378 = n17966 ;
  assign y9379 = n17973 ;
  assign y9380 = ~n17976 ;
  assign y9381 = n17979 ;
  assign y9382 = n17980 ;
  assign y9383 = ~n17981 ;
  assign y9384 = ~1'b0 ;
  assign y9385 = 1'b0 ;
  assign y9386 = ~1'b0 ;
  assign y9387 = ~n17985 ;
  assign y9388 = ~1'b0 ;
  assign y9389 = n17993 ;
  assign y9390 = n17994 ;
  assign y9391 = n17998 ;
  assign y9392 = n18001 ;
  assign y9393 = n18004 ;
  assign y9394 = n18010 ;
  assign y9395 = ~n18011 ;
  assign y9396 = ~n18012 ;
  assign y9397 = ~1'b0 ;
  assign y9398 = ~1'b0 ;
  assign y9399 = ~n18015 ;
  assign y9400 = ~n18016 ;
  assign y9401 = ~n18017 ;
  assign y9402 = n18019 ;
  assign y9403 = ~1'b0 ;
  assign y9404 = n18023 ;
  assign y9405 = n18024 ;
  assign y9406 = ~1'b0 ;
  assign y9407 = ~n18027 ;
  assign y9408 = ~1'b0 ;
  assign y9409 = ~1'b0 ;
  assign y9410 = n18031 ;
  assign y9411 = n18034 ;
  assign y9412 = n18039 ;
  assign y9413 = ~1'b0 ;
  assign y9414 = ~n18041 ;
  assign y9415 = n18046 ;
  assign y9416 = 1'b0 ;
  assign y9417 = ~n18055 ;
  assign y9418 = ~1'b0 ;
  assign y9419 = n18060 ;
  assign y9420 = ~n18064 ;
  assign y9421 = n18066 ;
  assign y9422 = ~1'b0 ;
  assign y9423 = n18067 ;
  assign y9424 = ~1'b0 ;
  assign y9425 = ~n18068 ;
  assign y9426 = ~n18070 ;
  assign y9427 = ~n18072 ;
  assign y9428 = n18073 ;
  assign y9429 = ~1'b0 ;
  assign y9430 = ~1'b0 ;
  assign y9431 = ~n5091 ;
  assign y9432 = ~n18079 ;
  assign y9433 = ~n18081 ;
  assign y9434 = ~n18085 ;
  assign y9435 = ~1'b0 ;
  assign y9436 = n18088 ;
  assign y9437 = n18090 ;
  assign y9438 = ~n18091 ;
  assign y9439 = ~1'b0 ;
  assign y9440 = 1'b0 ;
  assign y9441 = ~1'b0 ;
  assign y9442 = ~1'b0 ;
  assign y9443 = ~n18098 ;
  assign y9444 = 1'b0 ;
  assign y9445 = ~n18100 ;
  assign y9446 = ~n18102 ;
  assign y9447 = n18104 ;
  assign y9448 = n18109 ;
  assign y9449 = ~n18113 ;
  assign y9450 = n18115 ;
  assign y9451 = n18118 ;
  assign y9452 = ~1'b0 ;
  assign y9453 = 1'b0 ;
  assign y9454 = ~n18121 ;
  assign y9455 = n18126 ;
  assign y9456 = ~1'b0 ;
  assign y9457 = ~1'b0 ;
  assign y9458 = ~1'b0 ;
  assign y9459 = ~n18128 ;
  assign y9460 = ~n18131 ;
  assign y9461 = ~n18133 ;
  assign y9462 = ~n18134 ;
  assign y9463 = n18136 ;
  assign y9464 = n18137 ;
  assign y9465 = n8271 ;
  assign y9466 = ~n18139 ;
  assign y9467 = ~n18143 ;
  assign y9468 = n18145 ;
  assign y9469 = ~1'b0 ;
  assign y9470 = ~n13806 ;
  assign y9471 = n18147 ;
  assign y9472 = ~n18148 ;
  assign y9473 = ~n16810 ;
  assign y9474 = n18149 ;
  assign y9475 = x94 ;
  assign y9476 = n18153 ;
  assign y9477 = ~1'b0 ;
  assign y9478 = n18156 ;
  assign y9479 = n18161 ;
  assign y9480 = n3010 ;
  assign y9481 = 1'b0 ;
  assign y9482 = n18164 ;
  assign y9483 = ~1'b0 ;
  assign y9484 = ~1'b0 ;
  assign y9485 = ~1'b0 ;
  assign y9486 = ~1'b0 ;
  assign y9487 = ~1'b0 ;
  assign y9488 = ~n18170 ;
  assign y9489 = ~n18171 ;
  assign y9490 = ~n150 ;
  assign y9491 = ~1'b0 ;
  assign y9492 = ~n18174 ;
  assign y9493 = ~1'b0 ;
  assign y9494 = n18176 ;
  assign y9495 = ~1'b0 ;
  assign y9496 = ~1'b0 ;
  assign y9497 = n18177 ;
  assign y9498 = n18179 ;
  assign y9499 = n18180 ;
  assign y9500 = ~1'b0 ;
  assign y9501 = n18181 ;
  assign y9502 = n18182 ;
  assign y9503 = ~n18184 ;
  assign y9504 = n18185 ;
  assign y9505 = n18188 ;
  assign y9506 = ~n6139 ;
  assign y9507 = ~n18191 ;
  assign y9508 = ~n18193 ;
  assign y9509 = ~1'b0 ;
  assign y9510 = ~n18194 ;
  assign y9511 = ~1'b0 ;
  assign y9512 = ~n18195 ;
  assign y9513 = n18196 ;
  assign y9514 = ~n18198 ;
  assign y9515 = ~n18203 ;
  assign y9516 = n18205 ;
  assign y9517 = n18206 ;
  assign y9518 = ~n18207 ;
  assign y9519 = n18211 ;
  assign y9520 = n18212 ;
  assign y9521 = n18216 ;
  assign y9522 = ~n4541 ;
  assign y9523 = ~1'b0 ;
  assign y9524 = ~n18217 ;
  assign y9525 = ~1'b0 ;
  assign y9526 = n18219 ;
  assign y9527 = n18220 ;
  assign y9528 = n876 ;
  assign y9529 = ~n18224 ;
  assign y9530 = n18225 ;
  assign y9531 = ~n14610 ;
  assign y9532 = ~n18227 ;
  assign y9533 = n18229 ;
  assign y9534 = ~1'b0 ;
  assign y9535 = n18232 ;
  assign y9536 = ~1'b0 ;
  assign y9537 = n18234 ;
  assign y9538 = ~n18238 ;
  assign y9539 = n12709 ;
  assign y9540 = n18239 ;
  assign y9541 = n18244 ;
  assign y9542 = ~n18247 ;
  assign y9543 = ~1'b0 ;
  assign y9544 = ~n18248 ;
  assign y9545 = n18252 ;
  assign y9546 = ~1'b0 ;
  assign y9547 = n18255 ;
  assign y9548 = 1'b0 ;
  assign y9549 = ~1'b0 ;
  assign y9550 = ~1'b0 ;
  assign y9551 = n18258 ;
  assign y9552 = n4979 ;
  assign y9553 = n18259 ;
  assign y9554 = ~n18261 ;
  assign y9555 = n18262 ;
  assign y9556 = n18264 ;
  assign y9557 = ~1'b0 ;
  assign y9558 = ~1'b0 ;
  assign y9559 = n18265 ;
  assign y9560 = ~n18266 ;
  assign y9561 = n18268 ;
  assign y9562 = ~1'b0 ;
  assign y9563 = ~n18270 ;
  assign y9564 = ~n18272 ;
  assign y9565 = n18273 ;
  assign y9566 = n18274 ;
  assign y9567 = ~n18275 ;
  assign y9568 = ~n18280 ;
  assign y9569 = ~1'b0 ;
  assign y9570 = n18281 ;
  assign y9571 = ~1'b0 ;
  assign y9572 = ~1'b0 ;
  assign y9573 = 1'b0 ;
  assign y9574 = ~1'b0 ;
  assign y9575 = n18285 ;
  assign y9576 = 1'b0 ;
  assign y9577 = ~n18290 ;
  assign y9578 = ~1'b0 ;
  assign y9579 = ~n18291 ;
  assign y9580 = n18292 ;
  assign y9581 = n18293 ;
  assign y9582 = n18294 ;
  assign y9583 = ~n18299 ;
  assign y9584 = n18301 ;
  assign y9585 = n18303 ;
  assign y9586 = n18307 ;
  assign y9587 = ~n18309 ;
  assign y9588 = ~n18316 ;
  assign y9589 = ~n18319 ;
  assign y9590 = ~1'b0 ;
  assign y9591 = ~1'b0 ;
  assign y9592 = n18326 ;
  assign y9593 = n18328 ;
  assign y9594 = ~n18331 ;
  assign y9595 = ~n18334 ;
  assign y9596 = n18338 ;
  assign y9597 = ~n10109 ;
  assign y9598 = ~1'b0 ;
  assign y9599 = ~1'b0 ;
  assign y9600 = ~n18340 ;
  assign y9601 = ~n18341 ;
  assign y9602 = n18342 ;
  assign y9603 = ~1'b0 ;
  assign y9604 = ~1'b0 ;
  assign y9605 = n2235 ;
  assign y9606 = ~1'b0 ;
  assign y9607 = n18353 ;
  assign y9608 = ~1'b0 ;
  assign y9609 = ~n18354 ;
  assign y9610 = n18355 ;
  assign y9611 = n18356 ;
  assign y9612 = ~1'b0 ;
  assign y9613 = ~1'b0 ;
  assign y9614 = n18357 ;
  assign y9615 = ~n18359 ;
  assign y9616 = n18361 ;
  assign y9617 = ~n18362 ;
  assign y9618 = ~1'b0 ;
  assign y9619 = ~1'b0 ;
  assign y9620 = n18363 ;
  assign y9621 = ~n18364 ;
  assign y9622 = ~1'b0 ;
  assign y9623 = ~n18365 ;
  assign y9624 = ~1'b0 ;
  assign y9625 = n18368 ;
  assign y9626 = ~1'b0 ;
  assign y9627 = ~1'b0 ;
  assign y9628 = n18369 ;
  assign y9629 = ~n18371 ;
  assign y9630 = ~n18375 ;
  assign y9631 = n18380 ;
  assign y9632 = ~n18385 ;
  assign y9633 = n18390 ;
  assign y9634 = ~1'b0 ;
  assign y9635 = ~n18393 ;
  assign y9636 = ~n18394 ;
  assign y9637 = ~1'b0 ;
  assign y9638 = n18401 ;
  assign y9639 = ~n18404 ;
  assign y9640 = ~1'b0 ;
  assign y9641 = n18405 ;
  assign y9642 = 1'b0 ;
  assign y9643 = ~1'b0 ;
  assign y9644 = ~1'b0 ;
  assign y9645 = ~n18407 ;
  assign y9646 = ~1'b0 ;
  assign y9647 = n18410 ;
  assign y9648 = ~n18411 ;
  assign y9649 = n2635 ;
  assign y9650 = ~1'b0 ;
  assign y9651 = n18412 ;
  assign y9652 = ~n18415 ;
  assign y9653 = n18417 ;
  assign y9654 = ~n14387 ;
  assign y9655 = ~n18421 ;
  assign y9656 = ~n18423 ;
  assign y9657 = ~n18427 ;
  assign y9658 = ~n18430 ;
  assign y9659 = ~n18436 ;
  assign y9660 = ~n18438 ;
  assign y9661 = ~1'b0 ;
  assign y9662 = ~1'b0 ;
  assign y9663 = ~1'b0 ;
  assign y9664 = 1'b0 ;
  assign y9665 = ~n18439 ;
  assign y9666 = ~n18440 ;
  assign y9667 = ~1'b0 ;
  assign y9668 = ~1'b0 ;
  assign y9669 = ~1'b0 ;
  assign y9670 = n18442 ;
  assign y9671 = n18443 ;
  assign y9672 = ~1'b0 ;
  assign y9673 = n18444 ;
  assign y9674 = ~n18447 ;
  assign y9675 = ~n18448 ;
  assign y9676 = ~n18454 ;
  assign y9677 = ~n18455 ;
  assign y9678 = ~n18460 ;
  assign y9679 = ~n18462 ;
  assign y9680 = ~1'b0 ;
  assign y9681 = n18464 ;
  assign y9682 = ~n18469 ;
  assign y9683 = ~n18470 ;
  assign y9684 = ~n18473 ;
  assign y9685 = 1'b0 ;
  assign y9686 = ~n18474 ;
  assign y9687 = n11177 ;
  assign y9688 = n18477 ;
  assign y9689 = n18479 ;
  assign y9690 = n18481 ;
  assign y9691 = n18484 ;
  assign y9692 = ~1'b0 ;
  assign y9693 = ~1'b0 ;
  assign y9694 = ~1'b0 ;
  assign y9695 = ~n18487 ;
  assign y9696 = n18491 ;
  assign y9697 = ~1'b0 ;
  assign y9698 = n18493 ;
  assign y9699 = ~1'b0 ;
  assign y9700 = ~n18494 ;
  assign y9701 = n18499 ;
  assign y9702 = ~n18501 ;
  assign y9703 = ~n18504 ;
  assign y9704 = ~n18505 ;
  assign y9705 = n18510 ;
  assign y9706 = ~1'b0 ;
  assign y9707 = ~1'b0 ;
  assign y9708 = n18513 ;
  assign y9709 = ~n18515 ;
  assign y9710 = ~n18521 ;
  assign y9711 = n18540 ;
  assign y9712 = ~1'b0 ;
  assign y9713 = ~n18541 ;
  assign y9714 = ~n18544 ;
  assign y9715 = ~n18545 ;
  assign y9716 = ~1'b0 ;
  assign y9717 = ~n18552 ;
  assign y9718 = ~1'b0 ;
  assign y9719 = ~n18555 ;
  assign y9720 = ~n18556 ;
  assign y9721 = ~n18559 ;
  assign y9722 = n18560 ;
  assign y9723 = ~n18561 ;
  assign y9724 = n18562 ;
  assign y9725 = ~1'b0 ;
  assign y9726 = ~n18563 ;
  assign y9727 = n18564 ;
  assign y9728 = ~n18566 ;
  assign y9729 = ~n18567 ;
  assign y9730 = ~1'b0 ;
  assign y9731 = ~n18569 ;
  assign y9732 = ~1'b0 ;
  assign y9733 = ~n9666 ;
  assign y9734 = ~1'b0 ;
  assign y9735 = ~n18570 ;
  assign y9736 = ~1'b0 ;
  assign y9737 = ~1'b0 ;
  assign y9738 = n18573 ;
  assign y9739 = 1'b0 ;
  assign y9740 = 1'b0 ;
  assign y9741 = ~1'b0 ;
  assign y9742 = ~1'b0 ;
  assign y9743 = ~1'b0 ;
  assign y9744 = n18577 ;
  assign y9745 = n18581 ;
  assign y9746 = ~1'b0 ;
  assign y9747 = n18583 ;
  assign y9748 = ~1'b0 ;
  assign y9749 = ~n18585 ;
  assign y9750 = n18586 ;
  assign y9751 = ~n18588 ;
  assign y9752 = n18589 ;
  assign y9753 = ~n18591 ;
  assign y9754 = ~n18592 ;
  assign y9755 = 1'b0 ;
  assign y9756 = ~n18593 ;
  assign y9757 = ~n18597 ;
  assign y9758 = 1'b0 ;
  assign y9759 = ~1'b0 ;
  assign y9760 = n18600 ;
  assign y9761 = n18602 ;
  assign y9762 = ~n18603 ;
  assign y9763 = ~n18608 ;
  assign y9764 = n18609 ;
  assign y9765 = n18610 ;
  assign y9766 = ~n18611 ;
  assign y9767 = n18613 ;
  assign y9768 = n18614 ;
  assign y9769 = ~n18615 ;
  assign y9770 = ~1'b0 ;
  assign y9771 = ~n18616 ;
  assign y9772 = ~x102 ;
  assign y9773 = n18617 ;
  assign y9774 = ~n9192 ;
  assign y9775 = ~n18620 ;
  assign y9776 = ~n18622 ;
  assign y9777 = ~1'b0 ;
  assign y9778 = n18625 ;
  assign y9779 = ~1'b0 ;
  assign y9780 = ~1'b0 ;
  assign y9781 = ~1'b0 ;
  assign y9782 = n10191 ;
  assign y9783 = n13511 ;
  assign y9784 = ~n18627 ;
  assign y9785 = ~n18629 ;
  assign y9786 = n18631 ;
  assign y9787 = ~n18636 ;
  assign y9788 = n18639 ;
  assign y9789 = n18646 ;
  assign y9790 = n6021 ;
  assign y9791 = ~1'b0 ;
  assign y9792 = ~n18648 ;
  assign y9793 = n18650 ;
  assign y9794 = n18651 ;
  assign y9795 = ~1'b0 ;
  assign y9796 = n18652 ;
  assign y9797 = ~n18655 ;
  assign y9798 = 1'b0 ;
  assign y9799 = n18656 ;
  assign y9800 = ~n18657 ;
  assign y9801 = ~n18659 ;
  assign y9802 = n9396 ;
  assign y9803 = ~n18661 ;
  assign y9804 = ~n18666 ;
  assign y9805 = ~1'b0 ;
  assign y9806 = ~n18668 ;
  assign y9807 = ~n18673 ;
  assign y9808 = ~1'b0 ;
  assign y9809 = ~n18676 ;
  assign y9810 = ~1'b0 ;
  assign y9811 = ~n18677 ;
  assign y9812 = n18679 ;
  assign y9813 = ~1'b0 ;
  assign y9814 = n9528 ;
  assign y9815 = n18680 ;
  assign y9816 = n18682 ;
  assign y9817 = n18683 ;
  assign y9818 = ~n18685 ;
  assign y9819 = ~1'b0 ;
  assign y9820 = ~1'b0 ;
  assign y9821 = ~1'b0 ;
  assign y9822 = n18690 ;
  assign y9823 = ~1'b0 ;
  assign y9824 = n18695 ;
  assign y9825 = ~n18697 ;
  assign y9826 = ~1'b0 ;
  assign y9827 = ~1'b0 ;
  assign y9828 = n18699 ;
  assign y9829 = ~n18700 ;
  assign y9830 = ~n9768 ;
  assign y9831 = n18702 ;
  assign y9832 = ~n18703 ;
  assign y9833 = n18704 ;
  assign y9834 = n18706 ;
  assign y9835 = ~n18707 ;
  assign y9836 = ~1'b0 ;
  assign y9837 = ~1'b0 ;
  assign y9838 = n18708 ;
  assign y9839 = ~n18709 ;
  assign y9840 = n18711 ;
  assign y9841 = ~n18713 ;
  assign y9842 = n18715 ;
  assign y9843 = ~1'b0 ;
  assign y9844 = ~n18716 ;
  assign y9845 = ~1'b0 ;
  assign y9846 = n18718 ;
  assign y9847 = 1'b0 ;
  assign y9848 = ~1'b0 ;
  assign y9849 = n18720 ;
  assign y9850 = ~1'b0 ;
  assign y9851 = n18724 ;
  assign y9852 = ~1'b0 ;
  assign y9853 = ~n18725 ;
  assign y9854 = 1'b0 ;
  assign y9855 = ~n9467 ;
  assign y9856 = n792 ;
  assign y9857 = n18726 ;
  assign y9858 = ~n18735 ;
  assign y9859 = ~n18738 ;
  assign y9860 = n18739 ;
  assign y9861 = ~1'b0 ;
  assign y9862 = n18741 ;
  assign y9863 = n18743 ;
  assign y9864 = n18745 ;
  assign y9865 = ~1'b0 ;
  assign y9866 = ~1'b0 ;
  assign y9867 = ~n18746 ;
  assign y9868 = ~n18750 ;
  assign y9869 = ~n18752 ;
  assign y9870 = ~n18754 ;
  assign y9871 = n18757 ;
  assign y9872 = ~n13046 ;
  assign y9873 = ~n18758 ;
  assign y9874 = ~1'b0 ;
  assign y9875 = ~1'b0 ;
  assign y9876 = ~n18761 ;
  assign y9877 = ~n18763 ;
  assign y9878 = ~n18766 ;
  assign y9879 = ~n18770 ;
  assign y9880 = ~1'b0 ;
  assign y9881 = ~n18773 ;
  assign y9882 = ~n18774 ;
  assign y9883 = n18775 ;
  assign y9884 = ~1'b0 ;
  assign y9885 = ~1'b0 ;
  assign y9886 = ~n11947 ;
  assign y9887 = ~n12158 ;
  assign y9888 = n18776 ;
  assign y9889 = ~n18778 ;
  assign y9890 = ~n18783 ;
  assign y9891 = ~1'b0 ;
  assign y9892 = n18785 ;
  assign y9893 = n18787 ;
  assign y9894 = ~n18791 ;
  assign y9895 = n18792 ;
  assign y9896 = n18793 ;
  assign y9897 = n18794 ;
  assign y9898 = n18801 ;
  assign y9899 = n18802 ;
  assign y9900 = n18803 ;
  assign y9901 = ~n18804 ;
  assign y9902 = ~n18806 ;
  assign y9903 = n18808 ;
  assign y9904 = ~1'b0 ;
  assign y9905 = ~1'b0 ;
  assign y9906 = ~n18810 ;
  assign y9907 = ~1'b0 ;
  assign y9908 = ~n18811 ;
  assign y9909 = n18814 ;
  assign y9910 = ~1'b0 ;
  assign y9911 = ~n13580 ;
  assign y9912 = n18820 ;
  assign y9913 = n18822 ;
  assign y9914 = n1555 ;
  assign y9915 = ~1'b0 ;
  assign y9916 = ~n18823 ;
  assign y9917 = n1259 ;
  assign y9918 = ~n18828 ;
  assign y9919 = ~1'b0 ;
  assign y9920 = n18833 ;
  assign y9921 = ~1'b0 ;
  assign y9922 = ~n18834 ;
  assign y9923 = ~n18835 ;
  assign y9924 = ~n6568 ;
  assign y9925 = ~1'b0 ;
  assign y9926 = n18837 ;
  assign y9927 = ~1'b0 ;
  assign y9928 = ~1'b0 ;
  assign y9929 = ~n18838 ;
  assign y9930 = n10169 ;
  assign y9931 = ~n18839 ;
  assign y9932 = ~n18840 ;
  assign y9933 = n18841 ;
  assign y9934 = n18845 ;
  assign y9935 = ~n18847 ;
  assign y9936 = ~n18848 ;
  assign y9937 = n18851 ;
  assign y9938 = n18854 ;
  assign y9939 = n18858 ;
  assign y9940 = n18860 ;
  assign y9941 = ~n18861 ;
  assign y9942 = ~n4403 ;
  assign y9943 = n18862 ;
  assign y9944 = n18866 ;
  assign y9945 = n18867 ;
  assign y9946 = n18871 ;
  assign y9947 = ~n10875 ;
  assign y9948 = ~1'b0 ;
  assign y9949 = n18874 ;
  assign y9950 = ~1'b0 ;
  assign y9951 = ~1'b0 ;
  assign y9952 = ~n18877 ;
  assign y9953 = ~1'b0 ;
  assign y9954 = ~1'b0 ;
  assign y9955 = n18378 ;
  assign y9956 = ~1'b0 ;
  assign y9957 = n18880 ;
  assign y9958 = ~n18884 ;
  assign y9959 = ~1'b0 ;
  assign y9960 = n18886 ;
  assign y9961 = ~1'b0 ;
  assign y9962 = ~n18887 ;
  assign y9963 = n18888 ;
  assign y9964 = n18892 ;
  assign y9965 = ~1'b0 ;
  assign y9966 = n18896 ;
  assign y9967 = ~n18900 ;
  assign y9968 = n18903 ;
  assign y9969 = ~n18904 ;
  assign y9970 = ~1'b0 ;
  assign y9971 = n18908 ;
  assign y9972 = n18909 ;
  assign y9973 = ~1'b0 ;
  assign y9974 = ~1'b0 ;
  assign y9975 = ~1'b0 ;
  assign y9976 = n18926 ;
  assign y9977 = ~n18930 ;
  assign y9978 = ~n18934 ;
  assign y9979 = ~n7353 ;
  assign y9980 = ~n18937 ;
  assign y9981 = n3606 ;
  assign y9982 = ~1'b0 ;
  assign y9983 = ~1'b0 ;
  assign y9984 = ~n9865 ;
  assign y9985 = n18938 ;
  assign y9986 = n18940 ;
  assign y9987 = n18943 ;
  assign y9988 = n5524 ;
  assign y9989 = n18944 ;
  assign y9990 = ~n14441 ;
  assign y9991 = ~n18945 ;
  assign y9992 = n18946 ;
  assign y9993 = ~n18948 ;
  assign y9994 = ~n18951 ;
  assign y9995 = ~1'b0 ;
  assign y9996 = ~1'b0 ;
  assign y9997 = n18954 ;
  assign y9998 = n18955 ;
  assign y9999 = ~n18956 ;
  assign y10000 = ~1'b0 ;
  assign y10001 = n18958 ;
  assign y10002 = ~n18959 ;
  assign y10003 = n18960 ;
  assign y10004 = 1'b0 ;
  assign y10005 = ~n18962 ;
  assign y10006 = n18963 ;
  assign y10007 = ~n18964 ;
  assign y10008 = n18968 ;
  assign y10009 = n18970 ;
  assign y10010 = ~n18973 ;
  assign y10011 = ~1'b0 ;
  assign y10012 = ~n18975 ;
  assign y10013 = ~n18976 ;
  assign y10014 = n1535 ;
  assign y10015 = n18978 ;
  assign y10016 = ~n18979 ;
  assign y10017 = ~n12417 ;
  assign y10018 = n18980 ;
  assign y10019 = ~n13373 ;
  assign y10020 = ~1'b0 ;
  assign y10021 = ~n18981 ;
  assign y10022 = n18986 ;
  assign y10023 = n5011 ;
  assign y10024 = ~n18989 ;
  assign y10025 = ~n18991 ;
  assign y10026 = ~1'b0 ;
  assign y10027 = n18993 ;
  assign y10028 = ~n6899 ;
  assign y10029 = ~n4571 ;
  assign y10030 = ~1'b0 ;
  assign y10031 = 1'b0 ;
  assign y10032 = ~n18997 ;
  assign y10033 = ~n18999 ;
  assign y10034 = ~1'b0 ;
  assign y10035 = ~1'b0 ;
  assign y10036 = ~n19002 ;
  assign y10037 = ~1'b0 ;
  assign y10038 = 1'b0 ;
  assign y10039 = ~n19003 ;
  assign y10040 = 1'b0 ;
  assign y10041 = ~1'b0 ;
  assign y10042 = ~n19007 ;
  assign y10043 = ~n18719 ;
  assign y10044 = ~1'b0 ;
  assign y10045 = 1'b0 ;
  assign y10046 = n19008 ;
  assign y10047 = ~n19009 ;
  assign y10048 = n19010 ;
  assign y10049 = n8801 ;
  assign y10050 = n19011 ;
  assign y10051 = ~n19012 ;
  assign y10052 = ~n19019 ;
  assign y10053 = ~1'b0 ;
  assign y10054 = n11642 ;
  assign y10055 = ~n19020 ;
  assign y10056 = ~1'b0 ;
  assign y10057 = ~1'b0 ;
  assign y10058 = ~n19022 ;
  assign y10059 = ~1'b0 ;
  assign y10060 = ~1'b0 ;
  assign y10061 = ~1'b0 ;
  assign y10062 = ~1'b0 ;
  assign y10063 = ~n19026 ;
  assign y10064 = n19027 ;
  assign y10065 = ~1'b0 ;
  assign y10066 = n19029 ;
  assign y10067 = ~n19031 ;
  assign y10068 = n19034 ;
  assign y10069 = ~1'b0 ;
  assign y10070 = ~1'b0 ;
  assign y10071 = ~1'b0 ;
  assign y10072 = ~n19036 ;
  assign y10073 = ~1'b0 ;
  assign y10074 = ~n19040 ;
  assign y10075 = ~n6623 ;
  assign y10076 = n19042 ;
  assign y10077 = ~n19043 ;
  assign y10078 = ~1'b0 ;
  assign y10079 = ~n19046 ;
  assign y10080 = n19048 ;
  assign y10081 = n19053 ;
  assign y10082 = n19054 ;
  assign y10083 = n19060 ;
  assign y10084 = ~1'b0 ;
  assign y10085 = ~n19063 ;
  assign y10086 = ~1'b0 ;
  assign y10087 = n19069 ;
  assign y10088 = n19070 ;
  assign y10089 = n19074 ;
  assign y10090 = n15327 ;
  assign y10091 = ~1'b0 ;
  assign y10092 = ~1'b0 ;
  assign y10093 = ~1'b0 ;
  assign y10094 = ~1'b0 ;
  assign y10095 = ~n19076 ;
  assign y10096 = ~n8810 ;
  assign y10097 = ~n19077 ;
  assign y10098 = n19078 ;
  assign y10099 = ~n19086 ;
  assign y10100 = n19089 ;
  assign y10101 = ~n19091 ;
  assign y10102 = ~n19094 ;
  assign y10103 = ~n19095 ;
  assign y10104 = n3620 ;
  assign y10105 = n19096 ;
  assign y10106 = ~n19097 ;
  assign y10107 = ~n19098 ;
  assign y10108 = ~n19102 ;
  assign y10109 = ~n19104 ;
  assign y10110 = ~1'b0 ;
  assign y10111 = n19106 ;
  assign y10112 = ~1'b0 ;
  assign y10113 = n19109 ;
  assign y10114 = n19112 ;
  assign y10115 = ~n19113 ;
  assign y10116 = ~n19115 ;
  assign y10117 = ~n8062 ;
  assign y10118 = ~n8720 ;
  assign y10119 = ~n19121 ;
  assign y10120 = ~n5737 ;
  assign y10121 = n19128 ;
  assign y10122 = n19131 ;
  assign y10123 = ~1'b0 ;
  assign y10124 = ~1'b0 ;
  assign y10125 = n19132 ;
  assign y10126 = ~1'b0 ;
  assign y10127 = ~1'b0 ;
  assign y10128 = n19136 ;
  assign y10129 = 1'b0 ;
  assign y10130 = n563 ;
  assign y10131 = ~n19139 ;
  assign y10132 = ~n19140 ;
  assign y10133 = n19142 ;
  assign y10134 = ~n19143 ;
  assign y10135 = ~n19145 ;
  assign y10136 = n19149 ;
  assign y10137 = ~1'b0 ;
  assign y10138 = ~n19151 ;
  assign y10139 = ~1'b0 ;
  assign y10140 = ~n19152 ;
  assign y10141 = ~n19153 ;
  assign y10142 = ~n19155 ;
  assign y10143 = ~1'b0 ;
  assign y10144 = n19156 ;
  assign y10145 = ~1'b0 ;
  assign y10146 = n18932 ;
  assign y10147 = n19157 ;
  assign y10148 = ~n19158 ;
  assign y10149 = ~n19159 ;
  assign y10150 = n19161 ;
  assign y10151 = n19162 ;
  assign y10152 = n19163 ;
  assign y10153 = ~n19165 ;
  assign y10154 = ~n19166 ;
  assign y10155 = n6821 ;
  assign y10156 = ~n19169 ;
  assign y10157 = n19170 ;
  assign y10158 = ~n19171 ;
  assign y10159 = n19174 ;
  assign y10160 = n19178 ;
  assign y10161 = n19180 ;
  assign y10162 = ~n19181 ;
  assign y10163 = 1'b0 ;
  assign y10164 = ~n19183 ;
  assign y10165 = ~n19186 ;
  assign y10166 = ~1'b0 ;
  assign y10167 = ~n17857 ;
  assign y10168 = ~1'b0 ;
  assign y10169 = ~n19188 ;
  assign y10170 = ~n19190 ;
  assign y10171 = ~1'b0 ;
  assign y10172 = ~n19191 ;
  assign y10173 = ~n19193 ;
  assign y10174 = n19195 ;
  assign y10175 = n19196 ;
  assign y10176 = n19199 ;
  assign y10177 = n19201 ;
  assign y10178 = n19202 ;
  assign y10179 = n19203 ;
  assign y10180 = ~n19204 ;
  assign y10181 = ~n19207 ;
  assign y10182 = ~n19208 ;
  assign y10183 = ~1'b0 ;
  assign y10184 = n19210 ;
  assign y10185 = ~n19212 ;
  assign y10186 = ~n19217 ;
  assign y10187 = n19221 ;
  assign y10188 = ~1'b0 ;
  assign y10189 = ~n19222 ;
  assign y10190 = ~n19225 ;
  assign y10191 = n1720 ;
  assign y10192 = ~n19233 ;
  assign y10193 = ~1'b0 ;
  assign y10194 = ~1'b0 ;
  assign y10195 = n3943 ;
  assign y10196 = ~n19234 ;
  assign y10197 = ~n7612 ;
  assign y10198 = ~n19237 ;
  assign y10199 = n19239 ;
  assign y10200 = n14880 ;
  assign y10201 = ~n19242 ;
  assign y10202 = ~n19250 ;
  assign y10203 = n19251 ;
  assign y10204 = ~1'b0 ;
  assign y10205 = ~n17418 ;
  assign y10206 = ~1'b0 ;
  assign y10207 = ~n19256 ;
  assign y10208 = ~1'b0 ;
  assign y10209 = ~n19265 ;
  assign y10210 = ~1'b0 ;
  assign y10211 = n19267 ;
  assign y10212 = ~1'b0 ;
  assign y10213 = n19268 ;
  assign y10214 = ~1'b0 ;
  assign y10215 = ~1'b0 ;
  assign y10216 = n802 ;
  assign y10217 = ~n19269 ;
  assign y10218 = ~n19270 ;
  assign y10219 = n19271 ;
  assign y10220 = n19274 ;
  assign y10221 = n19275 ;
  assign y10222 = ~1'b0 ;
  assign y10223 = ~1'b0 ;
  assign y10224 = n19277 ;
  assign y10225 = ~1'b0 ;
  assign y10226 = n19278 ;
  assign y10227 = n19282 ;
  assign y10228 = n19284 ;
  assign y10229 = n11913 ;
  assign y10230 = n19288 ;
  assign y10231 = ~n19289 ;
  assign y10232 = ~n362 ;
  assign y10233 = ~n19290 ;
  assign y10234 = ~1'b0 ;
  assign y10235 = n19291 ;
  assign y10236 = n19292 ;
  assign y10237 = ~1'b0 ;
  assign y10238 = ~n19295 ;
  assign y10239 = n15949 ;
  assign y10240 = ~1'b0 ;
  assign y10241 = ~n1396 ;
  assign y10242 = ~n5991 ;
  assign y10243 = n19296 ;
  assign y10244 = ~n19300 ;
  assign y10245 = ~1'b0 ;
  assign y10246 = ~n19302 ;
  assign y10247 = n19304 ;
  assign y10248 = n19310 ;
  assign y10249 = n19312 ;
  assign y10250 = ~1'b0 ;
  assign y10251 = ~1'b0 ;
  assign y10252 = n19313 ;
  assign y10253 = n19314 ;
  assign y10254 = ~n19315 ;
  assign y10255 = ~1'b0 ;
  assign y10256 = ~1'b0 ;
  assign y10257 = n19316 ;
  assign y10258 = n19319 ;
  assign y10259 = ~n19328 ;
  assign y10260 = ~n19330 ;
  assign y10261 = ~1'b0 ;
  assign y10262 = ~n19331 ;
  assign y10263 = ~n19332 ;
  assign y10264 = n19334 ;
  assign y10265 = ~n19335 ;
  assign y10266 = ~n19336 ;
  assign y10267 = ~1'b0 ;
  assign y10268 = ~n4355 ;
  assign y10269 = ~n19339 ;
  assign y10270 = ~n19346 ;
  assign y10271 = n19348 ;
  assign y10272 = ~1'b0 ;
  assign y10273 = ~n3869 ;
  assign y10274 = ~n19349 ;
  assign y10275 = ~1'b0 ;
  assign y10276 = ~1'b0 ;
  assign y10277 = ~1'b0 ;
  assign y10278 = ~1'b0 ;
  assign y10279 = n3792 ;
  assign y10280 = ~n19351 ;
  assign y10281 = ~1'b0 ;
  assign y10282 = ~1'b0 ;
  assign y10283 = ~n19352 ;
  assign y10284 = ~1'b0 ;
  assign y10285 = n19356 ;
  assign y10286 = ~n19358 ;
  assign y10287 = ~n19360 ;
  assign y10288 = n19361 ;
  assign y10289 = n19362 ;
  assign y10290 = ~1'b0 ;
  assign y10291 = ~n19365 ;
  assign y10292 = ~n4141 ;
  assign y10293 = ~1'b0 ;
  assign y10294 = ~1'b0 ;
  assign y10295 = ~1'b0 ;
  assign y10296 = ~1'b0 ;
  assign y10297 = ~n19367 ;
  assign y10298 = ~n11577 ;
  assign y10299 = ~n19368 ;
  assign y10300 = ~1'b0 ;
  assign y10301 = ~1'b0 ;
  assign y10302 = n19371 ;
  assign y10303 = ~1'b0 ;
  assign y10304 = ~n19373 ;
  assign y10305 = n19374 ;
  assign y10306 = n19375 ;
  assign y10307 = ~n19376 ;
  assign y10308 = ~1'b0 ;
  assign y10309 = ~n19378 ;
  assign y10310 = n19379 ;
  assign y10311 = n19380 ;
  assign y10312 = n1970 ;
  assign y10313 = n19384 ;
  assign y10314 = n19385 ;
  assign y10315 = ~n19386 ;
  assign y10316 = n19387 ;
  assign y10317 = ~1'b0 ;
  assign y10318 = ~n19388 ;
  assign y10319 = n19389 ;
  assign y10320 = ~1'b0 ;
  assign y10321 = ~1'b0 ;
  assign y10322 = ~1'b0 ;
  assign y10323 = ~n19391 ;
  assign y10324 = n18631 ;
  assign y10325 = ~1'b0 ;
  assign y10326 = ~1'b0 ;
  assign y10327 = ~1'b0 ;
  assign y10328 = n19393 ;
  assign y10329 = ~n19394 ;
  assign y10330 = ~1'b0 ;
  assign y10331 = ~1'b0 ;
  assign y10332 = ~1'b0 ;
  assign y10333 = n19396 ;
  assign y10334 = n19401 ;
  assign y10335 = n19402 ;
  assign y10336 = ~n19407 ;
  assign y10337 = n19409 ;
  assign y10338 = n19410 ;
  assign y10339 = ~n19411 ;
  assign y10340 = ~n19414 ;
  assign y10341 = ~1'b0 ;
  assign y10342 = n19416 ;
  assign y10343 = n19421 ;
  assign y10344 = n19431 ;
  assign y10345 = ~n19434 ;
  assign y10346 = ~n19438 ;
  assign y10347 = ~1'b0 ;
  assign y10348 = ~n19440 ;
  assign y10349 = ~n19441 ;
  assign y10350 = ~n19442 ;
  assign y10351 = ~n19445 ;
  assign y10352 = ~n19446 ;
  assign y10353 = ~n19448 ;
  assign y10354 = ~1'b0 ;
  assign y10355 = ~1'b0 ;
  assign y10356 = ~n19452 ;
  assign y10357 = n19453 ;
  assign y10358 = n19454 ;
  assign y10359 = ~n19455 ;
  assign y10360 = ~1'b0 ;
  assign y10361 = ~n19457 ;
  assign y10362 = n19463 ;
  assign y10363 = ~n19464 ;
  assign y10364 = n19465 ;
  assign y10365 = ~n19468 ;
  assign y10366 = n4224 ;
  assign y10367 = ~n19471 ;
  assign y10368 = ~n19472 ;
  assign y10369 = ~1'b0 ;
  assign y10370 = ~n9847 ;
  assign y10371 = ~n1679 ;
  assign y10372 = ~1'b0 ;
  assign y10373 = n19474 ;
  assign y10374 = n19475 ;
  assign y10375 = ~1'b0 ;
  assign y10376 = ~n19478 ;
  assign y10377 = ~1'b0 ;
  assign y10378 = n19480 ;
  assign y10379 = ~1'b0 ;
  assign y10380 = n19482 ;
  assign y10381 = ~1'b0 ;
  assign y10382 = ~1'b0 ;
  assign y10383 = ~n19485 ;
  assign y10384 = n19487 ;
  assign y10385 = ~n19491 ;
  assign y10386 = n19493 ;
  assign y10387 = n19495 ;
  assign y10388 = ~1'b0 ;
  assign y10389 = ~1'b0 ;
  assign y10390 = ~1'b0 ;
  assign y10391 = n19497 ;
  assign y10392 = n794 ;
  assign y10393 = n19499 ;
  assign y10394 = ~1'b0 ;
  assign y10395 = 1'b0 ;
  assign y10396 = ~1'b0 ;
  assign y10397 = n19501 ;
  assign y10398 = ~1'b0 ;
  assign y10399 = ~n19502 ;
  assign y10400 = ~n19503 ;
  assign y10401 = ~1'b0 ;
  assign y10402 = n19509 ;
  assign y10403 = ~n19510 ;
  assign y10404 = ~n19512 ;
  assign y10405 = ~1'b0 ;
  assign y10406 = n19522 ;
  assign y10407 = ~n19524 ;
  assign y10408 = ~n19525 ;
  assign y10409 = ~1'b0 ;
  assign y10410 = ~1'b0 ;
  assign y10411 = n19529 ;
  assign y10412 = n13331 ;
  assign y10413 = n19530 ;
  assign y10414 = n19531 ;
  assign y10415 = n2821 ;
  assign y10416 = n19538 ;
  assign y10417 = ~n2607 ;
  assign y10418 = ~n19542 ;
  assign y10419 = ~1'b0 ;
  assign y10420 = n19543 ;
  assign y10421 = n19544 ;
  assign y10422 = ~1'b0 ;
  assign y10423 = ~1'b0 ;
  assign y10424 = n19547 ;
  assign y10425 = ~1'b0 ;
  assign y10426 = ~1'b0 ;
  assign y10427 = 1'b0 ;
  assign y10428 = ~1'b0 ;
  assign y10429 = n19553 ;
  assign y10430 = n1281 ;
  assign y10431 = ~1'b0 ;
  assign y10432 = n19555 ;
  assign y10433 = ~n19556 ;
  assign y10434 = ~1'b0 ;
  assign y10435 = n19557 ;
  assign y10436 = ~n19558 ;
  assign y10437 = n19559 ;
  assign y10438 = n19563 ;
  assign y10439 = ~1'b0 ;
  assign y10440 = n16032 ;
  assign y10441 = ~1'b0 ;
  assign y10442 = n19569 ;
  assign y10443 = ~n19570 ;
  assign y10444 = ~1'b0 ;
  assign y10445 = ~n19579 ;
  assign y10446 = n19580 ;
  assign y10447 = n7145 ;
  assign y10448 = ~1'b0 ;
  assign y10449 = n19583 ;
  assign y10450 = ~n16028 ;
  assign y10451 = n10775 ;
  assign y10452 = ~1'b0 ;
  assign y10453 = ~n19586 ;
  assign y10454 = n19589 ;
  assign y10455 = n19590 ;
  assign y10456 = ~n19595 ;
  assign y10457 = n19601 ;
  assign y10458 = ~n19607 ;
  assign y10459 = ~n19608 ;
  assign y10460 = n19609 ;
  assign y10461 = n19611 ;
  assign y10462 = ~1'b0 ;
  assign y10463 = ~n19613 ;
  assign y10464 = n19616 ;
  assign y10465 = ~n630 ;
  assign y10466 = ~n19621 ;
  assign y10467 = n10271 ;
  assign y10468 = ~n19622 ;
  assign y10469 = ~n19623 ;
  assign y10470 = n19624 ;
  assign y10471 = n19625 ;
  assign y10472 = ~1'b0 ;
  assign y10473 = n8452 ;
  assign y10474 = n4886 ;
  assign y10475 = ~n19629 ;
  assign y10476 = n19636 ;
  assign y10477 = ~n4522 ;
  assign y10478 = ~n19641 ;
  assign y10479 = n19642 ;
  assign y10480 = ~1'b0 ;
  assign y10481 = ~1'b0 ;
  assign y10482 = n19645 ;
  assign y10483 = ~1'b0 ;
  assign y10484 = ~n19647 ;
  assign y10485 = ~1'b0 ;
  assign y10486 = n19648 ;
  assign y10487 = ~n19649 ;
  assign y10488 = n19655 ;
  assign y10489 = ~n19657 ;
  assign y10490 = ~1'b0 ;
  assign y10491 = ~n1439 ;
  assign y10492 = n19659 ;
  assign y10493 = ~1'b0 ;
  assign y10494 = n19660 ;
  assign y10495 = n19662 ;
  assign y10496 = ~n19665 ;
  assign y10497 = n19676 ;
  assign y10498 = ~1'b0 ;
  assign y10499 = n19681 ;
  assign y10500 = ~1'b0 ;
  assign y10501 = ~n19683 ;
  assign y10502 = n19686 ;
  assign y10503 = ~n15400 ;
  assign y10504 = n19691 ;
  assign y10505 = ~1'b0 ;
  assign y10506 = ~1'b0 ;
  assign y10507 = n19692 ;
  assign y10508 = ~1'b0 ;
  assign y10509 = n19693 ;
  assign y10510 = n19694 ;
  assign y10511 = 1'b0 ;
  assign y10512 = ~n19696 ;
  assign y10513 = 1'b0 ;
  assign y10514 = ~n19697 ;
  assign y10515 = n19700 ;
  assign y10516 = ~n19702 ;
  assign y10517 = ~n19703 ;
  assign y10518 = n8003 ;
  assign y10519 = n19704 ;
  assign y10520 = ~n4870 ;
  assign y10521 = ~1'b0 ;
  assign y10522 = ~n19708 ;
  assign y10523 = n19711 ;
  assign y10524 = ~n19712 ;
  assign y10525 = ~n19713 ;
  assign y10526 = ~n19715 ;
  assign y10527 = 1'b0 ;
  assign y10528 = n19719 ;
  assign y10529 = n19720 ;
  assign y10530 = ~1'b0 ;
  assign y10531 = ~n19722 ;
  assign y10532 = ~n19724 ;
  assign y10533 = ~n19725 ;
  assign y10534 = ~n19728 ;
  assign y10535 = ~1'b0 ;
  assign y10536 = ~n19734 ;
  assign y10537 = ~1'b0 ;
  assign y10538 = ~1'b0 ;
  assign y10539 = ~1'b0 ;
  assign y10540 = ~n19735 ;
  assign y10541 = ~n19736 ;
  assign y10542 = n19737 ;
  assign y10543 = ~1'b0 ;
  assign y10544 = ~1'b0 ;
  assign y10545 = ~n19739 ;
  assign y10546 = ~1'b0 ;
  assign y10547 = ~1'b0 ;
  assign y10548 = ~1'b0 ;
  assign y10549 = ~n19740 ;
  assign y10550 = n19742 ;
  assign y10551 = ~n19747 ;
  assign y10552 = ~n3572 ;
  assign y10553 = ~n19749 ;
  assign y10554 = ~n11149 ;
  assign y10555 = ~n19751 ;
  assign y10556 = ~n19753 ;
  assign y10557 = n19756 ;
  assign y10558 = n19757 ;
  assign y10559 = ~n12336 ;
  assign y10560 = ~n19759 ;
  assign y10561 = n19165 ;
  assign y10562 = n19761 ;
  assign y10563 = ~n19763 ;
  assign y10564 = n19765 ;
  assign y10565 = ~n19768 ;
  assign y10566 = ~n19769 ;
  assign y10567 = ~1'b0 ;
  assign y10568 = ~n19771 ;
  assign y10569 = ~1'b0 ;
  assign y10570 = n19773 ;
  assign y10571 = ~n19775 ;
  assign y10572 = ~n4526 ;
  assign y10573 = n19778 ;
  assign y10574 = ~n19780 ;
  assign y10575 = n19784 ;
  assign y10576 = ~n19787 ;
  assign y10577 = ~n19791 ;
  assign y10578 = ~n19794 ;
  assign y10579 = ~n19795 ;
  assign y10580 = ~n19800 ;
  assign y10581 = ~n19806 ;
  assign y10582 = n19811 ;
  assign y10583 = ~1'b0 ;
  assign y10584 = n19814 ;
  assign y10585 = n19815 ;
  assign y10586 = ~n19822 ;
  assign y10587 = ~1'b0 ;
  assign y10588 = ~1'b0 ;
  assign y10589 = ~1'b0 ;
  assign y10590 = n19823 ;
  assign y10591 = ~n19824 ;
  assign y10592 = ~n19827 ;
  assign y10593 = ~n19828 ;
  assign y10594 = ~1'b0 ;
  assign y10595 = ~n19829 ;
  assign y10596 = ~n19831 ;
  assign y10597 = n19833 ;
  assign y10598 = ~n19835 ;
  assign y10599 = ~n19837 ;
  assign y10600 = n15002 ;
  assign y10601 = n19839 ;
  assign y10602 = ~n19840 ;
  assign y10603 = n19846 ;
  assign y10604 = ~1'b0 ;
  assign y10605 = ~1'b0 ;
  assign y10606 = ~1'b0 ;
  assign y10607 = n19848 ;
  assign y10608 = ~1'b0 ;
  assign y10609 = ~1'b0 ;
  assign y10610 = ~n19849 ;
  assign y10611 = ~1'b0 ;
  assign y10612 = n19852 ;
  assign y10613 = ~n18725 ;
  assign y10614 = ~n19854 ;
  assign y10615 = ~n19856 ;
  assign y10616 = ~1'b0 ;
  assign y10617 = n19857 ;
  assign y10618 = ~n19859 ;
  assign y10619 = ~n19864 ;
  assign y10620 = n1128 ;
  assign y10621 = ~n19866 ;
  assign y10622 = ~1'b0 ;
  assign y10623 = ~n19867 ;
  assign y10624 = n19870 ;
  assign y10625 = n19875 ;
  assign y10626 = n19876 ;
  assign y10627 = ~n19878 ;
  assign y10628 = ~n19879 ;
  assign y10629 = ~n19881 ;
  assign y10630 = n19882 ;
  assign y10631 = ~n19885 ;
  assign y10632 = ~1'b0 ;
  assign y10633 = n19887 ;
  assign y10634 = ~n19888 ;
  assign y10635 = ~n19890 ;
  assign y10636 = ~1'b0 ;
  assign y10637 = ~1'b0 ;
  assign y10638 = n19892 ;
  assign y10639 = ~n19894 ;
  assign y10640 = 1'b0 ;
  assign y10641 = ~1'b0 ;
  assign y10642 = ~n19898 ;
  assign y10643 = ~1'b0 ;
  assign y10644 = ~1'b0 ;
  assign y10645 = ~1'b0 ;
  assign y10646 = ~n19899 ;
  assign y10647 = n19905 ;
  assign y10648 = ~n19908 ;
  assign y10649 = ~n19909 ;
  assign y10650 = ~n19913 ;
  assign y10651 = n19919 ;
  assign y10652 = ~n8885 ;
  assign y10653 = ~n19921 ;
  assign y10654 = ~1'b0 ;
  assign y10655 = ~n19924 ;
  assign y10656 = ~n19928 ;
  assign y10657 = n16926 ;
  assign y10658 = ~1'b0 ;
  assign y10659 = ~n19931 ;
  assign y10660 = n19933 ;
  assign y10661 = ~n19942 ;
  assign y10662 = n19943 ;
  assign y10663 = ~n19944 ;
  assign y10664 = ~n19946 ;
  assign y10665 = ~n7408 ;
  assign y10666 = ~n19947 ;
  assign y10667 = n19950 ;
  assign y10668 = ~n19952 ;
  assign y10669 = n19954 ;
  assign y10670 = ~1'b0 ;
  assign y10671 = ~1'b0 ;
  assign y10672 = n19956 ;
  assign y10673 = ~1'b0 ;
  assign y10674 = ~n19962 ;
  assign y10675 = n10825 ;
  assign y10676 = ~1'b0 ;
  assign y10677 = n19964 ;
  assign y10678 = n19966 ;
  assign y10679 = n19967 ;
  assign y10680 = ~1'b0 ;
  assign y10681 = ~n19968 ;
  assign y10682 = ~n7100 ;
  assign y10683 = ~1'b0 ;
  assign y10684 = ~n19976 ;
  assign y10685 = n19978 ;
  assign y10686 = ~n19979 ;
  assign y10687 = ~n19980 ;
  assign y10688 = ~1'b0 ;
  assign y10689 = n19981 ;
  assign y10690 = ~n19982 ;
  assign y10691 = ~n19984 ;
  assign y10692 = ~1'b0 ;
  assign y10693 = ~n19987 ;
  assign y10694 = ~n19994 ;
  assign y10695 = ~n19998 ;
  assign y10696 = 1'b0 ;
  assign y10697 = ~n20008 ;
  assign y10698 = n14365 ;
  assign y10699 = ~1'b0 ;
  assign y10700 = ~n20009 ;
  assign y10701 = ~1'b0 ;
  assign y10702 = n20010 ;
  assign y10703 = ~n20011 ;
  assign y10704 = n20014 ;
  assign y10705 = ~n20034 ;
  assign y10706 = ~n20035 ;
  assign y10707 = ~n20038 ;
  assign y10708 = ~n20041 ;
  assign y10709 = n20042 ;
  assign y10710 = ~1'b0 ;
  assign y10711 = n20043 ;
  assign y10712 = ~n20044 ;
  assign y10713 = n20047 ;
  assign y10714 = n20049 ;
  assign y10715 = n20051 ;
  assign y10716 = ~1'b0 ;
  assign y10717 = ~n20052 ;
  assign y10718 = ~n20056 ;
  assign y10719 = n20057 ;
  assign y10720 = ~n20059 ;
  assign y10721 = ~1'b0 ;
  assign y10722 = n20060 ;
  assign y10723 = ~n20062 ;
  assign y10724 = ~1'b0 ;
  assign y10725 = ~1'b0 ;
  assign y10726 = ~n2062 ;
  assign y10727 = n20063 ;
  assign y10728 = ~1'b0 ;
  assign y10729 = n20066 ;
  assign y10730 = ~1'b0 ;
  assign y10731 = ~n20068 ;
  assign y10732 = n20069 ;
  assign y10733 = ~n20071 ;
  assign y10734 = ~1'b0 ;
  assign y10735 = ~n20074 ;
  assign y10736 = n20076 ;
  assign y10737 = ~1'b0 ;
  assign y10738 = ~n20077 ;
  assign y10739 = ~n20079 ;
  assign y10740 = ~n20081 ;
  assign y10741 = ~1'b0 ;
  assign y10742 = ~1'b0 ;
  assign y10743 = ~1'b0 ;
  assign y10744 = ~1'b0 ;
  assign y10745 = n20082 ;
  assign y10746 = ~n20086 ;
  assign y10747 = ~n20089 ;
  assign y10748 = ~n20092 ;
  assign y10749 = ~1'b0 ;
  assign y10750 = ~1'b0 ;
  assign y10751 = n20094 ;
  assign y10752 = ~1'b0 ;
  assign y10753 = ~n20095 ;
  assign y10754 = n20097 ;
  assign y10755 = ~1'b0 ;
  assign y10756 = ~n20098 ;
  assign y10757 = ~n17823 ;
  assign y10758 = ~1'b0 ;
  assign y10759 = ~1'b0 ;
  assign y10760 = ~n20099 ;
  assign y10761 = ~n20105 ;
  assign y10762 = ~n20106 ;
  assign y10763 = ~n20108 ;
  assign y10764 = ~n20111 ;
  assign y10765 = ~1'b0 ;
  assign y10766 = n20114 ;
  assign y10767 = ~1'b0 ;
  assign y10768 = ~1'b0 ;
  assign y10769 = ~1'b0 ;
  assign y10770 = n20120 ;
  assign y10771 = n20121 ;
  assign y10772 = ~n20122 ;
  assign y10773 = ~1'b0 ;
  assign y10774 = ~1'b0 ;
  assign y10775 = ~n20123 ;
  assign y10776 = ~n20125 ;
  assign y10777 = ~1'b0 ;
  assign y10778 = ~1'b0 ;
  assign y10779 = n20135 ;
  assign y10780 = ~1'b0 ;
  assign y10781 = ~1'b0 ;
  assign y10782 = n20136 ;
  assign y10783 = ~n20140 ;
  assign y10784 = ~n20145 ;
  assign y10785 = ~1'b0 ;
  assign y10786 = n20156 ;
  assign y10787 = ~n20162 ;
  assign y10788 = n20163 ;
  assign y10789 = ~1'b0 ;
  assign y10790 = ~1'b0 ;
  assign y10791 = ~1'b0 ;
  assign y10792 = ~1'b0 ;
  assign y10793 = n20165 ;
  assign y10794 = n20167 ;
  assign y10795 = n20168 ;
  assign y10796 = ~1'b0 ;
  assign y10797 = ~1'b0 ;
  assign y10798 = n20170 ;
  assign y10799 = ~n1424 ;
  assign y10800 = ~1'b0 ;
  assign y10801 = n16366 ;
  assign y10802 = ~1'b0 ;
  assign y10803 = n13523 ;
  assign y10804 = ~1'b0 ;
  assign y10805 = ~1'b0 ;
  assign y10806 = n11329 ;
  assign y10807 = ~n20173 ;
  assign y10808 = ~1'b0 ;
  assign y10809 = ~1'b0 ;
  assign y10810 = n20174 ;
  assign y10811 = ~n20177 ;
  assign y10812 = ~n20181 ;
  assign y10813 = n20184 ;
  assign y10814 = ~n20185 ;
  assign y10815 = n20187 ;
  assign y10816 = ~1'b0 ;
  assign y10817 = ~1'b0 ;
  assign y10818 = ~1'b0 ;
  assign y10819 = n20189 ;
  assign y10820 = ~n20194 ;
  assign y10821 = ~n20197 ;
  assign y10822 = ~n20198 ;
  assign y10823 = n20199 ;
  assign y10824 = n20200 ;
  assign y10825 = ~n20201 ;
  assign y10826 = ~1'b0 ;
  assign y10827 = ~n20204 ;
  assign y10828 = ~n20205 ;
  assign y10829 = ~n6841 ;
  assign y10830 = ~n593 ;
  assign y10831 = n20206 ;
  assign y10832 = ~n14248 ;
  assign y10833 = ~1'b0 ;
  assign y10834 = ~1'b0 ;
  assign y10835 = n20208 ;
  assign y10836 = ~n20213 ;
  assign y10837 = n20214 ;
  assign y10838 = ~n20216 ;
  assign y10839 = ~n20219 ;
  assign y10840 = ~1'b0 ;
  assign y10841 = n20220 ;
  assign y10842 = ~n20221 ;
  assign y10843 = n20222 ;
  assign y10844 = ~n20223 ;
  assign y10845 = n20224 ;
  assign y10846 = ~1'b0 ;
  assign y10847 = ~n8368 ;
  assign y10848 = ~1'b0 ;
  assign y10849 = ~n20228 ;
  assign y10850 = ~n1150 ;
  assign y10851 = n20242 ;
  assign y10852 = ~1'b0 ;
  assign y10853 = n20243 ;
  assign y10854 = ~n20246 ;
  assign y10855 = n20247 ;
  assign y10856 = ~1'b0 ;
  assign y10857 = n20248 ;
  assign y10858 = n20249 ;
  assign y10859 = 1'b0 ;
  assign y10860 = ~1'b0 ;
  assign y10861 = ~1'b0 ;
  assign y10862 = ~n20253 ;
  assign y10863 = ~n20258 ;
  assign y10864 = n20262 ;
  assign y10865 = ~1'b0 ;
  assign y10866 = n20263 ;
  assign y10867 = n20264 ;
  assign y10868 = n20266 ;
  assign y10869 = ~n20268 ;
  assign y10870 = ~1'b0 ;
  assign y10871 = n20272 ;
  assign y10872 = ~1'b0 ;
  assign y10873 = ~1'b0 ;
  assign y10874 = 1'b0 ;
  assign y10875 = ~n20273 ;
  assign y10876 = ~n20276 ;
  assign y10877 = n20279 ;
  assign y10878 = 1'b0 ;
  assign y10879 = n20283 ;
  assign y10880 = n20285 ;
  assign y10881 = n20287 ;
  assign y10882 = n20289 ;
  assign y10883 = n20290 ;
  assign y10884 = ~n20295 ;
  assign y10885 = ~n20296 ;
  assign y10886 = ~n20298 ;
  assign y10887 = n20299 ;
  assign y10888 = ~n20303 ;
  assign y10889 = ~1'b0 ;
  assign y10890 = n20307 ;
  assign y10891 = ~1'b0 ;
  assign y10892 = ~1'b0 ;
  assign y10893 = n20308 ;
  assign y10894 = n20309 ;
  assign y10895 = ~n20312 ;
  assign y10896 = ~n20313 ;
  assign y10897 = ~n20320 ;
  assign y10898 = n7444 ;
  assign y10899 = ~1'b0 ;
  assign y10900 = ~n20325 ;
  assign y10901 = ~n2412 ;
  assign y10902 = 1'b0 ;
  assign y10903 = ~n20326 ;
  assign y10904 = ~1'b0 ;
  assign y10905 = ~n20328 ;
  assign y10906 = ~1'b0 ;
  assign y10907 = ~1'b0 ;
  assign y10908 = n20333 ;
  assign y10909 = ~n20336 ;
  assign y10910 = ~n20340 ;
  assign y10911 = n20342 ;
  assign y10912 = n20343 ;
  assign y10913 = n20348 ;
  assign y10914 = n13539 ;
  assign y10915 = ~n20350 ;
  assign y10916 = n20355 ;
  assign y10917 = ~n20361 ;
  assign y10918 = ~1'b0 ;
  assign y10919 = ~n20368 ;
  assign y10920 = n20369 ;
  assign y10921 = ~n20371 ;
  assign y10922 = ~1'b0 ;
  assign y10923 = n20375 ;
  assign y10924 = ~1'b0 ;
  assign y10925 = ~1'b0 ;
  assign y10926 = ~1'b0 ;
  assign y10927 = ~1'b0 ;
  assign y10928 = ~1'b0 ;
  assign y10929 = ~n20376 ;
  assign y10930 = ~n20377 ;
  assign y10931 = n20380 ;
  assign y10932 = n20382 ;
  assign y10933 = ~1'b0 ;
  assign y10934 = ~n20384 ;
  assign y10935 = n20385 ;
  assign y10936 = n20387 ;
  assign y10937 = n20389 ;
  assign y10938 = ~n20390 ;
  assign y10939 = ~n20391 ;
  assign y10940 = ~1'b0 ;
  assign y10941 = ~n20394 ;
  assign y10942 = ~1'b0 ;
  assign y10943 = ~n20395 ;
  assign y10944 = ~n20398 ;
  assign y10945 = ~n20400 ;
  assign y10946 = ~1'b0 ;
  assign y10947 = n20401 ;
  assign y10948 = ~1'b0 ;
  assign y10949 = n20402 ;
  assign y10950 = ~n20405 ;
  assign y10951 = ~1'b0 ;
  assign y10952 = ~n8643 ;
  assign y10953 = n20407 ;
  assign y10954 = ~n20409 ;
  assign y10955 = n20412 ;
  assign y10956 = ~1'b0 ;
  assign y10957 = n20421 ;
  assign y10958 = ~n20422 ;
  assign y10959 = n2341 ;
  assign y10960 = ~n20425 ;
  assign y10961 = ~1'b0 ;
  assign y10962 = n20426 ;
  assign y10963 = ~1'b0 ;
  assign y10964 = n20428 ;
  assign y10965 = n20429 ;
  assign y10966 = n20433 ;
  assign y10967 = ~n3590 ;
  assign y10968 = ~1'b0 ;
  assign y10969 = ~1'b0 ;
  assign y10970 = ~n20434 ;
  assign y10971 = ~1'b0 ;
  assign y10972 = ~1'b0 ;
  assign y10973 = n20436 ;
  assign y10974 = ~n20438 ;
  assign y10975 = ~n20443 ;
  assign y10976 = ~n20444 ;
  assign y10977 = ~1'b0 ;
  assign y10978 = n20445 ;
  assign y10979 = ~n20448 ;
  assign y10980 = ~1'b0 ;
  assign y10981 = n20452 ;
  assign y10982 = n20454 ;
  assign y10983 = n20455 ;
  assign y10984 = ~n20456 ;
  assign y10985 = n20461 ;
  assign y10986 = n20462 ;
  assign y10987 = ~n20463 ;
  assign y10988 = ~1'b0 ;
  assign y10989 = n20467 ;
  assign y10990 = n20469 ;
  assign y10991 = ~1'b0 ;
  assign y10992 = n20471 ;
  assign y10993 = ~n20472 ;
  assign y10994 = n20473 ;
  assign y10995 = ~n9286 ;
  assign y10996 = ~n20475 ;
  assign y10997 = ~1'b0 ;
  assign y10998 = ~n4107 ;
  assign y10999 = ~1'b0 ;
  assign y11000 = n20476 ;
  assign y11001 = ~1'b0 ;
  assign y11002 = n20477 ;
  assign y11003 = ~n20479 ;
  assign y11004 = ~1'b0 ;
  assign y11005 = n20481 ;
  assign y11006 = ~1'b0 ;
  assign y11007 = ~1'b0 ;
  assign y11008 = ~n20482 ;
  assign y11009 = n20484 ;
  assign y11010 = n20486 ;
  assign y11011 = n20488 ;
  assign y11012 = ~1'b0 ;
  assign y11013 = n6643 ;
  assign y11014 = ~n20491 ;
  assign y11015 = ~n20492 ;
  assign y11016 = n20498 ;
  assign y11017 = n20500 ;
  assign y11018 = n20501 ;
  assign y11019 = ~1'b0 ;
  assign y11020 = ~n20503 ;
  assign y11021 = ~1'b0 ;
  assign y11022 = n1652 ;
  assign y11023 = ~n20506 ;
  assign y11024 = ~n20507 ;
  assign y11025 = ~n20508 ;
  assign y11026 = ~1'b0 ;
  assign y11027 = ~1'b0 ;
  assign y11028 = n20512 ;
  assign y11029 = ~1'b0 ;
  assign y11030 = ~1'b0 ;
  assign y11031 = ~n20514 ;
  assign y11032 = ~n20515 ;
  assign y11033 = ~1'b0 ;
  assign y11034 = ~n20516 ;
  assign y11035 = ~n20517 ;
  assign y11036 = ~n20518 ;
  assign y11037 = n20519 ;
  assign y11038 = n20523 ;
  assign y11039 = n20526 ;
  assign y11040 = n20530 ;
  assign y11041 = n20532 ;
  assign y11042 = n20534 ;
  assign y11043 = ~n20535 ;
  assign y11044 = n20536 ;
  assign y11045 = n20538 ;
  assign y11046 = ~1'b0 ;
  assign y11047 = n20541 ;
  assign y11048 = ~n20542 ;
  assign y11049 = ~n11404 ;
  assign y11050 = ~1'b0 ;
  assign y11051 = ~n20545 ;
  assign y11052 = ~1'b0 ;
  assign y11053 = n20547 ;
  assign y11054 = ~1'b0 ;
  assign y11055 = n20548 ;
  assign y11056 = ~n20551 ;
  assign y11057 = ~1'b0 ;
  assign y11058 = n20552 ;
  assign y11059 = n20559 ;
  assign y11060 = ~n20561 ;
  assign y11061 = ~n20563 ;
  assign y11062 = n20565 ;
  assign y11063 = ~1'b0 ;
  assign y11064 = n20568 ;
  assign y11065 = ~1'b0 ;
  assign y11066 = n20569 ;
  assign y11067 = n20575 ;
  assign y11068 = ~1'b0 ;
  assign y11069 = ~1'b0 ;
  assign y11070 = n20577 ;
  assign y11071 = n20579 ;
  assign y11072 = ~1'b0 ;
  assign y11073 = ~1'b0 ;
  assign y11074 = n6034 ;
  assign y11075 = ~n20580 ;
  assign y11076 = ~n20582 ;
  assign y11077 = ~1'b0 ;
  assign y11078 = ~n5002 ;
  assign y11079 = ~1'b0 ;
  assign y11080 = n20584 ;
  assign y11081 = ~n20588 ;
  assign y11082 = n20590 ;
  assign y11083 = n20593 ;
  assign y11084 = ~n20594 ;
  assign y11085 = ~n20596 ;
  assign y11086 = ~n20598 ;
  assign y11087 = ~1'b0 ;
  assign y11088 = ~n7241 ;
  assign y11089 = ~1'b0 ;
  assign y11090 = ~1'b0 ;
  assign y11091 = ~1'b0 ;
  assign y11092 = ~n20601 ;
  assign y11093 = n20603 ;
  assign y11094 = n20606 ;
  assign y11095 = n11237 ;
  assign y11096 = ~1'b0 ;
  assign y11097 = ~1'b0 ;
  assign y11098 = n20608 ;
  assign y11099 = ~n20611 ;
  assign y11100 = ~n20613 ;
  assign y11101 = n20614 ;
  assign y11102 = n20615 ;
  assign y11103 = n20618 ;
  assign y11104 = ~n648 ;
  assign y11105 = ~1'b0 ;
  assign y11106 = ~n11875 ;
  assign y11107 = n20619 ;
  assign y11108 = ~1'b0 ;
  assign y11109 = ~n20620 ;
  assign y11110 = ~1'b0 ;
  assign y11111 = ~n20623 ;
  assign y11112 = ~n11368 ;
  assign y11113 = ~n20624 ;
  assign y11114 = ~1'b0 ;
  assign y11115 = ~1'b0 ;
  assign y11116 = ~n20626 ;
  assign y11117 = n20627 ;
  assign y11118 = ~1'b0 ;
  assign y11119 = n20628 ;
  assign y11120 = ~n20629 ;
  assign y11121 = n20630 ;
  assign y11122 = n20631 ;
  assign y11123 = ~n17898 ;
  assign y11124 = ~1'b0 ;
  assign y11125 = 1'b0 ;
  assign y11126 = ~n20633 ;
  assign y11127 = n20634 ;
  assign y11128 = n20635 ;
  assign y11129 = n19071 ;
  assign y11130 = ~n20636 ;
  assign y11131 = n20640 ;
  assign y11132 = ~n20641 ;
  assign y11133 = ~n20643 ;
  assign y11134 = ~n20645 ;
  assign y11135 = ~n20647 ;
  assign y11136 = n20648 ;
  assign y11137 = n11351 ;
  assign y11138 = n20651 ;
  assign y11139 = ~n20654 ;
  assign y11140 = n3940 ;
  assign y11141 = ~1'b0 ;
  assign y11142 = ~1'b0 ;
  assign y11143 = ~1'b0 ;
  assign y11144 = ~n20662 ;
  assign y11145 = ~n20664 ;
  assign y11146 = n20668 ;
  assign y11147 = n20671 ;
  assign y11148 = ~n20673 ;
  assign y11149 = n20675 ;
  assign y11150 = n20677 ;
  assign y11151 = ~1'b0 ;
  assign y11152 = ~n20678 ;
  assign y11153 = ~n20682 ;
  assign y11154 = n20683 ;
  assign y11155 = ~n20686 ;
  assign y11156 = ~1'b0 ;
  assign y11157 = n1600 ;
  assign y11158 = ~n20689 ;
  assign y11159 = ~n20691 ;
  assign y11160 = ~1'b0 ;
  assign y11161 = ~n20692 ;
  assign y11162 = ~n20693 ;
  assign y11163 = ~n15131 ;
  assign y11164 = ~n20695 ;
  assign y11165 = ~n20696 ;
  assign y11166 = ~1'b0 ;
  assign y11167 = ~n20697 ;
  assign y11168 = n20699 ;
  assign y11169 = ~1'b0 ;
  assign y11170 = n1784 ;
  assign y11171 = ~n20701 ;
  assign y11172 = ~n8080 ;
  assign y11173 = ~1'b0 ;
  assign y11174 = ~1'b0 ;
  assign y11175 = ~n20706 ;
  assign y11176 = ~1'b0 ;
  assign y11177 = n20707 ;
  assign y11178 = ~n20709 ;
  assign y11179 = n20710 ;
  assign y11180 = n20715 ;
  assign y11181 = n20717 ;
  assign y11182 = n20718 ;
  assign y11183 = ~1'b0 ;
  assign y11184 = ~1'b0 ;
  assign y11185 = ~1'b0 ;
  assign y11186 = ~n20719 ;
  assign y11187 = ~n2434 ;
  assign y11188 = ~n20720 ;
  assign y11189 = ~n20722 ;
  assign y11190 = ~n20723 ;
  assign y11191 = n20724 ;
  assign y11192 = ~n20725 ;
  assign y11193 = n20729 ;
  assign y11194 = ~1'b0 ;
  assign y11195 = ~1'b0 ;
  assign y11196 = n20734 ;
  assign y11197 = n20736 ;
  assign y11198 = ~n20737 ;
  assign y11199 = n20738 ;
  assign y11200 = ~1'b0 ;
  assign y11201 = n20739 ;
  assign y11202 = ~n20741 ;
  assign y11203 = n19436 ;
  assign y11204 = ~1'b0 ;
  assign y11205 = ~n20745 ;
  assign y11206 = n20748 ;
  assign y11207 = 1'b0 ;
  assign y11208 = n20749 ;
  assign y11209 = ~n20751 ;
  assign y11210 = ~n20753 ;
  assign y11211 = ~1'b0 ;
  assign y11212 = ~1'b0 ;
  assign y11213 = ~n20757 ;
  assign y11214 = ~1'b0 ;
  assign y11215 = n13436 ;
  assign y11216 = ~n20759 ;
  assign y11217 = ~1'b0 ;
  assign y11218 = ~1'b0 ;
  assign y11219 = n20762 ;
  assign y11220 = ~1'b0 ;
  assign y11221 = ~n4440 ;
  assign y11222 = ~n18481 ;
  assign y11223 = n20763 ;
  assign y11224 = n20765 ;
  assign y11225 = 1'b0 ;
  assign y11226 = ~1'b0 ;
  assign y11227 = n20766 ;
  assign y11228 = ~n20771 ;
  assign y11229 = ~n20775 ;
  assign y11230 = ~n305 ;
  assign y11231 = ~n20777 ;
  assign y11232 = ~n20778 ;
  assign y11233 = ~n20781 ;
  assign y11234 = ~n20784 ;
  assign y11235 = ~1'b0 ;
  assign y11236 = ~1'b0 ;
  assign y11237 = ~1'b0 ;
  assign y11238 = n20785 ;
  assign y11239 = n11014 ;
  assign y11240 = 1'b0 ;
  assign y11241 = n20787 ;
  assign y11242 = ~n20789 ;
  assign y11243 = ~n20790 ;
  assign y11244 = n20791 ;
  assign y11245 = ~1'b0 ;
  assign y11246 = ~n20792 ;
  assign y11247 = ~1'b0 ;
  assign y11248 = ~1'b0 ;
  assign y11249 = n20795 ;
  assign y11250 = n20799 ;
  assign y11251 = ~n20800 ;
  assign y11252 = n20801 ;
  assign y11253 = ~1'b0 ;
  assign y11254 = ~n20805 ;
  assign y11255 = ~n4416 ;
  assign y11256 = 1'b0 ;
  assign y11257 = ~n20806 ;
  assign y11258 = n20808 ;
  assign y11259 = ~n20811 ;
  assign y11260 = n9178 ;
  assign y11261 = ~n20812 ;
  assign y11262 = ~1'b0 ;
  assign y11263 = ~n20813 ;
  assign y11264 = ~n20814 ;
  assign y11265 = ~1'b0 ;
  assign y11266 = ~n20817 ;
  assign y11267 = ~n20819 ;
  assign y11268 = ~n20820 ;
  assign y11269 = ~1'b0 ;
  assign y11270 = n20825 ;
  assign y11271 = n20826 ;
  assign y11272 = ~n20828 ;
  assign y11273 = n20829 ;
  assign y11274 = n20830 ;
  assign y11275 = ~1'b0 ;
  assign y11276 = n20831 ;
  assign y11277 = n20838 ;
  assign y11278 = ~n20839 ;
  assign y11279 = n20842 ;
  assign y11280 = ~n20844 ;
  assign y11281 = ~1'b0 ;
  assign y11282 = ~1'b0 ;
  assign y11283 = 1'b0 ;
  assign y11284 = ~1'b0 ;
  assign y11285 = ~1'b0 ;
  assign y11286 = ~n6386 ;
  assign y11287 = ~n20846 ;
  assign y11288 = ~n8062 ;
  assign y11289 = n20854 ;
  assign y11290 = n20856 ;
  assign y11291 = n20859 ;
  assign y11292 = ~1'b0 ;
  assign y11293 = ~n3726 ;
  assign y11294 = n20864 ;
  assign y11295 = n20866 ;
  assign y11296 = ~n20868 ;
  assign y11297 = ~n20872 ;
  assign y11298 = ~n20875 ;
  assign y11299 = ~n388 ;
  assign y11300 = ~1'b0 ;
  assign y11301 = ~1'b0 ;
  assign y11302 = ~n20878 ;
  assign y11303 = 1'b0 ;
  assign y11304 = n20880 ;
  assign y11305 = n20882 ;
  assign y11306 = ~n10699 ;
  assign y11307 = n20884 ;
  assign y11308 = n20886 ;
  assign y11309 = ~n20887 ;
  assign y11310 = ~n20888 ;
  assign y11311 = n20890 ;
  assign y11312 = n20891 ;
  assign y11313 = ~1'b0 ;
  assign y11314 = ~1'b0 ;
  assign y11315 = ~n20892 ;
  assign y11316 = ~n20893 ;
  assign y11317 = ~1'b0 ;
  assign y11318 = n20894 ;
  assign y11319 = n20898 ;
  assign y11320 = n20901 ;
  assign y11321 = ~n20903 ;
  assign y11322 = n20904 ;
  assign y11323 = n7851 ;
  assign y11324 = n20908 ;
  assign y11325 = ~1'b0 ;
  assign y11326 = 1'b0 ;
  assign y11327 = ~n8430 ;
  assign y11328 = ~n7019 ;
  assign y11329 = n20910 ;
  assign y11330 = n20915 ;
  assign y11331 = ~1'b0 ;
  assign y11332 = ~1'b0 ;
  assign y11333 = ~1'b0 ;
  assign y11334 = n20918 ;
  assign y11335 = n20920 ;
  assign y11336 = ~n20925 ;
  assign y11337 = ~n2278 ;
  assign y11338 = ~1'b0 ;
  assign y11339 = n20926 ;
  assign y11340 = ~n20929 ;
  assign y11341 = ~1'b0 ;
  assign y11342 = ~1'b0 ;
  assign y11343 = n20930 ;
  assign y11344 = n20932 ;
  assign y11345 = n20935 ;
  assign y11346 = ~1'b0 ;
  assign y11347 = ~1'b0 ;
  assign y11348 = n3904 ;
  assign y11349 = ~n20938 ;
  assign y11350 = n9876 ;
  assign y11351 = ~n20940 ;
  assign y11352 = ~n20942 ;
  assign y11353 = n20617 ;
  assign y11354 = ~1'b0 ;
  assign y11355 = ~1'b0 ;
  assign y11356 = ~n20945 ;
  assign y11357 = ~n20946 ;
  assign y11358 = ~1'b0 ;
  assign y11359 = ~1'b0 ;
  assign y11360 = n20950 ;
  assign y11361 = ~n20959 ;
  assign y11362 = ~1'b0 ;
  assign y11363 = ~n20960 ;
  assign y11364 = ~1'b0 ;
  assign y11365 = ~n20962 ;
  assign y11366 = ~1'b0 ;
  assign y11367 = ~n20964 ;
  assign y11368 = ~n20967 ;
  assign y11369 = n20968 ;
  assign y11370 = n20971 ;
  assign y11371 = ~1'b0 ;
  assign y11372 = n20972 ;
  assign y11373 = n20975 ;
  assign y11374 = n20977 ;
  assign y11375 = ~1'b0 ;
  assign y11376 = ~1'b0 ;
  assign y11377 = n20981 ;
  assign y11378 = n20982 ;
  assign y11379 = n20985 ;
  assign y11380 = ~1'b0 ;
  assign y11381 = ~1'b0 ;
  assign y11382 = ~n20987 ;
  assign y11383 = ~1'b0 ;
  assign y11384 = ~1'b0 ;
  assign y11385 = ~1'b0 ;
  assign y11386 = ~n20990 ;
  assign y11387 = ~1'b0 ;
  assign y11388 = ~n15176 ;
  assign y11389 = ~n20991 ;
  assign y11390 = ~n20993 ;
  assign y11391 = ~1'b0 ;
  assign y11392 = ~n1169 ;
  assign y11393 = n20994 ;
  assign y11394 = n20996 ;
  assign y11395 = n20997 ;
  assign y11396 = ~n21001 ;
  assign y11397 = ~n21002 ;
  assign y11398 = ~n20561 ;
  assign y11399 = n21008 ;
  assign y11400 = ~n21012 ;
  assign y11401 = ~1'b0 ;
  assign y11402 = ~n21015 ;
  assign y11403 = ~1'b0 ;
  assign y11404 = n21017 ;
  assign y11405 = n21019 ;
  assign y11406 = n21020 ;
  assign y11407 = ~1'b0 ;
  assign y11408 = n21021 ;
  assign y11409 = ~1'b0 ;
  assign y11410 = ~n21023 ;
  assign y11411 = ~1'b0 ;
  assign y11412 = n21024 ;
  assign y11413 = n4350 ;
  assign y11414 = ~n21027 ;
  assign y11415 = ~1'b0 ;
  assign y11416 = n6809 ;
  assign y11417 = n21029 ;
  assign y11418 = n21031 ;
  assign y11419 = ~1'b0 ;
  assign y11420 = ~n21033 ;
  assign y11421 = ~1'b0 ;
  assign y11422 = ~1'b0 ;
  assign y11423 = n21036 ;
  assign y11424 = ~n21037 ;
  assign y11425 = ~1'b0 ;
  assign y11426 = ~1'b0 ;
  assign y11427 = n21040 ;
  assign y11428 = ~1'b0 ;
  assign y11429 = n18067 ;
  assign y11430 = ~1'b0 ;
  assign y11431 = n21042 ;
  assign y11432 = ~n21045 ;
  assign y11433 = n21048 ;
  assign y11434 = n21049 ;
  assign y11435 = ~n21054 ;
  assign y11436 = ~1'b0 ;
  assign y11437 = ~n21058 ;
  assign y11438 = n1259 ;
  assign y11439 = ~n21059 ;
  assign y11440 = ~n21061 ;
  assign y11441 = ~1'b0 ;
  assign y11442 = ~n21065 ;
  assign y11443 = n21071 ;
  assign y11444 = n21075 ;
  assign y11445 = ~1'b0 ;
  assign y11446 = ~n21076 ;
  assign y11447 = ~n21077 ;
  assign y11448 = ~n21078 ;
  assign y11449 = ~n21079 ;
  assign y11450 = n21082 ;
  assign y11451 = ~1'b0 ;
  assign y11452 = n21084 ;
  assign y11453 = ~n21089 ;
  assign y11454 = n21090 ;
  assign y11455 = ~1'b0 ;
  assign y11456 = ~1'b0 ;
  assign y11457 = ~1'b0 ;
  assign y11458 = n21092 ;
  assign y11459 = ~1'b0 ;
  assign y11460 = ~1'b0 ;
  assign y11461 = n21094 ;
  assign y11462 = n21097 ;
  assign y11463 = ~n20084 ;
  assign y11464 = ~1'b0 ;
  assign y11465 = ~1'b0 ;
  assign y11466 = ~1'b0 ;
  assign y11467 = n21098 ;
  assign y11468 = ~1'b0 ;
  assign y11469 = n21101 ;
  assign y11470 = n21104 ;
  assign y11471 = ~1'b0 ;
  assign y11472 = ~n21109 ;
  assign y11473 = ~n21111 ;
  assign y11474 = ~n21112 ;
  assign y11475 = n21114 ;
  assign y11476 = ~n21117 ;
  assign y11477 = ~n21118 ;
  assign y11478 = ~n8543 ;
  assign y11479 = ~1'b0 ;
  assign y11480 = 1'b0 ;
  assign y11481 = ~n21119 ;
  assign y11482 = n21120 ;
  assign y11483 = 1'b0 ;
  assign y11484 = ~n21121 ;
  assign y11485 = ~1'b0 ;
  assign y11486 = ~n21123 ;
  assign y11487 = ~1'b0 ;
  assign y11488 = ~1'b0 ;
  assign y11489 = ~n21126 ;
  assign y11490 = ~n21128 ;
  assign y11491 = ~1'b0 ;
  assign y11492 = n21129 ;
  assign y11493 = n21131 ;
  assign y11494 = ~n21132 ;
  assign y11495 = ~n21133 ;
  assign y11496 = ~1'b0 ;
  assign y11497 = ~n21134 ;
  assign y11498 = ~1'b0 ;
  assign y11499 = n21136 ;
  assign y11500 = n21139 ;
  assign y11501 = n21141 ;
  assign y11502 = n21144 ;
  assign y11503 = ~1'b0 ;
  assign y11504 = ~1'b0 ;
  assign y11505 = ~n16974 ;
  assign y11506 = ~n21145 ;
  assign y11507 = ~n21147 ;
  assign y11508 = ~n21149 ;
  assign y11509 = ~1'b0 ;
  assign y11510 = ~1'b0 ;
  assign y11511 = ~1'b0 ;
  assign y11512 = ~1'b0 ;
  assign y11513 = n21150 ;
  assign y11514 = ~1'b0 ;
  assign y11515 = ~n21152 ;
  assign y11516 = n21154 ;
  assign y11517 = ~n21155 ;
  assign y11518 = n21158 ;
  assign y11519 = ~n21159 ;
  assign y11520 = n21161 ;
  assign y11521 = n20595 ;
  assign y11522 = n21164 ;
  assign y11523 = ~n2054 ;
  assign y11524 = n21166 ;
  assign y11525 = ~n21167 ;
  assign y11526 = ~n21169 ;
  assign y11527 = ~n21175 ;
  assign y11528 = ~1'b0 ;
  assign y11529 = n21176 ;
  assign y11530 = ~1'b0 ;
  assign y11531 = ~1'b0 ;
  assign y11532 = 1'b0 ;
  assign y11533 = n21181 ;
  assign y11534 = n21182 ;
  assign y11535 = 1'b0 ;
  assign y11536 = ~1'b0 ;
  assign y11537 = n21185 ;
  assign y11538 = ~1'b0 ;
  assign y11539 = n21188 ;
  assign y11540 = n21191 ;
  assign y11541 = n21192 ;
  assign y11542 = n21198 ;
  assign y11543 = n21199 ;
  assign y11544 = ~n21200 ;
  assign y11545 = ~1'b0 ;
  assign y11546 = ~1'b0 ;
  assign y11547 = ~1'b0 ;
  assign y11548 = ~n21202 ;
  assign y11549 = n21204 ;
  assign y11550 = ~1'b0 ;
  assign y11551 = n5431 ;
  assign y11552 = n21210 ;
  assign y11553 = ~1'b0 ;
  assign y11554 = ~1'b0 ;
  assign y11555 = 1'b0 ;
  assign y11556 = ~1'b0 ;
  assign y11557 = ~n21211 ;
  assign y11558 = ~n21212 ;
  assign y11559 = ~n21214 ;
  assign y11560 = ~1'b0 ;
  assign y11561 = ~1'b0 ;
  assign y11562 = n21215 ;
  assign y11563 = n21219 ;
  assign y11564 = ~1'b0 ;
  assign y11565 = n21221 ;
  assign y11566 = ~n21222 ;
  assign y11567 = n21224 ;
  assign y11568 = n7366 ;
  assign y11569 = n21225 ;
  assign y11570 = ~n21226 ;
  assign y11571 = ~1'b0 ;
  assign y11572 = n21228 ;
  assign y11573 = ~n21230 ;
  assign y11574 = 1'b0 ;
  assign y11575 = ~1'b0 ;
  assign y11576 = n21231 ;
  assign y11577 = n10880 ;
  assign y11578 = ~1'b0 ;
  assign y11579 = ~n7222 ;
  assign y11580 = ~1'b0 ;
  assign y11581 = ~n21232 ;
  assign y11582 = n21233 ;
  assign y11583 = n21234 ;
  assign y11584 = 1'b0 ;
  assign y11585 = ~n21238 ;
  assign y11586 = ~n21240 ;
  assign y11587 = ~1'b0 ;
  assign y11588 = ~1'b0 ;
  assign y11589 = n21241 ;
  assign y11590 = ~n21242 ;
  assign y11591 = n21243 ;
  assign y11592 = n21244 ;
  assign y11593 = ~n21247 ;
  assign y11594 = ~1'b0 ;
  assign y11595 = ~n21252 ;
  assign y11596 = ~1'b0 ;
  assign y11597 = n21258 ;
  assign y11598 = ~n21259 ;
  assign y11599 = ~1'b0 ;
  assign y11600 = ~n13170 ;
  assign y11601 = n1078 ;
  assign y11602 = n21260 ;
  assign y11603 = ~1'b0 ;
  assign y11604 = ~n21264 ;
  assign y11605 = ~n21266 ;
  assign y11606 = n21267 ;
  assign y11607 = n21270 ;
  assign y11608 = ~n21271 ;
  assign y11609 = ~1'b0 ;
  assign y11610 = n21275 ;
  assign y11611 = n21278 ;
  assign y11612 = ~n21283 ;
  assign y11613 = n21284 ;
  assign y11614 = ~n21288 ;
  assign y11615 = ~n2812 ;
  assign y11616 = n21289 ;
  assign y11617 = ~1'b0 ;
  assign y11618 = ~1'b0 ;
  assign y11619 = ~n21290 ;
  assign y11620 = ~1'b0 ;
  assign y11621 = ~n21300 ;
  assign y11622 = ~n21305 ;
  assign y11623 = n21315 ;
  assign y11624 = ~n21317 ;
  assign y11625 = ~1'b0 ;
  assign y11626 = ~1'b0 ;
  assign y11627 = ~n21318 ;
  assign y11628 = n21319 ;
  assign y11629 = ~1'b0 ;
  assign y11630 = n21327 ;
  assign y11631 = ~1'b0 ;
  assign y11632 = n21328 ;
  assign y11633 = n21330 ;
  assign y11634 = ~n21331 ;
  assign y11635 = ~1'b0 ;
  assign y11636 = ~1'b0 ;
  assign y11637 = ~1'b0 ;
  assign y11638 = 1'b0 ;
  assign y11639 = ~n21334 ;
  assign y11640 = n21335 ;
  assign y11641 = n21337 ;
  assign y11642 = ~n21342 ;
  assign y11643 = ~1'b0 ;
  assign y11644 = n21345 ;
  assign y11645 = ~1'b0 ;
  assign y11646 = ~n21349 ;
  assign y11647 = n21350 ;
  assign y11648 = n21356 ;
  assign y11649 = ~1'b0 ;
  assign y11650 = ~n21359 ;
  assign y11651 = ~n14321 ;
  assign y11652 = ~1'b0 ;
  assign y11653 = n21360 ;
  assign y11654 = ~1'b0 ;
  assign y11655 = n21361 ;
  assign y11656 = n21362 ;
  assign y11657 = ~n21363 ;
  assign y11658 = ~n14693 ;
  assign y11659 = ~1'b0 ;
  assign y11660 = ~1'b0 ;
  assign y11661 = ~n21365 ;
  assign y11662 = n21368 ;
  assign y11663 = ~1'b0 ;
  assign y11664 = n7192 ;
  assign y11665 = ~n21369 ;
  assign y11666 = ~n21371 ;
  assign y11667 = n21372 ;
  assign y11668 = n21374 ;
  assign y11669 = ~1'b0 ;
  assign y11670 = n21377 ;
  assign y11671 = ~1'b0 ;
  assign y11672 = n21387 ;
  assign y11673 = n21388 ;
  assign y11674 = n21389 ;
  assign y11675 = n21390 ;
  assign y11676 = ~n21393 ;
  assign y11677 = ~1'b0 ;
  assign y11678 = ~n13193 ;
  assign y11679 = n21395 ;
  assign y11680 = ~1'b0 ;
  assign y11681 = ~n21396 ;
  assign y11682 = ~1'b0 ;
  assign y11683 = ~1'b0 ;
  assign y11684 = n21397 ;
  assign y11685 = ~n21398 ;
  assign y11686 = ~n21404 ;
  assign y11687 = n21405 ;
  assign y11688 = n21406 ;
  assign y11689 = ~1'b0 ;
  assign y11690 = ~1'b0 ;
  assign y11691 = ~n17357 ;
  assign y11692 = n21408 ;
  assign y11693 = ~1'b0 ;
  assign y11694 = ~n21411 ;
  assign y11695 = ~n21412 ;
  assign y11696 = ~n21414 ;
  assign y11697 = ~n21422 ;
  assign y11698 = n21423 ;
  assign y11699 = ~n21424 ;
  assign y11700 = ~1'b0 ;
  assign y11701 = ~1'b0 ;
  assign y11702 = n21427 ;
  assign y11703 = ~n21430 ;
  assign y11704 = ~n21431 ;
  assign y11705 = ~1'b0 ;
  assign y11706 = ~n21432 ;
  assign y11707 = ~n21433 ;
  assign y11708 = ~n21436 ;
  assign y11709 = ~n21438 ;
  assign y11710 = ~1'b0 ;
  assign y11711 = ~1'b0 ;
  assign y11712 = ~n21441 ;
  assign y11713 = ~1'b0 ;
  assign y11714 = n21442 ;
  assign y11715 = ~n21444 ;
  assign y11716 = ~1'b0 ;
  assign y11717 = ~1'b0 ;
  assign y11718 = ~1'b0 ;
  assign y11719 = ~1'b0 ;
  assign y11720 = ~n21449 ;
  assign y11721 = ~1'b0 ;
  assign y11722 = ~1'b0 ;
  assign y11723 = n21452 ;
  assign y11724 = ~n21453 ;
  assign y11725 = ~n21455 ;
  assign y11726 = n21456 ;
  assign y11727 = n21462 ;
  assign y11728 = n21464 ;
  assign y11729 = n21470 ;
  assign y11730 = ~n21475 ;
  assign y11731 = n21477 ;
  assign y11732 = ~1'b0 ;
  assign y11733 = ~n21478 ;
  assign y11734 = n21480 ;
  assign y11735 = n21481 ;
  assign y11736 = ~n2066 ;
  assign y11737 = ~n21483 ;
  assign y11738 = ~n21484 ;
  assign y11739 = ~1'b0 ;
  assign y11740 = ~n21485 ;
  assign y11741 = n21487 ;
  assign y11742 = n21490 ;
  assign y11743 = n21494 ;
  assign y11744 = n21495 ;
  assign y11745 = n21496 ;
  assign y11746 = ~1'b0 ;
  assign y11747 = ~1'b0 ;
  assign y11748 = ~n21504 ;
  assign y11749 = n21511 ;
  assign y11750 = n21517 ;
  assign y11751 = n16585 ;
  assign y11752 = 1'b0 ;
  assign y11753 = ~n21518 ;
  assign y11754 = ~1'b0 ;
  assign y11755 = n21519 ;
  assign y11756 = ~1'b0 ;
  assign y11757 = ~1'b0 ;
  assign y11758 = ~n21520 ;
  assign y11759 = n21527 ;
  assign y11760 = ~n21530 ;
  assign y11761 = n21534 ;
  assign y11762 = ~1'b0 ;
  assign y11763 = ~n21535 ;
  assign y11764 = n21536 ;
  assign y11765 = ~1'b0 ;
  assign y11766 = ~1'b0 ;
  assign y11767 = n5622 ;
  assign y11768 = ~n21538 ;
  assign y11769 = ~n21539 ;
  assign y11770 = ~n21543 ;
  assign y11771 = 1'b0 ;
  assign y11772 = n21547 ;
  assign y11773 = ~1'b0 ;
  assign y11774 = ~1'b0 ;
  assign y11775 = n21553 ;
  assign y11776 = 1'b0 ;
  assign y11777 = n21554 ;
  assign y11778 = ~1'b0 ;
  assign y11779 = n21555 ;
  assign y11780 = ~1'b0 ;
  assign y11781 = ~1'b0 ;
  assign y11782 = ~1'b0 ;
  assign y11783 = ~1'b0 ;
  assign y11784 = ~n21556 ;
  assign y11785 = ~n21557 ;
  assign y11786 = ~n21558 ;
  assign y11787 = ~n21559 ;
  assign y11788 = n20801 ;
  assign y11789 = n21561 ;
  assign y11790 = n21565 ;
  assign y11791 = n21566 ;
  assign y11792 = ~n9000 ;
  assign y11793 = ~n21568 ;
  assign y11794 = ~1'b0 ;
  assign y11795 = ~n21571 ;
  assign y11796 = n9291 ;
  assign y11797 = n21573 ;
  assign y11798 = ~1'b0 ;
  assign y11799 = ~n21576 ;
  assign y11800 = ~n21579 ;
  assign y11801 = n10301 ;
  assign y11802 = ~1'b0 ;
  assign y11803 = ~1'b0 ;
  assign y11804 = ~n21580 ;
  assign y11805 = ~n21581 ;
  assign y11806 = n21582 ;
  assign y11807 = ~1'b0 ;
  assign y11808 = ~1'b0 ;
  assign y11809 = n21583 ;
  assign y11810 = ~1'b0 ;
  assign y11811 = n14576 ;
  assign y11812 = ~1'b0 ;
  assign y11813 = ~n14025 ;
  assign y11814 = ~n21585 ;
  assign y11815 = ~1'b0 ;
  assign y11816 = n21586 ;
  assign y11817 = ~1'b0 ;
  assign y11818 = ~1'b0 ;
  assign y11819 = ~n21587 ;
  assign y11820 = n21588 ;
  assign y11821 = ~1'b0 ;
  assign y11822 = ~1'b0 ;
  assign y11823 = ~n21589 ;
  assign y11824 = ~n1512 ;
  assign y11825 = ~n21593 ;
  assign y11826 = ~1'b0 ;
  assign y11827 = n7331 ;
  assign y11828 = n21594 ;
  assign y11829 = ~1'b0 ;
  assign y11830 = ~1'b0 ;
  assign y11831 = n21597 ;
  assign y11832 = n21600 ;
  assign y11833 = ~1'b0 ;
  assign y11834 = n21601 ;
  assign y11835 = n21602 ;
  assign y11836 = ~n21603 ;
  assign y11837 = ~1'b0 ;
  assign y11838 = ~n21605 ;
  assign y11839 = ~n21609 ;
  assign y11840 = ~n21612 ;
  assign y11841 = n21613 ;
  assign y11842 = ~n21618 ;
  assign y11843 = ~n21620 ;
  assign y11844 = n21626 ;
  assign y11845 = ~n21631 ;
  assign y11846 = ~1'b0 ;
  assign y11847 = 1'b0 ;
  assign y11848 = n21632 ;
  assign y11849 = n21633 ;
  assign y11850 = ~n21634 ;
  assign y11851 = ~n21636 ;
  assign y11852 = n21638 ;
  assign y11853 = n21639 ;
  assign y11854 = n21642 ;
  assign y11855 = ~n21644 ;
  assign y11856 = n21654 ;
  assign y11857 = ~1'b0 ;
  assign y11858 = ~1'b0 ;
  assign y11859 = ~1'b0 ;
  assign y11860 = n21656 ;
  assign y11861 = n21657 ;
  assign y11862 = n21658 ;
  assign y11863 = n21660 ;
  assign y11864 = ~1'b0 ;
  assign y11865 = ~n21666 ;
  assign y11866 = ~1'b0 ;
  assign y11867 = ~1'b0 ;
  assign y11868 = ~1'b0 ;
  assign y11869 = n21670 ;
  assign y11870 = 1'b0 ;
  assign y11871 = ~n3961 ;
  assign y11872 = n21680 ;
  assign y11873 = n21683 ;
  assign y11874 = ~1'b0 ;
  assign y11875 = ~1'b0 ;
  assign y11876 = ~n8468 ;
  assign y11877 = ~n21685 ;
  assign y11878 = ~n486 ;
  assign y11879 = n21688 ;
  assign y11880 = 1'b0 ;
  assign y11881 = n21690 ;
  assign y11882 = n21693 ;
  assign y11883 = n21695 ;
  assign y11884 = n21699 ;
  assign y11885 = n21700 ;
  assign y11886 = ~n21702 ;
  assign y11887 = ~n21704 ;
  assign y11888 = ~n21707 ;
  assign y11889 = ~1'b0 ;
  assign y11890 = n21710 ;
  assign y11891 = ~1'b0 ;
  assign y11892 = n21711 ;
  assign y11893 = ~1'b0 ;
  assign y11894 = n21713 ;
  assign y11895 = ~1'b0 ;
  assign y11896 = n21715 ;
  assign y11897 = ~1'b0 ;
  assign y11898 = n21717 ;
  assign y11899 = n21719 ;
  assign y11900 = n21722 ;
  assign y11901 = ~1'b0 ;
  assign y11902 = ~n21732 ;
  assign y11903 = n21737 ;
  assign y11904 = ~1'b0 ;
  assign y11905 = ~n21738 ;
  assign y11906 = ~1'b0 ;
  assign y11907 = n21740 ;
  assign y11908 = ~1'b0 ;
  assign y11909 = ~n21741 ;
  assign y11910 = ~n8023 ;
  assign y11911 = n21743 ;
  assign y11912 = ~1'b0 ;
  assign y11913 = ~n21744 ;
  assign y11914 = ~1'b0 ;
  assign y11915 = n12044 ;
  assign y11916 = ~n21752 ;
  assign y11917 = n21753 ;
  assign y11918 = ~n21754 ;
  assign y11919 = ~n21755 ;
  assign y11920 = ~n21756 ;
  assign y11921 = n21757 ;
  assign y11922 = 1'b0 ;
  assign y11923 = ~n21762 ;
  assign y11924 = ~n21765 ;
  assign y11925 = 1'b0 ;
  assign y11926 = ~n811 ;
  assign y11927 = ~1'b0 ;
  assign y11928 = ~n21766 ;
  assign y11929 = ~n21768 ;
  assign y11930 = ~1'b0 ;
  assign y11931 = ~1'b0 ;
  assign y11932 = ~1'b0 ;
  assign y11933 = ~1'b0 ;
  assign y11934 = n21771 ;
  assign y11935 = ~n21773 ;
  assign y11936 = ~1'b0 ;
  assign y11937 = ~n21778 ;
  assign y11938 = ~n21781 ;
  assign y11939 = n20727 ;
  assign y11940 = ~1'b0 ;
  assign y11941 = n21782 ;
  assign y11942 = ~n21784 ;
  assign y11943 = ~1'b0 ;
  assign y11944 = n1609 ;
  assign y11945 = ~n21790 ;
  assign y11946 = n21791 ;
  assign y11947 = n21792 ;
  assign y11948 = ~n21795 ;
  assign y11949 = ~n21796 ;
  assign y11950 = ~1'b0 ;
  assign y11951 = ~1'b0 ;
  assign y11952 = ~n21797 ;
  assign y11953 = ~1'b0 ;
  assign y11954 = ~n4012 ;
  assign y11955 = n21798 ;
  assign y11956 = n14091 ;
  assign y11957 = n21799 ;
  assign y11958 = ~1'b0 ;
  assign y11959 = ~1'b0 ;
  assign y11960 = ~n21802 ;
  assign y11961 = ~1'b0 ;
  assign y11962 = ~n21803 ;
  assign y11963 = ~1'b0 ;
  assign y11964 = ~1'b0 ;
  assign y11965 = n21805 ;
  assign y11966 = ~n21807 ;
  assign y11967 = ~n21808 ;
  assign y11968 = n21809 ;
  assign y11969 = ~1'b0 ;
  assign y11970 = n9242 ;
  assign y11971 = ~n21810 ;
  assign y11972 = n21811 ;
  assign y11973 = ~n21813 ;
  assign y11974 = n21815 ;
  assign y11975 = n21817 ;
  assign y11976 = n21818 ;
  assign y11977 = n21820 ;
  assign y11978 = ~1'b0 ;
  assign y11979 = ~1'b0 ;
  assign y11980 = n21821 ;
  assign y11981 = ~n21823 ;
  assign y11982 = ~n21825 ;
  assign y11983 = n21828 ;
  assign y11984 = 1'b0 ;
  assign y11985 = ~1'b0 ;
  assign y11986 = ~1'b0 ;
  assign y11987 = ~1'b0 ;
  assign y11988 = ~1'b0 ;
  assign y11989 = ~1'b0 ;
  assign y11990 = ~n21833 ;
  assign y11991 = ~n21834 ;
  assign y11992 = ~n21835 ;
  assign y11993 = ~n21836 ;
  assign y11994 = ~n21838 ;
  assign y11995 = n21839 ;
  assign y11996 = ~n21841 ;
  assign y11997 = n21844 ;
  assign y11998 = ~n21845 ;
  assign y11999 = n21847 ;
  assign y12000 = ~n21849 ;
  assign y12001 = n7465 ;
  assign y12002 = ~n21850 ;
  assign y12003 = n21854 ;
  assign y12004 = ~n21855 ;
  assign y12005 = n21858 ;
  assign y12006 = ~1'b0 ;
  assign y12007 = ~n21862 ;
  assign y12008 = ~n21865 ;
  assign y12009 = ~1'b0 ;
  assign y12010 = ~n21866 ;
  assign y12011 = n1247 ;
  assign y12012 = ~n21314 ;
  assign y12013 = ~n21867 ;
  assign y12014 = ~n21871 ;
  assign y12015 = ~1'b0 ;
  assign y12016 = ~n21874 ;
  assign y12017 = ~1'b0 ;
  assign y12018 = ~n21876 ;
  assign y12019 = n21877 ;
  assign y12020 = n21878 ;
  assign y12021 = ~n21879 ;
  assign y12022 = ~n21884 ;
  assign y12023 = ~1'b0 ;
  assign y12024 = ~n21885 ;
  assign y12025 = 1'b0 ;
  assign y12026 = ~1'b0 ;
  assign y12027 = ~1'b0 ;
  assign y12028 = n21887 ;
  assign y12029 = ~1'b0 ;
  assign y12030 = n21888 ;
  assign y12031 = n21889 ;
  assign y12032 = n21891 ;
  assign y12033 = ~1'b0 ;
  assign y12034 = ~n21892 ;
  assign y12035 = ~n21893 ;
  assign y12036 = ~n21897 ;
  assign y12037 = ~n21901 ;
  assign y12038 = n21902 ;
  assign y12039 = ~1'b0 ;
  assign y12040 = n21903 ;
  assign y12041 = ~n21907 ;
  assign y12042 = ~n11420 ;
  assign y12043 = ~1'b0 ;
  assign y12044 = ~n21908 ;
  assign y12045 = ~1'b0 ;
  assign y12046 = ~1'b0 ;
  assign y12047 = ~1'b0 ;
  assign y12048 = ~1'b0 ;
  assign y12049 = ~1'b0 ;
  assign y12050 = n21910 ;
  assign y12051 = n21912 ;
  assign y12052 = ~n21915 ;
  assign y12053 = ~n17353 ;
  assign y12054 = ~n21917 ;
  assign y12055 = ~n21920 ;
  assign y12056 = n21921 ;
  assign y12057 = ~1'b0 ;
  assign y12058 = ~1'b0 ;
  assign y12059 = n21922 ;
  assign y12060 = ~1'b0 ;
  assign y12061 = n21925 ;
  assign y12062 = ~n21927 ;
  assign y12063 = n21929 ;
  assign y12064 = ~1'b0 ;
  assign y12065 = n21931 ;
  assign y12066 = ~1'b0 ;
  assign y12067 = n21938 ;
  assign y12068 = n21942 ;
  assign y12069 = ~1'b0 ;
  assign y12070 = n21952 ;
  assign y12071 = ~n21961 ;
  assign y12072 = ~n21963 ;
  assign y12073 = n21966 ;
  assign y12074 = ~n21967 ;
  assign y12075 = ~1'b0 ;
  assign y12076 = ~n21968 ;
  assign y12077 = n21969 ;
  assign y12078 = ~n15759 ;
  assign y12079 = ~n21971 ;
  assign y12080 = n21972 ;
  assign y12081 = ~n21973 ;
  assign y12082 = ~n21974 ;
  assign y12083 = ~1'b0 ;
  assign y12084 = n21976 ;
  assign y12085 = ~n13786 ;
  assign y12086 = ~n16053 ;
  assign y12087 = 1'b0 ;
  assign y12088 = n21978 ;
  assign y12089 = ~n18305 ;
  assign y12090 = ~1'b0 ;
  assign y12091 = ~n21980 ;
  assign y12092 = ~n21982 ;
  assign y12093 = ~1'b0 ;
  assign y12094 = n21985 ;
  assign y12095 = n21986 ;
  assign y12096 = n21989 ;
  assign y12097 = ~n21990 ;
  assign y12098 = n21992 ;
  assign y12099 = n21995 ;
  assign y12100 = ~n7937 ;
  assign y12101 = n21996 ;
  assign y12102 = ~1'b0 ;
  assign y12103 = ~1'b0 ;
  assign y12104 = ~n21998 ;
  assign y12105 = ~1'b0 ;
  assign y12106 = n22002 ;
  assign y12107 = ~1'b0 ;
  assign y12108 = n22004 ;
  assign y12109 = ~1'b0 ;
  assign y12110 = ~n22008 ;
  assign y12111 = n22010 ;
  assign y12112 = ~n15012 ;
  assign y12113 = ~n22012 ;
  assign y12114 = ~n22014 ;
  assign y12115 = ~n22017 ;
  assign y12116 = n22019 ;
  assign y12117 = ~n22021 ;
  assign y12118 = ~n22025 ;
  assign y12119 = ~n22027 ;
  assign y12120 = ~n22028 ;
  assign y12121 = ~n22029 ;
  assign y12122 = n22034 ;
  assign y12123 = ~n22036 ;
  assign y12124 = ~n22038 ;
  assign y12125 = ~n22039 ;
  assign y12126 = ~n22042 ;
  assign y12127 = ~n22043 ;
  assign y12128 = ~1'b0 ;
  assign y12129 = ~n22044 ;
  assign y12130 = n22045 ;
  assign y12131 = ~1'b0 ;
  assign y12132 = ~n2912 ;
  assign y12133 = 1'b0 ;
  assign y12134 = n22046 ;
  assign y12135 = ~1'b0 ;
  assign y12136 = n22049 ;
  assign y12137 = n22051 ;
  assign y12138 = n22053 ;
  assign y12139 = ~1'b0 ;
  assign y12140 = ~n1425 ;
  assign y12141 = ~1'b0 ;
  assign y12142 = n22054 ;
  assign y12143 = ~1'b0 ;
  assign y12144 = ~n22058 ;
  assign y12145 = ~n22060 ;
  assign y12146 = ~n22061 ;
  assign y12147 = ~1'b0 ;
  assign y12148 = ~1'b0 ;
  assign y12149 = n14479 ;
  assign y12150 = ~n22065 ;
  assign y12151 = ~n22066 ;
  assign y12152 = ~1'b0 ;
  assign y12153 = ~1'b0 ;
  assign y12154 = ~1'b0 ;
  assign y12155 = ~n22067 ;
  assign y12156 = n22068 ;
  assign y12157 = ~1'b0 ;
  assign y12158 = n22069 ;
  assign y12159 = n10970 ;
  assign y12160 = ~1'b0 ;
  assign y12161 = n22072 ;
  assign y12162 = ~n22075 ;
  assign y12163 = ~n22078 ;
  assign y12164 = ~n7884 ;
  assign y12165 = ~n22081 ;
  assign y12166 = ~n22082 ;
  assign y12167 = ~1'b0 ;
  assign y12168 = ~n22084 ;
  assign y12169 = ~1'b0 ;
  assign y12170 = n22088 ;
  assign y12171 = n22089 ;
  assign y12172 = ~n22090 ;
  assign y12173 = ~1'b0 ;
  assign y12174 = ~n8895 ;
  assign y12175 = n22091 ;
  assign y12176 = ~n22092 ;
  assign y12177 = 1'b0 ;
  assign y12178 = n22093 ;
  assign y12179 = ~n22096 ;
  assign y12180 = ~n22098 ;
  assign y12181 = n2070 ;
  assign y12182 = n22100 ;
  assign y12183 = n13698 ;
  assign y12184 = n22104 ;
  assign y12185 = ~n22108 ;
  assign y12186 = ~1'b0 ;
  assign y12187 = ~n22110 ;
  assign y12188 = ~n4215 ;
  assign y12189 = ~n22111 ;
  assign y12190 = ~1'b0 ;
  assign y12191 = n22112 ;
  assign y12192 = n22118 ;
  assign y12193 = ~n22120 ;
  assign y12194 = ~n22127 ;
  assign y12195 = ~n3459 ;
  assign y12196 = ~n22128 ;
  assign y12197 = n22129 ;
  assign y12198 = ~n22130 ;
  assign y12199 = ~1'b0 ;
  assign y12200 = ~1'b0 ;
  assign y12201 = ~n22131 ;
  assign y12202 = ~n22135 ;
  assign y12203 = ~n22136 ;
  assign y12204 = ~n22138 ;
  assign y12205 = 1'b0 ;
  assign y12206 = ~1'b0 ;
  assign y12207 = ~n22141 ;
  assign y12208 = ~n22142 ;
  assign y12209 = ~n22144 ;
  assign y12210 = ~1'b0 ;
  assign y12211 = ~n22146 ;
  assign y12212 = ~1'b0 ;
  assign y12213 = ~n22150 ;
  assign y12214 = n22153 ;
  assign y12215 = n9320 ;
  assign y12216 = ~1'b0 ;
  assign y12217 = n22161 ;
  assign y12218 = ~1'b0 ;
  assign y12219 = ~n4632 ;
  assign y12220 = ~1'b0 ;
  assign y12221 = n22162 ;
  assign y12222 = n22164 ;
  assign y12223 = ~1'b0 ;
  assign y12224 = ~1'b0 ;
  assign y12225 = ~n22166 ;
  assign y12226 = n2718 ;
  assign y12227 = ~n22168 ;
  assign y12228 = ~n22170 ;
  assign y12229 = ~n22171 ;
  assign y12230 = ~n22173 ;
  assign y12231 = n22178 ;
  assign y12232 = ~n22180 ;
  assign y12233 = ~n22183 ;
  assign y12234 = ~1'b0 ;
  assign y12235 = n22186 ;
  assign y12236 = n22189 ;
  assign y12237 = ~n22202 ;
  assign y12238 = n22206 ;
  assign y12239 = n22210 ;
  assign y12240 = n22212 ;
  assign y12241 = ~n22216 ;
  assign y12242 = ~1'b0 ;
  assign y12243 = ~1'b0 ;
  assign y12244 = n22218 ;
  assign y12245 = ~n22221 ;
  assign y12246 = ~n22227 ;
  assign y12247 = ~n22229 ;
  assign y12248 = ~n22236 ;
  assign y12249 = n22241 ;
  assign y12250 = n22242 ;
  assign y12251 = ~n22243 ;
  assign y12252 = ~n22245 ;
  assign y12253 = ~n22249 ;
  assign y12254 = ~1'b0 ;
  assign y12255 = ~1'b0 ;
  assign y12256 = ~n22254 ;
  assign y12257 = ~n22255 ;
  assign y12258 = 1'b0 ;
  assign y12259 = ~1'b0 ;
  assign y12260 = ~n22260 ;
  assign y12261 = ~1'b0 ;
  assign y12262 = ~1'b0 ;
  assign y12263 = n22261 ;
  assign y12264 = ~n22263 ;
  assign y12265 = ~1'b0 ;
  assign y12266 = n22267 ;
  assign y12267 = n22269 ;
  assign y12268 = ~n8805 ;
  assign y12269 = ~1'b0 ;
  assign y12270 = n22271 ;
  assign y12271 = ~1'b0 ;
  assign y12272 = n22272 ;
  assign y12273 = n15681 ;
  assign y12274 = ~n22273 ;
  assign y12275 = ~1'b0 ;
  assign y12276 = n22274 ;
  assign y12277 = ~n22275 ;
  assign y12278 = ~n22276 ;
  assign y12279 = ~n22277 ;
  assign y12280 = ~1'b0 ;
  assign y12281 = n9151 ;
  assign y12282 = ~1'b0 ;
  assign y12283 = ~n22278 ;
  assign y12284 = ~n22282 ;
  assign y12285 = n22284 ;
  assign y12286 = ~1'b0 ;
  assign y12287 = ~1'b0 ;
  assign y12288 = ~n22288 ;
  assign y12289 = n22289 ;
  assign y12290 = ~1'b0 ;
  assign y12291 = ~n13024 ;
  assign y12292 = ~1'b0 ;
  assign y12293 = ~1'b0 ;
  assign y12294 = ~n22291 ;
  assign y12295 = ~n22292 ;
  assign y12296 = ~n22294 ;
  assign y12297 = ~1'b0 ;
  assign y12298 = ~n22298 ;
  assign y12299 = ~n22300 ;
  assign y12300 = ~1'b0 ;
  assign y12301 = ~1'b0 ;
  assign y12302 = ~n22302 ;
  assign y12303 = ~n22303 ;
  assign y12304 = n22307 ;
  assign y12305 = n22310 ;
  assign y12306 = ~n22313 ;
  assign y12307 = ~1'b0 ;
  assign y12308 = n22317 ;
  assign y12309 = n22319 ;
  assign y12310 = ~n22322 ;
  assign y12311 = n22323 ;
  assign y12312 = n22326 ;
  assign y12313 = ~n22327 ;
  assign y12314 = n22329 ;
  assign y12315 = n22330 ;
  assign y12316 = ~n22332 ;
  assign y12317 = n22339 ;
  assign y12318 = ~n22341 ;
  assign y12319 = ~1'b0 ;
  assign y12320 = 1'b0 ;
  assign y12321 = n22343 ;
  assign y12322 = n1679 ;
  assign y12323 = 1'b0 ;
  assign y12324 = n22346 ;
  assign y12325 = ~1'b0 ;
  assign y12326 = n3601 ;
  assign y12327 = ~1'b0 ;
  assign y12328 = ~n22347 ;
  assign y12329 = n22348 ;
  assign y12330 = ~n19661 ;
  assign y12331 = ~n22349 ;
  assign y12332 = n22351 ;
  assign y12333 = ~1'b0 ;
  assign y12334 = n22352 ;
  assign y12335 = ~1'b0 ;
  assign y12336 = ~n22353 ;
  assign y12337 = n22355 ;
  assign y12338 = n22358 ;
  assign y12339 = ~n22360 ;
  assign y12340 = ~n22362 ;
  assign y12341 = ~1'b0 ;
  assign y12342 = ~1'b0 ;
  assign y12343 = ~1'b0 ;
  assign y12344 = n18318 ;
  assign y12345 = n22365 ;
  assign y12346 = ~1'b0 ;
  assign y12347 = n22366 ;
  assign y12348 = ~n22370 ;
  assign y12349 = ~1'b0 ;
  assign y12350 = ~1'b0 ;
  assign y12351 = ~1'b0 ;
  assign y12352 = ~n2328 ;
  assign y12353 = n22371 ;
  assign y12354 = ~n22373 ;
  assign y12355 = n22375 ;
  assign y12356 = n22376 ;
  assign y12357 = ~n22377 ;
  assign y12358 = n14514 ;
  assign y12359 = n22378 ;
  assign y12360 = ~n16092 ;
  assign y12361 = n22381 ;
  assign y12362 = n22385 ;
  assign y12363 = 1'b0 ;
  assign y12364 = n22389 ;
  assign y12365 = ~n22396 ;
  assign y12366 = ~n22398 ;
  assign y12367 = n22399 ;
  assign y12368 = ~n22400 ;
  assign y12369 = ~1'b0 ;
  assign y12370 = ~n22402 ;
  assign y12371 = n22409 ;
  assign y12372 = n22411 ;
  assign y12373 = n22415 ;
  assign y12374 = n22416 ;
  assign y12375 = ~1'b0 ;
  assign y12376 = ~1'b0 ;
  assign y12377 = ~n3391 ;
  assign y12378 = n22418 ;
  assign y12379 = ~n22419 ;
  assign y12380 = ~1'b0 ;
  assign y12381 = ~1'b0 ;
  assign y12382 = ~1'b0 ;
  assign y12383 = ~1'b0 ;
  assign y12384 = ~1'b0 ;
  assign y12385 = n22420 ;
  assign y12386 = n22426 ;
  assign y12387 = n22427 ;
  assign y12388 = ~n22429 ;
  assign y12389 = ~1'b0 ;
  assign y12390 = n21106 ;
  assign y12391 = n22432 ;
  assign y12392 = ~1'b0 ;
  assign y12393 = n22434 ;
  assign y12394 = ~n22439 ;
  assign y12395 = ~n22440 ;
  assign y12396 = ~n22443 ;
  assign y12397 = ~n22445 ;
  assign y12398 = ~n22448 ;
  assign y12399 = n19459 ;
  assign y12400 = n22452 ;
  assign y12401 = ~n22455 ;
  assign y12402 = n2564 ;
  assign y12403 = ~1'b0 ;
  assign y12404 = ~n22458 ;
  assign y12405 = ~n22463 ;
  assign y12406 = ~1'b0 ;
  assign y12407 = ~n22467 ;
  assign y12408 = n22475 ;
  assign y12409 = ~n22476 ;
  assign y12410 = n22477 ;
  assign y12411 = 1'b0 ;
  assign y12412 = ~n22480 ;
  assign y12413 = ~1'b0 ;
  assign y12414 = ~n22483 ;
  assign y12415 = ~1'b0 ;
  assign y12416 = ~n6938 ;
  assign y12417 = n22484 ;
  assign y12418 = ~n22487 ;
  assign y12419 = n22489 ;
  assign y12420 = ~n22492 ;
  assign y12421 = n22496 ;
  assign y12422 = ~1'b0 ;
  assign y12423 = ~1'b0 ;
  assign y12424 = n22497 ;
  assign y12425 = ~1'b0 ;
  assign y12426 = ~n22499 ;
  assign y12427 = 1'b0 ;
  assign y12428 = n22502 ;
  assign y12429 = ~n22506 ;
  assign y12430 = ~1'b0 ;
  assign y12431 = n22508 ;
  assign y12432 = ~n22511 ;
  assign y12433 = ~n22512 ;
  assign y12434 = ~n12911 ;
  assign y12435 = 1'b0 ;
  assign y12436 = n22515 ;
  assign y12437 = ~1'b0 ;
  assign y12438 = n22516 ;
  assign y12439 = ~n16377 ;
  assign y12440 = n3193 ;
  assign y12441 = ~n22517 ;
  assign y12442 = n22520 ;
  assign y12443 = n22521 ;
  assign y12444 = ~1'b0 ;
  assign y12445 = n22522 ;
  assign y12446 = n645 ;
  assign y12447 = ~n22525 ;
  assign y12448 = ~n22526 ;
  assign y12449 = n22528 ;
  assign y12450 = ~n22529 ;
  assign y12451 = ~n22530 ;
  assign y12452 = ~n22531 ;
  assign y12453 = x34 ;
  assign y12454 = ~1'b0 ;
  assign y12455 = n22533 ;
  assign y12456 = ~n22536 ;
  assign y12457 = n22538 ;
  assign y12458 = ~n22540 ;
  assign y12459 = 1'b0 ;
  assign y12460 = ~n22541 ;
  assign y12461 = ~1'b0 ;
  assign y12462 = n22543 ;
  assign y12463 = ~1'b0 ;
  assign y12464 = ~1'b0 ;
  assign y12465 = ~n22544 ;
  assign y12466 = n12748 ;
  assign y12467 = ~n15223 ;
  assign y12468 = ~1'b0 ;
  assign y12469 = ~1'b0 ;
  assign y12470 = ~n22546 ;
  assign y12471 = ~n22548 ;
  assign y12472 = n22550 ;
  assign y12473 = ~n22553 ;
  assign y12474 = ~1'b0 ;
  assign y12475 = n22557 ;
  assign y12476 = ~1'b0 ;
  assign y12477 = n15736 ;
  assign y12478 = ~n22558 ;
  assign y12479 = ~n22560 ;
  assign y12480 = n22569 ;
  assign y12481 = ~1'b0 ;
  assign y12482 = ~n15404 ;
  assign y12483 = ~1'b0 ;
  assign y12484 = n3353 ;
  assign y12485 = n22570 ;
  assign y12486 = n22572 ;
  assign y12487 = ~n5576 ;
  assign y12488 = ~1'b0 ;
  assign y12489 = ~1'b0 ;
  assign y12490 = n22574 ;
  assign y12491 = n22576 ;
  assign y12492 = ~1'b0 ;
  assign y12493 = n4463 ;
  assign y12494 = n11228 ;
  assign y12495 = ~n22584 ;
  assign y12496 = n22587 ;
  assign y12497 = ~n22592 ;
  assign y12498 = ~n22595 ;
  assign y12499 = n22596 ;
  assign y12500 = n22599 ;
  assign y12501 = ~1'b0 ;
  assign y12502 = n22600 ;
  assign y12503 = ~1'b0 ;
  assign y12504 = n22601 ;
  assign y12505 = n22604 ;
  assign y12506 = n22606 ;
  assign y12507 = ~n22608 ;
  assign y12508 = ~n22609 ;
  assign y12509 = ~1'b0 ;
  assign y12510 = ~n22611 ;
  assign y12511 = n22613 ;
  assign y12512 = n22614 ;
  assign y12513 = ~n22615 ;
  assign y12514 = ~n14651 ;
  assign y12515 = ~1'b0 ;
  assign y12516 = n22616 ;
  assign y12517 = n10001 ;
  assign y12518 = ~1'b0 ;
  assign y12519 = n22618 ;
  assign y12520 = ~n22620 ;
  assign y12521 = n22624 ;
  assign y12522 = n22626 ;
  assign y12523 = ~n22627 ;
  assign y12524 = ~n22633 ;
  assign y12525 = ~1'b0 ;
  assign y12526 = ~1'b0 ;
  assign y12527 = ~1'b0 ;
  assign y12528 = ~n22634 ;
  assign y12529 = n22636 ;
  assign y12530 = ~1'b0 ;
  assign y12531 = ~n22638 ;
  assign y12532 = n22639 ;
  assign y12533 = n22640 ;
  assign y12534 = ~1'b0 ;
  assign y12535 = ~1'b0 ;
  assign y12536 = n22643 ;
  assign y12537 = ~n22644 ;
  assign y12538 = n22645 ;
  assign y12539 = ~n22648 ;
  assign y12540 = n22651 ;
  assign y12541 = ~1'b0 ;
  assign y12542 = ~1'b0 ;
  assign y12543 = n22652 ;
  assign y12544 = ~n22663 ;
  assign y12545 = ~n22666 ;
  assign y12546 = n6729 ;
  assign y12547 = ~n22673 ;
  assign y12548 = n22677 ;
  assign y12549 = ~n1819 ;
  assign y12550 = ~1'b0 ;
  assign y12551 = n22679 ;
  assign y12552 = ~n22680 ;
  assign y12553 = ~n22685 ;
  assign y12554 = ~n22689 ;
  assign y12555 = ~1'b0 ;
  assign y12556 = 1'b0 ;
  assign y12557 = ~1'b0 ;
  assign y12558 = ~n22690 ;
  assign y12559 = ~n22691 ;
  assign y12560 = 1'b0 ;
  assign y12561 = ~n22694 ;
  assign y12562 = ~n22695 ;
  assign y12563 = n22698 ;
  assign y12564 = ~n22700 ;
  assign y12565 = n12188 ;
  assign y12566 = n2973 ;
  assign y12567 = ~1'b0 ;
  assign y12568 = ~n22702 ;
  assign y12569 = ~1'b0 ;
  assign y12570 = ~n22711 ;
  assign y12571 = ~n22714 ;
  assign y12572 = ~n22715 ;
  assign y12573 = ~1'b0 ;
  assign y12574 = n22717 ;
  assign y12575 = ~1'b0 ;
  assign y12576 = ~1'b0 ;
  assign y12577 = ~1'b0 ;
  assign y12578 = ~1'b0 ;
  assign y12579 = ~n22719 ;
  assign y12580 = ~n22721 ;
  assign y12581 = n22727 ;
  assign y12582 = ~n22729 ;
  assign y12583 = n22730 ;
  assign y12584 = ~1'b0 ;
  assign y12585 = 1'b0 ;
  assign y12586 = n22734 ;
  assign y12587 = ~1'b0 ;
  assign y12588 = ~n22736 ;
  assign y12589 = ~n22739 ;
  assign y12590 = n22742 ;
  assign y12591 = ~1'b0 ;
  assign y12592 = ~n22744 ;
  assign y12593 = ~1'b0 ;
  assign y12594 = 1'b0 ;
  assign y12595 = n22745 ;
  assign y12596 = ~1'b0 ;
  assign y12597 = n22747 ;
  assign y12598 = n22748 ;
  assign y12599 = ~n22749 ;
  assign y12600 = n22750 ;
  assign y12601 = ~1'b0 ;
  assign y12602 = ~n22751 ;
  assign y12603 = ~1'b0 ;
  assign y12604 = ~n22752 ;
  assign y12605 = n22753 ;
  assign y12606 = ~1'b0 ;
  assign y12607 = ~1'b0 ;
  assign y12608 = ~1'b0 ;
  assign y12609 = ~n22756 ;
  assign y12610 = n22757 ;
  assign y12611 = n19521 ;
  assign y12612 = ~1'b0 ;
  assign y12613 = ~n17639 ;
  assign y12614 = ~n22759 ;
  assign y12615 = ~n22762 ;
  assign y12616 = ~1'b0 ;
  assign y12617 = n22763 ;
  assign y12618 = n22766 ;
  assign y12619 = n22768 ;
  assign y12620 = ~n22769 ;
  assign y12621 = n22770 ;
  assign y12622 = ~n22776 ;
  assign y12623 = ~1'b0 ;
  assign y12624 = ~1'b0 ;
  assign y12625 = n22778 ;
  assign y12626 = ~1'b0 ;
  assign y12627 = n22779 ;
  assign y12628 = ~1'b0 ;
  assign y12629 = ~1'b0 ;
  assign y12630 = n22783 ;
  assign y12631 = ~n22786 ;
  assign y12632 = ~n22788 ;
  assign y12633 = n22793 ;
  assign y12634 = n22795 ;
  assign y12635 = ~n22797 ;
  assign y12636 = n22800 ;
  assign y12637 = ~1'b0 ;
  assign y12638 = ~n22801 ;
  assign y12639 = n22802 ;
  assign y12640 = n22805 ;
  assign y12641 = ~n22807 ;
  assign y12642 = ~n22808 ;
  assign y12643 = ~1'b0 ;
  assign y12644 = ~1'b0 ;
  assign y12645 = ~n22809 ;
  assign y12646 = ~1'b0 ;
  assign y12647 = n22811 ;
  assign y12648 = ~n22813 ;
  assign y12649 = ~1'b0 ;
  assign y12650 = ~n22815 ;
  assign y12651 = n22818 ;
  assign y12652 = ~1'b0 ;
  assign y12653 = ~n22822 ;
  assign y12654 = n22823 ;
  assign y12655 = ~1'b0 ;
  assign y12656 = ~n22827 ;
  assign y12657 = n22833 ;
  assign y12658 = ~1'b0 ;
  assign y12659 = n22834 ;
  assign y12660 = ~n22835 ;
  assign y12661 = n22836 ;
  assign y12662 = ~n22838 ;
  assign y12663 = n22840 ;
  assign y12664 = n2635 ;
  assign y12665 = ~1'b0 ;
  assign y12666 = ~n22841 ;
  assign y12667 = ~1'b0 ;
  assign y12668 = n22843 ;
  assign y12669 = n22845 ;
  assign y12670 = ~n22846 ;
  assign y12671 = n1056 ;
  assign y12672 = ~n3056 ;
  assign y12673 = n22848 ;
  assign y12674 = ~1'b0 ;
  assign y12675 = n22850 ;
  assign y12676 = 1'b0 ;
  assign y12677 = n22854 ;
  assign y12678 = ~1'b0 ;
  assign y12679 = ~1'b0 ;
  assign y12680 = ~n22858 ;
  assign y12681 = ~n22860 ;
  assign y12682 = ~1'b0 ;
  assign y12683 = ~n22863 ;
  assign y12684 = n22865 ;
  assign y12685 = n22866 ;
  assign y12686 = ~1'b0 ;
  assign y12687 = ~n22870 ;
  assign y12688 = 1'b0 ;
  assign y12689 = n1465 ;
  assign y12690 = n22871 ;
  assign y12691 = n22873 ;
  assign y12692 = ~n22874 ;
  assign y12693 = ~n22879 ;
  assign y12694 = ~n22880 ;
  assign y12695 = ~n22887 ;
  assign y12696 = ~n22890 ;
  assign y12697 = ~1'b0 ;
  assign y12698 = ~n22892 ;
  assign y12699 = ~1'b0 ;
  assign y12700 = n10865 ;
  assign y12701 = ~n19896 ;
  assign y12702 = n22893 ;
  assign y12703 = ~n22896 ;
  assign y12704 = ~n22899 ;
  assign y12705 = ~n22900 ;
  assign y12706 = ~n22905 ;
  assign y12707 = ~1'b0 ;
  assign y12708 = ~1'b0 ;
  assign y12709 = ~1'b0 ;
  assign y12710 = n22909 ;
  assign y12711 = ~1'b0 ;
  assign y12712 = n22910 ;
  assign y12713 = ~1'b0 ;
  assign y12714 = ~n22911 ;
  assign y12715 = ~n22914 ;
  assign y12716 = ~1'b0 ;
  assign y12717 = n22916 ;
  assign y12718 = ~1'b0 ;
  assign y12719 = ~1'b0 ;
  assign y12720 = ~1'b0 ;
  assign y12721 = n4269 ;
  assign y12722 = ~n22917 ;
  assign y12723 = ~n22918 ;
  assign y12724 = ~1'b0 ;
  assign y12725 = n22920 ;
  assign y12726 = n22922 ;
  assign y12727 = ~n22923 ;
  assign y12728 = ~n22925 ;
  assign y12729 = ~n17421 ;
  assign y12730 = ~1'b0 ;
  assign y12731 = ~1'b0 ;
  assign y12732 = n22926 ;
  assign y12733 = ~1'b0 ;
  assign y12734 = ~1'b0 ;
  assign y12735 = ~1'b0 ;
  assign y12736 = ~n22927 ;
  assign y12737 = ~1'b0 ;
  assign y12738 = ~n22932 ;
  assign y12739 = ~n22933 ;
  assign y12740 = ~n22935 ;
  assign y12741 = ~n22937 ;
  assign y12742 = ~n22939 ;
  assign y12743 = ~n22940 ;
  assign y12744 = ~1'b0 ;
  assign y12745 = n22941 ;
  assign y12746 = ~1'b0 ;
  assign y12747 = ~n22945 ;
  assign y12748 = ~1'b0 ;
  assign y12749 = ~1'b0 ;
  assign y12750 = ~n22947 ;
  assign y12751 = ~1'b0 ;
  assign y12752 = ~n22948 ;
  assign y12753 = ~n22949 ;
  assign y12754 = n22951 ;
  assign y12755 = ~1'b0 ;
  assign y12756 = ~n22953 ;
  assign y12757 = ~1'b0 ;
  assign y12758 = n22955 ;
  assign y12759 = ~n22956 ;
  assign y12760 = ~1'b0 ;
  assign y12761 = ~1'b0 ;
  assign y12762 = ~n22957 ;
  assign y12763 = ~1'b0 ;
  assign y12764 = ~n22958 ;
  assign y12765 = n22959 ;
  assign y12766 = ~n22961 ;
  assign y12767 = n22962 ;
  assign y12768 = n2154 ;
  assign y12769 = ~1'b0 ;
  assign y12770 = ~n22964 ;
  assign y12771 = ~1'b0 ;
  assign y12772 = n22965 ;
  assign y12773 = ~n22970 ;
  assign y12774 = n22974 ;
  assign y12775 = n22975 ;
  assign y12776 = ~1'b0 ;
  assign y12777 = ~n22977 ;
  assign y12778 = ~1'b0 ;
  assign y12779 = ~1'b0 ;
  assign y12780 = n22979 ;
  assign y12781 = n22981 ;
  assign y12782 = n22983 ;
  assign y12783 = ~n22985 ;
  assign y12784 = ~1'b0 ;
  assign y12785 = ~1'b0 ;
  assign y12786 = ~1'b0 ;
  assign y12787 = ~1'b0 ;
  assign y12788 = n22986 ;
  assign y12789 = ~n22988 ;
  assign y12790 = ~n22989 ;
  assign y12791 = n3700 ;
  assign y12792 = ~n22990 ;
  assign y12793 = ~n13147 ;
  assign y12794 = ~n22992 ;
  assign y12795 = ~n22994 ;
  assign y12796 = ~1'b0 ;
  assign y12797 = ~1'b0 ;
  assign y12798 = ~1'b0 ;
  assign y12799 = ~n22064 ;
  assign y12800 = ~n22999 ;
  assign y12801 = n23001 ;
  assign y12802 = ~n23006 ;
  assign y12803 = n23008 ;
  assign y12804 = ~n981 ;
  assign y12805 = ~n23009 ;
  assign y12806 = ~n23010 ;
  assign y12807 = n23011 ;
  assign y12808 = n23013 ;
  assign y12809 = ~n23017 ;
  assign y12810 = ~n23018 ;
  assign y12811 = ~n23019 ;
  assign y12812 = ~n23024 ;
  assign y12813 = ~1'b0 ;
  assign y12814 = n23027 ;
  assign y12815 = n23028 ;
  assign y12816 = ~1'b0 ;
  assign y12817 = n2479 ;
  assign y12818 = ~n23033 ;
  assign y12819 = ~n23034 ;
  assign y12820 = n23035 ;
  assign y12821 = n23037 ;
  assign y12822 = n23039 ;
  assign y12823 = ~n23041 ;
  assign y12824 = ~n23043 ;
  assign y12825 = ~n23046 ;
  assign y12826 = n23047 ;
  assign y12827 = ~n14253 ;
  assign y12828 = n23049 ;
  assign y12829 = ~1'b0 ;
  assign y12830 = ~n23050 ;
  assign y12831 = n23051 ;
  assign y12832 = ~1'b0 ;
  assign y12833 = ~1'b0 ;
  assign y12834 = ~n23052 ;
  assign y12835 = ~1'b0 ;
  assign y12836 = ~n23054 ;
  assign y12837 = 1'b0 ;
  assign y12838 = ~1'b0 ;
  assign y12839 = n14935 ;
  assign y12840 = ~n23058 ;
  assign y12841 = n23059 ;
  assign y12842 = ~n23064 ;
  assign y12843 = ~1'b0 ;
  assign y12844 = n23066 ;
  assign y12845 = n18279 ;
  assign y12846 = n11420 ;
  assign y12847 = ~1'b0 ;
  assign y12848 = ~1'b0 ;
  assign y12849 = ~1'b0 ;
  assign y12850 = n23067 ;
  assign y12851 = n23074 ;
  assign y12852 = ~n23075 ;
  assign y12853 = n23081 ;
  assign y12854 = ~n23085 ;
  assign y12855 = ~1'b0 ;
  assign y12856 = n23086 ;
  assign y12857 = ~n14185 ;
  assign y12858 = ~n11704 ;
  assign y12859 = ~n23088 ;
  assign y12860 = ~1'b0 ;
  assign y12861 = n23093 ;
  assign y12862 = ~n23094 ;
  assign y12863 = n23096 ;
  assign y12864 = n23101 ;
  assign y12865 = ~n9529 ;
  assign y12866 = ~1'b0 ;
  assign y12867 = n23105 ;
  assign y12868 = ~n23106 ;
  assign y12869 = n23109 ;
  assign y12870 = n23111 ;
  assign y12871 = ~1'b0 ;
  assign y12872 = ~n23113 ;
  assign y12873 = n23116 ;
  assign y12874 = n23117 ;
  assign y12875 = ~1'b0 ;
  assign y12876 = n12573 ;
  assign y12877 = n4707 ;
  assign y12878 = n23118 ;
  assign y12879 = ~n23120 ;
  assign y12880 = ~1'b0 ;
  assign y12881 = n23122 ;
  assign y12882 = n20781 ;
  assign y12883 = n23123 ;
  assign y12884 = n23129 ;
  assign y12885 = n23131 ;
  assign y12886 = n23134 ;
  assign y12887 = n23135 ;
  assign y12888 = ~1'b0 ;
  assign y12889 = ~1'b0 ;
  assign y12890 = n23136 ;
  assign y12891 = n23138 ;
  assign y12892 = n23147 ;
  assign y12893 = n23149 ;
  assign y12894 = ~n23150 ;
  assign y12895 = ~n23152 ;
  assign y12896 = n23154 ;
  assign y12897 = n23160 ;
  assign y12898 = n23165 ;
  assign y12899 = ~n23168 ;
  assign y12900 = ~1'b0 ;
  assign y12901 = ~n23172 ;
  assign y12902 = ~1'b0 ;
  assign y12903 = ~n23174 ;
  assign y12904 = ~1'b0 ;
  assign y12905 = ~1'b0 ;
  assign y12906 = n23175 ;
  assign y12907 = ~1'b0 ;
  assign y12908 = n23176 ;
  assign y12909 = n23177 ;
  assign y12910 = 1'b0 ;
  assign y12911 = n23179 ;
  assign y12912 = ~n23186 ;
  assign y12913 = ~1'b0 ;
  assign y12914 = ~1'b0 ;
  assign y12915 = ~n150 ;
  assign y12916 = ~n23187 ;
  assign y12917 = ~n23189 ;
  assign y12918 = ~n12392 ;
  assign y12919 = n23191 ;
  assign y12920 = n12520 ;
  assign y12921 = n23193 ;
  assign y12922 = ~n23195 ;
  assign y12923 = n23198 ;
  assign y12924 = ~1'b0 ;
  assign y12925 = ~n23202 ;
  assign y12926 = n23204 ;
  assign y12927 = ~n15662 ;
  assign y12928 = ~1'b0 ;
  assign y12929 = n23205 ;
  assign y12930 = n23207 ;
  assign y12931 = n23208 ;
  assign y12932 = ~n23213 ;
  assign y12933 = 1'b0 ;
  assign y12934 = ~1'b0 ;
  assign y12935 = ~1'b0 ;
  assign y12936 = n23215 ;
  assign y12937 = ~n23216 ;
  assign y12938 = ~n23217 ;
  assign y12939 = ~n23218 ;
  assign y12940 = ~1'b0 ;
  assign y12941 = ~n23220 ;
  assign y12942 = n23221 ;
  assign y12943 = n23226 ;
  assign y12944 = ~1'b0 ;
  assign y12945 = ~1'b0 ;
  assign y12946 = ~n4884 ;
  assign y12947 = ~1'b0 ;
  assign y12948 = ~n23227 ;
  assign y12949 = ~n23228 ;
  assign y12950 = ~1'b0 ;
  assign y12951 = 1'b0 ;
  assign y12952 = n4793 ;
  assign y12953 = ~1'b0 ;
  assign y12954 = n23234 ;
  assign y12955 = ~n23235 ;
  assign y12956 = n23241 ;
  assign y12957 = n23244 ;
  assign y12958 = 1'b0 ;
  assign y12959 = ~n23246 ;
  assign y12960 = n5011 ;
  assign y12961 = ~1'b0 ;
  assign y12962 = ~1'b0 ;
  assign y12963 = ~1'b0 ;
  assign y12964 = n20900 ;
  assign y12965 = n15759 ;
  assign y12966 = ~n2330 ;
  assign y12967 = ~n23248 ;
  assign y12968 = ~n5966 ;
  assign y12969 = n3853 ;
  assign y12970 = ~n14694 ;
  assign y12971 = ~n23251 ;
  assign y12972 = ~1'b0 ;
  assign y12973 = ~n23256 ;
  assign y12974 = n23258 ;
  assign y12975 = ~1'b0 ;
  assign y12976 = ~1'b0 ;
  assign y12977 = ~1'b0 ;
  assign y12978 = n23260 ;
  assign y12979 = n23264 ;
  assign y12980 = n23266 ;
  assign y12981 = n5605 ;
  assign y12982 = ~1'b0 ;
  assign y12983 = n23267 ;
  assign y12984 = ~1'b0 ;
  assign y12985 = ~1'b0 ;
  assign y12986 = n23269 ;
  assign y12987 = n12735 ;
  assign y12988 = n4138 ;
  assign y12989 = n23270 ;
  assign y12990 = ~n23271 ;
  assign y12991 = n23273 ;
  assign y12992 = ~n23276 ;
  assign y12993 = ~n23279 ;
  assign y12994 = ~1'b0 ;
  assign y12995 = n23282 ;
  assign y12996 = n4931 ;
  assign y12997 = ~1'b0 ;
  assign y12998 = ~n23286 ;
  assign y12999 = ~n8847 ;
  assign y13000 = 1'b0 ;
  assign y13001 = n23287 ;
  assign y13002 = n23290 ;
  assign y13003 = n23291 ;
  assign y13004 = ~1'b0 ;
  assign y13005 = ~1'b0 ;
  assign y13006 = ~n23293 ;
  assign y13007 = ~1'b0 ;
  assign y13008 = n23295 ;
  assign y13009 = n2874 ;
  assign y13010 = 1'b0 ;
  assign y13011 = ~n23296 ;
  assign y13012 = ~n23297 ;
  assign y13013 = ~n23299 ;
  assign y13014 = n23300 ;
  assign y13015 = n23302 ;
  assign y13016 = n4266 ;
  assign y13017 = ~1'b0 ;
  assign y13018 = ~1'b0 ;
  assign y13019 = ~n23303 ;
  assign y13020 = ~n23304 ;
  assign y13021 = n23306 ;
  assign y13022 = ~n23308 ;
  assign y13023 = ~1'b0 ;
  assign y13024 = ~n23312 ;
  assign y13025 = n23313 ;
  assign y13026 = n23315 ;
  assign y13027 = ~n23318 ;
  assign y13028 = ~n23320 ;
  assign y13029 = 1'b0 ;
  assign y13030 = ~n23321 ;
  assign y13031 = n23325 ;
  assign y13032 = n23327 ;
  assign y13033 = n6850 ;
  assign y13034 = ~n23329 ;
  assign y13035 = n23331 ;
  assign y13036 = ~n23332 ;
  assign y13037 = ~1'b0 ;
  assign y13038 = ~1'b0 ;
  assign y13039 = n23336 ;
  assign y13040 = ~n23338 ;
  assign y13041 = n23340 ;
  assign y13042 = ~n3010 ;
  assign y13043 = n23341 ;
  assign y13044 = ~1'b0 ;
  assign y13045 = ~n11880 ;
  assign y13046 = ~n23342 ;
  assign y13047 = ~1'b0 ;
  assign y13048 = ~1'b0 ;
  assign y13049 = ~n6038 ;
  assign y13050 = ~n23345 ;
  assign y13051 = ~n755 ;
  assign y13052 = n23346 ;
  assign y13053 = n23348 ;
  assign y13054 = ~n23349 ;
  assign y13055 = ~1'b0 ;
  assign y13056 = ~1'b0 ;
  assign y13057 = n23350 ;
  assign y13058 = ~1'b0 ;
  assign y13059 = ~1'b0 ;
  assign y13060 = ~1'b0 ;
  assign y13061 = ~n23351 ;
  assign y13062 = ~n23356 ;
  assign y13063 = n23357 ;
  assign y13064 = 1'b0 ;
  assign y13065 = n23359 ;
  assign y13066 = ~n23361 ;
  assign y13067 = n23365 ;
  assign y13068 = ~1'b0 ;
  assign y13069 = n23367 ;
  assign y13070 = 1'b0 ;
  assign y13071 = n23370 ;
  assign y13072 = ~n23372 ;
  assign y13073 = ~n23373 ;
  assign y13074 = ~1'b0 ;
  assign y13075 = ~1'b0 ;
  assign y13076 = ~1'b0 ;
  assign y13077 = ~n23376 ;
  assign y13078 = n23377 ;
  assign y13079 = n9749 ;
  assign y13080 = ~n23380 ;
  assign y13081 = ~1'b0 ;
  assign y13082 = n23381 ;
  assign y13083 = ~n23383 ;
  assign y13084 = n23384 ;
  assign y13085 = n23386 ;
  assign y13086 = n23388 ;
  assign y13087 = ~n23390 ;
  assign y13088 = ~1'b0 ;
  assign y13089 = ~1'b0 ;
  assign y13090 = n23391 ;
  assign y13091 = n23394 ;
  assign y13092 = ~1'b0 ;
  assign y13093 = ~n23395 ;
  assign y13094 = ~n23396 ;
  assign y13095 = n3041 ;
  assign y13096 = ~1'b0 ;
  assign y13097 = ~n23401 ;
  assign y13098 = ~n23402 ;
  assign y13099 = ~n23404 ;
  assign y13100 = ~1'b0 ;
  assign y13101 = n23406 ;
  assign y13102 = n23407 ;
  assign y13103 = ~n23408 ;
  assign y13104 = ~1'b0 ;
  assign y13105 = ~n23409 ;
  assign y13106 = ~n23411 ;
  assign y13107 = ~n23415 ;
  assign y13108 = ~1'b0 ;
  assign y13109 = ~n5261 ;
  assign y13110 = ~n23416 ;
  assign y13111 = ~1'b0 ;
  assign y13112 = 1'b0 ;
  assign y13113 = ~n23418 ;
  assign y13114 = ~n23420 ;
  assign y13115 = ~n23421 ;
  assign y13116 = n23422 ;
  assign y13117 = ~n23424 ;
  assign y13118 = n5329 ;
  assign y13119 = n23426 ;
  assign y13120 = ~n5109 ;
  assign y13121 = ~1'b0 ;
  assign y13122 = ~n23427 ;
  assign y13123 = ~n23431 ;
  assign y13124 = ~1'b0 ;
  assign y13125 = ~n23432 ;
  assign y13126 = ~n23433 ;
  assign y13127 = n23435 ;
  assign y13128 = ~1'b0 ;
  assign y13129 = ~1'b0 ;
  assign y13130 = ~n23437 ;
  assign y13131 = n23441 ;
  assign y13132 = ~1'b0 ;
  assign y13133 = n23442 ;
  assign y13134 = ~1'b0 ;
  assign y13135 = ~n23446 ;
  assign y13136 = ~1'b0 ;
  assign y13137 = n23450 ;
  assign y13138 = n23451 ;
  assign y13139 = n23452 ;
  assign y13140 = ~1'b0 ;
  assign y13141 = ~n21786 ;
  assign y13142 = ~1'b0 ;
  assign y13143 = n23453 ;
  assign y13144 = ~1'b0 ;
  assign y13145 = ~1'b0 ;
  assign y13146 = ~1'b0 ;
  assign y13147 = ~n23455 ;
  assign y13148 = n23457 ;
  assign y13149 = ~n23458 ;
  assign y13150 = ~n23461 ;
  assign y13151 = n23463 ;
  assign y13152 = ~1'b0 ;
  assign y13153 = ~1'b0 ;
  assign y13154 = ~1'b0 ;
  assign y13155 = n23466 ;
  assign y13156 = ~1'b0 ;
  assign y13157 = ~1'b0 ;
  assign y13158 = ~n23468 ;
  assign y13159 = n23475 ;
  assign y13160 = ~n23476 ;
  assign y13161 = 1'b0 ;
  assign y13162 = 1'b0 ;
  assign y13163 = ~1'b0 ;
  assign y13164 = ~n23478 ;
  assign y13165 = ~n23479 ;
  assign y13166 = ~1'b0 ;
  assign y13167 = ~n23480 ;
  assign y13168 = ~n23483 ;
  assign y13169 = ~n2417 ;
  assign y13170 = ~n23484 ;
  assign y13171 = ~1'b0 ;
  assign y13172 = n23485 ;
  assign y13173 = n15791 ;
  assign y13174 = ~1'b0 ;
  assign y13175 = ~n23486 ;
  assign y13176 = n23488 ;
  assign y13177 = n23490 ;
  assign y13178 = ~1'b0 ;
  assign y13179 = n23491 ;
  assign y13180 = ~1'b0 ;
  assign y13181 = ~n1937 ;
  assign y13182 = ~1'b0 ;
  assign y13183 = ~n23492 ;
  assign y13184 = n23502 ;
  assign y13185 = ~1'b0 ;
  assign y13186 = ~1'b0 ;
  assign y13187 = n23504 ;
  assign y13188 = ~1'b0 ;
  assign y13189 = n23506 ;
  assign y13190 = ~n23510 ;
  assign y13191 = n23511 ;
  assign y13192 = ~1'b0 ;
  assign y13193 = ~1'b0 ;
  assign y13194 = ~n23513 ;
  assign y13195 = ~1'b0 ;
  assign y13196 = ~1'b0 ;
  assign y13197 = n23514 ;
  assign y13198 = ~n23516 ;
  assign y13199 = ~n23523 ;
  assign y13200 = ~n23524 ;
  assign y13201 = n23525 ;
  assign y13202 = n23528 ;
  assign y13203 = ~1'b0 ;
  assign y13204 = ~n23529 ;
  assign y13205 = n23531 ;
  assign y13206 = ~1'b0 ;
  assign y13207 = ~1'b0 ;
  assign y13208 = n23533 ;
  assign y13209 = n23535 ;
  assign y13210 = n23536 ;
  assign y13211 = n12355 ;
  assign y13212 = ~n23540 ;
  assign y13213 = ~1'b0 ;
  assign y13214 = n23542 ;
  assign y13215 = ~n23544 ;
  assign y13216 = n23546 ;
  assign y13217 = ~1'b0 ;
  assign y13218 = ~1'b0 ;
  assign y13219 = ~n21797 ;
  assign y13220 = ~1'b0 ;
  assign y13221 = ~n23549 ;
  assign y13222 = ~n23551 ;
  assign y13223 = ~n23552 ;
  assign y13224 = n23554 ;
  assign y13225 = ~n23557 ;
  assign y13226 = ~1'b0 ;
  assign y13227 = ~1'b0 ;
  assign y13228 = ~n23560 ;
  assign y13229 = n23563 ;
  assign y13230 = n23573 ;
  assign y13231 = ~n23577 ;
  assign y13232 = n23578 ;
  assign y13233 = ~n23579 ;
  assign y13234 = ~n23582 ;
  assign y13235 = n23585 ;
  assign y13236 = ~n23586 ;
  assign y13237 = ~n23588 ;
  assign y13238 = ~1'b0 ;
  assign y13239 = ~n10244 ;
  assign y13240 = ~1'b0 ;
  assign y13241 = ~1'b0 ;
  assign y13242 = n23591 ;
  assign y13243 = 1'b0 ;
  assign y13244 = ~n23593 ;
  assign y13245 = n23597 ;
  assign y13246 = ~1'b0 ;
  assign y13247 = ~1'b0 ;
  assign y13248 = ~1'b0 ;
  assign y13249 = ~1'b0 ;
  assign y13250 = ~n23599 ;
  assign y13251 = ~n3533 ;
  assign y13252 = ~n23601 ;
  assign y13253 = ~1'b0 ;
  assign y13254 = n23602 ;
  assign y13255 = ~n23607 ;
  assign y13256 = ~1'b0 ;
  assign y13257 = ~n23611 ;
  assign y13258 = n23612 ;
  assign y13259 = ~n14772 ;
  assign y13260 = n23617 ;
  assign y13261 = n21981 ;
  assign y13262 = ~n23619 ;
  assign y13263 = n23621 ;
  assign y13264 = n23622 ;
  assign y13265 = ~n23627 ;
  assign y13266 = n23629 ;
  assign y13267 = n23635 ;
  assign y13268 = n23636 ;
  assign y13269 = ~n23640 ;
  assign y13270 = ~1'b0 ;
  assign y13271 = 1'b0 ;
  assign y13272 = ~1'b0 ;
  assign y13273 = n23641 ;
  assign y13274 = ~1'b0 ;
  assign y13275 = ~n23644 ;
  assign y13276 = n23647 ;
  assign y13277 = ~1'b0 ;
  assign y13278 = ~n23648 ;
  assign y13279 = n13433 ;
  assign y13280 = n23649 ;
  assign y13281 = ~1'b0 ;
  assign y13282 = n23651 ;
  assign y13283 = n23652 ;
  assign y13284 = 1'b0 ;
  assign y13285 = n23654 ;
  assign y13286 = n23501 ;
  assign y13287 = ~n23656 ;
  assign y13288 = n23657 ;
  assign y13289 = ~1'b0 ;
  assign y13290 = ~1'b0 ;
  assign y13291 = ~n4586 ;
  assign y13292 = n23661 ;
  assign y13293 = ~1'b0 ;
  assign y13294 = n23664 ;
  assign y13295 = n23666 ;
  assign y13296 = ~n23671 ;
  assign y13297 = n23676 ;
  assign y13298 = ~n23681 ;
  assign y13299 = ~1'b0 ;
  assign y13300 = n23684 ;
  assign y13301 = n23690 ;
  assign y13302 = ~n23692 ;
  assign y13303 = n23693 ;
  assign y13304 = n23695 ;
  assign y13305 = n23701 ;
  assign y13306 = n23702 ;
  assign y13307 = ~n23703 ;
  assign y13308 = n23707 ;
  assign y13309 = ~n2743 ;
  assign y13310 = ~1'b0 ;
  assign y13311 = n23711 ;
  assign y13312 = ~1'b0 ;
  assign y13313 = ~n23712 ;
  assign y13314 = n23713 ;
  assign y13315 = 1'b0 ;
  assign y13316 = ~n23715 ;
  assign y13317 = n23722 ;
  assign y13318 = n23723 ;
  assign y13319 = ~n23725 ;
  assign y13320 = ~1'b0 ;
  assign y13321 = 1'b0 ;
  assign y13322 = ~n23726 ;
  assign y13323 = ~n23727 ;
  assign y13324 = ~n5062 ;
  assign y13325 = n672 ;
  assign y13326 = ~n23732 ;
  assign y13327 = ~n15508 ;
  assign y13328 = ~n23735 ;
  assign y13329 = ~n23737 ;
  assign y13330 = n23739 ;
  assign y13331 = ~1'b0 ;
  assign y13332 = ~1'b0 ;
  assign y13333 = ~1'b0 ;
  assign y13334 = ~n23741 ;
  assign y13335 = ~n23744 ;
  assign y13336 = ~n23746 ;
  assign y13337 = ~1'b0 ;
  assign y13338 = n23747 ;
  assign y13339 = ~1'b0 ;
  assign y13340 = ~1'b0 ;
  assign y13341 = ~n23749 ;
  assign y13342 = ~n23751 ;
  assign y13343 = ~n23755 ;
  assign y13344 = n23757 ;
  assign y13345 = n23758 ;
  assign y13346 = ~1'b0 ;
  assign y13347 = n23760 ;
  assign y13348 = n23769 ;
  assign y13349 = n23773 ;
  assign y13350 = ~1'b0 ;
  assign y13351 = n23774 ;
  assign y13352 = n2945 ;
  assign y13353 = ~n23779 ;
  assign y13354 = ~n23780 ;
  assign y13355 = ~n23782 ;
  assign y13356 = ~n23783 ;
  assign y13357 = ~n23785 ;
  assign y13358 = ~1'b0 ;
  assign y13359 = ~n23787 ;
  assign y13360 = n23790 ;
  assign y13361 = ~n23791 ;
  assign y13362 = ~n23792 ;
  assign y13363 = n23794 ;
  assign y13364 = ~n23795 ;
  assign y13365 = ~1'b0 ;
  assign y13366 = n14317 ;
  assign y13367 = ~1'b0 ;
  assign y13368 = ~n23798 ;
  assign y13369 = ~n23804 ;
  assign y13370 = ~n23806 ;
  assign y13371 = ~1'b0 ;
  assign y13372 = ~n23807 ;
  assign y13373 = ~n23810 ;
  assign y13374 = ~n23812 ;
  assign y13375 = n23814 ;
  assign y13376 = ~n23816 ;
  assign y13377 = ~1'b0 ;
  assign y13378 = ~n23818 ;
  assign y13379 = ~n21099 ;
  assign y13380 = ~1'b0 ;
  assign y13381 = n3877 ;
  assign y13382 = ~1'b0 ;
  assign y13383 = ~n23821 ;
  assign y13384 = n23822 ;
  assign y13385 = ~1'b0 ;
  assign y13386 = n23823 ;
  assign y13387 = ~n23827 ;
  assign y13388 = n23828 ;
  assign y13389 = n23829 ;
  assign y13390 = ~n23830 ;
  assign y13391 = ~1'b0 ;
  assign y13392 = ~1'b0 ;
  assign y13393 = ~1'b0 ;
  assign y13394 = n23832 ;
  assign y13395 = n23833 ;
  assign y13396 = ~1'b0 ;
  assign y13397 = ~n765 ;
  assign y13398 = ~1'b0 ;
  assign y13399 = ~n23835 ;
  assign y13400 = ~n23836 ;
  assign y13401 = ~1'b0 ;
  assign y13402 = ~n23838 ;
  assign y13403 = n23842 ;
  assign y13404 = ~n23849 ;
  assign y13405 = ~n23851 ;
  assign y13406 = ~n23854 ;
  assign y13407 = ~n23856 ;
  assign y13408 = ~n23858 ;
  assign y13409 = ~1'b0 ;
  assign y13410 = ~1'b0 ;
  assign y13411 = ~n23864 ;
  assign y13412 = n23867 ;
  assign y13413 = ~n23868 ;
  assign y13414 = ~n23869 ;
  assign y13415 = ~n23870 ;
  assign y13416 = ~n23871 ;
  assign y13417 = n5357 ;
  assign y13418 = n23872 ;
  assign y13419 = ~1'b0 ;
  assign y13420 = n23874 ;
  assign y13421 = ~1'b0 ;
  assign y13422 = n23875 ;
  assign y13423 = ~n430 ;
  assign y13424 = n23880 ;
  assign y13425 = n23882 ;
  assign y13426 = ~n23887 ;
  assign y13427 = ~n23888 ;
  assign y13428 = ~n23889 ;
  assign y13429 = ~1'b0 ;
  assign y13430 = ~n23892 ;
  assign y13431 = ~n23896 ;
  assign y13432 = ~1'b0 ;
  assign y13433 = ~1'b0 ;
  assign y13434 = ~n23898 ;
  assign y13435 = ~1'b0 ;
  assign y13436 = ~n23900 ;
  assign y13437 = ~1'b0 ;
  assign y13438 = n23901 ;
  assign y13439 = ~n23902 ;
  assign y13440 = ~1'b0 ;
  assign y13441 = ~n23908 ;
  assign y13442 = n23909 ;
  assign y13443 = ~1'b0 ;
  assign y13444 = ~n23910 ;
  assign y13445 = ~1'b0 ;
  assign y13446 = n23913 ;
  assign y13447 = ~n23914 ;
  assign y13448 = ~n23917 ;
  assign y13449 = ~n23919 ;
  assign y13450 = ~1'b0 ;
  assign y13451 = ~1'b0 ;
  assign y13452 = ~n23921 ;
  assign y13453 = ~1'b0 ;
  assign y13454 = ~n23928 ;
  assign y13455 = ~n23931 ;
  assign y13456 = n23933 ;
  assign y13457 = n23935 ;
  assign y13458 = n23936 ;
  assign y13459 = ~n23940 ;
  assign y13460 = n23941 ;
  assign y13461 = n23943 ;
  assign y13462 = ~n23945 ;
  assign y13463 = ~n23946 ;
  assign y13464 = ~n23949 ;
  assign y13465 = ~n23951 ;
  assign y13466 = n20757 ;
  assign y13467 = n23956 ;
  assign y13468 = ~n23957 ;
  assign y13469 = ~n23961 ;
  assign y13470 = n23962 ;
  assign y13471 = n21409 ;
  assign y13472 = n23963 ;
  assign y13473 = ~1'b0 ;
  assign y13474 = ~n23964 ;
  assign y13475 = ~1'b0 ;
  assign y13476 = ~1'b0 ;
  assign y13477 = ~n23966 ;
  assign y13478 = ~1'b0 ;
  assign y13479 = ~n23969 ;
  assign y13480 = ~1'b0 ;
  assign y13481 = ~n23970 ;
  assign y13482 = ~n23972 ;
  assign y13483 = n23975 ;
  assign y13484 = ~1'b0 ;
  assign y13485 = ~n23977 ;
  assign y13486 = ~1'b0 ;
  assign y13487 = n6862 ;
  assign y13488 = n23982 ;
  assign y13489 = n23984 ;
  assign y13490 = n23985 ;
  assign y13491 = ~1'b0 ;
  assign y13492 = ~n23987 ;
  assign y13493 = ~n23991 ;
  assign y13494 = n23994 ;
  assign y13495 = ~1'b0 ;
  assign y13496 = ~n23996 ;
  assign y13497 = ~n23997 ;
  assign y13498 = n24000 ;
  assign y13499 = ~1'b0 ;
  assign y13500 = ~n24003 ;
  assign y13501 = n24005 ;
  assign y13502 = ~n24007 ;
  assign y13503 = n24010 ;
  assign y13504 = n24012 ;
  assign y13505 = n24014 ;
  assign y13506 = ~1'b0 ;
  assign y13507 = ~n24016 ;
  assign y13508 = n24017 ;
  assign y13509 = n24021 ;
  assign y13510 = n8483 ;
  assign y13511 = n24025 ;
  assign y13512 = ~1'b0 ;
  assign y13513 = ~n24028 ;
  assign y13514 = n24029 ;
  assign y13515 = ~n5822 ;
  assign y13516 = ~n24030 ;
  assign y13517 = ~1'b0 ;
  assign y13518 = n24034 ;
  assign y13519 = n24035 ;
  assign y13520 = n24037 ;
  assign y13521 = n24041 ;
  assign y13522 = ~n24043 ;
  assign y13523 = ~n487 ;
  assign y13524 = n11892 ;
  assign y13525 = ~n24046 ;
  assign y13526 = n24047 ;
  assign y13527 = n24049 ;
  assign y13528 = ~1'b0 ;
  assign y13529 = n4786 ;
  assign y13530 = ~n24050 ;
  assign y13531 = ~n19957 ;
  assign y13532 = ~n2150 ;
  assign y13533 = n24054 ;
  assign y13534 = n24058 ;
  assign y13535 = n24059 ;
  assign y13536 = ~n24060 ;
  assign y13537 = n24061 ;
  assign y13538 = ~n9261 ;
  assign y13539 = ~1'b0 ;
  assign y13540 = ~n24063 ;
  assign y13541 = ~1'b0 ;
  assign y13542 = ~1'b0 ;
  assign y13543 = ~1'b0 ;
  assign y13544 = ~1'b0 ;
  assign y13545 = ~1'b0 ;
  assign y13546 = n24064 ;
  assign y13547 = ~n24066 ;
  assign y13548 = ~1'b0 ;
  assign y13549 = n24067 ;
  assign y13550 = ~1'b0 ;
  assign y13551 = ~1'b0 ;
  assign y13552 = ~1'b0 ;
  assign y13553 = n24074 ;
  assign y13554 = ~1'b0 ;
  assign y13555 = ~1'b0 ;
  assign y13556 = n24075 ;
  assign y13557 = ~n24076 ;
  assign y13558 = n24077 ;
  assign y13559 = ~1'b0 ;
  assign y13560 = n24080 ;
  assign y13561 = ~n4808 ;
  assign y13562 = ~1'b0 ;
  assign y13563 = n24081 ;
  assign y13564 = ~n24083 ;
  assign y13565 = n24084 ;
  assign y13566 = n24085 ;
  assign y13567 = n24089 ;
  assign y13568 = 1'b0 ;
  assign y13569 = n23644 ;
  assign y13570 = 1'b0 ;
  assign y13571 = ~n24090 ;
  assign y13572 = ~1'b0 ;
  assign y13573 = ~1'b0 ;
  assign y13574 = ~1'b0 ;
  assign y13575 = ~1'b0 ;
  assign y13576 = ~1'b0 ;
  assign y13577 = n24091 ;
  assign y13578 = n24092 ;
  assign y13579 = n24093 ;
  assign y13580 = ~1'b0 ;
  assign y13581 = ~n24095 ;
  assign y13582 = ~n24098 ;
  assign y13583 = ~1'b0 ;
  assign y13584 = 1'b0 ;
  assign y13585 = n24104 ;
  assign y13586 = ~n24109 ;
  assign y13587 = n24110 ;
  assign y13588 = ~1'b0 ;
  assign y13589 = n20560 ;
  assign y13590 = n4721 ;
  assign y13591 = n24115 ;
  assign y13592 = ~n24116 ;
  assign y13593 = ~1'b0 ;
  assign y13594 = ~n24119 ;
  assign y13595 = ~1'b0 ;
  assign y13596 = n24120 ;
  assign y13597 = ~n24121 ;
  assign y13598 = n24124 ;
  assign y13599 = ~n24126 ;
  assign y13600 = ~n24130 ;
  assign y13601 = ~n24132 ;
  assign y13602 = ~n24134 ;
  assign y13603 = n24138 ;
  assign y13604 = ~1'b0 ;
  assign y13605 = ~1'b0 ;
  assign y13606 = ~1'b0 ;
  assign y13607 = ~n24139 ;
  assign y13608 = n24140 ;
  assign y13609 = ~1'b0 ;
  assign y13610 = ~n24142 ;
  assign y13611 = 1'b0 ;
  assign y13612 = ~1'b0 ;
  assign y13613 = ~n24145 ;
  assign y13614 = n24146 ;
  assign y13615 = ~1'b0 ;
  assign y13616 = ~1'b0 ;
  assign y13617 = ~n24150 ;
  assign y13618 = n24152 ;
  assign y13619 = ~1'b0 ;
  assign y13620 = n24154 ;
  assign y13621 = n24156 ;
  assign y13622 = ~1'b0 ;
  assign y13623 = n24158 ;
  assign y13624 = ~1'b0 ;
  assign y13625 = ~1'b0 ;
  assign y13626 = ~n9901 ;
  assign y13627 = 1'b0 ;
  assign y13628 = ~n24161 ;
  assign y13629 = ~1'b0 ;
  assign y13630 = n24165 ;
  assign y13631 = n24166 ;
  assign y13632 = n24167 ;
  assign y13633 = ~n24172 ;
  assign y13634 = ~n24174 ;
  assign y13635 = ~n24175 ;
  assign y13636 = ~1'b0 ;
  assign y13637 = 1'b0 ;
  assign y13638 = n24176 ;
  assign y13639 = ~1'b0 ;
  assign y13640 = ~n24179 ;
  assign y13641 = ~n3429 ;
  assign y13642 = ~1'b0 ;
  assign y13643 = ~n24183 ;
  assign y13644 = ~n16788 ;
  assign y13645 = ~n10640 ;
  assign y13646 = ~n24186 ;
  assign y13647 = n24190 ;
  assign y13648 = ~n24191 ;
  assign y13649 = 1'b0 ;
  assign y13650 = ~1'b0 ;
  assign y13651 = ~n24192 ;
  assign y13652 = n24194 ;
  assign y13653 = ~1'b0 ;
  assign y13654 = n24198 ;
  assign y13655 = ~n24199 ;
  assign y13656 = ~n24201 ;
  assign y13657 = ~1'b0 ;
  assign y13658 = ~n24202 ;
  assign y13659 = ~1'b0 ;
  assign y13660 = n24203 ;
  assign y13661 = n24208 ;
  assign y13662 = n2945 ;
  assign y13663 = n24212 ;
  assign y13664 = ~1'b0 ;
  assign y13665 = ~1'b0 ;
  assign y13666 = n24213 ;
  assign y13667 = n24215 ;
  assign y13668 = n24217 ;
  assign y13669 = ~1'b0 ;
  assign y13670 = ~1'b0 ;
  assign y13671 = 1'b0 ;
  assign y13672 = n24218 ;
  assign y13673 = n24222 ;
  assign y13674 = n24227 ;
  assign y13675 = n24229 ;
  assign y13676 = n24232 ;
  assign y13677 = n24237 ;
  assign y13678 = ~1'b0 ;
  assign y13679 = ~n24239 ;
  assign y13680 = ~1'b0 ;
  assign y13681 = ~1'b0 ;
  assign y13682 = n24241 ;
  assign y13683 = ~1'b0 ;
  assign y13684 = ~n24244 ;
  assign y13685 = ~1'b0 ;
  assign y13686 = n24245 ;
  assign y13687 = n1370 ;
  assign y13688 = ~1'b0 ;
  assign y13689 = ~1'b0 ;
  assign y13690 = n24247 ;
  assign y13691 = ~n737 ;
  assign y13692 = ~n24248 ;
  assign y13693 = n24251 ;
  assign y13694 = ~1'b0 ;
  assign y13695 = ~1'b0 ;
  assign y13696 = ~n24254 ;
  assign y13697 = n24256 ;
  assign y13698 = n24257 ;
  assign y13699 = ~1'b0 ;
  assign y13700 = ~n24259 ;
  assign y13701 = ~n24263 ;
  assign y13702 = ~n24241 ;
  assign y13703 = ~n24268 ;
  assign y13704 = ~1'b0 ;
  assign y13705 = ~n24269 ;
  assign y13706 = ~1'b0 ;
  assign y13707 = ~1'b0 ;
  assign y13708 = n24272 ;
  assign y13709 = ~n24273 ;
  assign y13710 = n24276 ;
  assign y13711 = ~n3114 ;
  assign y13712 = ~1'b0 ;
  assign y13713 = n15341 ;
  assign y13714 = ~n11859 ;
  assign y13715 = ~n24280 ;
  assign y13716 = n24282 ;
  assign y13717 = ~1'b0 ;
  assign y13718 = ~n24284 ;
  assign y13719 = n20062 ;
  assign y13720 = ~n24285 ;
  assign y13721 = n24286 ;
  assign y13722 = ~n24288 ;
  assign y13723 = ~1'b0 ;
  assign y13724 = n19995 ;
  assign y13725 = ~n24289 ;
  assign y13726 = ~n24294 ;
  assign y13727 = ~1'b0 ;
  assign y13728 = ~n24296 ;
  assign y13729 = ~1'b0 ;
  assign y13730 = ~n24298 ;
  assign y13731 = ~1'b0 ;
  assign y13732 = ~1'b0 ;
  assign y13733 = ~1'b0 ;
  assign y13734 = ~1'b0 ;
  assign y13735 = ~1'b0 ;
  assign y13736 = ~n24299 ;
  assign y13737 = ~1'b0 ;
  assign y13738 = n24303 ;
  assign y13739 = ~1'b0 ;
  assign y13740 = n24307 ;
  assign y13741 = ~n24311 ;
  assign y13742 = n24317 ;
  assign y13743 = ~1'b0 ;
  assign y13744 = n24320 ;
  assign y13745 = ~n24322 ;
  assign y13746 = ~n24326 ;
  assign y13747 = n24327 ;
  assign y13748 = n24328 ;
  assign y13749 = n24331 ;
  assign y13750 = n24332 ;
  assign y13751 = ~1'b0 ;
endmodule
